Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_12x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A75: buffer std_logic
);
end x25_12x;

architecture x25_12x_behav of x25_12x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a768a,a772a,a773a,a774a,a778a,a779a,a783a,a784a,a785a,a786a,a790a,a791a,a795a,a796a,a797a,a801a,a802a,a806a,a807a,a808a,a809a,a810a,a814a,a815a,a819a,a820a,a821a,a825a,a826a,a830a,a831a,a832a,a833a,a837a,a838a,a842a,a843a,a844a,a848a,a849a,a853a,a854a,a855a,a856a,a857a,a858a,a862a,a863a,a867a,a868a,a869a,a873a,a874a,a878a,a879a,a880a,a881a,a885a,a886a,a890a,a891a,a892a,a896a,a897a,a901a,a902a,a903a,a904a,a905a,a909a,a910a,a914a,a915a,a916a,a920a,a921a,a925a,a926a,a927a,a928a,a932a,a933a,a937a,a938a,a939a,a943a,a944a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a958a,a959a,a963a,a964a,a965a,a969a,a970a,a974a,a975a,a976a,a977a,a981a,a982a,a986a,a987a,a988a,a992a,a993a,a997a,a998a,a999a,a1000a,a1001a,a1005a,a1006a,a1010a,a1011a,a1012a,a1016a,a1017a,a1021a,a1022a,a1023a,a1024a,a1028a,a1029a,a1033a,a1034a,a1035a,a1039a,a1040a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1053a,a1054a,a1058a,a1059a,a1060a,a1064a,a1065a,a1069a,a1070a,a1071a,a1072a,a1076a,a1077a,a1081a,a1082a,a1083a,a1087a,a1088a,a1092a,a1093a,a1094a,a1095a,a1096a,a1100a,a1101a,a1105a,a1106a,a1107a,a1111a,a1112a,a1116a,a1117a,a1118a,a1119a,a1123a,a1124a,a1128a,a1129a,a1130a,a1134a,a1135a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1149a,a1153a,a1154a,a1155a,a1159a,a1160a,a1164a,a1165a,a1166a,a1167a,a1171a,a1172a,a1176a,a1177a,a1178a,a1182a,a1183a,a1187a,a1188a,a1189a,a1190a,a1191a,a1195a,a1196a,a1200a,a1201a,a1202a,a1206a,a1207a,a1211a,a1212a,a1213a,a1214a,a1218a,a1219a,a1223a,a1224a,a1225a,a1229a,a1230a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1243a,a1244a,a1248a,a1249a,a1250a,a1254a,a1255a,a1259a,a1260a,a1261a,a1262a,a1266a,a1267a,a1271a,a1272a,a1273a,a1277a,a1278a,a1282a,a1283a,a1284a,a1285a,a1286a,a1290a,a1291a,a1295a,a1296a,a1297a,a1301a,a1302a,a1306a,a1307a,a1308a,a1309a,a1313a,a1314a,a1318a,a1319a,a1320a,a1324a,a1325a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1339a,a1340a,a1344a,a1345a,a1346a,a1350a,a1351a,a1355a,a1356a,a1357a,a1358a,a1362a,a1363a,a1367a,a1368a,a1369a,a1373a,a1374a,a1378a,a1379a,a1380a,a1381a,a1382a,a1386a,a1387a,a1391a,a1392a,a1393a,a1397a,a1398a,a1402a,a1403a,a1404a,a1405a,a1409a,a1410a,a1414a,a1415a,a1416a,a1420a,a1421a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1434a,a1435a,a1439a,a1440a,a1441a,a1445a,a1446a,a1450a,a1451a,a1452a,a1453a,a1457a,a1458a,a1462a,a1463a,a1464a,a1468a,a1469a,a1473a,a1474a,a1475a,a1476a,a1477a,a1481a,a1482a,a1486a,a1487a,a1488a,a1492a,a1493a,a1497a,a1498a,a1499a,a1500a,a1504a,a1505a,a1509a,a1510a,a1511a,a1515a,a1516a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1531a,a1535a,a1536a,a1537a,a1541a,a1542a,a1546a,a1547a,a1548a,a1549a,a1553a,a1554a,a1558a,a1559a,a1560a,a1564a,a1565a,a1569a,a1570a,a1571a,a1572a,a1573a,a1577a,a1578a,a1582a,a1583a,a1584a,a1588a,a1589a,a1593a,a1594a,a1595a,a1596a,a1600a,a1601a,a1605a,a1606a,a1607a,a1611a,a1612a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1625a,a1626a,a1630a,a1631a,a1632a,a1636a,a1637a,a1641a,a1642a,a1643a,a1644a,a1648a,a1649a,a1653a,a1654a,a1655a,a1659a,a1660a,a1664a,a1665a,a1666a,a1667a,a1668a,a1672a,a1673a,a1677a,a1678a,a1679a,a1683a,a1684a,a1688a,a1689a,a1690a,a1691a,a1695a,a1696a,a1700a,a1701a,a1702a,a1706a,a1707a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1721a,a1722a,a1726a,a1727a,a1728a,a1732a,a1733a,a1737a,a1738a,a1739a,a1740a,a1744a,a1745a,a1749a,a1750a,a1751a,a1755a,a1756a,a1760a,a1761a,a1762a,a1763a,a1764a,a1768a,a1769a,a1773a,a1774a,a1775a,a1779a,a1780a,a1784a,a1785a,a1786a,a1787a,a1791a,a1792a,a1796a,a1797a,a1798a,a1802a,a1803a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1816a,a1817a,a1821a,a1822a,a1823a,a1827a,a1828a,a1832a,a1833a,a1834a,a1835a,a1839a,a1840a,a1844a,a1845a,a1846a,a1850a,a1851a,a1855a,a1856a,a1857a,a1858a,a1859a,a1863a,a1864a,a1868a,a1869a,a1870a,a1874a,a1875a,a1879a,a1880a,a1881a,a1882a,a1886a,a1887a,a1891a,a1892a,a1893a,a1897a,a1898a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1913a,a1914a,a1918a,a1919a,a1920a,a1924a,a1925a,a1929a,a1930a,a1931a,a1932a,a1936a,a1937a,a1941a,a1942a,a1943a,a1947a,a1948a,a1952a,a1953a,a1954a,a1955a,a1956a,a1960a,a1961a,a1965a,a1966a,a1967a,a1971a,a1972a,a1976a,a1977a,a1978a,a1979a,a1983a,a1984a,a1988a,a1989a,a1990a,a1994a,a1995a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2008a,a2009a,a2013a,a2014a,a2015a,a2019a,a2020a,a2024a,a2025a,a2026a,a2027a,a2031a,a2032a,a2036a,a2037a,a2038a,a2042a,a2043a,a2047a,a2048a,a2049a,a2050a,a2051a,a2055a,a2056a,a2060a,a2061a,a2062a,a2066a,a2067a,a2071a,a2072a,a2073a,a2074a,a2078a,a2079a,a2083a,a2084a,a2085a,a2089a,a2090a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2104a,a2105a,a2109a,a2110a,a2111a,a2115a,a2116a,a2120a,a2121a,a2122a,a2123a,a2127a,a2128a,a2132a,a2133a,a2134a,a2138a,a2139a,a2143a,a2144a,a2145a,a2146a,a2147a,a2151a,a2152a,a2156a,a2157a,a2158a,a2162a,a2163a,a2167a,a2168a,a2169a,a2170a,a2174a,a2175a,a2179a,a2180a,a2181a,a2185a,a2186a,a2190a,a2191a,a2192a,a2193a,a2194a,a2195a,a2199a,a2200a,a2204a,a2205a,a2206a,a2210a,a2211a,a2215a,a2216a,a2217a,a2218a,a2222a,a2223a,a2227a,a2228a,a2229a,a2233a,a2234a,a2238a,a2239a,a2240a,a2241a,a2242a,a2246a,a2247a,a2251a,a2252a,a2253a,a2257a,a2258a,a2262a,a2263a,a2264a,a2265a,a2269a,a2270a,a2274a,a2275a,a2276a,a2280a,a2281a,a2285a,a2286a,a2287a,a2288a,a2289a,a2290a,a2291a,a2292a,a2293a,a2296a,a2299a,a2302a,a2305a,a2308a,a2312a,a2313a,a2316a,a2320a,a2321a,a2324a,a2328a,a2329a,a2332a,a2336a,a2337a,a2340a,a2344a,a2345a,a2349a,a2350a,a2354a,a2355a,a2359a,a2360a,a2364a,a2365a,a2369a,a2370a,a2374a,a2375a,a2379a,a2380a,a2384a,a2385a,a2389a,a2390a,a2394a,a2395a,a2399a,a2400a,a2404a,a2405a,a2409a,a2410a,a2414a,a2415a,a2419a,a2420a,a2424a,a2425a,a2429a,a2430a,a2434a,a2435a,a2439a,a2440a,a2444a,a2445a,a2449a,a2450a,a2453a,a2456a,a2457a,a2461a,a2462a,a2465a,a2468a,a2469a,a2473a,a2474a,a2477a,a2480a,a2481a,a2485a,a2486a,a2489a,a2492a,a2493a,a2497a,a2498a,a2501a,a2504a,a2505a,a2509a,a2510a,a2513a,a2516a,a2517a,a2521a,a2522a,a2525a,a2528a,a2529a,a2533a,a2534a,a2537a,a2540a,a2541a,a2545a,a2546a,a2549a,a2552a,a2553a,a2557a,a2558a,a2561a,a2564a,a2565a,a2569a,a2570a,a2573a,a2576a,a2577a,a2581a,a2582a,a2585a,a2588a,a2589a,a2593a,a2594a,a2597a,a2600a,a2601a,a2605a,a2606a,a2609a,a2612a,a2613a,a2617a,a2618a,a2621a,a2624a,a2625a,a2629a,a2630a,a2633a,a2636a,a2637a,a2641a,a2642a,a2645a,a2648a,a2649a,a2653a,a2654a,a2657a,a2660a,a2661a,a2665a,a2666a,a2669a,a2672a,a2673a,a2677a,a2678a,a2681a,a2684a,a2685a,a2689a,a2690a,a2693a,a2696a,a2697a,a2701a,a2702a,a2705a,a2708a,a2709a,a2713a,a2714a,a2717a,a2720a,a2721a,a2725a,a2726a,a2729a,a2732a,a2733a,a2737a,a2738a,a2741a,a2744a,a2745a,a2749a,a2750a,a2753a,a2756a,a2757a,a2761a,a2762a,a2765a,a2768a,a2769a,a2773a,a2774a,a2777a,a2780a,a2781a,a2784a,a2787a,a2788a,a2791a,a2794a,a2795a,a2798a,a2801a,a2802a,a2805a,a2808a,a2809a,a2812a,a2815a,a2816a,a2819a,a2822a,a2823a,a2826a,a2829a,a2830a,a2833a,a2836a,a2837a,a2840a,a2843a,a2844a,a2847a,a2850a,a2851a,a2854a,a2857a,a2858a,a2861a,a2864a,a2865a,a2868a,a2871a,a2872a,a2875a,a2878a,a2879a,a2882a,a2885a,a2886a,a2889a,a2892a,a2893a,a2896a,a2899a,a2900a,a2903a,a2906a,a2907a,a2910a,a2913a,a2914a,a2917a,a2920a,a2921a,a2924a,a2927a,a2928a,a2931a,a2934a,a2935a,a2938a,a2941a,a2942a,a2945a,a2948a,a2949a,a2952a,a2955a,a2956a,a2959a,a2962a,a2963a,a2966a,a2969a,a2970a,a2973a,a2976a,a2977a,a2980a,a2983a,a2984a,a2987a,a2990a,a2991a,a2994a,a2997a,a2998a,a3001a,a3004a,a3005a,a3008a,a3011a,a3012a,a3015a,a3018a,a3019a,a3022a,a3025a,a3026a,a3029a,a3032a,a3033a,a3036a,a3039a,a3040a,a3043a,a3046a,a3047a,a3050a,a3053a,a3054a,a3057a,a3060a,a3061a,a3064a,a3067a,a3068a,a3071a,a3074a,a3075a,a3078a,a3081a,a3082a,a3085a,a3088a,a3089a,a3092a,a3095a,a3096a,a3099a,a3102a,a3103a,a3106a,a3109a,a3110a,a3113a,a3116a,a3117a,a3120a,a3123a,a3124a,a3127a,a3130a,a3131a,a3134a,a3137a,a3138a,a3141a,a3144a,a3145a,a3148a,a3151a,a3152a,a3155a,a3158a,a3159a,a3162a,a3165a,a3166a,a3169a,a3172a,a3173a,a3176a,a3179a,a3180a,a3183a,a3186a,a3187a,a3190a,a3193a,a3194a,a3197a,a3200a,a3201a,a3204a,a3207a,a3208a,a3211a,a3214a,a3215a,a3218a,a3221a,a3222a,a3225a,a3228a,a3229a,a3232a,a3235a,a3236a,a3239a,a3242a,a3243a,a3246a,a3249a,a3250a,a3253a,a3256a,a3257a,a3260a,a3263a,a3264a,a3267a,a3270a,a3271a,a3274a,a3277a,a3278a,a3281a,a3284a,a3285a,a3288a,a3291a,a3292a,a3295a,a3298a,a3299a,a3302a,a3305a,a3306a,a3309a,a3312a,a3313a,a3316a,a3319a,a3320a,a3323a,a3326a,a3327a,a3330a,a3333a,a3334a,a3337a,a3340a,a3341a,a3344a,a3347a,a3348a,a3351a,a3354a,a3355a,a3358a,a3361a,a3362a,a3365a,a3368a,a3369a,a3372a,a3375a,a3376a,a3379a,a3382a,a3383a,a3386a,a3389a,a3390a,a3393a,a3396a,a3397a,a3400a,a3403a,a3404a,a3407a,a3410a,a3411a,a3414a,a3417a,a3418a,a3421a,a3424a,a3425a,a3428a,a3431a,a3432a,a3435a,a3438a,a3439a,a3442a,a3445a,a3446a,a3449a,a3452a,a3453a,a3456a,a3459a,a3460a,a3463a,a3466a,a3467a,a3470a,a3473a,a3474a,a3477a,a3480a,a3481a,a3484a,a3487a,a3488a,a3491a,a3494a,a3495a,a3498a,a3501a,a3502a,a3505a,a3508a,a3509a,a3512a,a3515a,a3516a,a3519a,a3522a,a3523a,a3526a,a3529a,a3530a,a3533a,a3536a,a3537a,a3540a,a3543a,a3544a,a3547a,a3550a,a3551a,a3554a,a3557a,a3558a,a3561a,a3564a,a3565a,a3568a,a3571a,a3572a,a3575a,a3578a,a3579a,a3582a,a3585a,a3586a,a3589a,a3592a,a3593a,a3596a,a3599a,a3600a,a3603a,a3606a,a3607a,a3610a,a3613a,a3614a,a3617a,a3620a,a3621a,a3624a,a3627a,a3628a,a3631a,a3634a,a3635a,a3638a,a3641a,a3642a,a3645a,a3648a,a3649a,a3652a,a3655a,a3656a,a3659a,a3662a,a3663a,a3666a,a3669a,a3670a,a3673a,a3676a,a3677a,a3680a,a3683a,a3684a,a3687a,a3690a,a3691a,a3694a,a3697a,a3698a,a3701a,a3704a,a3705a,a3708a,a3711a,a3712a,a3715a,a3718a,a3719a,a3722a,a3725a,a3726a,a3729a,a3732a,a3733a,a3736a,a3739a,a3740a,a3743a,a3746a,a3747a,a3750a,a3753a,a3754a,a3757a,a3760a,a3761a,a3764a,a3767a,a3768a,a3771a,a3774a,a3775a,a3778a,a3781a,a3782a,a3785a,a3788a,a3789a,a3792a,a3795a,a3796a,a3799a,a3802a,a3803a,a3806a,a3809a,a3810a,a3813a,a3816a,a3817a,a3820a,a3823a,a3824a,a3827a,a3830a,a3831a,a3834a,a3837a,a3838a,a3841a,a3844a,a3845a,a3848a,a3851a,a3852a,a3855a,a3858a,a3859a,a3862a,a3865a,a3866a,a3869a,a3872a,a3873a,a3876a,a3879a,a3880a,a3883a,a3886a,a3887a,a3890a,a3893a,a3894a,a3897a,a3900a,a3901a,a3904a,a3907a,a3908a,a3911a,a3914a,a3915a,a3918a,a3921a,a3922a,a3925a,a3928a,a3929a,a3932a,a3935a,a3936a,a3939a,a3942a,a3943a,a3946a,a3949a,a3950a,a3953a,a3956a,a3957a,a3960a,a3963a,a3964a,a3967a,a3971a,a3972a,a3973a,a3976a,a3979a,a3980a,a3983a,a3987a,a3988a,a3989a,a3992a,a3995a,a3996a,a3999a,a4003a,a4004a,a4005a,a4008a,a4011a,a4012a,a4015a,a4019a,a4020a,a4021a,a4024a,a4027a,a4028a,a4031a,a4035a,a4036a,a4037a,a4040a,a4043a,a4044a,a4047a,a4051a,a4052a,a4053a,a4056a,a4059a,a4060a,a4063a,a4067a,a4068a,a4069a,a4072a,a4075a,a4076a,a4079a,a4083a,a4084a,a4085a,a4088a,a4091a,a4092a,a4095a,a4099a,a4100a,a4101a,a4104a,a4107a,a4108a,a4111a,a4115a,a4116a,a4117a,a4120a,a4123a,a4124a,a4127a,a4131a,a4132a,a4133a,a4136a,a4139a,a4140a,a4143a,a4147a,a4148a,a4149a,a4152a,a4155a,a4156a,a4159a,a4163a,a4164a,a4165a,a4168a,a4171a,a4172a,a4175a,a4179a,a4180a,a4181a,a4184a,a4187a,a4188a,a4191a,a4195a,a4196a,a4197a,a4200a,a4203a,a4204a,a4207a,a4211a,a4212a,a4213a,a4216a,a4219a,a4220a,a4223a,a4227a,a4228a,a4229a,a4232a,a4235a,a4236a,a4239a,a4243a,a4244a,a4245a,a4248a,a4251a,a4252a,a4255a,a4259a,a4260a,a4261a,a4264a,a4267a,a4268a,a4271a,a4275a,a4276a,a4277a,a4280a,a4283a,a4284a,a4287a,a4291a,a4292a,a4293a,a4296a,a4299a,a4300a,a4303a,a4307a,a4308a,a4309a,a4312a,a4315a,a4316a,a4319a,a4323a,a4324a,a4325a,a4328a,a4331a,a4332a,a4335a,a4339a,a4340a,a4341a,a4344a,a4347a,a4348a,a4351a,a4355a,a4356a,a4357a,a4360a,a4363a,a4364a,a4367a,a4371a,a4372a,a4373a,a4376a,a4379a,a4380a,a4383a,a4387a,a4388a,a4389a,a4392a,a4395a,a4396a,a4399a,a4403a,a4404a,a4405a,a4408a,a4411a,a4412a,a4415a,a4419a,a4420a,a4421a,a4424a,a4427a,a4428a,a4431a,a4435a,a4436a,a4437a,a4440a,a4443a,a4444a,a4447a,a4451a,a4452a,a4453a,a4456a,a4459a,a4460a,a4463a,a4467a,a4468a,a4469a,a4472a,a4475a,a4476a,a4479a,a4483a,a4484a,a4485a,a4488a,a4491a,a4492a,a4495a,a4499a,a4500a,a4501a,a4504a,a4507a,a4508a,a4511a,a4515a,a4516a,a4517a,a4520a,a4523a,a4524a,a4527a,a4531a,a4532a,a4533a,a4536a,a4539a,a4540a,a4543a,a4547a,a4548a,a4549a,a4552a,a4555a,a4556a,a4559a,a4563a,a4564a,a4565a,a4568a,a4571a,a4572a,a4575a,a4579a,a4580a,a4581a,a4584a,a4587a,a4588a,a4591a,a4595a,a4596a,a4597a,a4600a,a4603a,a4604a,a4607a,a4611a,a4612a,a4613a,a4616a,a4619a,a4620a,a4623a,a4627a,a4628a,a4629a,a4632a,a4635a,a4636a,a4639a,a4643a,a4644a,a4645a,a4648a,a4651a,a4652a,a4655a,a4659a,a4660a,a4661a,a4664a,a4667a,a4668a,a4671a,a4675a,a4676a,a4677a,a4680a,a4683a,a4684a,a4687a,a4691a,a4692a,a4693a,a4696a,a4699a,a4700a,a4703a,a4707a,a4708a,a4709a,a4712a,a4715a,a4716a,a4719a,a4723a,a4724a,a4725a,a4728a,a4731a,a4732a,a4735a,a4739a,a4740a,a4741a,a4744a,a4747a,a4748a,a4751a,a4755a,a4756a,a4757a,a4760a,a4763a,a4764a,a4767a,a4771a,a4772a,a4773a,a4776a,a4779a,a4780a,a4783a,a4787a,a4788a,a4789a,a4792a,a4795a,a4796a,a4799a,a4803a,a4804a,a4805a,a4808a,a4811a,a4812a,a4815a,a4819a,a4820a,a4821a,a4824a,a4827a,a4828a,a4831a,a4835a,a4836a,a4837a,a4840a,a4843a,a4844a,a4847a,a4851a,a4852a,a4853a,a4856a,a4859a,a4860a,a4863a,a4867a,a4868a,a4869a,a4872a,a4875a,a4876a,a4879a,a4883a,a4884a,a4885a,a4888a,a4891a,a4892a,a4895a,a4899a,a4900a,a4901a,a4904a,a4907a,a4908a,a4911a,a4915a,a4916a,a4917a,a4920a,a4923a,a4924a,a4927a,a4931a,a4932a,a4933a,a4936a,a4939a,a4940a,a4943a,a4947a,a4948a,a4949a,a4952a,a4955a,a4956a,a4959a,a4963a,a4964a,a4965a,a4968a,a4971a,a4972a,a4975a,a4979a,a4980a,a4981a,a4984a,a4987a,a4988a,a4991a,a4995a,a4996a,a4997a,a5000a,a5003a,a5004a,a5007a,a5011a,a5012a,a5013a,a5016a,a5019a,a5020a,a5023a,a5027a,a5028a,a5029a,a5032a,a5035a,a5036a,a5039a,a5043a,a5044a,a5045a,a5048a,a5051a,a5052a,a5055a,a5059a,a5060a,a5061a,a5064a,a5067a,a5068a,a5071a,a5075a,a5076a,a5077a,a5080a,a5083a,a5084a,a5087a,a5091a,a5092a,a5093a,a5096a,a5099a,a5100a,a5103a,a5107a,a5108a,a5109a,a5112a,a5115a,a5116a,a5119a,a5123a,a5124a,a5125a,a5128a,a5131a,a5132a,a5135a,a5139a,a5140a,a5141a,a5144a,a5147a,a5148a,a5151a,a5155a,a5156a,a5157a,a5160a,a5163a,a5164a,a5167a,a5171a,a5172a,a5173a,a5176a,a5179a,a5180a,a5183a,a5187a,a5188a,a5189a,a5192a,a5195a,a5196a,a5199a,a5203a,a5204a,a5205a,a5208a,a5211a,a5212a,a5215a,a5219a,a5220a,a5221a,a5224a,a5227a,a5228a,a5231a,a5235a,a5236a,a5237a,a5240a,a5243a,a5244a,a5247a,a5251a,a5252a,a5253a,a5256a,a5259a,a5260a,a5263a,a5267a,a5268a,a5269a,a5272a,a5275a,a5276a,a5279a,a5283a,a5284a,a5285a,a5288a,a5291a,a5292a,a5295a,a5299a,a5300a,a5301a,a5304a,a5307a,a5308a,a5311a,a5315a,a5316a,a5317a,a5320a,a5323a,a5324a,a5327a,a5331a,a5332a,a5333a,a5336a,a5339a,a5340a,a5343a,a5347a,a5348a,a5349a,a5352a,a5355a,a5356a,a5359a,a5363a,a5364a,a5365a,a5368a,a5371a,a5372a,a5375a,a5379a,a5380a,a5381a,a5384a,a5387a,a5388a,a5391a,a5395a,a5396a,a5397a,a5400a,a5403a,a5404a,a5407a,a5411a,a5412a,a5413a,a5416a,a5419a,a5420a,a5423a,a5427a,a5428a,a5429a,a5432a,a5435a,a5436a,a5439a,a5443a,a5444a,a5445a,a5448a,a5451a,a5452a,a5455a,a5459a,a5460a,a5461a,a5464a,a5467a,a5468a,a5471a,a5475a,a5476a,a5477a,a5480a,a5483a,a5484a,a5487a,a5491a,a5492a,a5493a,a5496a,a5499a,a5500a,a5503a,a5507a,a5508a,a5509a,a5512a,a5515a,a5516a,a5519a,a5523a,a5524a,a5525a,a5528a,a5531a,a5532a,a5535a,a5539a,a5540a,a5541a,a5544a,a5547a,a5548a,a5551a,a5555a,a5556a,a5557a,a5560a,a5563a,a5564a,a5567a,a5571a,a5572a,a5573a,a5576a,a5579a,a5580a,a5583a,a5587a,a5588a,a5589a,a5592a,a5595a,a5596a,a5599a,a5603a,a5604a,a5605a,a5608a,a5611a,a5612a,a5615a,a5619a,a5620a,a5621a,a5624a,a5627a,a5628a,a5631a,a5635a,a5636a,a5637a,a5640a,a5643a,a5644a,a5647a,a5651a,a5652a,a5653a,a5656a,a5659a,a5660a,a5663a,a5667a,a5668a,a5669a,a5672a,a5675a,a5676a,a5679a,a5683a,a5684a,a5685a,a5688a,a5691a,a5692a,a5695a,a5699a,a5700a,a5701a,a5704a,a5707a,a5708a,a5711a,a5715a,a5716a,a5717a,a5720a,a5723a,a5724a,a5727a,a5731a,a5732a,a5733a,a5736a,a5739a,a5740a,a5743a,a5747a,a5748a,a5749a,a5752a,a5755a,a5756a,a5759a,a5763a,a5764a,a5765a,a5768a,a5771a,a5772a,a5775a,a5779a,a5780a,a5781a,a5784a,a5787a,a5788a,a5791a,a5795a,a5796a,a5797a,a5800a,a5803a,a5804a,a5807a,a5811a,a5812a,a5813a,a5816a,a5819a,a5820a,a5823a,a5827a,a5828a,a5829a,a5832a,a5835a,a5836a,a5839a,a5843a,a5844a,a5845a,a5848a,a5851a,a5852a,a5855a,a5859a,a5860a,a5861a,a5864a,a5867a,a5868a,a5871a,a5875a,a5876a,a5877a,a5880a,a5883a,a5884a,a5887a,a5891a,a5892a,a5893a,a5896a,a5899a,a5900a,a5903a,a5907a,a5908a,a5909a,a5912a,a5915a,a5916a,a5919a,a5923a,a5924a,a5925a,a5928a,a5931a,a5932a,a5935a,a5939a,a5940a,a5941a,a5944a,a5947a,a5948a,a5951a,a5955a,a5956a,a5957a,a5960a,a5963a,a5964a,a5967a,a5971a,a5972a,a5973a,a5976a,a5979a,a5980a,a5983a,a5987a,a5988a,a5989a,a5992a,a5995a,a5996a,a5999a,a6003a,a6004a,a6005a,a6008a,a6011a,a6012a,a6015a,a6019a,a6020a,a6021a,a6024a,a6027a,a6028a,a6031a,a6035a,a6036a,a6037a,a6040a,a6043a,a6044a,a6047a,a6051a,a6052a,a6053a,a6056a,a6059a,a6060a,a6063a,a6067a,a6068a,a6069a,a6072a,a6075a,a6076a,a6079a,a6083a,a6084a,a6085a,a6088a,a6091a,a6092a,a6095a,a6099a,a6100a,a6101a,a6104a,a6107a,a6108a,a6111a,a6115a,a6116a,a6117a,a6120a,a6123a,a6124a,a6127a,a6131a,a6132a,a6133a,a6136a,a6139a,a6140a,a6143a,a6147a,a6148a,a6149a,a6152a,a6155a,a6156a,a6159a,a6163a,a6164a,a6165a,a6168a,a6171a,a6172a,a6175a,a6179a,a6180a,a6181a,a6184a,a6187a,a6188a,a6191a,a6195a,a6196a,a6197a,a6200a,a6203a,a6204a,a6207a,a6211a,a6212a,a6213a,a6216a,a6219a,a6220a,a6223a,a6227a,a6228a,a6229a,a6232a,a6235a,a6236a,a6239a,a6243a,a6244a,a6245a,a6248a,a6251a,a6252a,a6255a,a6259a,a6260a,a6261a,a6264a,a6267a,a6268a,a6271a,a6275a,a6276a,a6277a,a6280a,a6283a,a6284a,a6287a,a6291a,a6292a,a6293a,a6296a,a6299a,a6300a,a6303a,a6307a,a6308a,a6309a,a6312a,a6315a,a6316a,a6319a,a6323a,a6324a,a6325a,a6328a,a6331a,a6332a,a6335a,a6339a,a6340a,a6341a,a6344a,a6347a,a6348a,a6351a,a6355a,a6356a,a6357a,a6360a,a6363a,a6364a,a6367a,a6371a,a6372a,a6373a,a6376a,a6379a,a6380a,a6383a,a6387a,a6388a,a6389a,a6392a,a6395a,a6396a,a6399a,a6403a,a6404a,a6405a,a6408a,a6411a,a6412a,a6415a,a6419a,a6420a,a6421a,a6424a,a6427a,a6428a,a6431a,a6435a,a6436a,a6437a,a6440a,a6443a,a6444a,a6447a,a6451a,a6452a,a6453a,a6456a,a6459a,a6460a,a6463a,a6467a,a6468a,a6469a,a6472a,a6475a,a6476a,a6479a,a6483a,a6484a,a6485a,a6488a,a6491a,a6492a,a6495a,a6499a,a6500a,a6501a,a6504a,a6507a,a6508a,a6511a,a6515a,a6516a,a6517a,a6520a,a6523a,a6524a,a6527a,a6531a,a6532a,a6533a,a6536a,a6539a,a6540a,a6543a,a6547a,a6548a,a6549a,a6552a,a6555a,a6556a,a6559a,a6563a,a6564a,a6565a,a6568a,a6571a,a6572a,a6575a,a6579a,a6580a,a6581a,a6584a,a6588a,a6589a,a6590a,a6593a,a6597a,a6598a,a6599a,a6602a,a6606a,a6607a,a6608a,a6611a,a6615a,a6616a,a6617a,a6620a,a6624a,a6625a,a6626a,a6629a,a6633a,a6634a,a6635a,a6638a,a6642a,a6643a,a6644a,a6647a,a6651a,a6652a,a6653a,a6656a,a6660a,a6661a,a6662a,a6665a,a6669a,a6670a,a6671a,a6674a,a6678a,a6679a,a6680a,a6683a,a6687a,a6688a,a6689a,a6692a,a6696a,a6697a,a6698a,a6701a,a6705a,a6706a,a6707a,a6710a,a6714a,a6715a,a6716a,a6719a,a6723a,a6724a,a6725a,a6728a,a6732a,a6733a,a6734a,a6737a,a6741a,a6742a,a6743a,a6746a,a6750a,a6751a,a6752a,a6755a,a6759a,a6760a,a6761a,a6764a,a6768a,a6769a,a6770a,a6773a,a6777a,a6778a,a6779a,a6782a,a6786a,a6787a,a6788a,a6791a,a6795a,a6796a,a6797a,a6800a,a6804a,a6805a,a6806a,a6809a,a6813a,a6814a,a6815a,a6818a,a6822a,a6823a,a6824a,a6827a,a6831a,a6832a,a6833a,a6836a,a6840a,a6841a,a6842a,a6845a,a6849a,a6850a,a6851a,a6854a,a6858a,a6859a,a6860a,a6863a,a6867a,a6868a,a6869a,a6872a,a6876a,a6877a,a6878a,a6881a,a6885a,a6886a,a6887a,a6890a,a6894a,a6895a,a6896a,a6899a,a6903a,a6904a,a6905a,a6908a,a6912a,a6913a,a6914a,a6917a,a6921a,a6922a,a6923a,a6926a,a6930a,a6931a,a6932a,a6935a,a6939a,a6940a,a6941a,a6944a,a6948a,a6949a,a6950a,a6953a,a6957a,a6958a,a6959a,a6962a,a6966a,a6967a,a6968a,a6971a,a6975a,a6976a,a6977a,a6980a,a6984a,a6985a,a6986a,a6989a,a6993a,a6994a,a6995a,a6998a,a7002a,a7003a,a7004a,a7007a,a7011a,a7012a,a7013a,a7016a,a7020a,a7021a,a7022a,a7025a,a7029a,a7030a,a7031a,a7034a,a7038a,a7039a,a7040a,a7043a,a7047a,a7048a,a7049a,a7052a,a7056a,a7057a,a7058a,a7061a,a7065a,a7066a,a7067a,a7070a,a7074a,a7075a,a7076a,a7079a,a7083a,a7084a,a7085a,a7088a,a7092a,a7093a,a7094a,a7097a,a7101a,a7102a,a7103a,a7106a,a7110a,a7111a,a7112a,a7115a,a7119a,a7120a,a7121a,a7124a,a7128a,a7129a,a7130a,a7133a,a7137a,a7138a,a7139a,a7142a,a7146a,a7147a,a7148a,a7151a,a7155a,a7156a,a7157a,a7160a,a7164a,a7165a,a7166a,a7169a,a7173a,a7174a,a7175a,a7178a,a7182a,a7183a,a7184a,a7187a,a7191a,a7192a,a7193a,a7196a,a7200a,a7201a,a7202a,a7205a,a7209a,a7210a,a7211a,a7214a,a7218a,a7219a,a7220a,a7223a,a7227a,a7228a,a7229a,a7232a,a7236a,a7237a,a7238a,a7241a,a7245a,a7246a,a7247a,a7250a,a7254a,a7255a,a7256a,a7259a,a7263a,a7264a,a7265a,a7268a,a7272a,a7273a,a7274a,a7277a,a7281a,a7282a,a7283a,a7286a,a7290a,a7291a,a7292a,a7295a,a7299a,a7300a,a7301a,a7304a,a7308a,a7309a,a7310a,a7313a,a7317a,a7318a,a7319a,a7322a,a7326a,a7327a,a7328a,a7331a,a7335a,a7336a,a7337a,a7340a,a7344a,a7345a,a7346a,a7349a,a7353a,a7354a,a7355a,a7358a,a7362a,a7363a,a7364a,a7367a,a7371a,a7372a,a7373a,a7376a,a7380a,a7381a,a7382a,a7385a,a7389a,a7390a,a7391a,a7394a,a7398a,a7399a,a7400a,a7403a,a7407a,a7408a,a7409a,a7412a,a7416a,a7417a,a7418a,a7421a,a7425a,a7426a,a7427a,a7430a,a7434a,a7435a,a7436a,a7439a,a7443a,a7444a,a7445a,a7448a,a7452a,a7453a,a7454a,a7457a,a7461a,a7462a,a7463a,a7466a,a7470a,a7471a,a7472a,a7475a,a7479a,a7480a,a7481a,a7484a,a7488a,a7489a,a7490a,a7493a,a7497a,a7498a,a7499a,a7502a,a7506a,a7507a,a7508a,a7511a,a7515a,a7516a,a7517a,a7520a,a7524a,a7525a,a7526a,a7529a,a7533a,a7534a,a7535a,a7538a,a7542a,a7543a,a7544a,a7547a,a7551a,a7552a,a7553a,a7556a,a7560a,a7561a,a7562a,a7565a,a7569a,a7570a,a7571a,a7574a,a7578a,a7579a,a7580a,a7583a,a7587a,a7588a,a7589a,a7592a,a7596a,a7597a,a7598a,a7601a,a7605a,a7606a,a7607a,a7610a,a7614a,a7615a,a7616a,a7619a,a7623a,a7624a,a7625a,a7628a,a7632a,a7633a,a7634a,a7637a,a7641a,a7642a,a7643a,a7646a,a7650a,a7651a,a7652a,a7655a,a7659a,a7660a,a7661a,a7664a,a7668a,a7669a,a7670a,a7673a,a7677a,a7678a,a7679a,a7682a,a7686a,a7687a,a7688a,a7691a,a7695a,a7696a,a7697a,a7700a,a7704a,a7705a,a7706a,a7709a,a7713a,a7714a,a7715a,a7718a,a7722a,a7723a,a7724a,a7727a,a7731a,a7732a,a7733a,a7736a,a7740a,a7741a,a7742a,a7745a,a7749a,a7750a,a7751a,a7754a,a7758a,a7759a,a7760a,a7763a,a7767a,a7768a,a7769a,a7772a,a7776a,a7777a,a7778a,a7781a,a7785a,a7786a,a7787a,a7790a,a7794a,a7795a,a7796a,a7799a,a7803a,a7804a,a7805a,a7808a,a7812a,a7813a,a7814a,a7817a,a7821a,a7822a,a7823a,a7826a,a7830a,a7831a,a7832a,a7835a,a7839a,a7840a,a7841a,a7844a,a7848a,a7849a,a7850a,a7853a,a7857a,a7858a,a7859a,a7862a,a7866a,a7867a,a7868a,a7871a,a7875a,a7876a,a7877a,a7880a,a7884a,a7885a,a7886a,a7889a,a7893a,a7894a,a7895a,a7898a,a7902a,a7903a,a7904a,a7907a,a7911a,a7912a,a7913a,a7916a,a7920a,a7921a,a7922a,a7925a,a7929a,a7930a,a7931a,a7934a,a7938a,a7939a,a7940a,a7943a,a7947a,a7948a,a7949a,a7952a,a7956a,a7957a,a7958a,a7961a,a7965a,a7966a,a7967a,a7970a,a7974a,a7975a,a7976a,a7979a,a7983a,a7984a,a7985a,a7988a,a7992a,a7993a,a7994a,a7997a,a8001a,a8002a,a8003a,a8006a,a8010a,a8011a,a8012a,a8015a,a8019a,a8020a,a8021a,a8024a,a8028a,a8029a,a8030a,a8033a,a8037a,a8038a,a8039a,a8042a,a8046a,a8047a,a8048a,a8051a,a8055a,a8056a,a8057a,a8060a,a8064a,a8065a,a8066a,a8069a,a8073a,a8074a,a8075a,a8078a,a8082a,a8083a,a8084a,a8087a,a8091a,a8092a,a8093a,a8096a,a8100a,a8101a,a8102a,a8105a,a8109a,a8110a,a8111a,a8114a,a8118a,a8119a,a8120a,a8123a,a8127a,a8128a,a8129a,a8132a,a8136a,a8137a,a8138a,a8141a,a8145a,a8146a,a8147a,a8150a,a8154a,a8155a,a8156a,a8159a,a8163a,a8164a,a8165a,a8168a,a8172a,a8173a,a8174a,a8177a,a8181a,a8182a,a8183a,a8186a,a8190a,a8191a,a8192a,a8195a,a8199a,a8200a,a8201a,a8204a,a8208a,a8209a,a8210a,a8213a,a8217a,a8218a,a8219a,a8222a,a8226a,a8227a,a8228a,a8231a,a8235a,a8236a,a8237a,a8240a,a8244a,a8245a,a8246a,a8249a,a8253a,a8254a,a8255a,a8258a,a8262a,a8263a,a8264a,a8267a,a8271a,a8272a,a8273a,a8276a,a8280a,a8281a,a8282a,a8285a,a8289a,a8290a,a8291a,a8294a,a8298a,a8299a,a8300a,a8303a,a8307a,a8308a,a8309a,a8312a,a8316a,a8317a,a8318a,a8321a,a8325a,a8326a,a8327a,a8330a,a8334a,a8335a,a8336a,a8339a,a8343a,a8344a,a8345a,a8348a,a8352a,a8353a,a8354a,a8357a,a8361a,a8362a,a8363a,a8366a,a8370a,a8371a,a8372a,a8375a,a8379a,a8380a,a8381a,a8384a,a8388a,a8389a,a8390a,a8393a,a8397a,a8398a,a8399a,a8402a,a8406a,a8407a,a8408a,a8411a,a8415a,a8416a,a8417a,a8420a,a8424a,a8425a,a8426a,a8429a,a8433a,a8434a,a8435a,a8438a,a8442a,a8443a,a8444a,a8447a,a8451a,a8452a,a8453a,a8456a,a8460a,a8461a,a8462a,a8465a,a8469a,a8470a,a8471a,a8474a,a8478a,a8479a,a8480a,a8483a,a8487a,a8488a,a8489a,a8492a,a8496a,a8497a,a8498a,a8501a,a8505a,a8506a,a8507a,a8510a,a8514a,a8515a,a8516a,a8519a,a8523a,a8524a,a8525a,a8528a,a8532a,a8533a,a8534a,a8537a,a8541a,a8542a,a8543a,a8546a,a8550a,a8551a,a8552a,a8555a,a8559a,a8560a,a8561a,a8564a,a8568a,a8569a,a8570a,a8573a,a8577a,a8578a,a8579a,a8582a,a8586a,a8587a,a8588a,a8591a,a8595a,a8596a,a8597a,a8600a,a8604a,a8605a,a8606a,a8609a,a8613a,a8614a,a8615a,a8618a,a8622a,a8623a,a8624a,a8627a,a8631a,a8632a,a8633a,a8636a,a8640a,a8641a,a8642a,a8645a,a8649a,a8650a,a8651a,a8654a,a8658a,a8659a,a8660a,a8663a,a8667a,a8668a,a8669a,a8672a,a8676a,a8677a,a8678a,a8681a,a8685a,a8686a,a8687a,a8690a,a8694a,a8695a,a8696a,a8699a,a8703a,a8704a,a8705a,a8708a,a8712a,a8713a,a8714a,a8717a,a8721a,a8722a,a8723a,a8726a,a8730a,a8731a,a8732a,a8735a,a8739a,a8740a,a8741a,a8744a,a8748a,a8749a,a8750a,a8753a,a8757a,a8758a,a8759a,a8762a,a8766a,a8767a,a8768a,a8771a,a8775a,a8776a,a8777a,a8780a,a8784a,a8785a,a8786a,a8789a,a8793a,a8794a,a8795a,a8798a,a8802a,a8803a,a8804a,a8807a,a8811a,a8812a,a8813a,a8816a,a8820a,a8821a,a8822a,a8825a,a8829a,a8830a,a8831a,a8834a,a8838a,a8839a,a8840a,a8843a,a8847a,a8848a,a8849a,a8852a,a8856a,a8857a,a8858a,a8861a,a8865a,a8866a,a8867a,a8870a,a8874a,a8875a,a8876a,a8879a,a8883a,a8884a,a8885a,a8888a,a8892a,a8893a,a8894a,a8897a,a8901a,a8902a,a8903a,a8906a,a8910a,a8911a,a8912a,a8915a,a8919a,a8920a,a8921a,a8924a,a8928a,a8929a,a8930a,a8933a,a8937a,a8938a,a8939a,a8942a,a8946a,a8947a,a8948a,a8951a,a8955a,a8956a,a8957a,a8960a,a8964a,a8965a,a8966a,a8969a,a8973a,a8974a,a8975a,a8978a,a8982a,a8983a,a8984a,a8987a,a8991a,a8992a,a8993a,a8996a,a9000a,a9001a,a9002a,a9005a,a9009a,a9010a,a9011a,a9014a,a9018a,a9019a,a9020a,a9023a,a9027a,a9028a,a9029a,a9032a,a9036a,a9037a,a9038a,a9041a,a9045a,a9046a,a9047a,a9050a,a9054a,a9055a,a9056a,a9059a,a9063a,a9064a,a9065a,a9068a,a9072a,a9073a,a9074a,a9077a,a9081a,a9082a,a9083a,a9086a,a9090a,a9091a,a9092a,a9095a,a9099a,a9100a,a9101a,a9104a,a9108a,a9109a,a9110a,a9113a,a9117a,a9118a,a9119a,a9122a,a9126a,a9127a,a9128a,a9131a,a9135a,a9136a,a9137a,a9140a,a9144a,a9145a,a9146a,a9149a,a9153a,a9154a,a9155a,a9158a,a9162a,a9163a,a9164a,a9167a,a9171a,a9172a,a9173a,a9176a,a9180a,a9181a,a9182a,a9185a,a9189a,a9190a,a9191a,a9194a,a9198a,a9199a,a9200a,a9203a,a9207a,a9208a,a9209a,a9212a,a9216a,a9217a,a9218a,a9221a,a9225a,a9226a,a9227a,a9230a,a9234a,a9235a,a9236a,a9239a,a9243a,a9244a,a9245a,a9248a,a9252a,a9253a,a9254a,a9257a,a9261a,a9262a,a9263a,a9266a,a9270a,a9271a,a9272a,a9275a,a9279a,a9280a,a9281a,a9284a,a9288a,a9289a,a9290a,a9293a,a9297a,a9298a,a9299a,a9302a,a9306a,a9307a,a9308a,a9311a,a9315a,a9316a,a9317a,a9320a,a9324a,a9325a,a9326a,a9329a,a9333a,a9334a,a9335a,a9338a,a9342a,a9343a,a9344a,a9347a,a9351a,a9352a,a9353a,a9356a,a9360a,a9361a,a9362a,a9365a,a9369a,a9370a,a9371a,a9374a,a9378a,a9379a,a9380a,a9383a,a9387a,a9388a,a9389a,a9392a,a9396a,a9397a,a9398a,a9401a,a9405a,a9406a,a9407a,a9410a,a9414a,a9415a,a9416a,a9419a,a9423a,a9424a,a9425a,a9428a,a9432a,a9433a,a9434a,a9437a,a9441a,a9442a,a9443a,a9446a,a9450a,a9451a,a9452a,a9455a,a9459a,a9460a,a9461a,a9464a,a9468a,a9469a,a9470a,a9473a,a9477a,a9478a,a9479a,a9482a,a9486a,a9487a,a9488a,a9491a,a9495a,a9496a,a9497a,a9500a,a9504a,a9505a,a9506a,a9509a,a9513a,a9514a,a9515a,a9518a,a9522a,a9523a,a9524a,a9527a,a9531a,a9532a,a9533a,a9536a,a9540a,a9541a,a9542a,a9545a,a9549a,a9550a,a9551a,a9554a,a9558a,a9559a,a9560a,a9563a,a9567a,a9568a,a9569a,a9572a,a9576a,a9577a,a9578a,a9581a,a9585a,a9586a,a9587a,a9590a,a9594a,a9595a,a9596a,a9599a,a9603a,a9604a,a9605a,a9608a,a9612a,a9613a,a9614a,a9617a,a9621a,a9622a,a9623a,a9626a,a9630a,a9631a,a9632a,a9635a,a9639a,a9640a,a9641a,a9644a,a9648a,a9649a,a9650a,a9653a,a9657a,a9658a,a9659a,a9662a,a9666a,a9667a,a9668a,a9671a,a9675a,a9676a,a9677a,a9680a,a9684a,a9685a,a9686a,a9689a,a9693a,a9694a,a9695a,a9698a,a9702a,a9703a,a9704a,a9707a,a9711a,a9712a,a9713a,a9716a,a9720a,a9721a,a9722a,a9725a,a9729a,a9730a,a9731a,a9734a,a9738a,a9739a,a9740a,a9743a,a9747a,a9748a,a9749a,a9752a,a9756a,a9757a,a9758a,a9761a,a9765a,a9766a,a9767a,a9770a,a9774a,a9775a,a9776a,a9779a,a9783a,a9784a,a9785a,a9788a,a9792a,a9793a,a9794a,a9797a,a9801a,a9802a,a9803a,a9806a,a9810a,a9811a,a9812a,a9815a,a9819a,a9820a,a9821a,a9824a,a9828a,a9829a,a9830a,a9833a,a9837a,a9838a,a9839a,a9842a,a9846a,a9847a,a9848a,a9851a,a9855a,a9856a,a9857a,a9860a,a9864a,a9865a,a9866a,a9869a,a9873a,a9874a,a9875a,a9878a,a9882a,a9883a,a9884a,a9887a,a9891a,a9892a,a9893a,a9896a,a9900a,a9901a,a9902a,a9905a,a9909a,a9910a,a9911a,a9914a,a9918a,a9919a,a9920a,a9923a,a9927a,a9928a,a9929a,a9932a,a9936a,a9937a,a9938a,a9941a,a9945a,a9946a,a9947a,a9950a,a9954a,a9955a,a9956a,a9959a,a9963a,a9964a,a9965a,a9968a,a9972a,a9973a,a9974a,a9977a,a9981a,a9982a,a9983a,a9986a,a9990a,a9991a,a9992a,a9995a,a9999a,a10000a,a10001a,a10004a,a10008a,a10009a,a10010a,a10013a,a10017a,a10018a,a10019a,a10022a,a10026a,a10027a,a10028a,a10031a,a10035a,a10036a,a10037a,a10040a,a10044a,a10045a,a10046a,a10049a,a10053a,a10054a,a10055a,a10058a,a10062a,a10063a,a10064a,a10067a,a10071a,a10072a,a10073a,a10076a,a10080a,a10081a,a10082a,a10085a,a10089a,a10090a,a10091a,a10094a,a10098a,a10099a,a10100a,a10103a,a10107a,a10108a,a10109a,a10112a,a10116a,a10117a,a10118a,a10121a,a10125a,a10126a,a10127a,a10130a,a10134a,a10135a,a10136a,a10139a,a10143a,a10144a,a10145a,a10148a,a10152a,a10153a,a10154a,a10157a,a10161a,a10162a,a10163a,a10166a,a10170a,a10171a,a10172a,a10175a,a10179a,a10180a,a10181a,a10184a,a10188a,a10189a,a10190a,a10193a,a10197a,a10198a,a10199a,a10202a,a10206a,a10207a,a10208a,a10211a,a10215a,a10216a,a10217a,a10220a,a10224a,a10225a,a10226a,a10229a,a10233a,a10234a,a10235a,a10238a,a10242a,a10243a,a10244a,a10247a,a10251a,a10252a,a10253a,a10256a,a10260a,a10261a,a10262a,a10265a,a10269a,a10270a,a10271a,a10274a,a10278a,a10279a,a10280a,a10283a,a10287a,a10288a,a10289a,a10292a,a10296a,a10297a,a10298a,a10301a,a10305a,a10306a,a10307a,a10310a,a10314a,a10315a,a10316a,a10319a,a10323a,a10324a,a10325a,a10328a,a10332a,a10333a,a10334a,a10338a,a10339a,a10343a,a10344a,a10345a,a10348a,a10352a,a10353a,a10354a,a10358a,a10359a,a10363a,a10364a,a10365a,a10368a,a10372a,a10373a,a10374a,a10378a,a10379a,a10383a,a10384a,a10385a,a10388a,a10392a,a10393a,a10394a,a10398a,a10399a,a10403a,a10404a,a10405a,a10408a,a10412a,a10413a,a10414a,a10418a,a10419a,a10423a,a10424a,a10425a,a10428a,a10432a,a10433a,a10434a,a10438a,a10439a,a10443a,a10444a,a10445a,a10448a,a10452a,a10453a,a10454a,a10458a,a10459a,a10463a,a10464a,a10465a,a10468a,a10472a,a10473a,a10474a,a10478a,a10479a,a10483a,a10484a,a10485a,a10488a,a10492a,a10493a,a10494a,a10498a,a10499a,a10503a,a10504a,a10505a,a10508a,a10512a,a10513a,a10514a,a10518a,a10519a,a10523a,a10524a,a10525a,a10528a,a10532a,a10533a,a10534a,a10538a,a10539a,a10543a,a10544a,a10545a,a10548a,a10552a,a10553a,a10554a,a10558a,a10559a,a10563a,a10564a,a10565a,a10568a,a10572a,a10573a,a10574a,a10578a,a10579a,a10583a,a10584a,a10585a,a10588a,a10592a,a10593a,a10594a,a10598a,a10599a,a10603a,a10604a,a10605a,a10608a,a10612a,a10613a,a10614a,a10618a,a10619a,a10623a,a10624a,a10625a,a10628a,a10632a,a10633a,a10634a,a10638a,a10639a,a10643a,a10644a,a10645a,a10648a,a10652a,a10653a,a10654a,a10658a,a10659a,a10663a,a10664a,a10665a,a10668a,a10672a,a10673a,a10674a,a10678a,a10679a,a10683a,a10684a,a10685a,a10688a,a10692a,a10693a,a10694a,a10698a,a10699a,a10703a,a10704a,a10705a,a10708a,a10712a,a10713a,a10714a,a10718a,a10719a,a10723a,a10724a,a10725a,a10728a,a10732a,a10733a,a10734a,a10738a,a10739a,a10743a,a10744a,a10745a,a10748a,a10752a,a10753a,a10754a,a10758a,a10759a,a10763a,a10764a,a10765a,a10768a,a10772a,a10773a,a10774a,a10778a,a10779a,a10783a,a10784a,a10785a,a10788a,a10792a,a10793a,a10794a,a10798a,a10799a,a10803a,a10804a,a10805a,a10808a,a10812a,a10813a,a10814a,a10818a,a10819a,a10823a,a10824a,a10825a,a10828a,a10832a,a10833a,a10834a,a10838a,a10839a,a10843a,a10844a,a10845a,a10848a,a10852a,a10853a,a10854a,a10858a,a10859a,a10863a,a10864a,a10865a,a10868a,a10872a,a10873a,a10874a,a10878a,a10879a,a10883a,a10884a,a10885a,a10888a,a10892a,a10893a,a10894a,a10898a,a10899a,a10903a,a10904a,a10905a,a10908a,a10912a,a10913a,a10914a,a10918a,a10919a,a10923a,a10924a,a10925a,a10928a,a10932a,a10933a,a10934a,a10938a,a10939a,a10943a,a10944a,a10945a,a10948a,a10952a,a10953a,a10954a,a10958a,a10959a,a10963a,a10964a,a10965a,a10968a,a10972a,a10973a,a10974a,a10978a,a10979a,a10983a,a10984a,a10985a,a10988a,a10992a,a10993a,a10994a,a10998a,a10999a,a11003a,a11004a,a11005a,a11008a,a11012a,a11013a,a11014a,a11018a,a11019a,a11023a,a11024a,a11025a,a11028a,a11032a,a11033a,a11034a,a11038a,a11039a,a11043a,a11044a,a11045a,a11048a,a11052a,a11053a,a11054a,a11058a,a11059a,a11063a,a11064a,a11065a,a11068a,a11072a,a11073a,a11074a,a11078a,a11079a,a11083a,a11084a,a11085a,a11088a,a11092a,a11093a,a11094a,a11098a,a11099a,a11103a,a11104a,a11105a,a11108a,a11112a,a11113a,a11114a,a11118a,a11119a,a11123a,a11124a,a11125a,a11128a,a11132a,a11133a,a11134a,a11138a,a11139a,a11143a,a11144a,a11145a,a11148a,a11152a,a11153a,a11154a,a11158a,a11159a,a11163a,a11164a,a11165a,a11168a,a11172a,a11173a,a11174a,a11178a,a11179a,a11183a,a11184a,a11185a,a11188a,a11192a,a11193a,a11194a,a11198a,a11199a,a11203a,a11204a,a11205a,a11208a,a11212a,a11213a,a11214a,a11218a,a11219a,a11223a,a11224a,a11225a,a11228a,a11232a,a11233a,a11234a,a11238a,a11239a,a11243a,a11244a,a11245a,a11248a,a11252a,a11253a,a11254a,a11258a,a11259a,a11263a,a11264a,a11265a,a11268a,a11272a,a11273a,a11274a,a11278a,a11279a,a11283a,a11284a,a11285a,a11288a,a11292a,a11293a,a11294a,a11298a,a11299a,a11303a,a11304a,a11305a,a11308a,a11312a,a11313a,a11314a,a11318a,a11319a,a11323a,a11324a,a11325a,a11328a,a11332a,a11333a,a11334a,a11338a,a11339a,a11343a,a11344a,a11345a,a11348a,a11352a,a11353a,a11354a,a11358a,a11359a,a11363a,a11364a,a11365a,a11368a,a11372a,a11373a,a11374a,a11378a,a11379a,a11383a,a11384a,a11385a,a11388a,a11392a,a11393a,a11394a,a11398a,a11399a,a11403a,a11404a,a11405a,a11408a,a11412a,a11413a,a11414a,a11418a,a11419a,a11423a,a11424a,a11425a,a11428a,a11432a,a11433a,a11434a,a11438a,a11439a,a11443a,a11444a,a11445a,a11448a,a11452a,a11453a,a11454a,a11458a,a11459a,a11463a,a11464a,a11465a,a11468a,a11472a,a11473a,a11474a,a11478a,a11479a,a11483a,a11484a,a11485a,a11488a,a11492a,a11493a,a11494a,a11498a,a11499a,a11503a,a11504a,a11505a,a11508a,a11512a,a11513a,a11514a,a11518a,a11519a,a11523a,a11524a,a11525a,a11528a,a11532a,a11533a,a11534a,a11538a,a11539a,a11543a,a11544a,a11545a,a11548a,a11552a,a11553a,a11554a,a11558a,a11559a,a11563a,a11564a,a11565a,a11568a,a11572a,a11573a,a11574a,a11578a,a11579a,a11583a,a11584a,a11585a,a11588a,a11592a,a11593a,a11594a,a11598a,a11599a,a11603a,a11604a,a11605a,a11608a,a11612a,a11613a,a11614a,a11618a,a11619a,a11623a,a11624a,a11625a,a11628a,a11632a,a11633a,a11634a,a11638a,a11639a,a11643a,a11644a,a11645a,a11648a,a11652a,a11653a,a11654a,a11658a,a11659a,a11663a,a11664a,a11665a,a11668a,a11672a,a11673a,a11674a,a11678a,a11679a,a11683a,a11684a,a11685a,a11688a,a11692a,a11693a,a11694a,a11698a,a11699a,a11703a,a11704a,a11705a,a11708a,a11712a,a11713a,a11714a,a11718a,a11719a,a11723a,a11724a,a11725a,a11728a,a11732a,a11733a,a11734a,a11738a,a11739a,a11743a,a11744a,a11745a,a11748a,a11752a,a11753a,a11754a,a11758a,a11759a,a11763a,a11764a,a11765a,a11768a,a11772a,a11773a,a11774a,a11778a,a11779a,a11783a,a11784a,a11785a,a11788a,a11792a,a11793a,a11794a,a11798a,a11799a,a11803a,a11804a,a11805a,a11808a,a11812a,a11813a,a11814a,a11818a,a11819a,a11823a,a11824a,a11825a,a11828a,a11832a,a11833a,a11834a,a11838a,a11839a,a11843a,a11844a,a11845a,a11848a,a11852a,a11853a,a11854a,a11858a,a11859a,a11863a,a11864a,a11865a,a11868a,a11872a,a11873a,a11874a,a11878a,a11879a,a11883a,a11884a,a11885a,a11888a,a11892a,a11893a,a11894a,a11898a,a11899a,a11903a,a11904a,a11905a,a11908a,a11912a,a11913a,a11914a,a11918a,a11919a,a11923a,a11924a,a11925a,a11928a,a11932a,a11933a,a11934a,a11938a,a11939a,a11943a,a11944a,a11945a,a11948a,a11952a,a11953a,a11954a,a11958a,a11959a,a11963a,a11964a,a11965a,a11968a,a11972a,a11973a,a11974a,a11978a,a11979a,a11983a,a11984a,a11985a,a11988a,a11992a,a11993a,a11994a,a11998a,a11999a,a12003a,a12004a,a12005a,a12008a,a12012a,a12013a,a12014a,a12018a,a12019a,a12023a,a12024a,a12025a,a12028a,a12032a,a12033a,a12034a,a12038a,a12039a,a12043a,a12044a,a12045a,a12048a,a12052a,a12053a,a12054a,a12058a,a12059a,a12063a,a12064a,a12065a,a12068a,a12072a,a12073a,a12074a,a12078a,a12079a,a12083a,a12084a,a12085a,a12088a,a12092a,a12093a,a12094a,a12098a,a12099a,a12103a,a12104a,a12105a,a12108a,a12112a,a12113a,a12114a,a12118a,a12119a,a12123a,a12124a,a12125a,a12128a,a12132a,a12133a,a12134a,a12138a,a12139a,a12143a,a12144a,a12145a,a12148a,a12152a,a12153a,a12154a,a12158a,a12159a,a12163a,a12164a,a12165a,a12168a,a12172a,a12173a,a12174a,a12178a,a12179a,a12183a,a12184a,a12185a,a12188a,a12192a,a12193a,a12194a,a12198a,a12199a,a12203a,a12204a,a12205a,a12208a,a12212a,a12213a,a12214a,a12218a,a12219a,a12223a,a12224a,a12225a,a12228a,a12232a,a12233a,a12234a,a12238a,a12239a,a12243a,a12244a,a12245a,a12248a,a12252a,a12253a,a12254a,a12258a,a12259a,a12263a,a12264a,a12265a,a12268a,a12272a,a12273a,a12274a,a12278a,a12279a,a12283a,a12284a,a12285a,a12288a,a12292a,a12293a,a12294a,a12298a,a12299a,a12303a,a12304a,a12305a,a12308a,a12312a,a12313a,a12314a,a12318a,a12319a,a12323a,a12324a,a12325a,a12328a,a12332a,a12333a,a12334a,a12338a,a12339a,a12343a,a12344a,a12345a,a12348a,a12352a,a12353a,a12354a,a12358a,a12359a,a12363a,a12364a,a12365a,a12368a,a12372a,a12373a,a12374a,a12378a,a12379a,a12383a,a12384a,a12385a,a12388a,a12392a,a12393a,a12394a,a12398a,a12399a,a12403a,a12404a,a12405a,a12408a,a12412a,a12413a,a12414a,a12418a,a12419a,a12423a,a12424a,a12425a,a12428a,a12432a,a12433a,a12434a,a12438a,a12439a,a12443a,a12444a,a12445a,a12448a,a12452a,a12453a,a12454a,a12458a,a12459a,a12463a,a12464a,a12465a,a12468a,a12472a,a12473a,a12474a,a12478a,a12479a,a12483a,a12484a,a12485a,a12488a,a12492a,a12493a,a12494a,a12498a,a12499a,a12503a,a12504a,a12505a,a12508a,a12512a,a12513a,a12514a,a12518a,a12519a,a12523a,a12524a,a12525a,a12528a,a12532a,a12533a,a12534a,a12538a,a12539a,a12543a,a12544a,a12545a,a12548a,a12552a,a12553a,a12554a,a12558a,a12559a,a12563a,a12564a,a12565a,a12568a,a12572a,a12573a,a12574a,a12578a,a12579a,a12583a,a12584a,a12585a,a12588a,a12592a,a12593a,a12594a,a12598a,a12599a,a12603a,a12604a,a12605a,a12608a,a12612a,a12613a,a12614a,a12618a,a12619a,a12623a,a12624a,a12625a,a12628a,a12632a,a12633a,a12634a,a12638a,a12639a,a12643a,a12644a,a12645a,a12648a,a12652a,a12653a,a12654a,a12658a,a12659a,a12663a,a12664a,a12665a,a12668a,a12672a,a12673a,a12674a,a12678a,a12679a,a12683a,a12684a,a12685a,a12688a,a12692a,a12693a,a12694a,a12698a,a12699a,a12703a,a12704a,a12705a,a12708a,a12712a,a12713a,a12714a,a12718a,a12719a,a12723a,a12724a,a12725a,a12728a,a12732a,a12733a,a12734a,a12738a,a12739a,a12743a,a12744a,a12745a,a12748a,a12752a,a12753a,a12754a,a12758a,a12759a,a12763a,a12764a,a12765a,a12768a,a12772a,a12773a,a12774a,a12778a,a12779a,a12783a,a12784a,a12785a,a12788a,a12792a,a12793a,a12794a,a12798a,a12799a,a12803a,a12804a,a12805a,a12808a,a12812a,a12813a,a12814a,a12818a,a12819a,a12823a,a12824a,a12825a,a12828a,a12832a,a12833a,a12834a,a12838a,a12839a,a12843a,a12844a,a12845a,a12848a,a12852a,a12853a,a12854a,a12858a,a12859a,a12863a,a12864a,a12865a,a12868a,a12872a,a12873a,a12874a,a12878a,a12879a,a12883a,a12884a,a12885a,a12888a,a12892a,a12893a,a12894a,a12898a,a12899a,a12903a,a12904a,a12905a,a12908a,a12912a,a12913a,a12914a,a12918a,a12919a,a12923a,a12924a,a12925a,a12928a,a12932a,a12933a,a12934a,a12938a,a12939a,a12943a,a12944a,a12945a,a12948a,a12952a,a12953a,a12954a,a12958a,a12959a,a12963a,a12964a,a12965a,a12968a,a12972a,a12973a,a12974a,a12978a,a12979a,a12983a,a12984a,a12985a,a12988a,a12992a,a12993a,a12994a,a12998a,a12999a,a13003a,a13004a,a13005a,a13008a,a13012a,a13013a,a13014a,a13018a,a13019a,a13023a,a13024a,a13025a,a13028a,a13032a,a13033a,a13034a,a13038a,a13039a,a13043a,a13044a,a13045a,a13048a,a13052a,a13053a,a13054a,a13058a,a13059a,a13063a,a13064a,a13065a,a13068a,a13072a,a13073a,a13074a,a13078a,a13079a,a13083a,a13084a,a13085a,a13088a,a13092a,a13093a,a13094a,a13098a,a13099a,a13103a,a13104a,a13105a,a13108a,a13112a,a13113a,a13114a,a13118a,a13119a,a13123a,a13124a,a13125a,a13128a,a13132a,a13133a,a13134a,a13138a,a13139a,a13143a,a13144a,a13145a,a13148a,a13152a,a13153a,a13154a,a13158a,a13159a,a13163a,a13164a,a13165a,a13168a,a13172a,a13173a,a13174a,a13178a,a13179a,a13183a,a13184a,a13185a,a13188a,a13192a,a13193a,a13194a,a13198a,a13199a,a13203a,a13204a,a13205a,a13208a,a13212a,a13213a,a13214a,a13218a,a13219a,a13223a,a13224a,a13225a,a13228a,a13232a,a13233a,a13234a,a13238a,a13239a,a13243a,a13244a,a13245a,a13248a,a13252a,a13253a,a13254a,a13258a,a13259a,a13263a,a13264a,a13265a,a13268a,a13272a,a13273a,a13274a,a13278a,a13279a,a13283a,a13284a,a13285a,a13288a,a13292a,a13293a,a13294a,a13298a,a13299a,a13303a,a13304a,a13305a,a13308a,a13312a,a13313a,a13314a,a13318a,a13319a,a13323a,a13324a,a13325a,a13328a,a13332a,a13333a,a13334a,a13338a,a13339a,a13343a,a13344a,a13345a,a13348a,a13352a,a13353a,a13354a,a13358a,a13359a,a13363a,a13364a,a13365a,a13368a,a13372a,a13373a,a13374a,a13378a,a13379a,a13383a,a13384a,a13385a,a13388a,a13392a,a13393a,a13394a,a13398a,a13399a,a13403a,a13404a,a13405a,a13408a,a13412a,a13413a,a13414a,a13418a,a13419a,a13423a,a13424a,a13425a,a13428a,a13432a,a13433a,a13434a,a13438a,a13439a,a13443a,a13444a,a13445a,a13448a,a13452a,a13453a,a13454a,a13458a,a13459a,a13463a,a13464a,a13465a,a13468a,a13472a,a13473a,a13474a,a13478a,a13479a,a13483a,a13484a,a13485a,a13488a,a13492a,a13493a,a13494a,a13498a,a13499a,a13503a,a13504a,a13505a,a13508a,a13512a,a13513a,a13514a,a13518a,a13519a,a13523a,a13524a,a13525a,a13528a,a13532a,a13533a,a13534a,a13538a,a13539a,a13543a,a13544a,a13545a,a13548a,a13552a,a13553a,a13554a,a13558a,a13559a,a13563a,a13564a,a13565a,a13568a,a13572a,a13573a,a13574a,a13578a,a13579a,a13583a,a13584a,a13585a,a13588a,a13592a,a13593a,a13594a,a13598a,a13599a,a13603a,a13604a,a13605a,a13608a,a13612a,a13613a,a13614a,a13618a,a13619a,a13623a,a13624a,a13625a,a13628a,a13632a,a13633a,a13634a,a13638a,a13639a,a13643a,a13644a,a13645a,a13648a,a13652a,a13653a,a13654a,a13658a,a13659a,a13663a,a13664a,a13665a,a13668a,a13672a,a13673a,a13674a,a13678a,a13679a,a13683a,a13684a,a13685a,a13689a,a13690a,a13694a,a13695a,a13696a,a13700a,a13701a,a13705a,a13706a,a13707a,a13711a,a13712a,a13716a,a13717a,a13718a,a13722a,a13723a,a13727a,a13728a,a13729a,a13733a,a13734a,a13738a,a13739a,a13740a,a13744a,a13745a,a13749a,a13750a,a13751a,a13755a,a13756a,a13760a,a13761a,a13762a,a13766a,a13767a,a13771a,a13772a,a13773a,a13777a,a13778a,a13782a,a13783a,a13784a,a13788a,a13789a,a13793a,a13794a,a13795a,a13799a,a13800a,a13804a,a13805a,a13806a,a13810a,a13811a,a13815a,a13816a,a13817a,a13821a,a13822a,a13826a,a13827a,a13828a,a13832a,a13833a,a13837a,a13838a,a13839a,a13843a,a13844a,a13848a,a13849a,a13850a,a13854a,a13855a,a13859a,a13860a,a13861a,a13865a,a13866a,a13870a,a13871a,a13872a,a13876a,a13877a,a13881a,a13882a,a13883a,a13887a,a13888a,a13892a,a13893a,a13894a,a13898a,a13899a,a13903a,a13904a,a13905a,a13909a,a13910a,a13914a,a13915a,a13916a,a13920a,a13921a,a13925a,a13926a,a13927a,a13931a,a13932a,a13936a,a13937a,a13938a,a13942a,a13943a,a13947a,a13948a,a13949a,a13953a,a13954a,a13958a,a13959a,a13960a,a13964a,a13965a,a13969a,a13970a,a13971a,a13975a,a13976a,a13980a,a13981a,a13982a,a13986a,a13987a,a13991a,a13992a,a13993a,a13997a,a13998a,a14002a,a14003a,a14004a,a14008a,a14009a,a14013a,a14014a,a14015a,a14019a,a14020a,a14024a,a14025a,a14026a,a14030a,a14031a,a14035a,a14036a,a14037a,a14041a,a14042a,a14046a,a14047a,a14048a,a14052a,a14053a,a14057a,a14058a,a14059a,a14063a,a14064a,a14068a,a14069a,a14070a,a14074a,a14075a,a14079a,a14080a,a14081a,a14085a,a14086a,a14090a,a14091a,a14092a,a14096a,a14097a,a14101a,a14102a,a14103a,a14107a,a14108a,a14112a,a14113a,a14114a,a14118a,a14119a,a14123a,a14124a,a14125a,a14129a,a14130a,a14134a,a14135a,a14136a,a14140a,a14141a,a14145a,a14146a,a14147a,a14151a,a14152a,a14156a,a14157a,a14158a,a14162a,a14163a,a14167a,a14168a,a14169a,a14173a,a14174a,a14178a,a14179a,a14180a,a14184a,a14185a,a14189a,a14190a,a14191a,a14195a,a14196a,a14200a,a14201a,a14202a,a14206a,a14207a,a14211a,a14212a,a14213a,a14217a,a14218a,a14222a,a14223a,a14224a,a14228a,a14229a,a14233a,a14234a,a14235a,a14239a,a14240a,a14244a,a14245a,a14246a,a14250a,a14251a,a14255a,a14256a,a14257a,a14261a,a14262a,a14266a,a14267a,a14268a,a14272a,a14273a,a14277a,a14278a,a14279a,a14283a,a14284a,a14288a,a14289a,a14290a,a14294a,a14295a,a14299a,a14300a,a14301a,a14305a,a14306a,a14310a,a14311a,a14312a,a14316a,a14317a,a14321a,a14322a,a14323a,a14327a,a14328a,a14332a,a14333a,a14334a,a14338a,a14339a,a14343a,a14344a,a14345a,a14349a,a14350a,a14354a,a14355a,a14356a,a14360a,a14361a,a14365a,a14366a,a14367a,a14371a,a14372a,a14376a,a14377a,a14378a,a14382a,a14383a,a14387a,a14388a,a14389a,a14393a,a14394a,a14398a,a14399a,a14400a,a14404a,a14405a,a14409a,a14410a,a14411a,a14415a,a14416a,a14420a,a14421a,a14422a,a14426a,a14427a,a14431a,a14432a,a14433a,a14437a,a14438a,a14442a,a14443a,a14444a,a14448a,a14449a,a14453a,a14454a,a14455a,a14459a,a14460a,a14464a,a14465a,a14466a,a14470a,a14471a,a14475a,a14476a,a14477a,a14481a,a14482a,a14486a,a14487a,a14488a,a14492a,a14493a,a14497a,a14498a,a14499a,a14503a,a14504a,a14508a,a14509a,a14510a,a14514a,a14515a,a14519a,a14520a,a14521a,a14525a,a14526a,a14530a,a14531a,a14532a,a14536a,a14537a,a14541a,a14542a,a14543a,a14547a,a14548a,a14552a,a14553a,a14554a,a14558a,a14559a,a14563a,a14564a,a14565a,a14569a,a14570a,a14574a,a14575a,a14576a,a14580a,a14581a,a14585a,a14586a,a14587a,a14591a,a14592a,a14596a,a14597a,a14598a,a14602a,a14603a,a14607a,a14608a,a14609a,a14613a,a14614a,a14618a,a14619a,a14620a,a14624a,a14625a,a14629a,a14630a,a14631a,a14635a,a14636a,a14640a,a14641a,a14642a,a14646a,a14647a,a14651a,a14652a,a14653a,a14657a,a14658a,a14662a,a14663a,a14664a,a14668a,a14669a,a14673a,a14674a,a14675a,a14679a,a14680a,a14684a,a14685a,a14686a,a14690a,a14691a,a14695a,a14696a,a14697a,a14701a,a14702a,a14706a,a14707a,a14708a,a14712a,a14713a,a14717a,a14718a,a14719a,a14723a,a14724a,a14728a,a14729a,a14730a,a14734a,a14735a,a14739a,a14740a,a14741a,a14745a,a14746a,a14750a,a14751a,a14752a,a14756a,a14757a,a14761a,a14762a,a14763a,a14767a,a14768a,a14772a,a14773a,a14774a,a14778a,a14779a,a14783a,a14784a,a14785a,a14789a,a14790a,a14794a,a14795a,a14796a,a14800a,a14801a,a14805a,a14806a,a14807a,a14811a,a14812a,a14816a,a14817a,a14818a,a14822a,a14823a,a14827a,a14828a,a14829a,a14833a,a14834a,a14838a,a14839a,a14840a,a14844a,a14845a,a14849a,a14850a,a14851a,a14855a,a14856a,a14860a,a14861a,a14862a,a14866a,a14867a,a14871a,a14872a,a14873a,a14877a,a14878a,a14882a,a14883a,a14884a,a14888a,a14889a,a14893a,a14894a,a14895a,a14899a,a14900a,a14904a,a14905a,a14906a,a14910a,a14911a,a14915a,a14916a,a14917a,a14921a,a14922a,a14926a,a14927a,a14928a,a14932a,a14933a,a14937a,a14938a,a14939a,a14943a,a14944a,a14948a,a14949a,a14950a,a14954a,a14955a,a14959a,a14960a,a14961a,a14965a,a14966a,a14970a,a14971a,a14972a,a14976a,a14977a,a14981a,a14982a,a14983a,a14987a,a14988a,a14992a,a14993a,a14994a,a14998a,a14999a,a15003a,a15004a,a15005a,a15009a,a15010a,a15014a,a15015a,a15016a,a15020a,a15021a,a15025a,a15026a,a15027a,a15031a,a15032a,a15036a,a15037a,a15038a,a15042a,a15043a,a15047a,a15048a,a15049a,a15053a,a15054a,a15058a,a15059a,a15060a,a15064a,a15065a,a15069a,a15070a,a15071a,a15075a,a15076a,a15080a,a15081a,a15082a,a15086a,a15087a,a15091a,a15092a,a15093a,a15097a,a15098a,a15102a,a15103a,a15104a,a15108a,a15109a,a15113a,a15114a,a15115a,a15119a,a15120a,a15124a,a15125a,a15126a,a15130a,a15131a,a15135a,a15136a,a15137a,a15141a,a15142a,a15146a,a15147a,a15148a,a15152a,a15153a,a15157a,a15158a,a15159a,a15163a,a15164a,a15168a,a15169a,a15170a,a15174a,a15175a,a15179a,a15180a,a15181a,a15185a,a15186a,a15190a,a15191a,a15192a,a15196a,a15197a,a15201a,a15202a,a15203a,a15207a,a15208a,a15212a,a15213a,a15214a,a15218a,a15219a,a15223a,a15224a,a15225a,a15229a,a15230a,a15234a,a15235a,a15236a,a15240a,a15241a,a15245a,a15246a,a15247a,a15251a,a15252a,a15256a,a15257a,a15258a,a15262a,a15263a,a15267a,a15268a,a15269a,a15273a,a15274a,a15278a,a15279a,a15280a,a15284a,a15285a,a15289a,a15290a,a15291a,a15295a,a15296a,a15300a,a15301a,a15302a,a15306a,a15307a,a15311a,a15312a,a15313a,a15317a,a15318a,a15322a,a15323a,a15324a,a15328a,a15329a,a15333a,a15334a,a15335a,a15339a,a15340a,a15344a,a15345a,a15346a,a15350a,a15351a,a15355a,a15356a,a15357a,a15361a,a15362a,a15366a,a15367a,a15368a,a15372a,a15373a,a15377a,a15378a,a15379a,a15383a,a15384a,a15388a,a15389a,a15390a,a15394a,a15395a,a15399a,a15400a,a15401a,a15405a,a15406a,a15410a,a15411a,a15412a,a15416a,a15417a,a15421a,a15422a,a15423a,a15427a,a15428a,a15432a,a15433a,a15434a,a15438a,a15439a,a15443a,a15444a,a15445a,a15449a,a15450a,a15454a,a15455a,a15456a,a15460a,a15461a,a15464a,a15467a,a15468a,a15469a,a15473a,a15474a,a15478a,a15479a,a15480a,a15484a,a15485a,a15488a,a15491a,a15492a,a15493a,a15497a,a15498a,a15502a,a15503a,a15504a,a15508a,a15509a,a15512a,a15515a,a15516a,a15517a,a15521a,a15522a,a15526a,a15527a,a15528a,a15532a,a15533a,a15536a,a15539a,a15540a,a15541a,a15545a,a15546a,a15550a,a15551a,a15552a,a15556a,a15557a,a15560a,a15563a,a15564a,a15565a,a15569a,a15570a,a15574a,a15575a,a15576a,a15580a,a15581a,a15584a,a15587a,a15588a,a15589a,a15593a,a15594a,a15598a,a15599a,a15600a,a15604a,a15605a,a15608a,a15611a,a15612a,a15613a,a15617a,a15618a,a15622a,a15623a,a15624a,a15628a,a15629a,a15632a,a15635a,a15636a,a15637a,a15641a,a15642a,a15646a,a15647a,a15648a,a15652a,a15653a,a15656a,a15659a,a15660a,a15661a,a15665a,a15666a,a15670a,a15671a,a15672a,a15676a,a15677a,a15680a,a15683a,a15684a,a15685a,a15689a,a15690a,a15694a,a15695a,a15696a,a15700a,a15701a,a15704a,a15707a,a15708a,a15709a,a15713a,a15714a,a15718a,a15719a,a15720a,a15724a,a15725a,a15728a,a15731a,a15732a,a15733a,a15737a,a15738a,a15742a,a15743a,a15744a,a15748a,a15749a,a15752a,a15755a,a15756a,a15757a,a15761a,a15762a,a15766a,a15767a,a15768a,a15772a,a15773a,a15776a,a15779a,a15780a,a15781a,a15785a,a15786a,a15790a,a15791a,a15792a,a15796a,a15797a,a15800a,a15803a,a15804a,a15805a,a15809a,a15810a,a15814a,a15815a,a15816a,a15820a,a15821a,a15824a,a15827a,a15828a,a15829a: std_logic;
begin

A75 <=( a2293a ) or ( a1528a );
 a1a <=( a15829a  and  a15816a );
 a2a <=( a15805a  and  a15792a );
 a3a <=( a15781a  and  a15768a );
 a4a <=( a15757a  and  a15744a );
 a5a <=( a15733a  and  a15720a );
 a6a <=( a15709a  and  a15696a );
 a7a <=( a15685a  and  a15672a );
 a8a <=( a15661a  and  a15648a );
 a9a <=( a15637a  and  a15624a );
 a10a <=( a15613a  and  a15600a );
 a11a <=( a15589a  and  a15576a );
 a12a <=( a15565a  and  a15552a );
 a13a <=( a15541a  and  a15528a );
 a14a <=( a15517a  and  a15504a );
 a15a <=( a15493a  and  a15480a );
 a16a <=( a15469a  and  a15456a );
 a17a <=( a15445a  and  a15434a );
 a18a <=( a15423a  and  a15412a );
 a19a <=( a15401a  and  a15390a );
 a20a <=( a15379a  and  a15368a );
 a21a <=( a15357a  and  a15346a );
 a22a <=( a15335a  and  a15324a );
 a23a <=( a15313a  and  a15302a );
 a24a <=( a15291a  and  a15280a );
 a25a <=( a15269a  and  a15258a );
 a26a <=( a15247a  and  a15236a );
 a27a <=( a15225a  and  a15214a );
 a28a <=( a15203a  and  a15192a );
 a29a <=( a15181a  and  a15170a );
 a30a <=( a15159a  and  a15148a );
 a31a <=( a15137a  and  a15126a );
 a32a <=( a15115a  and  a15104a );
 a33a <=( a15093a  and  a15082a );
 a34a <=( a15071a  and  a15060a );
 a35a <=( a15049a  and  a15038a );
 a36a <=( a15027a  and  a15016a );
 a37a <=( a15005a  and  a14994a );
 a38a <=( a14983a  and  a14972a );
 a39a <=( a14961a  and  a14950a );
 a40a <=( a14939a  and  a14928a );
 a41a <=( a14917a  and  a14906a );
 a42a <=( a14895a  and  a14884a );
 a43a <=( a14873a  and  a14862a );
 a44a <=( a14851a  and  a14840a );
 a45a <=( a14829a  and  a14818a );
 a46a <=( a14807a  and  a14796a );
 a47a <=( a14785a  and  a14774a );
 a48a <=( a14763a  and  a14752a );
 a49a <=( a14741a  and  a14730a );
 a50a <=( a14719a  and  a14708a );
 a51a <=( a14697a  and  a14686a );
 a52a <=( a14675a  and  a14664a );
 a53a <=( a14653a  and  a14642a );
 a54a <=( a14631a  and  a14620a );
 a55a <=( a14609a  and  a14598a );
 a56a <=( a14587a  and  a14576a );
 a57a <=( a14565a  and  a14554a );
 a58a <=( a14543a  and  a14532a );
 a59a <=( a14521a  and  a14510a );
 a60a <=( a14499a  and  a14488a );
 a61a <=( a14477a  and  a14466a );
 a62a <=( a14455a  and  a14444a );
 a63a <=( a14433a  and  a14422a );
 a64a <=( a14411a  and  a14400a );
 a65a <=( a14389a  and  a14378a );
 a66a <=( a14367a  and  a14356a );
 a67a <=( a14345a  and  a14334a );
 a68a <=( a14323a  and  a14312a );
 a69a <=( a14301a  and  a14290a );
 a70a <=( a14279a  and  a14268a );
 a71a <=( a14257a  and  a14246a );
 a72a <=( a14235a  and  a14224a );
 a73a <=( a14213a  and  a14202a );
 a74a <=( a14191a  and  a14180a );
 a75a <=( a14169a  and  a14158a );
 a76a <=( a14147a  and  a14136a );
 a77a <=( a14125a  and  a14114a );
 a78a <=( a14103a  and  a14092a );
 a79a <=( a14081a  and  a14070a );
 a80a <=( a14059a  and  a14048a );
 a81a <=( a14037a  and  a14026a );
 a82a <=( a14015a  and  a14004a );
 a83a <=( a13993a  and  a13982a );
 a84a <=( a13971a  and  a13960a );
 a85a <=( a13949a  and  a13938a );
 a86a <=( a13927a  and  a13916a );
 a87a <=( a13905a  and  a13894a );
 a88a <=( a13883a  and  a13872a );
 a89a <=( a13861a  and  a13850a );
 a90a <=( a13839a  and  a13828a );
 a91a <=( a13817a  and  a13806a );
 a92a <=( a13795a  and  a13784a );
 a93a <=( a13773a  and  a13762a );
 a94a <=( a13751a  and  a13740a );
 a95a <=( a13729a  and  a13718a );
 a96a <=( a13707a  and  a13696a );
 a97a <=( a13685a  and  a13674a );
 a98a <=( a13665a  and  a13654a );
 a99a <=( a13645a  and  a13634a );
 a100a <=( a13625a  and  a13614a );
 a101a <=( a13605a  and  a13594a );
 a102a <=( a13585a  and  a13574a );
 a103a <=( a13565a  and  a13554a );
 a104a <=( a13545a  and  a13534a );
 a105a <=( a13525a  and  a13514a );
 a106a <=( a13505a  and  a13494a );
 a107a <=( a13485a  and  a13474a );
 a108a <=( a13465a  and  a13454a );
 a109a <=( a13445a  and  a13434a );
 a110a <=( a13425a  and  a13414a );
 a111a <=( a13405a  and  a13394a );
 a112a <=( a13385a  and  a13374a );
 a113a <=( a13365a  and  a13354a );
 a114a <=( a13345a  and  a13334a );
 a115a <=( a13325a  and  a13314a );
 a116a <=( a13305a  and  a13294a );
 a117a <=( a13285a  and  a13274a );
 a118a <=( a13265a  and  a13254a );
 a119a <=( a13245a  and  a13234a );
 a120a <=( a13225a  and  a13214a );
 a121a <=( a13205a  and  a13194a );
 a122a <=( a13185a  and  a13174a );
 a123a <=( a13165a  and  a13154a );
 a124a <=( a13145a  and  a13134a );
 a125a <=( a13125a  and  a13114a );
 a126a <=( a13105a  and  a13094a );
 a127a <=( a13085a  and  a13074a );
 a128a <=( a13065a  and  a13054a );
 a129a <=( a13045a  and  a13034a );
 a130a <=( a13025a  and  a13014a );
 a131a <=( a13005a  and  a12994a );
 a132a <=( a12985a  and  a12974a );
 a133a <=( a12965a  and  a12954a );
 a134a <=( a12945a  and  a12934a );
 a135a <=( a12925a  and  a12914a );
 a136a <=( a12905a  and  a12894a );
 a137a <=( a12885a  and  a12874a );
 a138a <=( a12865a  and  a12854a );
 a139a <=( a12845a  and  a12834a );
 a140a <=( a12825a  and  a12814a );
 a141a <=( a12805a  and  a12794a );
 a142a <=( a12785a  and  a12774a );
 a143a <=( a12765a  and  a12754a );
 a144a <=( a12745a  and  a12734a );
 a145a <=( a12725a  and  a12714a );
 a146a <=( a12705a  and  a12694a );
 a147a <=( a12685a  and  a12674a );
 a148a <=( a12665a  and  a12654a );
 a149a <=( a12645a  and  a12634a );
 a150a <=( a12625a  and  a12614a );
 a151a <=( a12605a  and  a12594a );
 a152a <=( a12585a  and  a12574a );
 a153a <=( a12565a  and  a12554a );
 a154a <=( a12545a  and  a12534a );
 a155a <=( a12525a  and  a12514a );
 a156a <=( a12505a  and  a12494a );
 a157a <=( a12485a  and  a12474a );
 a158a <=( a12465a  and  a12454a );
 a159a <=( a12445a  and  a12434a );
 a160a <=( a12425a  and  a12414a );
 a161a <=( a12405a  and  a12394a );
 a162a <=( a12385a  and  a12374a );
 a163a <=( a12365a  and  a12354a );
 a164a <=( a12345a  and  a12334a );
 a165a <=( a12325a  and  a12314a );
 a166a <=( a12305a  and  a12294a );
 a167a <=( a12285a  and  a12274a );
 a168a <=( a12265a  and  a12254a );
 a169a <=( a12245a  and  a12234a );
 a170a <=( a12225a  and  a12214a );
 a171a <=( a12205a  and  a12194a );
 a172a <=( a12185a  and  a12174a );
 a173a <=( a12165a  and  a12154a );
 a174a <=( a12145a  and  a12134a );
 a175a <=( a12125a  and  a12114a );
 a176a <=( a12105a  and  a12094a );
 a177a <=( a12085a  and  a12074a );
 a178a <=( a12065a  and  a12054a );
 a179a <=( a12045a  and  a12034a );
 a180a <=( a12025a  and  a12014a );
 a181a <=( a12005a  and  a11994a );
 a182a <=( a11985a  and  a11974a );
 a183a <=( a11965a  and  a11954a );
 a184a <=( a11945a  and  a11934a );
 a185a <=( a11925a  and  a11914a );
 a186a <=( a11905a  and  a11894a );
 a187a <=( a11885a  and  a11874a );
 a188a <=( a11865a  and  a11854a );
 a189a <=( a11845a  and  a11834a );
 a190a <=( a11825a  and  a11814a );
 a191a <=( a11805a  and  a11794a );
 a192a <=( a11785a  and  a11774a );
 a193a <=( a11765a  and  a11754a );
 a194a <=( a11745a  and  a11734a );
 a195a <=( a11725a  and  a11714a );
 a196a <=( a11705a  and  a11694a );
 a197a <=( a11685a  and  a11674a );
 a198a <=( a11665a  and  a11654a );
 a199a <=( a11645a  and  a11634a );
 a200a <=( a11625a  and  a11614a );
 a201a <=( a11605a  and  a11594a );
 a202a <=( a11585a  and  a11574a );
 a203a <=( a11565a  and  a11554a );
 a204a <=( a11545a  and  a11534a );
 a205a <=( a11525a  and  a11514a );
 a206a <=( a11505a  and  a11494a );
 a207a <=( a11485a  and  a11474a );
 a208a <=( a11465a  and  a11454a );
 a209a <=( a11445a  and  a11434a );
 a210a <=( a11425a  and  a11414a );
 a211a <=( a11405a  and  a11394a );
 a212a <=( a11385a  and  a11374a );
 a213a <=( a11365a  and  a11354a );
 a214a <=( a11345a  and  a11334a );
 a215a <=( a11325a  and  a11314a );
 a216a <=( a11305a  and  a11294a );
 a217a <=( a11285a  and  a11274a );
 a218a <=( a11265a  and  a11254a );
 a219a <=( a11245a  and  a11234a );
 a220a <=( a11225a  and  a11214a );
 a221a <=( a11205a  and  a11194a );
 a222a <=( a11185a  and  a11174a );
 a223a <=( a11165a  and  a11154a );
 a224a <=( a11145a  and  a11134a );
 a225a <=( a11125a  and  a11114a );
 a226a <=( a11105a  and  a11094a );
 a227a <=( a11085a  and  a11074a );
 a228a <=( a11065a  and  a11054a );
 a229a <=( a11045a  and  a11034a );
 a230a <=( a11025a  and  a11014a );
 a231a <=( a11005a  and  a10994a );
 a232a <=( a10985a  and  a10974a );
 a233a <=( a10965a  and  a10954a );
 a234a <=( a10945a  and  a10934a );
 a235a <=( a10925a  and  a10914a );
 a236a <=( a10905a  and  a10894a );
 a237a <=( a10885a  and  a10874a );
 a238a <=( a10865a  and  a10854a );
 a239a <=( a10845a  and  a10834a );
 a240a <=( a10825a  and  a10814a );
 a241a <=( a10805a  and  a10794a );
 a242a <=( a10785a  and  a10774a );
 a243a <=( a10765a  and  a10754a );
 a244a <=( a10745a  and  a10734a );
 a245a <=( a10725a  and  a10714a );
 a246a <=( a10705a  and  a10694a );
 a247a <=( a10685a  and  a10674a );
 a248a <=( a10665a  and  a10654a );
 a249a <=( a10645a  and  a10634a );
 a250a <=( a10625a  and  a10614a );
 a251a <=( a10605a  and  a10594a );
 a252a <=( a10585a  and  a10574a );
 a253a <=( a10565a  and  a10554a );
 a254a <=( a10545a  and  a10534a );
 a255a <=( a10525a  and  a10514a );
 a256a <=( a10505a  and  a10494a );
 a257a <=( a10485a  and  a10474a );
 a258a <=( a10465a  and  a10454a );
 a259a <=( a10445a  and  a10434a );
 a260a <=( a10425a  and  a10414a );
 a261a <=( a10405a  and  a10394a );
 a262a <=( a10385a  and  a10374a );
 a263a <=( a10365a  and  a10354a );
 a264a <=( a10345a  and  a10334a );
 a265a <=( a10325a  and  a10316a );
 a266a <=( a10307a  and  a10298a );
 a267a <=( a10289a  and  a10280a );
 a268a <=( a10271a  and  a10262a );
 a269a <=( a10253a  and  a10244a );
 a270a <=( a10235a  and  a10226a );
 a271a <=( a10217a  and  a10208a );
 a272a <=( a10199a  and  a10190a );
 a273a <=( a10181a  and  a10172a );
 a274a <=( a10163a  and  a10154a );
 a275a <=( a10145a  and  a10136a );
 a276a <=( a10127a  and  a10118a );
 a277a <=( a10109a  and  a10100a );
 a278a <=( a10091a  and  a10082a );
 a279a <=( a10073a  and  a10064a );
 a280a <=( a10055a  and  a10046a );
 a281a <=( a10037a  and  a10028a );
 a282a <=( a10019a  and  a10010a );
 a283a <=( a10001a  and  a9992a );
 a284a <=( a9983a  and  a9974a );
 a285a <=( a9965a  and  a9956a );
 a286a <=( a9947a  and  a9938a );
 a287a <=( a9929a  and  a9920a );
 a288a <=( a9911a  and  a9902a );
 a289a <=( a9893a  and  a9884a );
 a290a <=( a9875a  and  a9866a );
 a291a <=( a9857a  and  a9848a );
 a292a <=( a9839a  and  a9830a );
 a293a <=( a9821a  and  a9812a );
 a294a <=( a9803a  and  a9794a );
 a295a <=( a9785a  and  a9776a );
 a296a <=( a9767a  and  a9758a );
 a297a <=( a9749a  and  a9740a );
 a298a <=( a9731a  and  a9722a );
 a299a <=( a9713a  and  a9704a );
 a300a <=( a9695a  and  a9686a );
 a301a <=( a9677a  and  a9668a );
 a302a <=( a9659a  and  a9650a );
 a303a <=( a9641a  and  a9632a );
 a304a <=( a9623a  and  a9614a );
 a305a <=( a9605a  and  a9596a );
 a306a <=( a9587a  and  a9578a );
 a307a <=( a9569a  and  a9560a );
 a308a <=( a9551a  and  a9542a );
 a309a <=( a9533a  and  a9524a );
 a310a <=( a9515a  and  a9506a );
 a311a <=( a9497a  and  a9488a );
 a312a <=( a9479a  and  a9470a );
 a313a <=( a9461a  and  a9452a );
 a314a <=( a9443a  and  a9434a );
 a315a <=( a9425a  and  a9416a );
 a316a <=( a9407a  and  a9398a );
 a317a <=( a9389a  and  a9380a );
 a318a <=( a9371a  and  a9362a );
 a319a <=( a9353a  and  a9344a );
 a320a <=( a9335a  and  a9326a );
 a321a <=( a9317a  and  a9308a );
 a322a <=( a9299a  and  a9290a );
 a323a <=( a9281a  and  a9272a );
 a324a <=( a9263a  and  a9254a );
 a325a <=( a9245a  and  a9236a );
 a326a <=( a9227a  and  a9218a );
 a327a <=( a9209a  and  a9200a );
 a328a <=( a9191a  and  a9182a );
 a329a <=( a9173a  and  a9164a );
 a330a <=( a9155a  and  a9146a );
 a331a <=( a9137a  and  a9128a );
 a332a <=( a9119a  and  a9110a );
 a333a <=( a9101a  and  a9092a );
 a334a <=( a9083a  and  a9074a );
 a335a <=( a9065a  and  a9056a );
 a336a <=( a9047a  and  a9038a );
 a337a <=( a9029a  and  a9020a );
 a338a <=( a9011a  and  a9002a );
 a339a <=( a8993a  and  a8984a );
 a340a <=( a8975a  and  a8966a );
 a341a <=( a8957a  and  a8948a );
 a342a <=( a8939a  and  a8930a );
 a343a <=( a8921a  and  a8912a );
 a344a <=( a8903a  and  a8894a );
 a345a <=( a8885a  and  a8876a );
 a346a <=( a8867a  and  a8858a );
 a347a <=( a8849a  and  a8840a );
 a348a <=( a8831a  and  a8822a );
 a349a <=( a8813a  and  a8804a );
 a350a <=( a8795a  and  a8786a );
 a351a <=( a8777a  and  a8768a );
 a352a <=( a8759a  and  a8750a );
 a353a <=( a8741a  and  a8732a );
 a354a <=( a8723a  and  a8714a );
 a355a <=( a8705a  and  a8696a );
 a356a <=( a8687a  and  a8678a );
 a357a <=( a8669a  and  a8660a );
 a358a <=( a8651a  and  a8642a );
 a359a <=( a8633a  and  a8624a );
 a360a <=( a8615a  and  a8606a );
 a361a <=( a8597a  and  a8588a );
 a362a <=( a8579a  and  a8570a );
 a363a <=( a8561a  and  a8552a );
 a364a <=( a8543a  and  a8534a );
 a365a <=( a8525a  and  a8516a );
 a366a <=( a8507a  and  a8498a );
 a367a <=( a8489a  and  a8480a );
 a368a <=( a8471a  and  a8462a );
 a369a <=( a8453a  and  a8444a );
 a370a <=( a8435a  and  a8426a );
 a371a <=( a8417a  and  a8408a );
 a372a <=( a8399a  and  a8390a );
 a373a <=( a8381a  and  a8372a );
 a374a <=( a8363a  and  a8354a );
 a375a <=( a8345a  and  a8336a );
 a376a <=( a8327a  and  a8318a );
 a377a <=( a8309a  and  a8300a );
 a378a <=( a8291a  and  a8282a );
 a379a <=( a8273a  and  a8264a );
 a380a <=( a8255a  and  a8246a );
 a381a <=( a8237a  and  a8228a );
 a382a <=( a8219a  and  a8210a );
 a383a <=( a8201a  and  a8192a );
 a384a <=( a8183a  and  a8174a );
 a385a <=( a8165a  and  a8156a );
 a386a <=( a8147a  and  a8138a );
 a387a <=( a8129a  and  a8120a );
 a388a <=( a8111a  and  a8102a );
 a389a <=( a8093a  and  a8084a );
 a390a <=( a8075a  and  a8066a );
 a391a <=( a8057a  and  a8048a );
 a392a <=( a8039a  and  a8030a );
 a393a <=( a8021a  and  a8012a );
 a394a <=( a8003a  and  a7994a );
 a395a <=( a7985a  and  a7976a );
 a396a <=( a7967a  and  a7958a );
 a397a <=( a7949a  and  a7940a );
 a398a <=( a7931a  and  a7922a );
 a399a <=( a7913a  and  a7904a );
 a400a <=( a7895a  and  a7886a );
 a401a <=( a7877a  and  a7868a );
 a402a <=( a7859a  and  a7850a );
 a403a <=( a7841a  and  a7832a );
 a404a <=( a7823a  and  a7814a );
 a405a <=( a7805a  and  a7796a );
 a406a <=( a7787a  and  a7778a );
 a407a <=( a7769a  and  a7760a );
 a408a <=( a7751a  and  a7742a );
 a409a <=( a7733a  and  a7724a );
 a410a <=( a7715a  and  a7706a );
 a411a <=( a7697a  and  a7688a );
 a412a <=( a7679a  and  a7670a );
 a413a <=( a7661a  and  a7652a );
 a414a <=( a7643a  and  a7634a );
 a415a <=( a7625a  and  a7616a );
 a416a <=( a7607a  and  a7598a );
 a417a <=( a7589a  and  a7580a );
 a418a <=( a7571a  and  a7562a );
 a419a <=( a7553a  and  a7544a );
 a420a <=( a7535a  and  a7526a );
 a421a <=( a7517a  and  a7508a );
 a422a <=( a7499a  and  a7490a );
 a423a <=( a7481a  and  a7472a );
 a424a <=( a7463a  and  a7454a );
 a425a <=( a7445a  and  a7436a );
 a426a <=( a7427a  and  a7418a );
 a427a <=( a7409a  and  a7400a );
 a428a <=( a7391a  and  a7382a );
 a429a <=( a7373a  and  a7364a );
 a430a <=( a7355a  and  a7346a );
 a431a <=( a7337a  and  a7328a );
 a432a <=( a7319a  and  a7310a );
 a433a <=( a7301a  and  a7292a );
 a434a <=( a7283a  and  a7274a );
 a435a <=( a7265a  and  a7256a );
 a436a <=( a7247a  and  a7238a );
 a437a <=( a7229a  and  a7220a );
 a438a <=( a7211a  and  a7202a );
 a439a <=( a7193a  and  a7184a );
 a440a <=( a7175a  and  a7166a );
 a441a <=( a7157a  and  a7148a );
 a442a <=( a7139a  and  a7130a );
 a443a <=( a7121a  and  a7112a );
 a444a <=( a7103a  and  a7094a );
 a445a <=( a7085a  and  a7076a );
 a446a <=( a7067a  and  a7058a );
 a447a <=( a7049a  and  a7040a );
 a448a <=( a7031a  and  a7022a );
 a449a <=( a7013a  and  a7004a );
 a450a <=( a6995a  and  a6986a );
 a451a <=( a6977a  and  a6968a );
 a452a <=( a6959a  and  a6950a );
 a453a <=( a6941a  and  a6932a );
 a454a <=( a6923a  and  a6914a );
 a455a <=( a6905a  and  a6896a );
 a456a <=( a6887a  and  a6878a );
 a457a <=( a6869a  and  a6860a );
 a458a <=( a6851a  and  a6842a );
 a459a <=( a6833a  and  a6824a );
 a460a <=( a6815a  and  a6806a );
 a461a <=( a6797a  and  a6788a );
 a462a <=( a6779a  and  a6770a );
 a463a <=( a6761a  and  a6752a );
 a464a <=( a6743a  and  a6734a );
 a465a <=( a6725a  and  a6716a );
 a466a <=( a6707a  and  a6698a );
 a467a <=( a6689a  and  a6680a );
 a468a <=( a6671a  and  a6662a );
 a469a <=( a6653a  and  a6644a );
 a470a <=( a6635a  and  a6626a );
 a471a <=( a6617a  and  a6608a );
 a472a <=( a6599a  and  a6590a );
 a473a <=( a6581a  and  a6572a );
 a474a <=( a6565a  and  a6556a );
 a475a <=( a6549a  and  a6540a );
 a476a <=( a6533a  and  a6524a );
 a477a <=( a6517a  and  a6508a );
 a478a <=( a6501a  and  a6492a );
 a479a <=( a6485a  and  a6476a );
 a480a <=( a6469a  and  a6460a );
 a481a <=( a6453a  and  a6444a );
 a482a <=( a6437a  and  a6428a );
 a483a <=( a6421a  and  a6412a );
 a484a <=( a6405a  and  a6396a );
 a485a <=( a6389a  and  a6380a );
 a486a <=( a6373a  and  a6364a );
 a487a <=( a6357a  and  a6348a );
 a488a <=( a6341a  and  a6332a );
 a489a <=( a6325a  and  a6316a );
 a490a <=( a6309a  and  a6300a );
 a491a <=( a6293a  and  a6284a );
 a492a <=( a6277a  and  a6268a );
 a493a <=( a6261a  and  a6252a );
 a494a <=( a6245a  and  a6236a );
 a495a <=( a6229a  and  a6220a );
 a496a <=( a6213a  and  a6204a );
 a497a <=( a6197a  and  a6188a );
 a498a <=( a6181a  and  a6172a );
 a499a <=( a6165a  and  a6156a );
 a500a <=( a6149a  and  a6140a );
 a501a <=( a6133a  and  a6124a );
 a502a <=( a6117a  and  a6108a );
 a503a <=( a6101a  and  a6092a );
 a504a <=( a6085a  and  a6076a );
 a505a <=( a6069a  and  a6060a );
 a506a <=( a6053a  and  a6044a );
 a507a <=( a6037a  and  a6028a );
 a508a <=( a6021a  and  a6012a );
 a509a <=( a6005a  and  a5996a );
 a510a <=( a5989a  and  a5980a );
 a511a <=( a5973a  and  a5964a );
 a512a <=( a5957a  and  a5948a );
 a513a <=( a5941a  and  a5932a );
 a514a <=( a5925a  and  a5916a );
 a515a <=( a5909a  and  a5900a );
 a516a <=( a5893a  and  a5884a );
 a517a <=( a5877a  and  a5868a );
 a518a <=( a5861a  and  a5852a );
 a519a <=( a5845a  and  a5836a );
 a520a <=( a5829a  and  a5820a );
 a521a <=( a5813a  and  a5804a );
 a522a <=( a5797a  and  a5788a );
 a523a <=( a5781a  and  a5772a );
 a524a <=( a5765a  and  a5756a );
 a525a <=( a5749a  and  a5740a );
 a526a <=( a5733a  and  a5724a );
 a527a <=( a5717a  and  a5708a );
 a528a <=( a5701a  and  a5692a );
 a529a <=( a5685a  and  a5676a );
 a530a <=( a5669a  and  a5660a );
 a531a <=( a5653a  and  a5644a );
 a532a <=( a5637a  and  a5628a );
 a533a <=( a5621a  and  a5612a );
 a534a <=( a5605a  and  a5596a );
 a535a <=( a5589a  and  a5580a );
 a536a <=( a5573a  and  a5564a );
 a537a <=( a5557a  and  a5548a );
 a538a <=( a5541a  and  a5532a );
 a539a <=( a5525a  and  a5516a );
 a540a <=( a5509a  and  a5500a );
 a541a <=( a5493a  and  a5484a );
 a542a <=( a5477a  and  a5468a );
 a543a <=( a5461a  and  a5452a );
 a544a <=( a5445a  and  a5436a );
 a545a <=( a5429a  and  a5420a );
 a546a <=( a5413a  and  a5404a );
 a547a <=( a5397a  and  a5388a );
 a548a <=( a5381a  and  a5372a );
 a549a <=( a5365a  and  a5356a );
 a550a <=( a5349a  and  a5340a );
 a551a <=( a5333a  and  a5324a );
 a552a <=( a5317a  and  a5308a );
 a553a <=( a5301a  and  a5292a );
 a554a <=( a5285a  and  a5276a );
 a555a <=( a5269a  and  a5260a );
 a556a <=( a5253a  and  a5244a );
 a557a <=( a5237a  and  a5228a );
 a558a <=( a5221a  and  a5212a );
 a559a <=( a5205a  and  a5196a );
 a560a <=( a5189a  and  a5180a );
 a561a <=( a5173a  and  a5164a );
 a562a <=( a5157a  and  a5148a );
 a563a <=( a5141a  and  a5132a );
 a564a <=( a5125a  and  a5116a );
 a565a <=( a5109a  and  a5100a );
 a566a <=( a5093a  and  a5084a );
 a567a <=( a5077a  and  a5068a );
 a568a <=( a5061a  and  a5052a );
 a569a <=( a5045a  and  a5036a );
 a570a <=( a5029a  and  a5020a );
 a571a <=( a5013a  and  a5004a );
 a572a <=( a4997a  and  a4988a );
 a573a <=( a4981a  and  a4972a );
 a574a <=( a4965a  and  a4956a );
 a575a <=( a4949a  and  a4940a );
 a576a <=( a4933a  and  a4924a );
 a577a <=( a4917a  and  a4908a );
 a578a <=( a4901a  and  a4892a );
 a579a <=( a4885a  and  a4876a );
 a580a <=( a4869a  and  a4860a );
 a581a <=( a4853a  and  a4844a );
 a582a <=( a4837a  and  a4828a );
 a583a <=( a4821a  and  a4812a );
 a584a <=( a4805a  and  a4796a );
 a585a <=( a4789a  and  a4780a );
 a586a <=( a4773a  and  a4764a );
 a587a <=( a4757a  and  a4748a );
 a588a <=( a4741a  and  a4732a );
 a589a <=( a4725a  and  a4716a );
 a590a <=( a4709a  and  a4700a );
 a591a <=( a4693a  and  a4684a );
 a592a <=( a4677a  and  a4668a );
 a593a <=( a4661a  and  a4652a );
 a594a <=( a4645a  and  a4636a );
 a595a <=( a4629a  and  a4620a );
 a596a <=( a4613a  and  a4604a );
 a597a <=( a4597a  and  a4588a );
 a598a <=( a4581a  and  a4572a );
 a599a <=( a4565a  and  a4556a );
 a600a <=( a4549a  and  a4540a );
 a601a <=( a4533a  and  a4524a );
 a602a <=( a4517a  and  a4508a );
 a603a <=( a4501a  and  a4492a );
 a604a <=( a4485a  and  a4476a );
 a605a <=( a4469a  and  a4460a );
 a606a <=( a4453a  and  a4444a );
 a607a <=( a4437a  and  a4428a );
 a608a <=( a4421a  and  a4412a );
 a609a <=( a4405a  and  a4396a );
 a610a <=( a4389a  and  a4380a );
 a611a <=( a4373a  and  a4364a );
 a612a <=( a4357a  and  a4348a );
 a613a <=( a4341a  and  a4332a );
 a614a <=( a4325a  and  a4316a );
 a615a <=( a4309a  and  a4300a );
 a616a <=( a4293a  and  a4284a );
 a617a <=( a4277a  and  a4268a );
 a618a <=( a4261a  and  a4252a );
 a619a <=( a4245a  and  a4236a );
 a620a <=( a4229a  and  a4220a );
 a621a <=( a4213a  and  a4204a );
 a622a <=( a4197a  and  a4188a );
 a623a <=( a4181a  and  a4172a );
 a624a <=( a4165a  and  a4156a );
 a625a <=( a4149a  and  a4140a );
 a626a <=( a4133a  and  a4124a );
 a627a <=( a4117a  and  a4108a );
 a628a <=( a4101a  and  a4092a );
 a629a <=( a4085a  and  a4076a );
 a630a <=( a4069a  and  a4060a );
 a631a <=( a4053a  and  a4044a );
 a632a <=( a4037a  and  a4028a );
 a633a <=( a4021a  and  a4012a );
 a634a <=( a4005a  and  a3996a );
 a635a <=( a3989a  and  a3980a );
 a636a <=( a3973a  and  a3964a );
 a637a <=( a3957a  and  a3950a );
 a638a <=( a3943a  and  a3936a );
 a639a <=( a3929a  and  a3922a );
 a640a <=( a3915a  and  a3908a );
 a641a <=( a3901a  and  a3894a );
 a642a <=( a3887a  and  a3880a );
 a643a <=( a3873a  and  a3866a );
 a644a <=( a3859a  and  a3852a );
 a645a <=( a3845a  and  a3838a );
 a646a <=( a3831a  and  a3824a );
 a647a <=( a3817a  and  a3810a );
 a648a <=( a3803a  and  a3796a );
 a649a <=( a3789a  and  a3782a );
 a650a <=( a3775a  and  a3768a );
 a651a <=( a3761a  and  a3754a );
 a652a <=( a3747a  and  a3740a );
 a653a <=( a3733a  and  a3726a );
 a654a <=( a3719a  and  a3712a );
 a655a <=( a3705a  and  a3698a );
 a656a <=( a3691a  and  a3684a );
 a657a <=( a3677a  and  a3670a );
 a658a <=( a3663a  and  a3656a );
 a659a <=( a3649a  and  a3642a );
 a660a <=( a3635a  and  a3628a );
 a661a <=( a3621a  and  a3614a );
 a662a <=( a3607a  and  a3600a );
 a663a <=( a3593a  and  a3586a );
 a664a <=( a3579a  and  a3572a );
 a665a <=( a3565a  and  a3558a );
 a666a <=( a3551a  and  a3544a );
 a667a <=( a3537a  and  a3530a );
 a668a <=( a3523a  and  a3516a );
 a669a <=( a3509a  and  a3502a );
 a670a <=( a3495a  and  a3488a );
 a671a <=( a3481a  and  a3474a );
 a672a <=( a3467a  and  a3460a );
 a673a <=( a3453a  and  a3446a );
 a674a <=( a3439a  and  a3432a );
 a675a <=( a3425a  and  a3418a );
 a676a <=( a3411a  and  a3404a );
 a677a <=( a3397a  and  a3390a );
 a678a <=( a3383a  and  a3376a );
 a679a <=( a3369a  and  a3362a );
 a680a <=( a3355a  and  a3348a );
 a681a <=( a3341a  and  a3334a );
 a682a <=( a3327a  and  a3320a );
 a683a <=( a3313a  and  a3306a );
 a684a <=( a3299a  and  a3292a );
 a685a <=( a3285a  and  a3278a );
 a686a <=( a3271a  and  a3264a );
 a687a <=( a3257a  and  a3250a );
 a688a <=( a3243a  and  a3236a );
 a689a <=( a3229a  and  a3222a );
 a690a <=( a3215a  and  a3208a );
 a691a <=( a3201a  and  a3194a );
 a692a <=( a3187a  and  a3180a );
 a693a <=( a3173a  and  a3166a );
 a694a <=( a3159a  and  a3152a );
 a695a <=( a3145a  and  a3138a );
 a696a <=( a3131a  and  a3124a );
 a697a <=( a3117a  and  a3110a );
 a698a <=( a3103a  and  a3096a );
 a699a <=( a3089a  and  a3082a );
 a700a <=( a3075a  and  a3068a );
 a701a <=( a3061a  and  a3054a );
 a702a <=( a3047a  and  a3040a );
 a703a <=( a3033a  and  a3026a );
 a704a <=( a3019a  and  a3012a );
 a705a <=( a3005a  and  a2998a );
 a706a <=( a2991a  and  a2984a );
 a707a <=( a2977a  and  a2970a );
 a708a <=( a2963a  and  a2956a );
 a709a <=( a2949a  and  a2942a );
 a710a <=( a2935a  and  a2928a );
 a711a <=( a2921a  and  a2914a );
 a712a <=( a2907a  and  a2900a );
 a713a <=( a2893a  and  a2886a );
 a714a <=( a2879a  and  a2872a );
 a715a <=( a2865a  and  a2858a );
 a716a <=( a2851a  and  a2844a );
 a717a <=( a2837a  and  a2830a );
 a718a <=( a2823a  and  a2816a );
 a719a <=( a2809a  and  a2802a );
 a720a <=( a2795a  and  a2788a );
 a721a <=( a2781a  and  a2774a );
 a722a <=( a2769a  and  a2762a );
 a723a <=( a2757a  and  a2750a );
 a724a <=( a2745a  and  a2738a );
 a725a <=( a2733a  and  a2726a );
 a726a <=( a2721a  and  a2714a );
 a727a <=( a2709a  and  a2702a );
 a728a <=( a2697a  and  a2690a );
 a729a <=( a2685a  and  a2678a );
 a730a <=( a2673a  and  a2666a );
 a731a <=( a2661a  and  a2654a );
 a732a <=( a2649a  and  a2642a );
 a733a <=( a2637a  and  a2630a );
 a734a <=( a2625a  and  a2618a );
 a735a <=( a2613a  and  a2606a );
 a736a <=( a2601a  and  a2594a );
 a737a <=( a2589a  and  a2582a );
 a738a <=( a2577a  and  a2570a );
 a739a <=( a2565a  and  a2558a );
 a740a <=( a2553a  and  a2546a );
 a741a <=( a2541a  and  a2534a );
 a742a <=( a2529a  and  a2522a );
 a743a <=( a2517a  and  a2510a );
 a744a <=( a2505a  and  a2498a );
 a745a <=( a2493a  and  a2486a );
 a746a <=( a2481a  and  a2474a );
 a747a <=( a2469a  and  a2462a );
 a748a <=( a2457a  and  a2450a );
 a749a <=( a2445a  and  a2440a );
 a750a <=( a2435a  and  a2430a );
 a751a <=( a2425a  and  a2420a );
 a752a <=( a2415a  and  a2410a );
 a753a <=( a2405a  and  a2400a );
 a754a <=( a2395a  and  a2390a );
 a755a <=( a2385a  and  a2380a );
 a756a <=( a2375a  and  a2370a );
 a757a <=( a2365a  and  a2360a );
 a758a <=( a2355a  and  a2350a );
 a759a <=( a2345a  and  a2340a );
 a760a <=( a2337a  and  a2332a );
 a761a <=( a2329a  and  a2324a );
 a762a <=( a2321a  and  a2316a );
 a763a <=( a2313a  and  a2308a );
 a764a <=( a2305a  and  a2302a );
 a765a <=( a2299a  and  a2296a );
 a768a <=( a764a ) or ( a765a );
 a772a <=( a761a ) or ( a762a );
 a773a <=( a763a ) or ( a772a );
 a774a <=( a773a ) or ( a768a );
 a778a <=( a758a ) or ( a759a );
 a779a <=( a760a ) or ( a778a );
 a783a <=( a755a ) or ( a756a );
 a784a <=( a757a ) or ( a783a );
 a785a <=( a784a ) or ( a779a );
 a786a <=( a785a ) or ( a774a );
 a790a <=( a752a ) or ( a753a );
 a791a <=( a754a ) or ( a790a );
 a795a <=( a749a ) or ( a750a );
 a796a <=( a751a ) or ( a795a );
 a797a <=( a796a ) or ( a791a );
 a801a <=( a746a ) or ( a747a );
 a802a <=( a748a ) or ( a801a );
 a806a <=( a743a ) or ( a744a );
 a807a <=( a745a ) or ( a806a );
 a808a <=( a807a ) or ( a802a );
 a809a <=( a808a ) or ( a797a );
 a810a <=( a809a ) or ( a786a );
 a814a <=( a740a ) or ( a741a );
 a815a <=( a742a ) or ( a814a );
 a819a <=( a737a ) or ( a738a );
 a820a <=( a739a ) or ( a819a );
 a821a <=( a820a ) or ( a815a );
 a825a <=( a734a ) or ( a735a );
 a826a <=( a736a ) or ( a825a );
 a830a <=( a731a ) or ( a732a );
 a831a <=( a733a ) or ( a830a );
 a832a <=( a831a ) or ( a826a );
 a833a <=( a832a ) or ( a821a );
 a837a <=( a728a ) or ( a729a );
 a838a <=( a730a ) or ( a837a );
 a842a <=( a725a ) or ( a726a );
 a843a <=( a727a ) or ( a842a );
 a844a <=( a843a ) or ( a838a );
 a848a <=( a722a ) or ( a723a );
 a849a <=( a724a ) or ( a848a );
 a853a <=( a719a ) or ( a720a );
 a854a <=( a721a ) or ( a853a );
 a855a <=( a854a ) or ( a849a );
 a856a <=( a855a ) or ( a844a );
 a857a <=( a856a ) or ( a833a );
 a858a <=( a857a ) or ( a810a );
 a862a <=( a716a ) or ( a717a );
 a863a <=( a718a ) or ( a862a );
 a867a <=( a713a ) or ( a714a );
 a868a <=( a715a ) or ( a867a );
 a869a <=( a868a ) or ( a863a );
 a873a <=( a710a ) or ( a711a );
 a874a <=( a712a ) or ( a873a );
 a878a <=( a707a ) or ( a708a );
 a879a <=( a709a ) or ( a878a );
 a880a <=( a879a ) or ( a874a );
 a881a <=( a880a ) or ( a869a );
 a885a <=( a704a ) or ( a705a );
 a886a <=( a706a ) or ( a885a );
 a890a <=( a701a ) or ( a702a );
 a891a <=( a703a ) or ( a890a );
 a892a <=( a891a ) or ( a886a );
 a896a <=( a698a ) or ( a699a );
 a897a <=( a700a ) or ( a896a );
 a901a <=( a695a ) or ( a696a );
 a902a <=( a697a ) or ( a901a );
 a903a <=( a902a ) or ( a897a );
 a904a <=( a903a ) or ( a892a );
 a905a <=( a904a ) or ( a881a );
 a909a <=( a692a ) or ( a693a );
 a910a <=( a694a ) or ( a909a );
 a914a <=( a689a ) or ( a690a );
 a915a <=( a691a ) or ( a914a );
 a916a <=( a915a ) or ( a910a );
 a920a <=( a686a ) or ( a687a );
 a921a <=( a688a ) or ( a920a );
 a925a <=( a683a ) or ( a684a );
 a926a <=( a685a ) or ( a925a );
 a927a <=( a926a ) or ( a921a );
 a928a <=( a927a ) or ( a916a );
 a932a <=( a680a ) or ( a681a );
 a933a <=( a682a ) or ( a932a );
 a937a <=( a677a ) or ( a678a );
 a938a <=( a679a ) or ( a937a );
 a939a <=( a938a ) or ( a933a );
 a943a <=( a674a ) or ( a675a );
 a944a <=( a676a ) or ( a943a );
 a948a <=( a671a ) or ( a672a );
 a949a <=( a673a ) or ( a948a );
 a950a <=( a949a ) or ( a944a );
 a951a <=( a950a ) or ( a939a );
 a952a <=( a951a ) or ( a928a );
 a953a <=( a952a ) or ( a905a );
 a954a <=( a953a ) or ( a858a );
 a958a <=( a668a ) or ( a669a );
 a959a <=( a670a ) or ( a958a );
 a963a <=( a665a ) or ( a666a );
 a964a <=( a667a ) or ( a963a );
 a965a <=( a964a ) or ( a959a );
 a969a <=( a662a ) or ( a663a );
 a970a <=( a664a ) or ( a969a );
 a974a <=( a659a ) or ( a660a );
 a975a <=( a661a ) or ( a974a );
 a976a <=( a975a ) or ( a970a );
 a977a <=( a976a ) or ( a965a );
 a981a <=( a656a ) or ( a657a );
 a982a <=( a658a ) or ( a981a );
 a986a <=( a653a ) or ( a654a );
 a987a <=( a655a ) or ( a986a );
 a988a <=( a987a ) or ( a982a );
 a992a <=( a650a ) or ( a651a );
 a993a <=( a652a ) or ( a992a );
 a997a <=( a647a ) or ( a648a );
 a998a <=( a649a ) or ( a997a );
 a999a <=( a998a ) or ( a993a );
 a1000a <=( a999a ) or ( a988a );
 a1001a <=( a1000a ) or ( a977a );
 a1005a <=( a644a ) or ( a645a );
 a1006a <=( a646a ) or ( a1005a );
 a1010a <=( a641a ) or ( a642a );
 a1011a <=( a643a ) or ( a1010a );
 a1012a <=( a1011a ) or ( a1006a );
 a1016a <=( a638a ) or ( a639a );
 a1017a <=( a640a ) or ( a1016a );
 a1021a <=( a635a ) or ( a636a );
 a1022a <=( a637a ) or ( a1021a );
 a1023a <=( a1022a ) or ( a1017a );
 a1024a <=( a1023a ) or ( a1012a );
 a1028a <=( a632a ) or ( a633a );
 a1029a <=( a634a ) or ( a1028a );
 a1033a <=( a629a ) or ( a630a );
 a1034a <=( a631a ) or ( a1033a );
 a1035a <=( a1034a ) or ( a1029a );
 a1039a <=( a626a ) or ( a627a );
 a1040a <=( a628a ) or ( a1039a );
 a1044a <=( a623a ) or ( a624a );
 a1045a <=( a625a ) or ( a1044a );
 a1046a <=( a1045a ) or ( a1040a );
 a1047a <=( a1046a ) or ( a1035a );
 a1048a <=( a1047a ) or ( a1024a );
 a1049a <=( a1048a ) or ( a1001a );
 a1053a <=( a620a ) or ( a621a );
 a1054a <=( a622a ) or ( a1053a );
 a1058a <=( a617a ) or ( a618a );
 a1059a <=( a619a ) or ( a1058a );
 a1060a <=( a1059a ) or ( a1054a );
 a1064a <=( a614a ) or ( a615a );
 a1065a <=( a616a ) or ( a1064a );
 a1069a <=( a611a ) or ( a612a );
 a1070a <=( a613a ) or ( a1069a );
 a1071a <=( a1070a ) or ( a1065a );
 a1072a <=( a1071a ) or ( a1060a );
 a1076a <=( a608a ) or ( a609a );
 a1077a <=( a610a ) or ( a1076a );
 a1081a <=( a605a ) or ( a606a );
 a1082a <=( a607a ) or ( a1081a );
 a1083a <=( a1082a ) or ( a1077a );
 a1087a <=( a602a ) or ( a603a );
 a1088a <=( a604a ) or ( a1087a );
 a1092a <=( a599a ) or ( a600a );
 a1093a <=( a601a ) or ( a1092a );
 a1094a <=( a1093a ) or ( a1088a );
 a1095a <=( a1094a ) or ( a1083a );
 a1096a <=( a1095a ) or ( a1072a );
 a1100a <=( a596a ) or ( a597a );
 a1101a <=( a598a ) or ( a1100a );
 a1105a <=( a593a ) or ( a594a );
 a1106a <=( a595a ) or ( a1105a );
 a1107a <=( a1106a ) or ( a1101a );
 a1111a <=( a590a ) or ( a591a );
 a1112a <=( a592a ) or ( a1111a );
 a1116a <=( a587a ) or ( a588a );
 a1117a <=( a589a ) or ( a1116a );
 a1118a <=( a1117a ) or ( a1112a );
 a1119a <=( a1118a ) or ( a1107a );
 a1123a <=( a584a ) or ( a585a );
 a1124a <=( a586a ) or ( a1123a );
 a1128a <=( a581a ) or ( a582a );
 a1129a <=( a583a ) or ( a1128a );
 a1130a <=( a1129a ) or ( a1124a );
 a1134a <=( a578a ) or ( a579a );
 a1135a <=( a580a ) or ( a1134a );
 a1139a <=( a575a ) or ( a576a );
 a1140a <=( a577a ) or ( a1139a );
 a1141a <=( a1140a ) or ( a1135a );
 a1142a <=( a1141a ) or ( a1130a );
 a1143a <=( a1142a ) or ( a1119a );
 a1144a <=( a1143a ) or ( a1096a );
 a1145a <=( a1144a ) or ( a1049a );
 a1146a <=( a1145a ) or ( a954a );
 a1149a <=( a573a ) or ( a574a );
 a1153a <=( a570a ) or ( a571a );
 a1154a <=( a572a ) or ( a1153a );
 a1155a <=( a1154a ) or ( a1149a );
 a1159a <=( a567a ) or ( a568a );
 a1160a <=( a569a ) or ( a1159a );
 a1164a <=( a564a ) or ( a565a );
 a1165a <=( a566a ) or ( a1164a );
 a1166a <=( a1165a ) or ( a1160a );
 a1167a <=( a1166a ) or ( a1155a );
 a1171a <=( a561a ) or ( a562a );
 a1172a <=( a563a ) or ( a1171a );
 a1176a <=( a558a ) or ( a559a );
 a1177a <=( a560a ) or ( a1176a );
 a1178a <=( a1177a ) or ( a1172a );
 a1182a <=( a555a ) or ( a556a );
 a1183a <=( a557a ) or ( a1182a );
 a1187a <=( a552a ) or ( a553a );
 a1188a <=( a554a ) or ( a1187a );
 a1189a <=( a1188a ) or ( a1183a );
 a1190a <=( a1189a ) or ( a1178a );
 a1191a <=( a1190a ) or ( a1167a );
 a1195a <=( a549a ) or ( a550a );
 a1196a <=( a551a ) or ( a1195a );
 a1200a <=( a546a ) or ( a547a );
 a1201a <=( a548a ) or ( a1200a );
 a1202a <=( a1201a ) or ( a1196a );
 a1206a <=( a543a ) or ( a544a );
 a1207a <=( a545a ) or ( a1206a );
 a1211a <=( a540a ) or ( a541a );
 a1212a <=( a542a ) or ( a1211a );
 a1213a <=( a1212a ) or ( a1207a );
 a1214a <=( a1213a ) or ( a1202a );
 a1218a <=( a537a ) or ( a538a );
 a1219a <=( a539a ) or ( a1218a );
 a1223a <=( a534a ) or ( a535a );
 a1224a <=( a536a ) or ( a1223a );
 a1225a <=( a1224a ) or ( a1219a );
 a1229a <=( a531a ) or ( a532a );
 a1230a <=( a533a ) or ( a1229a );
 a1234a <=( a528a ) or ( a529a );
 a1235a <=( a530a ) or ( a1234a );
 a1236a <=( a1235a ) or ( a1230a );
 a1237a <=( a1236a ) or ( a1225a );
 a1238a <=( a1237a ) or ( a1214a );
 a1239a <=( a1238a ) or ( a1191a );
 a1243a <=( a525a ) or ( a526a );
 a1244a <=( a527a ) or ( a1243a );
 a1248a <=( a522a ) or ( a523a );
 a1249a <=( a524a ) or ( a1248a );
 a1250a <=( a1249a ) or ( a1244a );
 a1254a <=( a519a ) or ( a520a );
 a1255a <=( a521a ) or ( a1254a );
 a1259a <=( a516a ) or ( a517a );
 a1260a <=( a518a ) or ( a1259a );
 a1261a <=( a1260a ) or ( a1255a );
 a1262a <=( a1261a ) or ( a1250a );
 a1266a <=( a513a ) or ( a514a );
 a1267a <=( a515a ) or ( a1266a );
 a1271a <=( a510a ) or ( a511a );
 a1272a <=( a512a ) or ( a1271a );
 a1273a <=( a1272a ) or ( a1267a );
 a1277a <=( a507a ) or ( a508a );
 a1278a <=( a509a ) or ( a1277a );
 a1282a <=( a504a ) or ( a505a );
 a1283a <=( a506a ) or ( a1282a );
 a1284a <=( a1283a ) or ( a1278a );
 a1285a <=( a1284a ) or ( a1273a );
 a1286a <=( a1285a ) or ( a1262a );
 a1290a <=( a501a ) or ( a502a );
 a1291a <=( a503a ) or ( a1290a );
 a1295a <=( a498a ) or ( a499a );
 a1296a <=( a500a ) or ( a1295a );
 a1297a <=( a1296a ) or ( a1291a );
 a1301a <=( a495a ) or ( a496a );
 a1302a <=( a497a ) or ( a1301a );
 a1306a <=( a492a ) or ( a493a );
 a1307a <=( a494a ) or ( a1306a );
 a1308a <=( a1307a ) or ( a1302a );
 a1309a <=( a1308a ) or ( a1297a );
 a1313a <=( a489a ) or ( a490a );
 a1314a <=( a491a ) or ( a1313a );
 a1318a <=( a486a ) or ( a487a );
 a1319a <=( a488a ) or ( a1318a );
 a1320a <=( a1319a ) or ( a1314a );
 a1324a <=( a483a ) or ( a484a );
 a1325a <=( a485a ) or ( a1324a );
 a1329a <=( a480a ) or ( a481a );
 a1330a <=( a482a ) or ( a1329a );
 a1331a <=( a1330a ) or ( a1325a );
 a1332a <=( a1331a ) or ( a1320a );
 a1333a <=( a1332a ) or ( a1309a );
 a1334a <=( a1333a ) or ( a1286a );
 a1335a <=( a1334a ) or ( a1239a );
 a1339a <=( a477a ) or ( a478a );
 a1340a <=( a479a ) or ( a1339a );
 a1344a <=( a474a ) or ( a475a );
 a1345a <=( a476a ) or ( a1344a );
 a1346a <=( a1345a ) or ( a1340a );
 a1350a <=( a471a ) or ( a472a );
 a1351a <=( a473a ) or ( a1350a );
 a1355a <=( a468a ) or ( a469a );
 a1356a <=( a470a ) or ( a1355a );
 a1357a <=( a1356a ) or ( a1351a );
 a1358a <=( a1357a ) or ( a1346a );
 a1362a <=( a465a ) or ( a466a );
 a1363a <=( a467a ) or ( a1362a );
 a1367a <=( a462a ) or ( a463a );
 a1368a <=( a464a ) or ( a1367a );
 a1369a <=( a1368a ) or ( a1363a );
 a1373a <=( a459a ) or ( a460a );
 a1374a <=( a461a ) or ( a1373a );
 a1378a <=( a456a ) or ( a457a );
 a1379a <=( a458a ) or ( a1378a );
 a1380a <=( a1379a ) or ( a1374a );
 a1381a <=( a1380a ) or ( a1369a );
 a1382a <=( a1381a ) or ( a1358a );
 a1386a <=( a453a ) or ( a454a );
 a1387a <=( a455a ) or ( a1386a );
 a1391a <=( a450a ) or ( a451a );
 a1392a <=( a452a ) or ( a1391a );
 a1393a <=( a1392a ) or ( a1387a );
 a1397a <=( a447a ) or ( a448a );
 a1398a <=( a449a ) or ( a1397a );
 a1402a <=( a444a ) or ( a445a );
 a1403a <=( a446a ) or ( a1402a );
 a1404a <=( a1403a ) or ( a1398a );
 a1405a <=( a1404a ) or ( a1393a );
 a1409a <=( a441a ) or ( a442a );
 a1410a <=( a443a ) or ( a1409a );
 a1414a <=( a438a ) or ( a439a );
 a1415a <=( a440a ) or ( a1414a );
 a1416a <=( a1415a ) or ( a1410a );
 a1420a <=( a435a ) or ( a436a );
 a1421a <=( a437a ) or ( a1420a );
 a1425a <=( a432a ) or ( a433a );
 a1426a <=( a434a ) or ( a1425a );
 a1427a <=( a1426a ) or ( a1421a );
 a1428a <=( a1427a ) or ( a1416a );
 a1429a <=( a1428a ) or ( a1405a );
 a1430a <=( a1429a ) or ( a1382a );
 a1434a <=( a429a ) or ( a430a );
 a1435a <=( a431a ) or ( a1434a );
 a1439a <=( a426a ) or ( a427a );
 a1440a <=( a428a ) or ( a1439a );
 a1441a <=( a1440a ) or ( a1435a );
 a1445a <=( a423a ) or ( a424a );
 a1446a <=( a425a ) or ( a1445a );
 a1450a <=( a420a ) or ( a421a );
 a1451a <=( a422a ) or ( a1450a );
 a1452a <=( a1451a ) or ( a1446a );
 a1453a <=( a1452a ) or ( a1441a );
 a1457a <=( a417a ) or ( a418a );
 a1458a <=( a419a ) or ( a1457a );
 a1462a <=( a414a ) or ( a415a );
 a1463a <=( a416a ) or ( a1462a );
 a1464a <=( a1463a ) or ( a1458a );
 a1468a <=( a411a ) or ( a412a );
 a1469a <=( a413a ) or ( a1468a );
 a1473a <=( a408a ) or ( a409a );
 a1474a <=( a410a ) or ( a1473a );
 a1475a <=( a1474a ) or ( a1469a );
 a1476a <=( a1475a ) or ( a1464a );
 a1477a <=( a1476a ) or ( a1453a );
 a1481a <=( a405a ) or ( a406a );
 a1482a <=( a407a ) or ( a1481a );
 a1486a <=( a402a ) or ( a403a );
 a1487a <=( a404a ) or ( a1486a );
 a1488a <=( a1487a ) or ( a1482a );
 a1492a <=( a399a ) or ( a400a );
 a1493a <=( a401a ) or ( a1492a );
 a1497a <=( a396a ) or ( a397a );
 a1498a <=( a398a ) or ( a1497a );
 a1499a <=( a1498a ) or ( a1493a );
 a1500a <=( a1499a ) or ( a1488a );
 a1504a <=( a393a ) or ( a394a );
 a1505a <=( a395a ) or ( a1504a );
 a1509a <=( a390a ) or ( a391a );
 a1510a <=( a392a ) or ( a1509a );
 a1511a <=( a1510a ) or ( a1505a );
 a1515a <=( a387a ) or ( a388a );
 a1516a <=( a389a ) or ( a1515a );
 a1520a <=( a384a ) or ( a385a );
 a1521a <=( a386a ) or ( a1520a );
 a1522a <=( a1521a ) or ( a1516a );
 a1523a <=( a1522a ) or ( a1511a );
 a1524a <=( a1523a ) or ( a1500a );
 a1525a <=( a1524a ) or ( a1477a );
 a1526a <=( a1525a ) or ( a1430a );
 a1527a <=( a1526a ) or ( a1335a );
 a1528a <=( a1527a ) or ( a1146a );
 a1531a <=( a382a ) or ( a383a );
 a1535a <=( a379a ) or ( a380a );
 a1536a <=( a381a ) or ( a1535a );
 a1537a <=( a1536a ) or ( a1531a );
 a1541a <=( a376a ) or ( a377a );
 a1542a <=( a378a ) or ( a1541a );
 a1546a <=( a373a ) or ( a374a );
 a1547a <=( a375a ) or ( a1546a );
 a1548a <=( a1547a ) or ( a1542a );
 a1549a <=( a1548a ) or ( a1537a );
 a1553a <=( a370a ) or ( a371a );
 a1554a <=( a372a ) or ( a1553a );
 a1558a <=( a367a ) or ( a368a );
 a1559a <=( a369a ) or ( a1558a );
 a1560a <=( a1559a ) or ( a1554a );
 a1564a <=( a364a ) or ( a365a );
 a1565a <=( a366a ) or ( a1564a );
 a1569a <=( a361a ) or ( a362a );
 a1570a <=( a363a ) or ( a1569a );
 a1571a <=( a1570a ) or ( a1565a );
 a1572a <=( a1571a ) or ( a1560a );
 a1573a <=( a1572a ) or ( a1549a );
 a1577a <=( a358a ) or ( a359a );
 a1578a <=( a360a ) or ( a1577a );
 a1582a <=( a355a ) or ( a356a );
 a1583a <=( a357a ) or ( a1582a );
 a1584a <=( a1583a ) or ( a1578a );
 a1588a <=( a352a ) or ( a353a );
 a1589a <=( a354a ) or ( a1588a );
 a1593a <=( a349a ) or ( a350a );
 a1594a <=( a351a ) or ( a1593a );
 a1595a <=( a1594a ) or ( a1589a );
 a1596a <=( a1595a ) or ( a1584a );
 a1600a <=( a346a ) or ( a347a );
 a1601a <=( a348a ) or ( a1600a );
 a1605a <=( a343a ) or ( a344a );
 a1606a <=( a345a ) or ( a1605a );
 a1607a <=( a1606a ) or ( a1601a );
 a1611a <=( a340a ) or ( a341a );
 a1612a <=( a342a ) or ( a1611a );
 a1616a <=( a337a ) or ( a338a );
 a1617a <=( a339a ) or ( a1616a );
 a1618a <=( a1617a ) or ( a1612a );
 a1619a <=( a1618a ) or ( a1607a );
 a1620a <=( a1619a ) or ( a1596a );
 a1621a <=( a1620a ) or ( a1573a );
 a1625a <=( a334a ) or ( a335a );
 a1626a <=( a336a ) or ( a1625a );
 a1630a <=( a331a ) or ( a332a );
 a1631a <=( a333a ) or ( a1630a );
 a1632a <=( a1631a ) or ( a1626a );
 a1636a <=( a328a ) or ( a329a );
 a1637a <=( a330a ) or ( a1636a );
 a1641a <=( a325a ) or ( a326a );
 a1642a <=( a327a ) or ( a1641a );
 a1643a <=( a1642a ) or ( a1637a );
 a1644a <=( a1643a ) or ( a1632a );
 a1648a <=( a322a ) or ( a323a );
 a1649a <=( a324a ) or ( a1648a );
 a1653a <=( a319a ) or ( a320a );
 a1654a <=( a321a ) or ( a1653a );
 a1655a <=( a1654a ) or ( a1649a );
 a1659a <=( a316a ) or ( a317a );
 a1660a <=( a318a ) or ( a1659a );
 a1664a <=( a313a ) or ( a314a );
 a1665a <=( a315a ) or ( a1664a );
 a1666a <=( a1665a ) or ( a1660a );
 a1667a <=( a1666a ) or ( a1655a );
 a1668a <=( a1667a ) or ( a1644a );
 a1672a <=( a310a ) or ( a311a );
 a1673a <=( a312a ) or ( a1672a );
 a1677a <=( a307a ) or ( a308a );
 a1678a <=( a309a ) or ( a1677a );
 a1679a <=( a1678a ) or ( a1673a );
 a1683a <=( a304a ) or ( a305a );
 a1684a <=( a306a ) or ( a1683a );
 a1688a <=( a301a ) or ( a302a );
 a1689a <=( a303a ) or ( a1688a );
 a1690a <=( a1689a ) or ( a1684a );
 a1691a <=( a1690a ) or ( a1679a );
 a1695a <=( a298a ) or ( a299a );
 a1696a <=( a300a ) or ( a1695a );
 a1700a <=( a295a ) or ( a296a );
 a1701a <=( a297a ) or ( a1700a );
 a1702a <=( a1701a ) or ( a1696a );
 a1706a <=( a292a ) or ( a293a );
 a1707a <=( a294a ) or ( a1706a );
 a1711a <=( a289a ) or ( a290a );
 a1712a <=( a291a ) or ( a1711a );
 a1713a <=( a1712a ) or ( a1707a );
 a1714a <=( a1713a ) or ( a1702a );
 a1715a <=( a1714a ) or ( a1691a );
 a1716a <=( a1715a ) or ( a1668a );
 a1717a <=( a1716a ) or ( a1621a );
 a1721a <=( a286a ) or ( a287a );
 a1722a <=( a288a ) or ( a1721a );
 a1726a <=( a283a ) or ( a284a );
 a1727a <=( a285a ) or ( a1726a );
 a1728a <=( a1727a ) or ( a1722a );
 a1732a <=( a280a ) or ( a281a );
 a1733a <=( a282a ) or ( a1732a );
 a1737a <=( a277a ) or ( a278a );
 a1738a <=( a279a ) or ( a1737a );
 a1739a <=( a1738a ) or ( a1733a );
 a1740a <=( a1739a ) or ( a1728a );
 a1744a <=( a274a ) or ( a275a );
 a1745a <=( a276a ) or ( a1744a );
 a1749a <=( a271a ) or ( a272a );
 a1750a <=( a273a ) or ( a1749a );
 a1751a <=( a1750a ) or ( a1745a );
 a1755a <=( a268a ) or ( a269a );
 a1756a <=( a270a ) or ( a1755a );
 a1760a <=( a265a ) or ( a266a );
 a1761a <=( a267a ) or ( a1760a );
 a1762a <=( a1761a ) or ( a1756a );
 a1763a <=( a1762a ) or ( a1751a );
 a1764a <=( a1763a ) or ( a1740a );
 a1768a <=( a262a ) or ( a263a );
 a1769a <=( a264a ) or ( a1768a );
 a1773a <=( a259a ) or ( a260a );
 a1774a <=( a261a ) or ( a1773a );
 a1775a <=( a1774a ) or ( a1769a );
 a1779a <=( a256a ) or ( a257a );
 a1780a <=( a258a ) or ( a1779a );
 a1784a <=( a253a ) or ( a254a );
 a1785a <=( a255a ) or ( a1784a );
 a1786a <=( a1785a ) or ( a1780a );
 a1787a <=( a1786a ) or ( a1775a );
 a1791a <=( a250a ) or ( a251a );
 a1792a <=( a252a ) or ( a1791a );
 a1796a <=( a247a ) or ( a248a );
 a1797a <=( a249a ) or ( a1796a );
 a1798a <=( a1797a ) or ( a1792a );
 a1802a <=( a244a ) or ( a245a );
 a1803a <=( a246a ) or ( a1802a );
 a1807a <=( a241a ) or ( a242a );
 a1808a <=( a243a ) or ( a1807a );
 a1809a <=( a1808a ) or ( a1803a );
 a1810a <=( a1809a ) or ( a1798a );
 a1811a <=( a1810a ) or ( a1787a );
 a1812a <=( a1811a ) or ( a1764a );
 a1816a <=( a238a ) or ( a239a );
 a1817a <=( a240a ) or ( a1816a );
 a1821a <=( a235a ) or ( a236a );
 a1822a <=( a237a ) or ( a1821a );
 a1823a <=( a1822a ) or ( a1817a );
 a1827a <=( a232a ) or ( a233a );
 a1828a <=( a234a ) or ( a1827a );
 a1832a <=( a229a ) or ( a230a );
 a1833a <=( a231a ) or ( a1832a );
 a1834a <=( a1833a ) or ( a1828a );
 a1835a <=( a1834a ) or ( a1823a );
 a1839a <=( a226a ) or ( a227a );
 a1840a <=( a228a ) or ( a1839a );
 a1844a <=( a223a ) or ( a224a );
 a1845a <=( a225a ) or ( a1844a );
 a1846a <=( a1845a ) or ( a1840a );
 a1850a <=( a220a ) or ( a221a );
 a1851a <=( a222a ) or ( a1850a );
 a1855a <=( a217a ) or ( a218a );
 a1856a <=( a219a ) or ( a1855a );
 a1857a <=( a1856a ) or ( a1851a );
 a1858a <=( a1857a ) or ( a1846a );
 a1859a <=( a1858a ) or ( a1835a );
 a1863a <=( a214a ) or ( a215a );
 a1864a <=( a216a ) or ( a1863a );
 a1868a <=( a211a ) or ( a212a );
 a1869a <=( a213a ) or ( a1868a );
 a1870a <=( a1869a ) or ( a1864a );
 a1874a <=( a208a ) or ( a209a );
 a1875a <=( a210a ) or ( a1874a );
 a1879a <=( a205a ) or ( a206a );
 a1880a <=( a207a ) or ( a1879a );
 a1881a <=( a1880a ) or ( a1875a );
 a1882a <=( a1881a ) or ( a1870a );
 a1886a <=( a202a ) or ( a203a );
 a1887a <=( a204a ) or ( a1886a );
 a1891a <=( a199a ) or ( a200a );
 a1892a <=( a201a ) or ( a1891a );
 a1893a <=( a1892a ) or ( a1887a );
 a1897a <=( a196a ) or ( a197a );
 a1898a <=( a198a ) or ( a1897a );
 a1902a <=( a193a ) or ( a194a );
 a1903a <=( a195a ) or ( a1902a );
 a1904a <=( a1903a ) or ( a1898a );
 a1905a <=( a1904a ) or ( a1893a );
 a1906a <=( a1905a ) or ( a1882a );
 a1907a <=( a1906a ) or ( a1859a );
 a1908a <=( a1907a ) or ( a1812a );
 a1909a <=( a1908a ) or ( a1717a );
 a1913a <=( a190a ) or ( a191a );
 a1914a <=( a192a ) or ( a1913a );
 a1918a <=( a187a ) or ( a188a );
 a1919a <=( a189a ) or ( a1918a );
 a1920a <=( a1919a ) or ( a1914a );
 a1924a <=( a184a ) or ( a185a );
 a1925a <=( a186a ) or ( a1924a );
 a1929a <=( a181a ) or ( a182a );
 a1930a <=( a183a ) or ( a1929a );
 a1931a <=( a1930a ) or ( a1925a );
 a1932a <=( a1931a ) or ( a1920a );
 a1936a <=( a178a ) or ( a179a );
 a1937a <=( a180a ) or ( a1936a );
 a1941a <=( a175a ) or ( a176a );
 a1942a <=( a177a ) or ( a1941a );
 a1943a <=( a1942a ) or ( a1937a );
 a1947a <=( a172a ) or ( a173a );
 a1948a <=( a174a ) or ( a1947a );
 a1952a <=( a169a ) or ( a170a );
 a1953a <=( a171a ) or ( a1952a );
 a1954a <=( a1953a ) or ( a1948a );
 a1955a <=( a1954a ) or ( a1943a );
 a1956a <=( a1955a ) or ( a1932a );
 a1960a <=( a166a ) or ( a167a );
 a1961a <=( a168a ) or ( a1960a );
 a1965a <=( a163a ) or ( a164a );
 a1966a <=( a165a ) or ( a1965a );
 a1967a <=( a1966a ) or ( a1961a );
 a1971a <=( a160a ) or ( a161a );
 a1972a <=( a162a ) or ( a1971a );
 a1976a <=( a157a ) or ( a158a );
 a1977a <=( a159a ) or ( a1976a );
 a1978a <=( a1977a ) or ( a1972a );
 a1979a <=( a1978a ) or ( a1967a );
 a1983a <=( a154a ) or ( a155a );
 a1984a <=( a156a ) or ( a1983a );
 a1988a <=( a151a ) or ( a152a );
 a1989a <=( a153a ) or ( a1988a );
 a1990a <=( a1989a ) or ( a1984a );
 a1994a <=( a148a ) or ( a149a );
 a1995a <=( a150a ) or ( a1994a );
 a1999a <=( a145a ) or ( a146a );
 a2000a <=( a147a ) or ( a1999a );
 a2001a <=( a2000a ) or ( a1995a );
 a2002a <=( a2001a ) or ( a1990a );
 a2003a <=( a2002a ) or ( a1979a );
 a2004a <=( a2003a ) or ( a1956a );
 a2008a <=( a142a ) or ( a143a );
 a2009a <=( a144a ) or ( a2008a );
 a2013a <=( a139a ) or ( a140a );
 a2014a <=( a141a ) or ( a2013a );
 a2015a <=( a2014a ) or ( a2009a );
 a2019a <=( a136a ) or ( a137a );
 a2020a <=( a138a ) or ( a2019a );
 a2024a <=( a133a ) or ( a134a );
 a2025a <=( a135a ) or ( a2024a );
 a2026a <=( a2025a ) or ( a2020a );
 a2027a <=( a2026a ) or ( a2015a );
 a2031a <=( a130a ) or ( a131a );
 a2032a <=( a132a ) or ( a2031a );
 a2036a <=( a127a ) or ( a128a );
 a2037a <=( a129a ) or ( a2036a );
 a2038a <=( a2037a ) or ( a2032a );
 a2042a <=( a124a ) or ( a125a );
 a2043a <=( a126a ) or ( a2042a );
 a2047a <=( a121a ) or ( a122a );
 a2048a <=( a123a ) or ( a2047a );
 a2049a <=( a2048a ) or ( a2043a );
 a2050a <=( a2049a ) or ( a2038a );
 a2051a <=( a2050a ) or ( a2027a );
 a2055a <=( a118a ) or ( a119a );
 a2056a <=( a120a ) or ( a2055a );
 a2060a <=( a115a ) or ( a116a );
 a2061a <=( a117a ) or ( a2060a );
 a2062a <=( a2061a ) or ( a2056a );
 a2066a <=( a112a ) or ( a113a );
 a2067a <=( a114a ) or ( a2066a );
 a2071a <=( a109a ) or ( a110a );
 a2072a <=( a111a ) or ( a2071a );
 a2073a <=( a2072a ) or ( a2067a );
 a2074a <=( a2073a ) or ( a2062a );
 a2078a <=( a106a ) or ( a107a );
 a2079a <=( a108a ) or ( a2078a );
 a2083a <=( a103a ) or ( a104a );
 a2084a <=( a105a ) or ( a2083a );
 a2085a <=( a2084a ) or ( a2079a );
 a2089a <=( a100a ) or ( a101a );
 a2090a <=( a102a ) or ( a2089a );
 a2094a <=( a97a ) or ( a98a );
 a2095a <=( a99a ) or ( a2094a );
 a2096a <=( a2095a ) or ( a2090a );
 a2097a <=( a2096a ) or ( a2085a );
 a2098a <=( a2097a ) or ( a2074a );
 a2099a <=( a2098a ) or ( a2051a );
 a2100a <=( a2099a ) or ( a2004a );
 a2104a <=( a94a ) or ( a95a );
 a2105a <=( a96a ) or ( a2104a );
 a2109a <=( a91a ) or ( a92a );
 a2110a <=( a93a ) or ( a2109a );
 a2111a <=( a2110a ) or ( a2105a );
 a2115a <=( a88a ) or ( a89a );
 a2116a <=( a90a ) or ( a2115a );
 a2120a <=( a85a ) or ( a86a );
 a2121a <=( a87a ) or ( a2120a );
 a2122a <=( a2121a ) or ( a2116a );
 a2123a <=( a2122a ) or ( a2111a );
 a2127a <=( a82a ) or ( a83a );
 a2128a <=( a84a ) or ( a2127a );
 a2132a <=( a79a ) or ( a80a );
 a2133a <=( a81a ) or ( a2132a );
 a2134a <=( a2133a ) or ( a2128a );
 a2138a <=( a76a ) or ( a77a );
 a2139a <=( a78a ) or ( a2138a );
 a2143a <=( a73a ) or ( a74a );
 a2144a <=( a75a ) or ( a2143a );
 a2145a <=( a2144a ) or ( a2139a );
 a2146a <=( a2145a ) or ( a2134a );
 a2147a <=( a2146a ) or ( a2123a );
 a2151a <=( a70a ) or ( a71a );
 a2152a <=( a72a ) or ( a2151a );
 a2156a <=( a67a ) or ( a68a );
 a2157a <=( a69a ) or ( a2156a );
 a2158a <=( a2157a ) or ( a2152a );
 a2162a <=( a64a ) or ( a65a );
 a2163a <=( a66a ) or ( a2162a );
 a2167a <=( a61a ) or ( a62a );
 a2168a <=( a63a ) or ( a2167a );
 a2169a <=( a2168a ) or ( a2163a );
 a2170a <=( a2169a ) or ( a2158a );
 a2174a <=( a58a ) or ( a59a );
 a2175a <=( a60a ) or ( a2174a );
 a2179a <=( a55a ) or ( a56a );
 a2180a <=( a57a ) or ( a2179a );
 a2181a <=( a2180a ) or ( a2175a );
 a2185a <=( a52a ) or ( a53a );
 a2186a <=( a54a ) or ( a2185a );
 a2190a <=( a49a ) or ( a50a );
 a2191a <=( a51a ) or ( a2190a );
 a2192a <=( a2191a ) or ( a2186a );
 a2193a <=( a2192a ) or ( a2181a );
 a2194a <=( a2193a ) or ( a2170a );
 a2195a <=( a2194a ) or ( a2147a );
 a2199a <=( a46a ) or ( a47a );
 a2200a <=( a48a ) or ( a2199a );
 a2204a <=( a43a ) or ( a44a );
 a2205a <=( a45a ) or ( a2204a );
 a2206a <=( a2205a ) or ( a2200a );
 a2210a <=( a40a ) or ( a41a );
 a2211a <=( a42a ) or ( a2210a );
 a2215a <=( a37a ) or ( a38a );
 a2216a <=( a39a ) or ( a2215a );
 a2217a <=( a2216a ) or ( a2211a );
 a2218a <=( a2217a ) or ( a2206a );
 a2222a <=( a34a ) or ( a35a );
 a2223a <=( a36a ) or ( a2222a );
 a2227a <=( a31a ) or ( a32a );
 a2228a <=( a33a ) or ( a2227a );
 a2229a <=( a2228a ) or ( a2223a );
 a2233a <=( a28a ) or ( a29a );
 a2234a <=( a30a ) or ( a2233a );
 a2238a <=( a25a ) or ( a26a );
 a2239a <=( a27a ) or ( a2238a );
 a2240a <=( a2239a ) or ( a2234a );
 a2241a <=( a2240a ) or ( a2229a );
 a2242a <=( a2241a ) or ( a2218a );
 a2246a <=( a22a ) or ( a23a );
 a2247a <=( a24a ) or ( a2246a );
 a2251a <=( a19a ) or ( a20a );
 a2252a <=( a21a ) or ( a2251a );
 a2253a <=( a2252a ) or ( a2247a );
 a2257a <=( a16a ) or ( a17a );
 a2258a <=( a18a ) or ( a2257a );
 a2262a <=( a13a ) or ( a14a );
 a2263a <=( a15a ) or ( a2262a );
 a2264a <=( a2263a ) or ( a2258a );
 a2265a <=( a2264a ) or ( a2253a );
 a2269a <=( a10a ) or ( a11a );
 a2270a <=( a12a ) or ( a2269a );
 a2274a <=( a7a ) or ( a8a );
 a2275a <=( a9a ) or ( a2274a );
 a2276a <=( a2275a ) or ( a2270a );
 a2280a <=( a4a ) or ( a5a );
 a2281a <=( a6a ) or ( a2280a );
 a2285a <=( a1a ) or ( a2a );
 a2286a <=( a3a ) or ( a2285a );
 a2287a <=( a2286a ) or ( a2281a );
 a2288a <=( a2287a ) or ( a2276a );
 a2289a <=( a2288a ) or ( a2265a );
 a2290a <=( a2289a ) or ( a2242a );
 a2291a <=( a2290a ) or ( a2195a );
 a2292a <=( a2291a ) or ( a2100a );
 a2293a <=( a2292a ) or ( a1909a );
 a2296a <=( (not A167)  and  (not A169) );
 a2299a <=( A202  and  (not A166) );
 a2302a <=( (not A169)  and  (not A170) );
 a2305a <=( A202  and  (not A168) );
 a2308a <=( (not A167)  and  (not A169) );
 a2312a <=( A201  and  A199 );
 a2313a <=( (not A166)  and  a2312a );
 a2316a <=( (not A167)  and  (not A169) );
 a2320a <=( A201  and  A200 );
 a2321a <=( (not A166)  and  a2320a );
 a2324a <=( (not A168)  and  (not A169) );
 a2328a <=( A202  and  A166 );
 a2329a <=( A167  and  a2328a );
 a2332a <=( (not A169)  and  (not A170) );
 a2336a <=( A201  and  A199 );
 a2337a <=( (not A168)  and  a2336a );
 a2340a <=( (not A169)  and  (not A170) );
 a2344a <=( A201  and  A200 );
 a2345a <=( (not A168)  and  a2344a );
 a2349a <=( (not A202)  and  (not A201) );
 a2350a <=( A169  and  a2349a );
 a2354a <=( A301  and  A235 );
 a2355a <=( (not A203)  and  a2354a );
 a2359a <=( (not A202)  and  (not A201) );
 a2360a <=( A169  and  a2359a );
 a2364a <=( A268  and  A235 );
 a2365a <=( (not A203)  and  a2364a );
 a2369a <=( (not A200)  and  (not A199) );
 a2370a <=( A169  and  a2369a );
 a2374a <=( A301  and  A235 );
 a2375a <=( (not A202)  and  a2374a );
 a2379a <=( (not A200)  and  (not A199) );
 a2380a <=( A169  and  a2379a );
 a2384a <=( A268  and  A235 );
 a2385a <=( (not A202)  and  a2384a );
 a2389a <=( (not A166)  and  (not A167) );
 a2390a <=( (not A169)  and  a2389a );
 a2394a <=( A203  and  A200 );
 a2395a <=( (not A199)  and  a2394a );
 a2399a <=( (not A166)  and  (not A167) );
 a2400a <=( (not A169)  and  a2399a );
 a2404a <=( A203  and  (not A200) );
 a2405a <=( A199  and  a2404a );
 a2409a <=( A167  and  (not A168) );
 a2410a <=( (not A169)  and  a2409a );
 a2414a <=( A201  and  A199 );
 a2415a <=( A166  and  a2414a );
 a2419a <=( A167  and  (not A168) );
 a2420a <=( (not A169)  and  a2419a );
 a2424a <=( A201  and  A200 );
 a2425a <=( A166  and  a2424a );
 a2429a <=( (not A168)  and  (not A169) );
 a2430a <=( (not A170)  and  a2429a );
 a2434a <=( A203  and  A200 );
 a2435a <=( (not A199)  and  a2434a );
 a2439a <=( (not A168)  and  (not A169) );
 a2440a <=( (not A170)  and  a2439a );
 a2444a <=( A203  and  (not A200) );
 a2445a <=( A199  and  a2444a );
 a2449a <=( (not A201)  and  A166 );
 a2450a <=( A168  and  a2449a );
 a2453a <=( (not A203)  and  (not A202) );
 a2456a <=( A301  and  A235 );
 a2457a <=( a2456a  and  a2453a );
 a2461a <=( (not A201)  and  A166 );
 a2462a <=( A168  and  a2461a );
 a2465a <=( (not A203)  and  (not A202) );
 a2468a <=( A268  and  A235 );
 a2469a <=( a2468a  and  a2465a );
 a2473a <=( (not A199)  and  A166 );
 a2474a <=( A168  and  a2473a );
 a2477a <=( (not A202)  and  (not A200) );
 a2480a <=( A301  and  A235 );
 a2481a <=( a2480a  and  a2477a );
 a2485a <=( (not A199)  and  A166 );
 a2486a <=( A168  and  a2485a );
 a2489a <=( (not A202)  and  (not A200) );
 a2492a <=( A268  and  A235 );
 a2493a <=( a2492a  and  a2489a );
 a2497a <=( (not A201)  and  A167 );
 a2498a <=( A168  and  a2497a );
 a2501a <=( (not A203)  and  (not A202) );
 a2504a <=( A301  and  A235 );
 a2505a <=( a2504a  and  a2501a );
 a2509a <=( (not A201)  and  A167 );
 a2510a <=( A168  and  a2509a );
 a2513a <=( (not A203)  and  (not A202) );
 a2516a <=( A268  and  A235 );
 a2517a <=( a2516a  and  a2513a );
 a2521a <=( (not A199)  and  A167 );
 a2522a <=( A168  and  a2521a );
 a2525a <=( (not A202)  and  (not A200) );
 a2528a <=( A301  and  A235 );
 a2529a <=( a2528a  and  a2525a );
 a2533a <=( (not A199)  and  A167 );
 a2534a <=( A168  and  a2533a );
 a2537a <=( (not A202)  and  (not A200) );
 a2540a <=( A268  and  A235 );
 a2541a <=( a2540a  and  a2537a );
 a2545a <=( (not A202)  and  (not A201) );
 a2546a <=( A169  and  a2545a );
 a2549a <=( A235  and  (not A203) );
 a2552a <=( A300  and  A299 );
 a2553a <=( a2552a  and  a2549a );
 a2557a <=( (not A202)  and  (not A201) );
 a2558a <=( A169  and  a2557a );
 a2561a <=( A235  and  (not A203) );
 a2564a <=( A300  and  A298 );
 a2565a <=( a2564a  and  a2561a );
 a2569a <=( (not A202)  and  (not A201) );
 a2570a <=( A169  and  a2569a );
 a2573a <=( A235  and  (not A203) );
 a2576a <=( A267  and  A265 );
 a2577a <=( a2576a  and  a2573a );
 a2581a <=( (not A202)  and  (not A201) );
 a2582a <=( A169  and  a2581a );
 a2585a <=( A235  and  (not A203) );
 a2588a <=( A267  and  A266 );
 a2589a <=( a2588a  and  a2585a );
 a2593a <=( (not A202)  and  (not A201) );
 a2594a <=( A169  and  a2593a );
 a2597a <=( A232  and  (not A203) );
 a2600a <=( A301  and  A234 );
 a2601a <=( a2600a  and  a2597a );
 a2605a <=( (not A202)  and  (not A201) );
 a2606a <=( A169  and  a2605a );
 a2609a <=( A232  and  (not A203) );
 a2612a <=( A268  and  A234 );
 a2613a <=( a2612a  and  a2609a );
 a2617a <=( (not A202)  and  (not A201) );
 a2618a <=( A169  and  a2617a );
 a2621a <=( A233  and  (not A203) );
 a2624a <=( A301  and  A234 );
 a2625a <=( a2624a  and  a2621a );
 a2629a <=( (not A202)  and  (not A201) );
 a2630a <=( A169  and  a2629a );
 a2633a <=( A233  and  (not A203) );
 a2636a <=( A268  and  A234 );
 a2637a <=( a2636a  and  a2633a );
 a2641a <=( A200  and  A199 );
 a2642a <=( A169  and  a2641a );
 a2645a <=( (not A202)  and  (not A201) );
 a2648a <=( A301  and  A235 );
 a2649a <=( a2648a  and  a2645a );
 a2653a <=( A200  and  A199 );
 a2654a <=( A169  and  a2653a );
 a2657a <=( (not A202)  and  (not A201) );
 a2660a <=( A268  and  A235 );
 a2661a <=( a2660a  and  a2657a );
 a2665a <=( (not A200)  and  (not A199) );
 a2666a <=( A169  and  a2665a );
 a2669a <=( A235  and  (not A202) );
 a2672a <=( A300  and  A299 );
 a2673a <=( a2672a  and  a2669a );
 a2677a <=( (not A200)  and  (not A199) );
 a2678a <=( A169  and  a2677a );
 a2681a <=( A235  and  (not A202) );
 a2684a <=( A300  and  A298 );
 a2685a <=( a2684a  and  a2681a );
 a2689a <=( (not A200)  and  (not A199) );
 a2690a <=( A169  and  a2689a );
 a2693a <=( A235  and  (not A202) );
 a2696a <=( A267  and  A265 );
 a2697a <=( a2696a  and  a2693a );
 a2701a <=( (not A200)  and  (not A199) );
 a2702a <=( A169  and  a2701a );
 a2705a <=( A235  and  (not A202) );
 a2708a <=( A267  and  A266 );
 a2709a <=( a2708a  and  a2705a );
 a2713a <=( (not A200)  and  (not A199) );
 a2714a <=( A169  and  a2713a );
 a2717a <=( A232  and  (not A202) );
 a2720a <=( A301  and  A234 );
 a2721a <=( a2720a  and  a2717a );
 a2725a <=( (not A200)  and  (not A199) );
 a2726a <=( A169  and  a2725a );
 a2729a <=( A232  and  (not A202) );
 a2732a <=( A268  and  A234 );
 a2733a <=( a2732a  and  a2729a );
 a2737a <=( (not A200)  and  (not A199) );
 a2738a <=( A169  and  a2737a );
 a2741a <=( A233  and  (not A202) );
 a2744a <=( A301  and  A234 );
 a2745a <=( a2744a  and  a2741a );
 a2749a <=( (not A200)  and  (not A199) );
 a2750a <=( A169  and  a2749a );
 a2753a <=( A233  and  (not A202) );
 a2756a <=( A268  and  A234 );
 a2757a <=( a2756a  and  a2753a );
 a2761a <=( A167  and  (not A168) );
 a2762a <=( (not A169)  and  a2761a );
 a2765a <=( (not A199)  and  A166 );
 a2768a <=( A203  and  A200 );
 a2769a <=( a2768a  and  a2765a );
 a2773a <=( A167  and  (not A168) );
 a2774a <=( (not A169)  and  a2773a );
 a2777a <=( A199  and  A166 );
 a2780a <=( A203  and  (not A200) );
 a2781a <=( a2780a  and  a2777a );
 a2784a <=( A166  and  A168 );
 a2787a <=( (not A202)  and  (not A201) );
 a2788a <=( a2787a  and  a2784a );
 a2791a <=( A235  and  (not A203) );
 a2794a <=( A300  and  A299 );
 a2795a <=( a2794a  and  a2791a );
 a2798a <=( A166  and  A168 );
 a2801a <=( (not A202)  and  (not A201) );
 a2802a <=( a2801a  and  a2798a );
 a2805a <=( A235  and  (not A203) );
 a2808a <=( A300  and  A298 );
 a2809a <=( a2808a  and  a2805a );
 a2812a <=( A166  and  A168 );
 a2815a <=( (not A202)  and  (not A201) );
 a2816a <=( a2815a  and  a2812a );
 a2819a <=( A235  and  (not A203) );
 a2822a <=( A267  and  A265 );
 a2823a <=( a2822a  and  a2819a );
 a2826a <=( A166  and  A168 );
 a2829a <=( (not A202)  and  (not A201) );
 a2830a <=( a2829a  and  a2826a );
 a2833a <=( A235  and  (not A203) );
 a2836a <=( A267  and  A266 );
 a2837a <=( a2836a  and  a2833a );
 a2840a <=( A166  and  A168 );
 a2843a <=( (not A202)  and  (not A201) );
 a2844a <=( a2843a  and  a2840a );
 a2847a <=( A232  and  (not A203) );
 a2850a <=( A301  and  A234 );
 a2851a <=( a2850a  and  a2847a );
 a2854a <=( A166  and  A168 );
 a2857a <=( (not A202)  and  (not A201) );
 a2858a <=( a2857a  and  a2854a );
 a2861a <=( A232  and  (not A203) );
 a2864a <=( A268  and  A234 );
 a2865a <=( a2864a  and  a2861a );
 a2868a <=( A166  and  A168 );
 a2871a <=( (not A202)  and  (not A201) );
 a2872a <=( a2871a  and  a2868a );
 a2875a <=( A233  and  (not A203) );
 a2878a <=( A301  and  A234 );
 a2879a <=( a2878a  and  a2875a );
 a2882a <=( A166  and  A168 );
 a2885a <=( (not A202)  and  (not A201) );
 a2886a <=( a2885a  and  a2882a );
 a2889a <=( A233  and  (not A203) );
 a2892a <=( A268  and  A234 );
 a2893a <=( a2892a  and  a2889a );
 a2896a <=( A166  and  A168 );
 a2899a <=( A200  and  A199 );
 a2900a <=( a2899a  and  a2896a );
 a2903a <=( (not A202)  and  (not A201) );
 a2906a <=( A301  and  A235 );
 a2907a <=( a2906a  and  a2903a );
 a2910a <=( A166  and  A168 );
 a2913a <=( A200  and  A199 );
 a2914a <=( a2913a  and  a2910a );
 a2917a <=( (not A202)  and  (not A201) );
 a2920a <=( A268  and  A235 );
 a2921a <=( a2920a  and  a2917a );
 a2924a <=( A166  and  A168 );
 a2927a <=( (not A200)  and  (not A199) );
 a2928a <=( a2927a  and  a2924a );
 a2931a <=( A235  and  (not A202) );
 a2934a <=( A300  and  A299 );
 a2935a <=( a2934a  and  a2931a );
 a2938a <=( A166  and  A168 );
 a2941a <=( (not A200)  and  (not A199) );
 a2942a <=( a2941a  and  a2938a );
 a2945a <=( A235  and  (not A202) );
 a2948a <=( A300  and  A298 );
 a2949a <=( a2948a  and  a2945a );
 a2952a <=( A166  and  A168 );
 a2955a <=( (not A200)  and  (not A199) );
 a2956a <=( a2955a  and  a2952a );
 a2959a <=( A235  and  (not A202) );
 a2962a <=( A267  and  A265 );
 a2963a <=( a2962a  and  a2959a );
 a2966a <=( A166  and  A168 );
 a2969a <=( (not A200)  and  (not A199) );
 a2970a <=( a2969a  and  a2966a );
 a2973a <=( A235  and  (not A202) );
 a2976a <=( A267  and  A266 );
 a2977a <=( a2976a  and  a2973a );
 a2980a <=( A166  and  A168 );
 a2983a <=( (not A200)  and  (not A199) );
 a2984a <=( a2983a  and  a2980a );
 a2987a <=( A232  and  (not A202) );
 a2990a <=( A301  and  A234 );
 a2991a <=( a2990a  and  a2987a );
 a2994a <=( A166  and  A168 );
 a2997a <=( (not A200)  and  (not A199) );
 a2998a <=( a2997a  and  a2994a );
 a3001a <=( A232  and  (not A202) );
 a3004a <=( A268  and  A234 );
 a3005a <=( a3004a  and  a3001a );
 a3008a <=( A166  and  A168 );
 a3011a <=( (not A200)  and  (not A199) );
 a3012a <=( a3011a  and  a3008a );
 a3015a <=( A233  and  (not A202) );
 a3018a <=( A301  and  A234 );
 a3019a <=( a3018a  and  a3015a );
 a3022a <=( A166  and  A168 );
 a3025a <=( (not A200)  and  (not A199) );
 a3026a <=( a3025a  and  a3022a );
 a3029a <=( A233  and  (not A202) );
 a3032a <=( A268  and  A234 );
 a3033a <=( a3032a  and  a3029a );
 a3036a <=( A167  and  A168 );
 a3039a <=( (not A202)  and  (not A201) );
 a3040a <=( a3039a  and  a3036a );
 a3043a <=( A235  and  (not A203) );
 a3046a <=( A300  and  A299 );
 a3047a <=( a3046a  and  a3043a );
 a3050a <=( A167  and  A168 );
 a3053a <=( (not A202)  and  (not A201) );
 a3054a <=( a3053a  and  a3050a );
 a3057a <=( A235  and  (not A203) );
 a3060a <=( A300  and  A298 );
 a3061a <=( a3060a  and  a3057a );
 a3064a <=( A167  and  A168 );
 a3067a <=( (not A202)  and  (not A201) );
 a3068a <=( a3067a  and  a3064a );
 a3071a <=( A235  and  (not A203) );
 a3074a <=( A267  and  A265 );
 a3075a <=( a3074a  and  a3071a );
 a3078a <=( A167  and  A168 );
 a3081a <=( (not A202)  and  (not A201) );
 a3082a <=( a3081a  and  a3078a );
 a3085a <=( A235  and  (not A203) );
 a3088a <=( A267  and  A266 );
 a3089a <=( a3088a  and  a3085a );
 a3092a <=( A167  and  A168 );
 a3095a <=( (not A202)  and  (not A201) );
 a3096a <=( a3095a  and  a3092a );
 a3099a <=( A232  and  (not A203) );
 a3102a <=( A301  and  A234 );
 a3103a <=( a3102a  and  a3099a );
 a3106a <=( A167  and  A168 );
 a3109a <=( (not A202)  and  (not A201) );
 a3110a <=( a3109a  and  a3106a );
 a3113a <=( A232  and  (not A203) );
 a3116a <=( A268  and  A234 );
 a3117a <=( a3116a  and  a3113a );
 a3120a <=( A167  and  A168 );
 a3123a <=( (not A202)  and  (not A201) );
 a3124a <=( a3123a  and  a3120a );
 a3127a <=( A233  and  (not A203) );
 a3130a <=( A301  and  A234 );
 a3131a <=( a3130a  and  a3127a );
 a3134a <=( A167  and  A168 );
 a3137a <=( (not A202)  and  (not A201) );
 a3138a <=( a3137a  and  a3134a );
 a3141a <=( A233  and  (not A203) );
 a3144a <=( A268  and  A234 );
 a3145a <=( a3144a  and  a3141a );
 a3148a <=( A167  and  A168 );
 a3151a <=( A200  and  A199 );
 a3152a <=( a3151a  and  a3148a );
 a3155a <=( (not A202)  and  (not A201) );
 a3158a <=( A301  and  A235 );
 a3159a <=( a3158a  and  a3155a );
 a3162a <=( A167  and  A168 );
 a3165a <=( A200  and  A199 );
 a3166a <=( a3165a  and  a3162a );
 a3169a <=( (not A202)  and  (not A201) );
 a3172a <=( A268  and  A235 );
 a3173a <=( a3172a  and  a3169a );
 a3176a <=( A167  and  A168 );
 a3179a <=( (not A200)  and  (not A199) );
 a3180a <=( a3179a  and  a3176a );
 a3183a <=( A235  and  (not A202) );
 a3186a <=( A300  and  A299 );
 a3187a <=( a3186a  and  a3183a );
 a3190a <=( A167  and  A168 );
 a3193a <=( (not A200)  and  (not A199) );
 a3194a <=( a3193a  and  a3190a );
 a3197a <=( A235  and  (not A202) );
 a3200a <=( A300  and  A298 );
 a3201a <=( a3200a  and  a3197a );
 a3204a <=( A167  and  A168 );
 a3207a <=( (not A200)  and  (not A199) );
 a3208a <=( a3207a  and  a3204a );
 a3211a <=( A235  and  (not A202) );
 a3214a <=( A267  and  A265 );
 a3215a <=( a3214a  and  a3211a );
 a3218a <=( A167  and  A168 );
 a3221a <=( (not A200)  and  (not A199) );
 a3222a <=( a3221a  and  a3218a );
 a3225a <=( A235  and  (not A202) );
 a3228a <=( A267  and  A266 );
 a3229a <=( a3228a  and  a3225a );
 a3232a <=( A167  and  A168 );
 a3235a <=( (not A200)  and  (not A199) );
 a3236a <=( a3235a  and  a3232a );
 a3239a <=( A232  and  (not A202) );
 a3242a <=( A301  and  A234 );
 a3243a <=( a3242a  and  a3239a );
 a3246a <=( A167  and  A168 );
 a3249a <=( (not A200)  and  (not A199) );
 a3250a <=( a3249a  and  a3246a );
 a3253a <=( A232  and  (not A202) );
 a3256a <=( A268  and  A234 );
 a3257a <=( a3256a  and  a3253a );
 a3260a <=( A167  and  A168 );
 a3263a <=( (not A200)  and  (not A199) );
 a3264a <=( a3263a  and  a3260a );
 a3267a <=( A233  and  (not A202) );
 a3270a <=( A301  and  A234 );
 a3271a <=( a3270a  and  a3267a );
 a3274a <=( A167  and  A168 );
 a3277a <=( (not A200)  and  (not A199) );
 a3278a <=( a3277a  and  a3274a );
 a3281a <=( A233  and  (not A202) );
 a3284a <=( A268  and  A234 );
 a3285a <=( a3284a  and  a3281a );
 a3288a <=( A167  and  A170 );
 a3291a <=( (not A201)  and  (not A166) );
 a3292a <=( a3291a  and  a3288a );
 a3295a <=( (not A203)  and  (not A202) );
 a3298a <=( A301  and  A235 );
 a3299a <=( a3298a  and  a3295a );
 a3302a <=( A167  and  A170 );
 a3305a <=( (not A201)  and  (not A166) );
 a3306a <=( a3305a  and  a3302a );
 a3309a <=( (not A203)  and  (not A202) );
 a3312a <=( A268  and  A235 );
 a3313a <=( a3312a  and  a3309a );
 a3316a <=( A167  and  A170 );
 a3319a <=( (not A199)  and  (not A166) );
 a3320a <=( a3319a  and  a3316a );
 a3323a <=( (not A202)  and  (not A200) );
 a3326a <=( A301  and  A235 );
 a3327a <=( a3326a  and  a3323a );
 a3330a <=( A167  and  A170 );
 a3333a <=( (not A199)  and  (not A166) );
 a3334a <=( a3333a  and  a3330a );
 a3337a <=( (not A202)  and  (not A200) );
 a3340a <=( A268  and  A235 );
 a3341a <=( a3340a  and  a3337a );
 a3344a <=( (not A167)  and  A170 );
 a3347a <=( (not A201)  and  A166 );
 a3348a <=( a3347a  and  a3344a );
 a3351a <=( (not A203)  and  (not A202) );
 a3354a <=( A301  and  A235 );
 a3355a <=( a3354a  and  a3351a );
 a3358a <=( (not A167)  and  A170 );
 a3361a <=( (not A201)  and  A166 );
 a3362a <=( a3361a  and  a3358a );
 a3365a <=( (not A203)  and  (not A202) );
 a3368a <=( A268  and  A235 );
 a3369a <=( a3368a  and  a3365a );
 a3372a <=( (not A167)  and  A170 );
 a3375a <=( (not A199)  and  A166 );
 a3376a <=( a3375a  and  a3372a );
 a3379a <=( (not A202)  and  (not A200) );
 a3382a <=( A301  and  A235 );
 a3383a <=( a3382a  and  a3379a );
 a3386a <=( (not A167)  and  A170 );
 a3389a <=( (not A199)  and  A166 );
 a3390a <=( a3389a  and  a3386a );
 a3393a <=( (not A202)  and  (not A200) );
 a3396a <=( A268  and  A235 );
 a3397a <=( a3396a  and  a3393a );
 a3400a <=( (not A201)  and  A169 );
 a3403a <=( (not A203)  and  (not A202) );
 a3404a <=( a3403a  and  a3400a );
 a3407a <=( A298  and  A235 );
 a3410a <=( A302  and  (not A299) );
 a3411a <=( a3410a  and  a3407a );
 a3414a <=( (not A201)  and  A169 );
 a3417a <=( (not A203)  and  (not A202) );
 a3418a <=( a3417a  and  a3414a );
 a3421a <=( (not A298)  and  A235 );
 a3424a <=( A302  and  A299 );
 a3425a <=( a3424a  and  a3421a );
 a3428a <=( (not A201)  and  A169 );
 a3431a <=( (not A203)  and  (not A202) );
 a3432a <=( a3431a  and  a3428a );
 a3435a <=( (not A265)  and  A235 );
 a3438a <=( A269  and  A266 );
 a3439a <=( a3438a  and  a3435a );
 a3442a <=( (not A201)  and  A169 );
 a3445a <=( (not A203)  and  (not A202) );
 a3446a <=( a3445a  and  a3442a );
 a3449a <=( A265  and  A235 );
 a3452a <=( A269  and  (not A266) );
 a3453a <=( a3452a  and  a3449a );
 a3456a <=( (not A201)  and  A169 );
 a3459a <=( (not A203)  and  (not A202) );
 a3460a <=( a3459a  and  a3456a );
 a3463a <=( A234  and  A232 );
 a3466a <=( A300  and  A299 );
 a3467a <=( a3466a  and  a3463a );
 a3470a <=( (not A201)  and  A169 );
 a3473a <=( (not A203)  and  (not A202) );
 a3474a <=( a3473a  and  a3470a );
 a3477a <=( A234  and  A232 );
 a3480a <=( A300  and  A298 );
 a3481a <=( a3480a  and  a3477a );
 a3484a <=( (not A201)  and  A169 );
 a3487a <=( (not A203)  and  (not A202) );
 a3488a <=( a3487a  and  a3484a );
 a3491a <=( A234  and  A232 );
 a3494a <=( A267  and  A265 );
 a3495a <=( a3494a  and  a3491a );
 a3498a <=( (not A201)  and  A169 );
 a3501a <=( (not A203)  and  (not A202) );
 a3502a <=( a3501a  and  a3498a );
 a3505a <=( A234  and  A232 );
 a3508a <=( A267  and  A266 );
 a3509a <=( a3508a  and  a3505a );
 a3512a <=( (not A201)  and  A169 );
 a3515a <=( (not A203)  and  (not A202) );
 a3516a <=( a3515a  and  a3512a );
 a3519a <=( A234  and  A233 );
 a3522a <=( A300  and  A299 );
 a3523a <=( a3522a  and  a3519a );
 a3526a <=( (not A201)  and  A169 );
 a3529a <=( (not A203)  and  (not A202) );
 a3530a <=( a3529a  and  a3526a );
 a3533a <=( A234  and  A233 );
 a3536a <=( A300  and  A298 );
 a3537a <=( a3536a  and  a3533a );
 a3540a <=( (not A201)  and  A169 );
 a3543a <=( (not A203)  and  (not A202) );
 a3544a <=( a3543a  and  a3540a );
 a3547a <=( A234  and  A233 );
 a3550a <=( A267  and  A265 );
 a3551a <=( a3550a  and  a3547a );
 a3554a <=( (not A201)  and  A169 );
 a3557a <=( (not A203)  and  (not A202) );
 a3558a <=( a3557a  and  a3554a );
 a3561a <=( A234  and  A233 );
 a3564a <=( A267  and  A266 );
 a3565a <=( a3564a  and  a3561a );
 a3568a <=( (not A201)  and  A169 );
 a3571a <=( (not A203)  and  (not A202) );
 a3572a <=( a3571a  and  a3568a );
 a3575a <=( A233  and  (not A232) );
 a3578a <=( A301  and  A236 );
 a3579a <=( a3578a  and  a3575a );
 a3582a <=( (not A201)  and  A169 );
 a3585a <=( (not A203)  and  (not A202) );
 a3586a <=( a3585a  and  a3582a );
 a3589a <=( A233  and  (not A232) );
 a3592a <=( A268  and  A236 );
 a3593a <=( a3592a  and  a3589a );
 a3596a <=( (not A201)  and  A169 );
 a3599a <=( (not A203)  and  (not A202) );
 a3600a <=( a3599a  and  a3596a );
 a3603a <=( (not A233)  and  A232 );
 a3606a <=( A301  and  A236 );
 a3607a <=( a3606a  and  a3603a );
 a3610a <=( (not A201)  and  A169 );
 a3613a <=( (not A203)  and  (not A202) );
 a3614a <=( a3613a  and  a3610a );
 a3617a <=( (not A233)  and  A232 );
 a3620a <=( A268  and  A236 );
 a3621a <=( a3620a  and  a3617a );
 a3624a <=( A199  and  A169 );
 a3627a <=( (not A201)  and  A200 );
 a3628a <=( a3627a  and  a3624a );
 a3631a <=( A235  and  (not A202) );
 a3634a <=( A300  and  A299 );
 a3635a <=( a3634a  and  a3631a );
 a3638a <=( A199  and  A169 );
 a3641a <=( (not A201)  and  A200 );
 a3642a <=( a3641a  and  a3638a );
 a3645a <=( A235  and  (not A202) );
 a3648a <=( A300  and  A298 );
 a3649a <=( a3648a  and  a3645a );
 a3652a <=( A199  and  A169 );
 a3655a <=( (not A201)  and  A200 );
 a3656a <=( a3655a  and  a3652a );
 a3659a <=( A235  and  (not A202) );
 a3662a <=( A267  and  A265 );
 a3663a <=( a3662a  and  a3659a );
 a3666a <=( A199  and  A169 );
 a3669a <=( (not A201)  and  A200 );
 a3670a <=( a3669a  and  a3666a );
 a3673a <=( A235  and  (not A202) );
 a3676a <=( A267  and  A266 );
 a3677a <=( a3676a  and  a3673a );
 a3680a <=( A199  and  A169 );
 a3683a <=( (not A201)  and  A200 );
 a3684a <=( a3683a  and  a3680a );
 a3687a <=( A232  and  (not A202) );
 a3690a <=( A301  and  A234 );
 a3691a <=( a3690a  and  a3687a );
 a3694a <=( A199  and  A169 );
 a3697a <=( (not A201)  and  A200 );
 a3698a <=( a3697a  and  a3694a );
 a3701a <=( A232  and  (not A202) );
 a3704a <=( A268  and  A234 );
 a3705a <=( a3704a  and  a3701a );
 a3708a <=( A199  and  A169 );
 a3711a <=( (not A201)  and  A200 );
 a3712a <=( a3711a  and  a3708a );
 a3715a <=( A233  and  (not A202) );
 a3718a <=( A301  and  A234 );
 a3719a <=( a3718a  and  a3715a );
 a3722a <=( A199  and  A169 );
 a3725a <=( (not A201)  and  A200 );
 a3726a <=( a3725a  and  a3722a );
 a3729a <=( A233  and  (not A202) );
 a3732a <=( A268  and  A234 );
 a3733a <=( a3732a  and  a3729a );
 a3736a <=( (not A199)  and  A169 );
 a3739a <=( (not A202)  and  (not A200) );
 a3740a <=( a3739a  and  a3736a );
 a3743a <=( A298  and  A235 );
 a3746a <=( A302  and  (not A299) );
 a3747a <=( a3746a  and  a3743a );
 a3750a <=( (not A199)  and  A169 );
 a3753a <=( (not A202)  and  (not A200) );
 a3754a <=( a3753a  and  a3750a );
 a3757a <=( (not A298)  and  A235 );
 a3760a <=( A302  and  A299 );
 a3761a <=( a3760a  and  a3757a );
 a3764a <=( (not A199)  and  A169 );
 a3767a <=( (not A202)  and  (not A200) );
 a3768a <=( a3767a  and  a3764a );
 a3771a <=( (not A265)  and  A235 );
 a3774a <=( A269  and  A266 );
 a3775a <=( a3774a  and  a3771a );
 a3778a <=( (not A199)  and  A169 );
 a3781a <=( (not A202)  and  (not A200) );
 a3782a <=( a3781a  and  a3778a );
 a3785a <=( A265  and  A235 );
 a3788a <=( A269  and  (not A266) );
 a3789a <=( a3788a  and  a3785a );
 a3792a <=( (not A199)  and  A169 );
 a3795a <=( (not A202)  and  (not A200) );
 a3796a <=( a3795a  and  a3792a );
 a3799a <=( A234  and  A232 );
 a3802a <=( A300  and  A299 );
 a3803a <=( a3802a  and  a3799a );
 a3806a <=( (not A199)  and  A169 );
 a3809a <=( (not A202)  and  (not A200) );
 a3810a <=( a3809a  and  a3806a );
 a3813a <=( A234  and  A232 );
 a3816a <=( A300  and  A298 );
 a3817a <=( a3816a  and  a3813a );
 a3820a <=( (not A199)  and  A169 );
 a3823a <=( (not A202)  and  (not A200) );
 a3824a <=( a3823a  and  a3820a );
 a3827a <=( A234  and  A232 );
 a3830a <=( A267  and  A265 );
 a3831a <=( a3830a  and  a3827a );
 a3834a <=( (not A199)  and  A169 );
 a3837a <=( (not A202)  and  (not A200) );
 a3838a <=( a3837a  and  a3834a );
 a3841a <=( A234  and  A232 );
 a3844a <=( A267  and  A266 );
 a3845a <=( a3844a  and  a3841a );
 a3848a <=( (not A199)  and  A169 );
 a3851a <=( (not A202)  and  (not A200) );
 a3852a <=( a3851a  and  a3848a );
 a3855a <=( A234  and  A233 );
 a3858a <=( A300  and  A299 );
 a3859a <=( a3858a  and  a3855a );
 a3862a <=( (not A199)  and  A169 );
 a3865a <=( (not A202)  and  (not A200) );
 a3866a <=( a3865a  and  a3862a );
 a3869a <=( A234  and  A233 );
 a3872a <=( A300  and  A298 );
 a3873a <=( a3872a  and  a3869a );
 a3876a <=( (not A199)  and  A169 );
 a3879a <=( (not A202)  and  (not A200) );
 a3880a <=( a3879a  and  a3876a );
 a3883a <=( A234  and  A233 );
 a3886a <=( A267  and  A265 );
 a3887a <=( a3886a  and  a3883a );
 a3890a <=( (not A199)  and  A169 );
 a3893a <=( (not A202)  and  (not A200) );
 a3894a <=( a3893a  and  a3890a );
 a3897a <=( A234  and  A233 );
 a3900a <=( A267  and  A266 );
 a3901a <=( a3900a  and  a3897a );
 a3904a <=( (not A199)  and  A169 );
 a3907a <=( (not A202)  and  (not A200) );
 a3908a <=( a3907a  and  a3904a );
 a3911a <=( A233  and  (not A232) );
 a3914a <=( A301  and  A236 );
 a3915a <=( a3914a  and  a3911a );
 a3918a <=( (not A199)  and  A169 );
 a3921a <=( (not A202)  and  (not A200) );
 a3922a <=( a3921a  and  a3918a );
 a3925a <=( A233  and  (not A232) );
 a3928a <=( A268  and  A236 );
 a3929a <=( a3928a  and  a3925a );
 a3932a <=( (not A199)  and  A169 );
 a3935a <=( (not A202)  and  (not A200) );
 a3936a <=( a3935a  and  a3932a );
 a3939a <=( (not A233)  and  A232 );
 a3942a <=( A301  and  A236 );
 a3943a <=( a3942a  and  a3939a );
 a3946a <=( (not A199)  and  A169 );
 a3949a <=( (not A202)  and  (not A200) );
 a3950a <=( a3949a  and  a3946a );
 a3953a <=( (not A233)  and  A232 );
 a3956a <=( A268  and  A236 );
 a3957a <=( a3956a  and  a3953a );
 a3960a <=( A166  and  A168 );
 a3963a <=( (not A202)  and  (not A201) );
 a3964a <=( a3963a  and  a3960a );
 a3967a <=( A235  and  (not A203) );
 a3971a <=( A302  and  (not A299) );
 a3972a <=( A298  and  a3971a );
 a3973a <=( a3972a  and  a3967a );
 a3976a <=( A166  and  A168 );
 a3979a <=( (not A202)  and  (not A201) );
 a3980a <=( a3979a  and  a3976a );
 a3983a <=( A235  and  (not A203) );
 a3987a <=( A302  and  A299 );
 a3988a <=( (not A298)  and  a3987a );
 a3989a <=( a3988a  and  a3983a );
 a3992a <=( A166  and  A168 );
 a3995a <=( (not A202)  and  (not A201) );
 a3996a <=( a3995a  and  a3992a );
 a3999a <=( A235  and  (not A203) );
 a4003a <=( A269  and  A266 );
 a4004a <=( (not A265)  and  a4003a );
 a4005a <=( a4004a  and  a3999a );
 a4008a <=( A166  and  A168 );
 a4011a <=( (not A202)  and  (not A201) );
 a4012a <=( a4011a  and  a4008a );
 a4015a <=( A235  and  (not A203) );
 a4019a <=( A269  and  (not A266) );
 a4020a <=( A265  and  a4019a );
 a4021a <=( a4020a  and  a4015a );
 a4024a <=( A166  and  A168 );
 a4027a <=( (not A202)  and  (not A201) );
 a4028a <=( a4027a  and  a4024a );
 a4031a <=( A232  and  (not A203) );
 a4035a <=( A300  and  A299 );
 a4036a <=( A234  and  a4035a );
 a4037a <=( a4036a  and  a4031a );
 a4040a <=( A166  and  A168 );
 a4043a <=( (not A202)  and  (not A201) );
 a4044a <=( a4043a  and  a4040a );
 a4047a <=( A232  and  (not A203) );
 a4051a <=( A300  and  A298 );
 a4052a <=( A234  and  a4051a );
 a4053a <=( a4052a  and  a4047a );
 a4056a <=( A166  and  A168 );
 a4059a <=( (not A202)  and  (not A201) );
 a4060a <=( a4059a  and  a4056a );
 a4063a <=( A232  and  (not A203) );
 a4067a <=( A267  and  A265 );
 a4068a <=( A234  and  a4067a );
 a4069a <=( a4068a  and  a4063a );
 a4072a <=( A166  and  A168 );
 a4075a <=( (not A202)  and  (not A201) );
 a4076a <=( a4075a  and  a4072a );
 a4079a <=( A232  and  (not A203) );
 a4083a <=( A267  and  A266 );
 a4084a <=( A234  and  a4083a );
 a4085a <=( a4084a  and  a4079a );
 a4088a <=( A166  and  A168 );
 a4091a <=( (not A202)  and  (not A201) );
 a4092a <=( a4091a  and  a4088a );
 a4095a <=( A233  and  (not A203) );
 a4099a <=( A300  and  A299 );
 a4100a <=( A234  and  a4099a );
 a4101a <=( a4100a  and  a4095a );
 a4104a <=( A166  and  A168 );
 a4107a <=( (not A202)  and  (not A201) );
 a4108a <=( a4107a  and  a4104a );
 a4111a <=( A233  and  (not A203) );
 a4115a <=( A300  and  A298 );
 a4116a <=( A234  and  a4115a );
 a4117a <=( a4116a  and  a4111a );
 a4120a <=( A166  and  A168 );
 a4123a <=( (not A202)  and  (not A201) );
 a4124a <=( a4123a  and  a4120a );
 a4127a <=( A233  and  (not A203) );
 a4131a <=( A267  and  A265 );
 a4132a <=( A234  and  a4131a );
 a4133a <=( a4132a  and  a4127a );
 a4136a <=( A166  and  A168 );
 a4139a <=( (not A202)  and  (not A201) );
 a4140a <=( a4139a  and  a4136a );
 a4143a <=( A233  and  (not A203) );
 a4147a <=( A267  and  A266 );
 a4148a <=( A234  and  a4147a );
 a4149a <=( a4148a  and  a4143a );
 a4152a <=( A166  and  A168 );
 a4155a <=( (not A202)  and  (not A201) );
 a4156a <=( a4155a  and  a4152a );
 a4159a <=( (not A232)  and  (not A203) );
 a4163a <=( A301  and  A236 );
 a4164a <=( A233  and  a4163a );
 a4165a <=( a4164a  and  a4159a );
 a4168a <=( A166  and  A168 );
 a4171a <=( (not A202)  and  (not A201) );
 a4172a <=( a4171a  and  a4168a );
 a4175a <=( (not A232)  and  (not A203) );
 a4179a <=( A268  and  A236 );
 a4180a <=( A233  and  a4179a );
 a4181a <=( a4180a  and  a4175a );
 a4184a <=( A166  and  A168 );
 a4187a <=( (not A202)  and  (not A201) );
 a4188a <=( a4187a  and  a4184a );
 a4191a <=( A232  and  (not A203) );
 a4195a <=( A301  and  A236 );
 a4196a <=( (not A233)  and  a4195a );
 a4197a <=( a4196a  and  a4191a );
 a4200a <=( A166  and  A168 );
 a4203a <=( (not A202)  and  (not A201) );
 a4204a <=( a4203a  and  a4200a );
 a4207a <=( A232  and  (not A203) );
 a4211a <=( A268  and  A236 );
 a4212a <=( (not A233)  and  a4211a );
 a4213a <=( a4212a  and  a4207a );
 a4216a <=( A166  and  A168 );
 a4219a <=( A200  and  A199 );
 a4220a <=( a4219a  and  a4216a );
 a4223a <=( (not A202)  and  (not A201) );
 a4227a <=( A300  and  A299 );
 a4228a <=( A235  and  a4227a );
 a4229a <=( a4228a  and  a4223a );
 a4232a <=( A166  and  A168 );
 a4235a <=( A200  and  A199 );
 a4236a <=( a4235a  and  a4232a );
 a4239a <=( (not A202)  and  (not A201) );
 a4243a <=( A300  and  A298 );
 a4244a <=( A235  and  a4243a );
 a4245a <=( a4244a  and  a4239a );
 a4248a <=( A166  and  A168 );
 a4251a <=( A200  and  A199 );
 a4252a <=( a4251a  and  a4248a );
 a4255a <=( (not A202)  and  (not A201) );
 a4259a <=( A267  and  A265 );
 a4260a <=( A235  and  a4259a );
 a4261a <=( a4260a  and  a4255a );
 a4264a <=( A166  and  A168 );
 a4267a <=( A200  and  A199 );
 a4268a <=( a4267a  and  a4264a );
 a4271a <=( (not A202)  and  (not A201) );
 a4275a <=( A267  and  A266 );
 a4276a <=( A235  and  a4275a );
 a4277a <=( a4276a  and  a4271a );
 a4280a <=( A166  and  A168 );
 a4283a <=( A200  and  A199 );
 a4284a <=( a4283a  and  a4280a );
 a4287a <=( (not A202)  and  (not A201) );
 a4291a <=( A301  and  A234 );
 a4292a <=( A232  and  a4291a );
 a4293a <=( a4292a  and  a4287a );
 a4296a <=( A166  and  A168 );
 a4299a <=( A200  and  A199 );
 a4300a <=( a4299a  and  a4296a );
 a4303a <=( (not A202)  and  (not A201) );
 a4307a <=( A268  and  A234 );
 a4308a <=( A232  and  a4307a );
 a4309a <=( a4308a  and  a4303a );
 a4312a <=( A166  and  A168 );
 a4315a <=( A200  and  A199 );
 a4316a <=( a4315a  and  a4312a );
 a4319a <=( (not A202)  and  (not A201) );
 a4323a <=( A301  and  A234 );
 a4324a <=( A233  and  a4323a );
 a4325a <=( a4324a  and  a4319a );
 a4328a <=( A166  and  A168 );
 a4331a <=( A200  and  A199 );
 a4332a <=( a4331a  and  a4328a );
 a4335a <=( (not A202)  and  (not A201) );
 a4339a <=( A268  and  A234 );
 a4340a <=( A233  and  a4339a );
 a4341a <=( a4340a  and  a4335a );
 a4344a <=( A166  and  A168 );
 a4347a <=( (not A200)  and  (not A199) );
 a4348a <=( a4347a  and  a4344a );
 a4351a <=( A235  and  (not A202) );
 a4355a <=( A302  and  (not A299) );
 a4356a <=( A298  and  a4355a );
 a4357a <=( a4356a  and  a4351a );
 a4360a <=( A166  and  A168 );
 a4363a <=( (not A200)  and  (not A199) );
 a4364a <=( a4363a  and  a4360a );
 a4367a <=( A235  and  (not A202) );
 a4371a <=( A302  and  A299 );
 a4372a <=( (not A298)  and  a4371a );
 a4373a <=( a4372a  and  a4367a );
 a4376a <=( A166  and  A168 );
 a4379a <=( (not A200)  and  (not A199) );
 a4380a <=( a4379a  and  a4376a );
 a4383a <=( A235  and  (not A202) );
 a4387a <=( A269  and  A266 );
 a4388a <=( (not A265)  and  a4387a );
 a4389a <=( a4388a  and  a4383a );
 a4392a <=( A166  and  A168 );
 a4395a <=( (not A200)  and  (not A199) );
 a4396a <=( a4395a  and  a4392a );
 a4399a <=( A235  and  (not A202) );
 a4403a <=( A269  and  (not A266) );
 a4404a <=( A265  and  a4403a );
 a4405a <=( a4404a  and  a4399a );
 a4408a <=( A166  and  A168 );
 a4411a <=( (not A200)  and  (not A199) );
 a4412a <=( a4411a  and  a4408a );
 a4415a <=( A232  and  (not A202) );
 a4419a <=( A300  and  A299 );
 a4420a <=( A234  and  a4419a );
 a4421a <=( a4420a  and  a4415a );
 a4424a <=( A166  and  A168 );
 a4427a <=( (not A200)  and  (not A199) );
 a4428a <=( a4427a  and  a4424a );
 a4431a <=( A232  and  (not A202) );
 a4435a <=( A300  and  A298 );
 a4436a <=( A234  and  a4435a );
 a4437a <=( a4436a  and  a4431a );
 a4440a <=( A166  and  A168 );
 a4443a <=( (not A200)  and  (not A199) );
 a4444a <=( a4443a  and  a4440a );
 a4447a <=( A232  and  (not A202) );
 a4451a <=( A267  and  A265 );
 a4452a <=( A234  and  a4451a );
 a4453a <=( a4452a  and  a4447a );
 a4456a <=( A166  and  A168 );
 a4459a <=( (not A200)  and  (not A199) );
 a4460a <=( a4459a  and  a4456a );
 a4463a <=( A232  and  (not A202) );
 a4467a <=( A267  and  A266 );
 a4468a <=( A234  and  a4467a );
 a4469a <=( a4468a  and  a4463a );
 a4472a <=( A166  and  A168 );
 a4475a <=( (not A200)  and  (not A199) );
 a4476a <=( a4475a  and  a4472a );
 a4479a <=( A233  and  (not A202) );
 a4483a <=( A300  and  A299 );
 a4484a <=( A234  and  a4483a );
 a4485a <=( a4484a  and  a4479a );
 a4488a <=( A166  and  A168 );
 a4491a <=( (not A200)  and  (not A199) );
 a4492a <=( a4491a  and  a4488a );
 a4495a <=( A233  and  (not A202) );
 a4499a <=( A300  and  A298 );
 a4500a <=( A234  and  a4499a );
 a4501a <=( a4500a  and  a4495a );
 a4504a <=( A166  and  A168 );
 a4507a <=( (not A200)  and  (not A199) );
 a4508a <=( a4507a  and  a4504a );
 a4511a <=( A233  and  (not A202) );
 a4515a <=( A267  and  A265 );
 a4516a <=( A234  and  a4515a );
 a4517a <=( a4516a  and  a4511a );
 a4520a <=( A166  and  A168 );
 a4523a <=( (not A200)  and  (not A199) );
 a4524a <=( a4523a  and  a4520a );
 a4527a <=( A233  and  (not A202) );
 a4531a <=( A267  and  A266 );
 a4532a <=( A234  and  a4531a );
 a4533a <=( a4532a  and  a4527a );
 a4536a <=( A166  and  A168 );
 a4539a <=( (not A200)  and  (not A199) );
 a4540a <=( a4539a  and  a4536a );
 a4543a <=( (not A232)  and  (not A202) );
 a4547a <=( A301  and  A236 );
 a4548a <=( A233  and  a4547a );
 a4549a <=( a4548a  and  a4543a );
 a4552a <=( A166  and  A168 );
 a4555a <=( (not A200)  and  (not A199) );
 a4556a <=( a4555a  and  a4552a );
 a4559a <=( (not A232)  and  (not A202) );
 a4563a <=( A268  and  A236 );
 a4564a <=( A233  and  a4563a );
 a4565a <=( a4564a  and  a4559a );
 a4568a <=( A166  and  A168 );
 a4571a <=( (not A200)  and  (not A199) );
 a4572a <=( a4571a  and  a4568a );
 a4575a <=( A232  and  (not A202) );
 a4579a <=( A301  and  A236 );
 a4580a <=( (not A233)  and  a4579a );
 a4581a <=( a4580a  and  a4575a );
 a4584a <=( A166  and  A168 );
 a4587a <=( (not A200)  and  (not A199) );
 a4588a <=( a4587a  and  a4584a );
 a4591a <=( A232  and  (not A202) );
 a4595a <=( A268  and  A236 );
 a4596a <=( (not A233)  and  a4595a );
 a4597a <=( a4596a  and  a4591a );
 a4600a <=( A167  and  A168 );
 a4603a <=( (not A202)  and  (not A201) );
 a4604a <=( a4603a  and  a4600a );
 a4607a <=( A235  and  (not A203) );
 a4611a <=( A302  and  (not A299) );
 a4612a <=( A298  and  a4611a );
 a4613a <=( a4612a  and  a4607a );
 a4616a <=( A167  and  A168 );
 a4619a <=( (not A202)  and  (not A201) );
 a4620a <=( a4619a  and  a4616a );
 a4623a <=( A235  and  (not A203) );
 a4627a <=( A302  and  A299 );
 a4628a <=( (not A298)  and  a4627a );
 a4629a <=( a4628a  and  a4623a );
 a4632a <=( A167  and  A168 );
 a4635a <=( (not A202)  and  (not A201) );
 a4636a <=( a4635a  and  a4632a );
 a4639a <=( A235  and  (not A203) );
 a4643a <=( A269  and  A266 );
 a4644a <=( (not A265)  and  a4643a );
 a4645a <=( a4644a  and  a4639a );
 a4648a <=( A167  and  A168 );
 a4651a <=( (not A202)  and  (not A201) );
 a4652a <=( a4651a  and  a4648a );
 a4655a <=( A235  and  (not A203) );
 a4659a <=( A269  and  (not A266) );
 a4660a <=( A265  and  a4659a );
 a4661a <=( a4660a  and  a4655a );
 a4664a <=( A167  and  A168 );
 a4667a <=( (not A202)  and  (not A201) );
 a4668a <=( a4667a  and  a4664a );
 a4671a <=( A232  and  (not A203) );
 a4675a <=( A300  and  A299 );
 a4676a <=( A234  and  a4675a );
 a4677a <=( a4676a  and  a4671a );
 a4680a <=( A167  and  A168 );
 a4683a <=( (not A202)  and  (not A201) );
 a4684a <=( a4683a  and  a4680a );
 a4687a <=( A232  and  (not A203) );
 a4691a <=( A300  and  A298 );
 a4692a <=( A234  and  a4691a );
 a4693a <=( a4692a  and  a4687a );
 a4696a <=( A167  and  A168 );
 a4699a <=( (not A202)  and  (not A201) );
 a4700a <=( a4699a  and  a4696a );
 a4703a <=( A232  and  (not A203) );
 a4707a <=( A267  and  A265 );
 a4708a <=( A234  and  a4707a );
 a4709a <=( a4708a  and  a4703a );
 a4712a <=( A167  and  A168 );
 a4715a <=( (not A202)  and  (not A201) );
 a4716a <=( a4715a  and  a4712a );
 a4719a <=( A232  and  (not A203) );
 a4723a <=( A267  and  A266 );
 a4724a <=( A234  and  a4723a );
 a4725a <=( a4724a  and  a4719a );
 a4728a <=( A167  and  A168 );
 a4731a <=( (not A202)  and  (not A201) );
 a4732a <=( a4731a  and  a4728a );
 a4735a <=( A233  and  (not A203) );
 a4739a <=( A300  and  A299 );
 a4740a <=( A234  and  a4739a );
 a4741a <=( a4740a  and  a4735a );
 a4744a <=( A167  and  A168 );
 a4747a <=( (not A202)  and  (not A201) );
 a4748a <=( a4747a  and  a4744a );
 a4751a <=( A233  and  (not A203) );
 a4755a <=( A300  and  A298 );
 a4756a <=( A234  and  a4755a );
 a4757a <=( a4756a  and  a4751a );
 a4760a <=( A167  and  A168 );
 a4763a <=( (not A202)  and  (not A201) );
 a4764a <=( a4763a  and  a4760a );
 a4767a <=( A233  and  (not A203) );
 a4771a <=( A267  and  A265 );
 a4772a <=( A234  and  a4771a );
 a4773a <=( a4772a  and  a4767a );
 a4776a <=( A167  and  A168 );
 a4779a <=( (not A202)  and  (not A201) );
 a4780a <=( a4779a  and  a4776a );
 a4783a <=( A233  and  (not A203) );
 a4787a <=( A267  and  A266 );
 a4788a <=( A234  and  a4787a );
 a4789a <=( a4788a  and  a4783a );
 a4792a <=( A167  and  A168 );
 a4795a <=( (not A202)  and  (not A201) );
 a4796a <=( a4795a  and  a4792a );
 a4799a <=( (not A232)  and  (not A203) );
 a4803a <=( A301  and  A236 );
 a4804a <=( A233  and  a4803a );
 a4805a <=( a4804a  and  a4799a );
 a4808a <=( A167  and  A168 );
 a4811a <=( (not A202)  and  (not A201) );
 a4812a <=( a4811a  and  a4808a );
 a4815a <=( (not A232)  and  (not A203) );
 a4819a <=( A268  and  A236 );
 a4820a <=( A233  and  a4819a );
 a4821a <=( a4820a  and  a4815a );
 a4824a <=( A167  and  A168 );
 a4827a <=( (not A202)  and  (not A201) );
 a4828a <=( a4827a  and  a4824a );
 a4831a <=( A232  and  (not A203) );
 a4835a <=( A301  and  A236 );
 a4836a <=( (not A233)  and  a4835a );
 a4837a <=( a4836a  and  a4831a );
 a4840a <=( A167  and  A168 );
 a4843a <=( (not A202)  and  (not A201) );
 a4844a <=( a4843a  and  a4840a );
 a4847a <=( A232  and  (not A203) );
 a4851a <=( A268  and  A236 );
 a4852a <=( (not A233)  and  a4851a );
 a4853a <=( a4852a  and  a4847a );
 a4856a <=( A167  and  A168 );
 a4859a <=( A200  and  A199 );
 a4860a <=( a4859a  and  a4856a );
 a4863a <=( (not A202)  and  (not A201) );
 a4867a <=( A300  and  A299 );
 a4868a <=( A235  and  a4867a );
 a4869a <=( a4868a  and  a4863a );
 a4872a <=( A167  and  A168 );
 a4875a <=( A200  and  A199 );
 a4876a <=( a4875a  and  a4872a );
 a4879a <=( (not A202)  and  (not A201) );
 a4883a <=( A300  and  A298 );
 a4884a <=( A235  and  a4883a );
 a4885a <=( a4884a  and  a4879a );
 a4888a <=( A167  and  A168 );
 a4891a <=( A200  and  A199 );
 a4892a <=( a4891a  and  a4888a );
 a4895a <=( (not A202)  and  (not A201) );
 a4899a <=( A267  and  A265 );
 a4900a <=( A235  and  a4899a );
 a4901a <=( a4900a  and  a4895a );
 a4904a <=( A167  and  A168 );
 a4907a <=( A200  and  A199 );
 a4908a <=( a4907a  and  a4904a );
 a4911a <=( (not A202)  and  (not A201) );
 a4915a <=( A267  and  A266 );
 a4916a <=( A235  and  a4915a );
 a4917a <=( a4916a  and  a4911a );
 a4920a <=( A167  and  A168 );
 a4923a <=( A200  and  A199 );
 a4924a <=( a4923a  and  a4920a );
 a4927a <=( (not A202)  and  (not A201) );
 a4931a <=( A301  and  A234 );
 a4932a <=( A232  and  a4931a );
 a4933a <=( a4932a  and  a4927a );
 a4936a <=( A167  and  A168 );
 a4939a <=( A200  and  A199 );
 a4940a <=( a4939a  and  a4936a );
 a4943a <=( (not A202)  and  (not A201) );
 a4947a <=( A268  and  A234 );
 a4948a <=( A232  and  a4947a );
 a4949a <=( a4948a  and  a4943a );
 a4952a <=( A167  and  A168 );
 a4955a <=( A200  and  A199 );
 a4956a <=( a4955a  and  a4952a );
 a4959a <=( (not A202)  and  (not A201) );
 a4963a <=( A301  and  A234 );
 a4964a <=( A233  and  a4963a );
 a4965a <=( a4964a  and  a4959a );
 a4968a <=( A167  and  A168 );
 a4971a <=( A200  and  A199 );
 a4972a <=( a4971a  and  a4968a );
 a4975a <=( (not A202)  and  (not A201) );
 a4979a <=( A268  and  A234 );
 a4980a <=( A233  and  a4979a );
 a4981a <=( a4980a  and  a4975a );
 a4984a <=( A167  and  A168 );
 a4987a <=( (not A200)  and  (not A199) );
 a4988a <=( a4987a  and  a4984a );
 a4991a <=( A235  and  (not A202) );
 a4995a <=( A302  and  (not A299) );
 a4996a <=( A298  and  a4995a );
 a4997a <=( a4996a  and  a4991a );
 a5000a <=( A167  and  A168 );
 a5003a <=( (not A200)  and  (not A199) );
 a5004a <=( a5003a  and  a5000a );
 a5007a <=( A235  and  (not A202) );
 a5011a <=( A302  and  A299 );
 a5012a <=( (not A298)  and  a5011a );
 a5013a <=( a5012a  and  a5007a );
 a5016a <=( A167  and  A168 );
 a5019a <=( (not A200)  and  (not A199) );
 a5020a <=( a5019a  and  a5016a );
 a5023a <=( A235  and  (not A202) );
 a5027a <=( A269  and  A266 );
 a5028a <=( (not A265)  and  a5027a );
 a5029a <=( a5028a  and  a5023a );
 a5032a <=( A167  and  A168 );
 a5035a <=( (not A200)  and  (not A199) );
 a5036a <=( a5035a  and  a5032a );
 a5039a <=( A235  and  (not A202) );
 a5043a <=( A269  and  (not A266) );
 a5044a <=( A265  and  a5043a );
 a5045a <=( a5044a  and  a5039a );
 a5048a <=( A167  and  A168 );
 a5051a <=( (not A200)  and  (not A199) );
 a5052a <=( a5051a  and  a5048a );
 a5055a <=( A232  and  (not A202) );
 a5059a <=( A300  and  A299 );
 a5060a <=( A234  and  a5059a );
 a5061a <=( a5060a  and  a5055a );
 a5064a <=( A167  and  A168 );
 a5067a <=( (not A200)  and  (not A199) );
 a5068a <=( a5067a  and  a5064a );
 a5071a <=( A232  and  (not A202) );
 a5075a <=( A300  and  A298 );
 a5076a <=( A234  and  a5075a );
 a5077a <=( a5076a  and  a5071a );
 a5080a <=( A167  and  A168 );
 a5083a <=( (not A200)  and  (not A199) );
 a5084a <=( a5083a  and  a5080a );
 a5087a <=( A232  and  (not A202) );
 a5091a <=( A267  and  A265 );
 a5092a <=( A234  and  a5091a );
 a5093a <=( a5092a  and  a5087a );
 a5096a <=( A167  and  A168 );
 a5099a <=( (not A200)  and  (not A199) );
 a5100a <=( a5099a  and  a5096a );
 a5103a <=( A232  and  (not A202) );
 a5107a <=( A267  and  A266 );
 a5108a <=( A234  and  a5107a );
 a5109a <=( a5108a  and  a5103a );
 a5112a <=( A167  and  A168 );
 a5115a <=( (not A200)  and  (not A199) );
 a5116a <=( a5115a  and  a5112a );
 a5119a <=( A233  and  (not A202) );
 a5123a <=( A300  and  A299 );
 a5124a <=( A234  and  a5123a );
 a5125a <=( a5124a  and  a5119a );
 a5128a <=( A167  and  A168 );
 a5131a <=( (not A200)  and  (not A199) );
 a5132a <=( a5131a  and  a5128a );
 a5135a <=( A233  and  (not A202) );
 a5139a <=( A300  and  A298 );
 a5140a <=( A234  and  a5139a );
 a5141a <=( a5140a  and  a5135a );
 a5144a <=( A167  and  A168 );
 a5147a <=( (not A200)  and  (not A199) );
 a5148a <=( a5147a  and  a5144a );
 a5151a <=( A233  and  (not A202) );
 a5155a <=( A267  and  A265 );
 a5156a <=( A234  and  a5155a );
 a5157a <=( a5156a  and  a5151a );
 a5160a <=( A167  and  A168 );
 a5163a <=( (not A200)  and  (not A199) );
 a5164a <=( a5163a  and  a5160a );
 a5167a <=( A233  and  (not A202) );
 a5171a <=( A267  and  A266 );
 a5172a <=( A234  and  a5171a );
 a5173a <=( a5172a  and  a5167a );
 a5176a <=( A167  and  A168 );
 a5179a <=( (not A200)  and  (not A199) );
 a5180a <=( a5179a  and  a5176a );
 a5183a <=( (not A232)  and  (not A202) );
 a5187a <=( A301  and  A236 );
 a5188a <=( A233  and  a5187a );
 a5189a <=( a5188a  and  a5183a );
 a5192a <=( A167  and  A168 );
 a5195a <=( (not A200)  and  (not A199) );
 a5196a <=( a5195a  and  a5192a );
 a5199a <=( (not A232)  and  (not A202) );
 a5203a <=( A268  and  A236 );
 a5204a <=( A233  and  a5203a );
 a5205a <=( a5204a  and  a5199a );
 a5208a <=( A167  and  A168 );
 a5211a <=( (not A200)  and  (not A199) );
 a5212a <=( a5211a  and  a5208a );
 a5215a <=( A232  and  (not A202) );
 a5219a <=( A301  and  A236 );
 a5220a <=( (not A233)  and  a5219a );
 a5221a <=( a5220a  and  a5215a );
 a5224a <=( A167  and  A168 );
 a5227a <=( (not A200)  and  (not A199) );
 a5228a <=( a5227a  and  a5224a );
 a5231a <=( A232  and  (not A202) );
 a5235a <=( A268  and  A236 );
 a5236a <=( (not A233)  and  a5235a );
 a5237a <=( a5236a  and  a5231a );
 a5240a <=( A167  and  A170 );
 a5243a <=( (not A201)  and  (not A166) );
 a5244a <=( a5243a  and  a5240a );
 a5247a <=( (not A203)  and  (not A202) );
 a5251a <=( A300  and  A299 );
 a5252a <=( A235  and  a5251a );
 a5253a <=( a5252a  and  a5247a );
 a5256a <=( A167  and  A170 );
 a5259a <=( (not A201)  and  (not A166) );
 a5260a <=( a5259a  and  a5256a );
 a5263a <=( (not A203)  and  (not A202) );
 a5267a <=( A300  and  A298 );
 a5268a <=( A235  and  a5267a );
 a5269a <=( a5268a  and  a5263a );
 a5272a <=( A167  and  A170 );
 a5275a <=( (not A201)  and  (not A166) );
 a5276a <=( a5275a  and  a5272a );
 a5279a <=( (not A203)  and  (not A202) );
 a5283a <=( A267  and  A265 );
 a5284a <=( A235  and  a5283a );
 a5285a <=( a5284a  and  a5279a );
 a5288a <=( A167  and  A170 );
 a5291a <=( (not A201)  and  (not A166) );
 a5292a <=( a5291a  and  a5288a );
 a5295a <=( (not A203)  and  (not A202) );
 a5299a <=( A267  and  A266 );
 a5300a <=( A235  and  a5299a );
 a5301a <=( a5300a  and  a5295a );
 a5304a <=( A167  and  A170 );
 a5307a <=( (not A201)  and  (not A166) );
 a5308a <=( a5307a  and  a5304a );
 a5311a <=( (not A203)  and  (not A202) );
 a5315a <=( A301  and  A234 );
 a5316a <=( A232  and  a5315a );
 a5317a <=( a5316a  and  a5311a );
 a5320a <=( A167  and  A170 );
 a5323a <=( (not A201)  and  (not A166) );
 a5324a <=( a5323a  and  a5320a );
 a5327a <=( (not A203)  and  (not A202) );
 a5331a <=( A268  and  A234 );
 a5332a <=( A232  and  a5331a );
 a5333a <=( a5332a  and  a5327a );
 a5336a <=( A167  and  A170 );
 a5339a <=( (not A201)  and  (not A166) );
 a5340a <=( a5339a  and  a5336a );
 a5343a <=( (not A203)  and  (not A202) );
 a5347a <=( A301  and  A234 );
 a5348a <=( A233  and  a5347a );
 a5349a <=( a5348a  and  a5343a );
 a5352a <=( A167  and  A170 );
 a5355a <=( (not A201)  and  (not A166) );
 a5356a <=( a5355a  and  a5352a );
 a5359a <=( (not A203)  and  (not A202) );
 a5363a <=( A268  and  A234 );
 a5364a <=( A233  and  a5363a );
 a5365a <=( a5364a  and  a5359a );
 a5368a <=( A167  and  A170 );
 a5371a <=( A199  and  (not A166) );
 a5372a <=( a5371a  and  a5368a );
 a5375a <=( (not A201)  and  A200 );
 a5379a <=( A301  and  A235 );
 a5380a <=( (not A202)  and  a5379a );
 a5381a <=( a5380a  and  a5375a );
 a5384a <=( A167  and  A170 );
 a5387a <=( A199  and  (not A166) );
 a5388a <=( a5387a  and  a5384a );
 a5391a <=( (not A201)  and  A200 );
 a5395a <=( A268  and  A235 );
 a5396a <=( (not A202)  and  a5395a );
 a5397a <=( a5396a  and  a5391a );
 a5400a <=( A167  and  A170 );
 a5403a <=( (not A199)  and  (not A166) );
 a5404a <=( a5403a  and  a5400a );
 a5407a <=( (not A202)  and  (not A200) );
 a5411a <=( A300  and  A299 );
 a5412a <=( A235  and  a5411a );
 a5413a <=( a5412a  and  a5407a );
 a5416a <=( A167  and  A170 );
 a5419a <=( (not A199)  and  (not A166) );
 a5420a <=( a5419a  and  a5416a );
 a5423a <=( (not A202)  and  (not A200) );
 a5427a <=( A300  and  A298 );
 a5428a <=( A235  and  a5427a );
 a5429a <=( a5428a  and  a5423a );
 a5432a <=( A167  and  A170 );
 a5435a <=( (not A199)  and  (not A166) );
 a5436a <=( a5435a  and  a5432a );
 a5439a <=( (not A202)  and  (not A200) );
 a5443a <=( A267  and  A265 );
 a5444a <=( A235  and  a5443a );
 a5445a <=( a5444a  and  a5439a );
 a5448a <=( A167  and  A170 );
 a5451a <=( (not A199)  and  (not A166) );
 a5452a <=( a5451a  and  a5448a );
 a5455a <=( (not A202)  and  (not A200) );
 a5459a <=( A267  and  A266 );
 a5460a <=( A235  and  a5459a );
 a5461a <=( a5460a  and  a5455a );
 a5464a <=( A167  and  A170 );
 a5467a <=( (not A199)  and  (not A166) );
 a5468a <=( a5467a  and  a5464a );
 a5471a <=( (not A202)  and  (not A200) );
 a5475a <=( A301  and  A234 );
 a5476a <=( A232  and  a5475a );
 a5477a <=( a5476a  and  a5471a );
 a5480a <=( A167  and  A170 );
 a5483a <=( (not A199)  and  (not A166) );
 a5484a <=( a5483a  and  a5480a );
 a5487a <=( (not A202)  and  (not A200) );
 a5491a <=( A268  and  A234 );
 a5492a <=( A232  and  a5491a );
 a5493a <=( a5492a  and  a5487a );
 a5496a <=( A167  and  A170 );
 a5499a <=( (not A199)  and  (not A166) );
 a5500a <=( a5499a  and  a5496a );
 a5503a <=( (not A202)  and  (not A200) );
 a5507a <=( A301  and  A234 );
 a5508a <=( A233  and  a5507a );
 a5509a <=( a5508a  and  a5503a );
 a5512a <=( A167  and  A170 );
 a5515a <=( (not A199)  and  (not A166) );
 a5516a <=( a5515a  and  a5512a );
 a5519a <=( (not A202)  and  (not A200) );
 a5523a <=( A268  and  A234 );
 a5524a <=( A233  and  a5523a );
 a5525a <=( a5524a  and  a5519a );
 a5528a <=( (not A167)  and  A170 );
 a5531a <=( (not A201)  and  A166 );
 a5532a <=( a5531a  and  a5528a );
 a5535a <=( (not A203)  and  (not A202) );
 a5539a <=( A300  and  A299 );
 a5540a <=( A235  and  a5539a );
 a5541a <=( a5540a  and  a5535a );
 a5544a <=( (not A167)  and  A170 );
 a5547a <=( (not A201)  and  A166 );
 a5548a <=( a5547a  and  a5544a );
 a5551a <=( (not A203)  and  (not A202) );
 a5555a <=( A300  and  A298 );
 a5556a <=( A235  and  a5555a );
 a5557a <=( a5556a  and  a5551a );
 a5560a <=( (not A167)  and  A170 );
 a5563a <=( (not A201)  and  A166 );
 a5564a <=( a5563a  and  a5560a );
 a5567a <=( (not A203)  and  (not A202) );
 a5571a <=( A267  and  A265 );
 a5572a <=( A235  and  a5571a );
 a5573a <=( a5572a  and  a5567a );
 a5576a <=( (not A167)  and  A170 );
 a5579a <=( (not A201)  and  A166 );
 a5580a <=( a5579a  and  a5576a );
 a5583a <=( (not A203)  and  (not A202) );
 a5587a <=( A267  and  A266 );
 a5588a <=( A235  and  a5587a );
 a5589a <=( a5588a  and  a5583a );
 a5592a <=( (not A167)  and  A170 );
 a5595a <=( (not A201)  and  A166 );
 a5596a <=( a5595a  and  a5592a );
 a5599a <=( (not A203)  and  (not A202) );
 a5603a <=( A301  and  A234 );
 a5604a <=( A232  and  a5603a );
 a5605a <=( a5604a  and  a5599a );
 a5608a <=( (not A167)  and  A170 );
 a5611a <=( (not A201)  and  A166 );
 a5612a <=( a5611a  and  a5608a );
 a5615a <=( (not A203)  and  (not A202) );
 a5619a <=( A268  and  A234 );
 a5620a <=( A232  and  a5619a );
 a5621a <=( a5620a  and  a5615a );
 a5624a <=( (not A167)  and  A170 );
 a5627a <=( (not A201)  and  A166 );
 a5628a <=( a5627a  and  a5624a );
 a5631a <=( (not A203)  and  (not A202) );
 a5635a <=( A301  and  A234 );
 a5636a <=( A233  and  a5635a );
 a5637a <=( a5636a  and  a5631a );
 a5640a <=( (not A167)  and  A170 );
 a5643a <=( (not A201)  and  A166 );
 a5644a <=( a5643a  and  a5640a );
 a5647a <=( (not A203)  and  (not A202) );
 a5651a <=( A268  and  A234 );
 a5652a <=( A233  and  a5651a );
 a5653a <=( a5652a  and  a5647a );
 a5656a <=( (not A167)  and  A170 );
 a5659a <=( A199  and  A166 );
 a5660a <=( a5659a  and  a5656a );
 a5663a <=( (not A201)  and  A200 );
 a5667a <=( A301  and  A235 );
 a5668a <=( (not A202)  and  a5667a );
 a5669a <=( a5668a  and  a5663a );
 a5672a <=( (not A167)  and  A170 );
 a5675a <=( A199  and  A166 );
 a5676a <=( a5675a  and  a5672a );
 a5679a <=( (not A201)  and  A200 );
 a5683a <=( A268  and  A235 );
 a5684a <=( (not A202)  and  a5683a );
 a5685a <=( a5684a  and  a5679a );
 a5688a <=( (not A167)  and  A170 );
 a5691a <=( (not A199)  and  A166 );
 a5692a <=( a5691a  and  a5688a );
 a5695a <=( (not A202)  and  (not A200) );
 a5699a <=( A300  and  A299 );
 a5700a <=( A235  and  a5699a );
 a5701a <=( a5700a  and  a5695a );
 a5704a <=( (not A167)  and  A170 );
 a5707a <=( (not A199)  and  A166 );
 a5708a <=( a5707a  and  a5704a );
 a5711a <=( (not A202)  and  (not A200) );
 a5715a <=( A300  and  A298 );
 a5716a <=( A235  and  a5715a );
 a5717a <=( a5716a  and  a5711a );
 a5720a <=( (not A167)  and  A170 );
 a5723a <=( (not A199)  and  A166 );
 a5724a <=( a5723a  and  a5720a );
 a5727a <=( (not A202)  and  (not A200) );
 a5731a <=( A267  and  A265 );
 a5732a <=( A235  and  a5731a );
 a5733a <=( a5732a  and  a5727a );
 a5736a <=( (not A167)  and  A170 );
 a5739a <=( (not A199)  and  A166 );
 a5740a <=( a5739a  and  a5736a );
 a5743a <=( (not A202)  and  (not A200) );
 a5747a <=( A267  and  A266 );
 a5748a <=( A235  and  a5747a );
 a5749a <=( a5748a  and  a5743a );
 a5752a <=( (not A167)  and  A170 );
 a5755a <=( (not A199)  and  A166 );
 a5756a <=( a5755a  and  a5752a );
 a5759a <=( (not A202)  and  (not A200) );
 a5763a <=( A301  and  A234 );
 a5764a <=( A232  and  a5763a );
 a5765a <=( a5764a  and  a5759a );
 a5768a <=( (not A167)  and  A170 );
 a5771a <=( (not A199)  and  A166 );
 a5772a <=( a5771a  and  a5768a );
 a5775a <=( (not A202)  and  (not A200) );
 a5779a <=( A268  and  A234 );
 a5780a <=( A232  and  a5779a );
 a5781a <=( a5780a  and  a5775a );
 a5784a <=( (not A167)  and  A170 );
 a5787a <=( (not A199)  and  A166 );
 a5788a <=( a5787a  and  a5784a );
 a5791a <=( (not A202)  and  (not A200) );
 a5795a <=( A301  and  A234 );
 a5796a <=( A233  and  a5795a );
 a5797a <=( a5796a  and  a5791a );
 a5800a <=( (not A167)  and  A170 );
 a5803a <=( (not A199)  and  A166 );
 a5804a <=( a5803a  and  a5800a );
 a5807a <=( (not A202)  and  (not A200) );
 a5811a <=( A268  and  A234 );
 a5812a <=( A233  and  a5811a );
 a5813a <=( a5812a  and  a5807a );
 a5816a <=( (not A201)  and  A169 );
 a5819a <=( (not A203)  and  (not A202) );
 a5820a <=( a5819a  and  a5816a );
 a5823a <=( A234  and  A232 );
 a5827a <=( A302  and  (not A299) );
 a5828a <=( A298  and  a5827a );
 a5829a <=( a5828a  and  a5823a );
 a5832a <=( (not A201)  and  A169 );
 a5835a <=( (not A203)  and  (not A202) );
 a5836a <=( a5835a  and  a5832a );
 a5839a <=( A234  and  A232 );
 a5843a <=( A302  and  A299 );
 a5844a <=( (not A298)  and  a5843a );
 a5845a <=( a5844a  and  a5839a );
 a5848a <=( (not A201)  and  A169 );
 a5851a <=( (not A203)  and  (not A202) );
 a5852a <=( a5851a  and  a5848a );
 a5855a <=( A234  and  A232 );
 a5859a <=( A269  and  A266 );
 a5860a <=( (not A265)  and  a5859a );
 a5861a <=( a5860a  and  a5855a );
 a5864a <=( (not A201)  and  A169 );
 a5867a <=( (not A203)  and  (not A202) );
 a5868a <=( a5867a  and  a5864a );
 a5871a <=( A234  and  A232 );
 a5875a <=( A269  and  (not A266) );
 a5876a <=( A265  and  a5875a );
 a5877a <=( a5876a  and  a5871a );
 a5880a <=( (not A201)  and  A169 );
 a5883a <=( (not A203)  and  (not A202) );
 a5884a <=( a5883a  and  a5880a );
 a5887a <=( A234  and  A233 );
 a5891a <=( A302  and  (not A299) );
 a5892a <=( A298  and  a5891a );
 a5893a <=( a5892a  and  a5887a );
 a5896a <=( (not A201)  and  A169 );
 a5899a <=( (not A203)  and  (not A202) );
 a5900a <=( a5899a  and  a5896a );
 a5903a <=( A234  and  A233 );
 a5907a <=( A302  and  A299 );
 a5908a <=( (not A298)  and  a5907a );
 a5909a <=( a5908a  and  a5903a );
 a5912a <=( (not A201)  and  A169 );
 a5915a <=( (not A203)  and  (not A202) );
 a5916a <=( a5915a  and  a5912a );
 a5919a <=( A234  and  A233 );
 a5923a <=( A269  and  A266 );
 a5924a <=( (not A265)  and  a5923a );
 a5925a <=( a5924a  and  a5919a );
 a5928a <=( (not A201)  and  A169 );
 a5931a <=( (not A203)  and  (not A202) );
 a5932a <=( a5931a  and  a5928a );
 a5935a <=( A234  and  A233 );
 a5939a <=( A269  and  (not A266) );
 a5940a <=( A265  and  a5939a );
 a5941a <=( a5940a  and  a5935a );
 a5944a <=( (not A201)  and  A169 );
 a5947a <=( (not A203)  and  (not A202) );
 a5948a <=( a5947a  and  a5944a );
 a5951a <=( A233  and  (not A232) );
 a5955a <=( A300  and  A299 );
 a5956a <=( A236  and  a5955a );
 a5957a <=( a5956a  and  a5951a );
 a5960a <=( (not A201)  and  A169 );
 a5963a <=( (not A203)  and  (not A202) );
 a5964a <=( a5963a  and  a5960a );
 a5967a <=( A233  and  (not A232) );
 a5971a <=( A300  and  A298 );
 a5972a <=( A236  and  a5971a );
 a5973a <=( a5972a  and  a5967a );
 a5976a <=( (not A201)  and  A169 );
 a5979a <=( (not A203)  and  (not A202) );
 a5980a <=( a5979a  and  a5976a );
 a5983a <=( A233  and  (not A232) );
 a5987a <=( A267  and  A265 );
 a5988a <=( A236  and  a5987a );
 a5989a <=( a5988a  and  a5983a );
 a5992a <=( (not A201)  and  A169 );
 a5995a <=( (not A203)  and  (not A202) );
 a5996a <=( a5995a  and  a5992a );
 a5999a <=( A233  and  (not A232) );
 a6003a <=( A267  and  A266 );
 a6004a <=( A236  and  a6003a );
 a6005a <=( a6004a  and  a5999a );
 a6008a <=( (not A201)  and  A169 );
 a6011a <=( (not A203)  and  (not A202) );
 a6012a <=( a6011a  and  a6008a );
 a6015a <=( (not A233)  and  A232 );
 a6019a <=( A300  and  A299 );
 a6020a <=( A236  and  a6019a );
 a6021a <=( a6020a  and  a6015a );
 a6024a <=( (not A201)  and  A169 );
 a6027a <=( (not A203)  and  (not A202) );
 a6028a <=( a6027a  and  a6024a );
 a6031a <=( (not A233)  and  A232 );
 a6035a <=( A300  and  A298 );
 a6036a <=( A236  and  a6035a );
 a6037a <=( a6036a  and  a6031a );
 a6040a <=( (not A201)  and  A169 );
 a6043a <=( (not A203)  and  (not A202) );
 a6044a <=( a6043a  and  a6040a );
 a6047a <=( (not A233)  and  A232 );
 a6051a <=( A267  and  A265 );
 a6052a <=( A236  and  a6051a );
 a6053a <=( a6052a  and  a6047a );
 a6056a <=( (not A201)  and  A169 );
 a6059a <=( (not A203)  and  (not A202) );
 a6060a <=( a6059a  and  a6056a );
 a6063a <=( (not A233)  and  A232 );
 a6067a <=( A267  and  A266 );
 a6068a <=( A236  and  a6067a );
 a6069a <=( a6068a  and  a6063a );
 a6072a <=( A199  and  A169 );
 a6075a <=( (not A201)  and  A200 );
 a6076a <=( a6075a  and  a6072a );
 a6079a <=( A235  and  (not A202) );
 a6083a <=( A302  and  (not A299) );
 a6084a <=( A298  and  a6083a );
 a6085a <=( a6084a  and  a6079a );
 a6088a <=( A199  and  A169 );
 a6091a <=( (not A201)  and  A200 );
 a6092a <=( a6091a  and  a6088a );
 a6095a <=( A235  and  (not A202) );
 a6099a <=( A302  and  A299 );
 a6100a <=( (not A298)  and  a6099a );
 a6101a <=( a6100a  and  a6095a );
 a6104a <=( A199  and  A169 );
 a6107a <=( (not A201)  and  A200 );
 a6108a <=( a6107a  and  a6104a );
 a6111a <=( A235  and  (not A202) );
 a6115a <=( A269  and  A266 );
 a6116a <=( (not A265)  and  a6115a );
 a6117a <=( a6116a  and  a6111a );
 a6120a <=( A199  and  A169 );
 a6123a <=( (not A201)  and  A200 );
 a6124a <=( a6123a  and  a6120a );
 a6127a <=( A235  and  (not A202) );
 a6131a <=( A269  and  (not A266) );
 a6132a <=( A265  and  a6131a );
 a6133a <=( a6132a  and  a6127a );
 a6136a <=( A199  and  A169 );
 a6139a <=( (not A201)  and  A200 );
 a6140a <=( a6139a  and  a6136a );
 a6143a <=( A232  and  (not A202) );
 a6147a <=( A300  and  A299 );
 a6148a <=( A234  and  a6147a );
 a6149a <=( a6148a  and  a6143a );
 a6152a <=( A199  and  A169 );
 a6155a <=( (not A201)  and  A200 );
 a6156a <=( a6155a  and  a6152a );
 a6159a <=( A232  and  (not A202) );
 a6163a <=( A300  and  A298 );
 a6164a <=( A234  and  a6163a );
 a6165a <=( a6164a  and  a6159a );
 a6168a <=( A199  and  A169 );
 a6171a <=( (not A201)  and  A200 );
 a6172a <=( a6171a  and  a6168a );
 a6175a <=( A232  and  (not A202) );
 a6179a <=( A267  and  A265 );
 a6180a <=( A234  and  a6179a );
 a6181a <=( a6180a  and  a6175a );
 a6184a <=( A199  and  A169 );
 a6187a <=( (not A201)  and  A200 );
 a6188a <=( a6187a  and  a6184a );
 a6191a <=( A232  and  (not A202) );
 a6195a <=( A267  and  A266 );
 a6196a <=( A234  and  a6195a );
 a6197a <=( a6196a  and  a6191a );
 a6200a <=( A199  and  A169 );
 a6203a <=( (not A201)  and  A200 );
 a6204a <=( a6203a  and  a6200a );
 a6207a <=( A233  and  (not A202) );
 a6211a <=( A300  and  A299 );
 a6212a <=( A234  and  a6211a );
 a6213a <=( a6212a  and  a6207a );
 a6216a <=( A199  and  A169 );
 a6219a <=( (not A201)  and  A200 );
 a6220a <=( a6219a  and  a6216a );
 a6223a <=( A233  and  (not A202) );
 a6227a <=( A300  and  A298 );
 a6228a <=( A234  and  a6227a );
 a6229a <=( a6228a  and  a6223a );
 a6232a <=( A199  and  A169 );
 a6235a <=( (not A201)  and  A200 );
 a6236a <=( a6235a  and  a6232a );
 a6239a <=( A233  and  (not A202) );
 a6243a <=( A267  and  A265 );
 a6244a <=( A234  and  a6243a );
 a6245a <=( a6244a  and  a6239a );
 a6248a <=( A199  and  A169 );
 a6251a <=( (not A201)  and  A200 );
 a6252a <=( a6251a  and  a6248a );
 a6255a <=( A233  and  (not A202) );
 a6259a <=( A267  and  A266 );
 a6260a <=( A234  and  a6259a );
 a6261a <=( a6260a  and  a6255a );
 a6264a <=( A199  and  A169 );
 a6267a <=( (not A201)  and  A200 );
 a6268a <=( a6267a  and  a6264a );
 a6271a <=( (not A232)  and  (not A202) );
 a6275a <=( A301  and  A236 );
 a6276a <=( A233  and  a6275a );
 a6277a <=( a6276a  and  a6271a );
 a6280a <=( A199  and  A169 );
 a6283a <=( (not A201)  and  A200 );
 a6284a <=( a6283a  and  a6280a );
 a6287a <=( (not A232)  and  (not A202) );
 a6291a <=( A268  and  A236 );
 a6292a <=( A233  and  a6291a );
 a6293a <=( a6292a  and  a6287a );
 a6296a <=( A199  and  A169 );
 a6299a <=( (not A201)  and  A200 );
 a6300a <=( a6299a  and  a6296a );
 a6303a <=( A232  and  (not A202) );
 a6307a <=( A301  and  A236 );
 a6308a <=( (not A233)  and  a6307a );
 a6309a <=( a6308a  and  a6303a );
 a6312a <=( A199  and  A169 );
 a6315a <=( (not A201)  and  A200 );
 a6316a <=( a6315a  and  a6312a );
 a6319a <=( A232  and  (not A202) );
 a6323a <=( A268  and  A236 );
 a6324a <=( (not A233)  and  a6323a );
 a6325a <=( a6324a  and  a6319a );
 a6328a <=( (not A199)  and  A169 );
 a6331a <=( (not A202)  and  (not A200) );
 a6332a <=( a6331a  and  a6328a );
 a6335a <=( A234  and  A232 );
 a6339a <=( A302  and  (not A299) );
 a6340a <=( A298  and  a6339a );
 a6341a <=( a6340a  and  a6335a );
 a6344a <=( (not A199)  and  A169 );
 a6347a <=( (not A202)  and  (not A200) );
 a6348a <=( a6347a  and  a6344a );
 a6351a <=( A234  and  A232 );
 a6355a <=( A302  and  A299 );
 a6356a <=( (not A298)  and  a6355a );
 a6357a <=( a6356a  and  a6351a );
 a6360a <=( (not A199)  and  A169 );
 a6363a <=( (not A202)  and  (not A200) );
 a6364a <=( a6363a  and  a6360a );
 a6367a <=( A234  and  A232 );
 a6371a <=( A269  and  A266 );
 a6372a <=( (not A265)  and  a6371a );
 a6373a <=( a6372a  and  a6367a );
 a6376a <=( (not A199)  and  A169 );
 a6379a <=( (not A202)  and  (not A200) );
 a6380a <=( a6379a  and  a6376a );
 a6383a <=( A234  and  A232 );
 a6387a <=( A269  and  (not A266) );
 a6388a <=( A265  and  a6387a );
 a6389a <=( a6388a  and  a6383a );
 a6392a <=( (not A199)  and  A169 );
 a6395a <=( (not A202)  and  (not A200) );
 a6396a <=( a6395a  and  a6392a );
 a6399a <=( A234  and  A233 );
 a6403a <=( A302  and  (not A299) );
 a6404a <=( A298  and  a6403a );
 a6405a <=( a6404a  and  a6399a );
 a6408a <=( (not A199)  and  A169 );
 a6411a <=( (not A202)  and  (not A200) );
 a6412a <=( a6411a  and  a6408a );
 a6415a <=( A234  and  A233 );
 a6419a <=( A302  and  A299 );
 a6420a <=( (not A298)  and  a6419a );
 a6421a <=( a6420a  and  a6415a );
 a6424a <=( (not A199)  and  A169 );
 a6427a <=( (not A202)  and  (not A200) );
 a6428a <=( a6427a  and  a6424a );
 a6431a <=( A234  and  A233 );
 a6435a <=( A269  and  A266 );
 a6436a <=( (not A265)  and  a6435a );
 a6437a <=( a6436a  and  a6431a );
 a6440a <=( (not A199)  and  A169 );
 a6443a <=( (not A202)  and  (not A200) );
 a6444a <=( a6443a  and  a6440a );
 a6447a <=( A234  and  A233 );
 a6451a <=( A269  and  (not A266) );
 a6452a <=( A265  and  a6451a );
 a6453a <=( a6452a  and  a6447a );
 a6456a <=( (not A199)  and  A169 );
 a6459a <=( (not A202)  and  (not A200) );
 a6460a <=( a6459a  and  a6456a );
 a6463a <=( A233  and  (not A232) );
 a6467a <=( A300  and  A299 );
 a6468a <=( A236  and  a6467a );
 a6469a <=( a6468a  and  a6463a );
 a6472a <=( (not A199)  and  A169 );
 a6475a <=( (not A202)  and  (not A200) );
 a6476a <=( a6475a  and  a6472a );
 a6479a <=( A233  and  (not A232) );
 a6483a <=( A300  and  A298 );
 a6484a <=( A236  and  a6483a );
 a6485a <=( a6484a  and  a6479a );
 a6488a <=( (not A199)  and  A169 );
 a6491a <=( (not A202)  and  (not A200) );
 a6492a <=( a6491a  and  a6488a );
 a6495a <=( A233  and  (not A232) );
 a6499a <=( A267  and  A265 );
 a6500a <=( A236  and  a6499a );
 a6501a <=( a6500a  and  a6495a );
 a6504a <=( (not A199)  and  A169 );
 a6507a <=( (not A202)  and  (not A200) );
 a6508a <=( a6507a  and  a6504a );
 a6511a <=( A233  and  (not A232) );
 a6515a <=( A267  and  A266 );
 a6516a <=( A236  and  a6515a );
 a6517a <=( a6516a  and  a6511a );
 a6520a <=( (not A199)  and  A169 );
 a6523a <=( (not A202)  and  (not A200) );
 a6524a <=( a6523a  and  a6520a );
 a6527a <=( (not A233)  and  A232 );
 a6531a <=( A300  and  A299 );
 a6532a <=( A236  and  a6531a );
 a6533a <=( a6532a  and  a6527a );
 a6536a <=( (not A199)  and  A169 );
 a6539a <=( (not A202)  and  (not A200) );
 a6540a <=( a6539a  and  a6536a );
 a6543a <=( (not A233)  and  A232 );
 a6547a <=( A300  and  A298 );
 a6548a <=( A236  and  a6547a );
 a6549a <=( a6548a  and  a6543a );
 a6552a <=( (not A199)  and  A169 );
 a6555a <=( (not A202)  and  (not A200) );
 a6556a <=( a6555a  and  a6552a );
 a6559a <=( (not A233)  and  A232 );
 a6563a <=( A267  and  A265 );
 a6564a <=( A236  and  a6563a );
 a6565a <=( a6564a  and  a6559a );
 a6568a <=( (not A199)  and  A169 );
 a6571a <=( (not A202)  and  (not A200) );
 a6572a <=( a6571a  and  a6568a );
 a6575a <=( (not A233)  and  A232 );
 a6579a <=( A267  and  A266 );
 a6580a <=( A236  and  a6579a );
 a6581a <=( a6580a  and  a6575a );
 a6584a <=( A166  and  A168 );
 a6588a <=( (not A203)  and  (not A202) );
 a6589a <=( (not A201)  and  a6588a );
 a6590a <=( a6589a  and  a6584a );
 a6593a <=( A234  and  A232 );
 a6597a <=( A302  and  (not A299) );
 a6598a <=( A298  and  a6597a );
 a6599a <=( a6598a  and  a6593a );
 a6602a <=( A166  and  A168 );
 a6606a <=( (not A203)  and  (not A202) );
 a6607a <=( (not A201)  and  a6606a );
 a6608a <=( a6607a  and  a6602a );
 a6611a <=( A234  and  A232 );
 a6615a <=( A302  and  A299 );
 a6616a <=( (not A298)  and  a6615a );
 a6617a <=( a6616a  and  a6611a );
 a6620a <=( A166  and  A168 );
 a6624a <=( (not A203)  and  (not A202) );
 a6625a <=( (not A201)  and  a6624a );
 a6626a <=( a6625a  and  a6620a );
 a6629a <=( A234  and  A232 );
 a6633a <=( A269  and  A266 );
 a6634a <=( (not A265)  and  a6633a );
 a6635a <=( a6634a  and  a6629a );
 a6638a <=( A166  and  A168 );
 a6642a <=( (not A203)  and  (not A202) );
 a6643a <=( (not A201)  and  a6642a );
 a6644a <=( a6643a  and  a6638a );
 a6647a <=( A234  and  A232 );
 a6651a <=( A269  and  (not A266) );
 a6652a <=( A265  and  a6651a );
 a6653a <=( a6652a  and  a6647a );
 a6656a <=( A166  and  A168 );
 a6660a <=( (not A203)  and  (not A202) );
 a6661a <=( (not A201)  and  a6660a );
 a6662a <=( a6661a  and  a6656a );
 a6665a <=( A234  and  A233 );
 a6669a <=( A302  and  (not A299) );
 a6670a <=( A298  and  a6669a );
 a6671a <=( a6670a  and  a6665a );
 a6674a <=( A166  and  A168 );
 a6678a <=( (not A203)  and  (not A202) );
 a6679a <=( (not A201)  and  a6678a );
 a6680a <=( a6679a  and  a6674a );
 a6683a <=( A234  and  A233 );
 a6687a <=( A302  and  A299 );
 a6688a <=( (not A298)  and  a6687a );
 a6689a <=( a6688a  and  a6683a );
 a6692a <=( A166  and  A168 );
 a6696a <=( (not A203)  and  (not A202) );
 a6697a <=( (not A201)  and  a6696a );
 a6698a <=( a6697a  and  a6692a );
 a6701a <=( A234  and  A233 );
 a6705a <=( A269  and  A266 );
 a6706a <=( (not A265)  and  a6705a );
 a6707a <=( a6706a  and  a6701a );
 a6710a <=( A166  and  A168 );
 a6714a <=( (not A203)  and  (not A202) );
 a6715a <=( (not A201)  and  a6714a );
 a6716a <=( a6715a  and  a6710a );
 a6719a <=( A234  and  A233 );
 a6723a <=( A269  and  (not A266) );
 a6724a <=( A265  and  a6723a );
 a6725a <=( a6724a  and  a6719a );
 a6728a <=( A166  and  A168 );
 a6732a <=( (not A203)  and  (not A202) );
 a6733a <=( (not A201)  and  a6732a );
 a6734a <=( a6733a  and  a6728a );
 a6737a <=( A233  and  (not A232) );
 a6741a <=( A300  and  A299 );
 a6742a <=( A236  and  a6741a );
 a6743a <=( a6742a  and  a6737a );
 a6746a <=( A166  and  A168 );
 a6750a <=( (not A203)  and  (not A202) );
 a6751a <=( (not A201)  and  a6750a );
 a6752a <=( a6751a  and  a6746a );
 a6755a <=( A233  and  (not A232) );
 a6759a <=( A300  and  A298 );
 a6760a <=( A236  and  a6759a );
 a6761a <=( a6760a  and  a6755a );
 a6764a <=( A166  and  A168 );
 a6768a <=( (not A203)  and  (not A202) );
 a6769a <=( (not A201)  and  a6768a );
 a6770a <=( a6769a  and  a6764a );
 a6773a <=( A233  and  (not A232) );
 a6777a <=( A267  and  A265 );
 a6778a <=( A236  and  a6777a );
 a6779a <=( a6778a  and  a6773a );
 a6782a <=( A166  and  A168 );
 a6786a <=( (not A203)  and  (not A202) );
 a6787a <=( (not A201)  and  a6786a );
 a6788a <=( a6787a  and  a6782a );
 a6791a <=( A233  and  (not A232) );
 a6795a <=( A267  and  A266 );
 a6796a <=( A236  and  a6795a );
 a6797a <=( a6796a  and  a6791a );
 a6800a <=( A166  and  A168 );
 a6804a <=( (not A203)  and  (not A202) );
 a6805a <=( (not A201)  and  a6804a );
 a6806a <=( a6805a  and  a6800a );
 a6809a <=( (not A233)  and  A232 );
 a6813a <=( A300  and  A299 );
 a6814a <=( A236  and  a6813a );
 a6815a <=( a6814a  and  a6809a );
 a6818a <=( A166  and  A168 );
 a6822a <=( (not A203)  and  (not A202) );
 a6823a <=( (not A201)  and  a6822a );
 a6824a <=( a6823a  and  a6818a );
 a6827a <=( (not A233)  and  A232 );
 a6831a <=( A300  and  A298 );
 a6832a <=( A236  and  a6831a );
 a6833a <=( a6832a  and  a6827a );
 a6836a <=( A166  and  A168 );
 a6840a <=( (not A203)  and  (not A202) );
 a6841a <=( (not A201)  and  a6840a );
 a6842a <=( a6841a  and  a6836a );
 a6845a <=( (not A233)  and  A232 );
 a6849a <=( A267  and  A265 );
 a6850a <=( A236  and  a6849a );
 a6851a <=( a6850a  and  a6845a );
 a6854a <=( A166  and  A168 );
 a6858a <=( (not A203)  and  (not A202) );
 a6859a <=( (not A201)  and  a6858a );
 a6860a <=( a6859a  and  a6854a );
 a6863a <=( (not A233)  and  A232 );
 a6867a <=( A267  and  A266 );
 a6868a <=( A236  and  a6867a );
 a6869a <=( a6868a  and  a6863a );
 a6872a <=( A166  and  A168 );
 a6876a <=( (not A201)  and  A200 );
 a6877a <=( A199  and  a6876a );
 a6878a <=( a6877a  and  a6872a );
 a6881a <=( A235  and  (not A202) );
 a6885a <=( A302  and  (not A299) );
 a6886a <=( A298  and  a6885a );
 a6887a <=( a6886a  and  a6881a );
 a6890a <=( A166  and  A168 );
 a6894a <=( (not A201)  and  A200 );
 a6895a <=( A199  and  a6894a );
 a6896a <=( a6895a  and  a6890a );
 a6899a <=( A235  and  (not A202) );
 a6903a <=( A302  and  A299 );
 a6904a <=( (not A298)  and  a6903a );
 a6905a <=( a6904a  and  a6899a );
 a6908a <=( A166  and  A168 );
 a6912a <=( (not A201)  and  A200 );
 a6913a <=( A199  and  a6912a );
 a6914a <=( a6913a  and  a6908a );
 a6917a <=( A235  and  (not A202) );
 a6921a <=( A269  and  A266 );
 a6922a <=( (not A265)  and  a6921a );
 a6923a <=( a6922a  and  a6917a );
 a6926a <=( A166  and  A168 );
 a6930a <=( (not A201)  and  A200 );
 a6931a <=( A199  and  a6930a );
 a6932a <=( a6931a  and  a6926a );
 a6935a <=( A235  and  (not A202) );
 a6939a <=( A269  and  (not A266) );
 a6940a <=( A265  and  a6939a );
 a6941a <=( a6940a  and  a6935a );
 a6944a <=( A166  and  A168 );
 a6948a <=( (not A201)  and  A200 );
 a6949a <=( A199  and  a6948a );
 a6950a <=( a6949a  and  a6944a );
 a6953a <=( A232  and  (not A202) );
 a6957a <=( A300  and  A299 );
 a6958a <=( A234  and  a6957a );
 a6959a <=( a6958a  and  a6953a );
 a6962a <=( A166  and  A168 );
 a6966a <=( (not A201)  and  A200 );
 a6967a <=( A199  and  a6966a );
 a6968a <=( a6967a  and  a6962a );
 a6971a <=( A232  and  (not A202) );
 a6975a <=( A300  and  A298 );
 a6976a <=( A234  and  a6975a );
 a6977a <=( a6976a  and  a6971a );
 a6980a <=( A166  and  A168 );
 a6984a <=( (not A201)  and  A200 );
 a6985a <=( A199  and  a6984a );
 a6986a <=( a6985a  and  a6980a );
 a6989a <=( A232  and  (not A202) );
 a6993a <=( A267  and  A265 );
 a6994a <=( A234  and  a6993a );
 a6995a <=( a6994a  and  a6989a );
 a6998a <=( A166  and  A168 );
 a7002a <=( (not A201)  and  A200 );
 a7003a <=( A199  and  a7002a );
 a7004a <=( a7003a  and  a6998a );
 a7007a <=( A232  and  (not A202) );
 a7011a <=( A267  and  A266 );
 a7012a <=( A234  and  a7011a );
 a7013a <=( a7012a  and  a7007a );
 a7016a <=( A166  and  A168 );
 a7020a <=( (not A201)  and  A200 );
 a7021a <=( A199  and  a7020a );
 a7022a <=( a7021a  and  a7016a );
 a7025a <=( A233  and  (not A202) );
 a7029a <=( A300  and  A299 );
 a7030a <=( A234  and  a7029a );
 a7031a <=( a7030a  and  a7025a );
 a7034a <=( A166  and  A168 );
 a7038a <=( (not A201)  and  A200 );
 a7039a <=( A199  and  a7038a );
 a7040a <=( a7039a  and  a7034a );
 a7043a <=( A233  and  (not A202) );
 a7047a <=( A300  and  A298 );
 a7048a <=( A234  and  a7047a );
 a7049a <=( a7048a  and  a7043a );
 a7052a <=( A166  and  A168 );
 a7056a <=( (not A201)  and  A200 );
 a7057a <=( A199  and  a7056a );
 a7058a <=( a7057a  and  a7052a );
 a7061a <=( A233  and  (not A202) );
 a7065a <=( A267  and  A265 );
 a7066a <=( A234  and  a7065a );
 a7067a <=( a7066a  and  a7061a );
 a7070a <=( A166  and  A168 );
 a7074a <=( (not A201)  and  A200 );
 a7075a <=( A199  and  a7074a );
 a7076a <=( a7075a  and  a7070a );
 a7079a <=( A233  and  (not A202) );
 a7083a <=( A267  and  A266 );
 a7084a <=( A234  and  a7083a );
 a7085a <=( a7084a  and  a7079a );
 a7088a <=( A166  and  A168 );
 a7092a <=( (not A201)  and  A200 );
 a7093a <=( A199  and  a7092a );
 a7094a <=( a7093a  and  a7088a );
 a7097a <=( (not A232)  and  (not A202) );
 a7101a <=( A301  and  A236 );
 a7102a <=( A233  and  a7101a );
 a7103a <=( a7102a  and  a7097a );
 a7106a <=( A166  and  A168 );
 a7110a <=( (not A201)  and  A200 );
 a7111a <=( A199  and  a7110a );
 a7112a <=( a7111a  and  a7106a );
 a7115a <=( (not A232)  and  (not A202) );
 a7119a <=( A268  and  A236 );
 a7120a <=( A233  and  a7119a );
 a7121a <=( a7120a  and  a7115a );
 a7124a <=( A166  and  A168 );
 a7128a <=( (not A201)  and  A200 );
 a7129a <=( A199  and  a7128a );
 a7130a <=( a7129a  and  a7124a );
 a7133a <=( A232  and  (not A202) );
 a7137a <=( A301  and  A236 );
 a7138a <=( (not A233)  and  a7137a );
 a7139a <=( a7138a  and  a7133a );
 a7142a <=( A166  and  A168 );
 a7146a <=( (not A201)  and  A200 );
 a7147a <=( A199  and  a7146a );
 a7148a <=( a7147a  and  a7142a );
 a7151a <=( A232  and  (not A202) );
 a7155a <=( A268  and  A236 );
 a7156a <=( (not A233)  and  a7155a );
 a7157a <=( a7156a  and  a7151a );
 a7160a <=( A166  and  A168 );
 a7164a <=( (not A202)  and  (not A200) );
 a7165a <=( (not A199)  and  a7164a );
 a7166a <=( a7165a  and  a7160a );
 a7169a <=( A234  and  A232 );
 a7173a <=( A302  and  (not A299) );
 a7174a <=( A298  and  a7173a );
 a7175a <=( a7174a  and  a7169a );
 a7178a <=( A166  and  A168 );
 a7182a <=( (not A202)  and  (not A200) );
 a7183a <=( (not A199)  and  a7182a );
 a7184a <=( a7183a  and  a7178a );
 a7187a <=( A234  and  A232 );
 a7191a <=( A302  and  A299 );
 a7192a <=( (not A298)  and  a7191a );
 a7193a <=( a7192a  and  a7187a );
 a7196a <=( A166  and  A168 );
 a7200a <=( (not A202)  and  (not A200) );
 a7201a <=( (not A199)  and  a7200a );
 a7202a <=( a7201a  and  a7196a );
 a7205a <=( A234  and  A232 );
 a7209a <=( A269  and  A266 );
 a7210a <=( (not A265)  and  a7209a );
 a7211a <=( a7210a  and  a7205a );
 a7214a <=( A166  and  A168 );
 a7218a <=( (not A202)  and  (not A200) );
 a7219a <=( (not A199)  and  a7218a );
 a7220a <=( a7219a  and  a7214a );
 a7223a <=( A234  and  A232 );
 a7227a <=( A269  and  (not A266) );
 a7228a <=( A265  and  a7227a );
 a7229a <=( a7228a  and  a7223a );
 a7232a <=( A166  and  A168 );
 a7236a <=( (not A202)  and  (not A200) );
 a7237a <=( (not A199)  and  a7236a );
 a7238a <=( a7237a  and  a7232a );
 a7241a <=( A234  and  A233 );
 a7245a <=( A302  and  (not A299) );
 a7246a <=( A298  and  a7245a );
 a7247a <=( a7246a  and  a7241a );
 a7250a <=( A166  and  A168 );
 a7254a <=( (not A202)  and  (not A200) );
 a7255a <=( (not A199)  and  a7254a );
 a7256a <=( a7255a  and  a7250a );
 a7259a <=( A234  and  A233 );
 a7263a <=( A302  and  A299 );
 a7264a <=( (not A298)  and  a7263a );
 a7265a <=( a7264a  and  a7259a );
 a7268a <=( A166  and  A168 );
 a7272a <=( (not A202)  and  (not A200) );
 a7273a <=( (not A199)  and  a7272a );
 a7274a <=( a7273a  and  a7268a );
 a7277a <=( A234  and  A233 );
 a7281a <=( A269  and  A266 );
 a7282a <=( (not A265)  and  a7281a );
 a7283a <=( a7282a  and  a7277a );
 a7286a <=( A166  and  A168 );
 a7290a <=( (not A202)  and  (not A200) );
 a7291a <=( (not A199)  and  a7290a );
 a7292a <=( a7291a  and  a7286a );
 a7295a <=( A234  and  A233 );
 a7299a <=( A269  and  (not A266) );
 a7300a <=( A265  and  a7299a );
 a7301a <=( a7300a  and  a7295a );
 a7304a <=( A166  and  A168 );
 a7308a <=( (not A202)  and  (not A200) );
 a7309a <=( (not A199)  and  a7308a );
 a7310a <=( a7309a  and  a7304a );
 a7313a <=( A233  and  (not A232) );
 a7317a <=( A300  and  A299 );
 a7318a <=( A236  and  a7317a );
 a7319a <=( a7318a  and  a7313a );
 a7322a <=( A166  and  A168 );
 a7326a <=( (not A202)  and  (not A200) );
 a7327a <=( (not A199)  and  a7326a );
 a7328a <=( a7327a  and  a7322a );
 a7331a <=( A233  and  (not A232) );
 a7335a <=( A300  and  A298 );
 a7336a <=( A236  and  a7335a );
 a7337a <=( a7336a  and  a7331a );
 a7340a <=( A166  and  A168 );
 a7344a <=( (not A202)  and  (not A200) );
 a7345a <=( (not A199)  and  a7344a );
 a7346a <=( a7345a  and  a7340a );
 a7349a <=( A233  and  (not A232) );
 a7353a <=( A267  and  A265 );
 a7354a <=( A236  and  a7353a );
 a7355a <=( a7354a  and  a7349a );
 a7358a <=( A166  and  A168 );
 a7362a <=( (not A202)  and  (not A200) );
 a7363a <=( (not A199)  and  a7362a );
 a7364a <=( a7363a  and  a7358a );
 a7367a <=( A233  and  (not A232) );
 a7371a <=( A267  and  A266 );
 a7372a <=( A236  and  a7371a );
 a7373a <=( a7372a  and  a7367a );
 a7376a <=( A166  and  A168 );
 a7380a <=( (not A202)  and  (not A200) );
 a7381a <=( (not A199)  and  a7380a );
 a7382a <=( a7381a  and  a7376a );
 a7385a <=( (not A233)  and  A232 );
 a7389a <=( A300  and  A299 );
 a7390a <=( A236  and  a7389a );
 a7391a <=( a7390a  and  a7385a );
 a7394a <=( A166  and  A168 );
 a7398a <=( (not A202)  and  (not A200) );
 a7399a <=( (not A199)  and  a7398a );
 a7400a <=( a7399a  and  a7394a );
 a7403a <=( (not A233)  and  A232 );
 a7407a <=( A300  and  A298 );
 a7408a <=( A236  and  a7407a );
 a7409a <=( a7408a  and  a7403a );
 a7412a <=( A166  and  A168 );
 a7416a <=( (not A202)  and  (not A200) );
 a7417a <=( (not A199)  and  a7416a );
 a7418a <=( a7417a  and  a7412a );
 a7421a <=( (not A233)  and  A232 );
 a7425a <=( A267  and  A265 );
 a7426a <=( A236  and  a7425a );
 a7427a <=( a7426a  and  a7421a );
 a7430a <=( A166  and  A168 );
 a7434a <=( (not A202)  and  (not A200) );
 a7435a <=( (not A199)  and  a7434a );
 a7436a <=( a7435a  and  a7430a );
 a7439a <=( (not A233)  and  A232 );
 a7443a <=( A267  and  A266 );
 a7444a <=( A236  and  a7443a );
 a7445a <=( a7444a  and  a7439a );
 a7448a <=( A167  and  A168 );
 a7452a <=( (not A203)  and  (not A202) );
 a7453a <=( (not A201)  and  a7452a );
 a7454a <=( a7453a  and  a7448a );
 a7457a <=( A234  and  A232 );
 a7461a <=( A302  and  (not A299) );
 a7462a <=( A298  and  a7461a );
 a7463a <=( a7462a  and  a7457a );
 a7466a <=( A167  and  A168 );
 a7470a <=( (not A203)  and  (not A202) );
 a7471a <=( (not A201)  and  a7470a );
 a7472a <=( a7471a  and  a7466a );
 a7475a <=( A234  and  A232 );
 a7479a <=( A302  and  A299 );
 a7480a <=( (not A298)  and  a7479a );
 a7481a <=( a7480a  and  a7475a );
 a7484a <=( A167  and  A168 );
 a7488a <=( (not A203)  and  (not A202) );
 a7489a <=( (not A201)  and  a7488a );
 a7490a <=( a7489a  and  a7484a );
 a7493a <=( A234  and  A232 );
 a7497a <=( A269  and  A266 );
 a7498a <=( (not A265)  and  a7497a );
 a7499a <=( a7498a  and  a7493a );
 a7502a <=( A167  and  A168 );
 a7506a <=( (not A203)  and  (not A202) );
 a7507a <=( (not A201)  and  a7506a );
 a7508a <=( a7507a  and  a7502a );
 a7511a <=( A234  and  A232 );
 a7515a <=( A269  and  (not A266) );
 a7516a <=( A265  and  a7515a );
 a7517a <=( a7516a  and  a7511a );
 a7520a <=( A167  and  A168 );
 a7524a <=( (not A203)  and  (not A202) );
 a7525a <=( (not A201)  and  a7524a );
 a7526a <=( a7525a  and  a7520a );
 a7529a <=( A234  and  A233 );
 a7533a <=( A302  and  (not A299) );
 a7534a <=( A298  and  a7533a );
 a7535a <=( a7534a  and  a7529a );
 a7538a <=( A167  and  A168 );
 a7542a <=( (not A203)  and  (not A202) );
 a7543a <=( (not A201)  and  a7542a );
 a7544a <=( a7543a  and  a7538a );
 a7547a <=( A234  and  A233 );
 a7551a <=( A302  and  A299 );
 a7552a <=( (not A298)  and  a7551a );
 a7553a <=( a7552a  and  a7547a );
 a7556a <=( A167  and  A168 );
 a7560a <=( (not A203)  and  (not A202) );
 a7561a <=( (not A201)  and  a7560a );
 a7562a <=( a7561a  and  a7556a );
 a7565a <=( A234  and  A233 );
 a7569a <=( A269  and  A266 );
 a7570a <=( (not A265)  and  a7569a );
 a7571a <=( a7570a  and  a7565a );
 a7574a <=( A167  and  A168 );
 a7578a <=( (not A203)  and  (not A202) );
 a7579a <=( (not A201)  and  a7578a );
 a7580a <=( a7579a  and  a7574a );
 a7583a <=( A234  and  A233 );
 a7587a <=( A269  and  (not A266) );
 a7588a <=( A265  and  a7587a );
 a7589a <=( a7588a  and  a7583a );
 a7592a <=( A167  and  A168 );
 a7596a <=( (not A203)  and  (not A202) );
 a7597a <=( (not A201)  and  a7596a );
 a7598a <=( a7597a  and  a7592a );
 a7601a <=( A233  and  (not A232) );
 a7605a <=( A300  and  A299 );
 a7606a <=( A236  and  a7605a );
 a7607a <=( a7606a  and  a7601a );
 a7610a <=( A167  and  A168 );
 a7614a <=( (not A203)  and  (not A202) );
 a7615a <=( (not A201)  and  a7614a );
 a7616a <=( a7615a  and  a7610a );
 a7619a <=( A233  and  (not A232) );
 a7623a <=( A300  and  A298 );
 a7624a <=( A236  and  a7623a );
 a7625a <=( a7624a  and  a7619a );
 a7628a <=( A167  and  A168 );
 a7632a <=( (not A203)  and  (not A202) );
 a7633a <=( (not A201)  and  a7632a );
 a7634a <=( a7633a  and  a7628a );
 a7637a <=( A233  and  (not A232) );
 a7641a <=( A267  and  A265 );
 a7642a <=( A236  and  a7641a );
 a7643a <=( a7642a  and  a7637a );
 a7646a <=( A167  and  A168 );
 a7650a <=( (not A203)  and  (not A202) );
 a7651a <=( (not A201)  and  a7650a );
 a7652a <=( a7651a  and  a7646a );
 a7655a <=( A233  and  (not A232) );
 a7659a <=( A267  and  A266 );
 a7660a <=( A236  and  a7659a );
 a7661a <=( a7660a  and  a7655a );
 a7664a <=( A167  and  A168 );
 a7668a <=( (not A203)  and  (not A202) );
 a7669a <=( (not A201)  and  a7668a );
 a7670a <=( a7669a  and  a7664a );
 a7673a <=( (not A233)  and  A232 );
 a7677a <=( A300  and  A299 );
 a7678a <=( A236  and  a7677a );
 a7679a <=( a7678a  and  a7673a );
 a7682a <=( A167  and  A168 );
 a7686a <=( (not A203)  and  (not A202) );
 a7687a <=( (not A201)  and  a7686a );
 a7688a <=( a7687a  and  a7682a );
 a7691a <=( (not A233)  and  A232 );
 a7695a <=( A300  and  A298 );
 a7696a <=( A236  and  a7695a );
 a7697a <=( a7696a  and  a7691a );
 a7700a <=( A167  and  A168 );
 a7704a <=( (not A203)  and  (not A202) );
 a7705a <=( (not A201)  and  a7704a );
 a7706a <=( a7705a  and  a7700a );
 a7709a <=( (not A233)  and  A232 );
 a7713a <=( A267  and  A265 );
 a7714a <=( A236  and  a7713a );
 a7715a <=( a7714a  and  a7709a );
 a7718a <=( A167  and  A168 );
 a7722a <=( (not A203)  and  (not A202) );
 a7723a <=( (not A201)  and  a7722a );
 a7724a <=( a7723a  and  a7718a );
 a7727a <=( (not A233)  and  A232 );
 a7731a <=( A267  and  A266 );
 a7732a <=( A236  and  a7731a );
 a7733a <=( a7732a  and  a7727a );
 a7736a <=( A167  and  A168 );
 a7740a <=( (not A201)  and  A200 );
 a7741a <=( A199  and  a7740a );
 a7742a <=( a7741a  and  a7736a );
 a7745a <=( A235  and  (not A202) );
 a7749a <=( A302  and  (not A299) );
 a7750a <=( A298  and  a7749a );
 a7751a <=( a7750a  and  a7745a );
 a7754a <=( A167  and  A168 );
 a7758a <=( (not A201)  and  A200 );
 a7759a <=( A199  and  a7758a );
 a7760a <=( a7759a  and  a7754a );
 a7763a <=( A235  and  (not A202) );
 a7767a <=( A302  and  A299 );
 a7768a <=( (not A298)  and  a7767a );
 a7769a <=( a7768a  and  a7763a );
 a7772a <=( A167  and  A168 );
 a7776a <=( (not A201)  and  A200 );
 a7777a <=( A199  and  a7776a );
 a7778a <=( a7777a  and  a7772a );
 a7781a <=( A235  and  (not A202) );
 a7785a <=( A269  and  A266 );
 a7786a <=( (not A265)  and  a7785a );
 a7787a <=( a7786a  and  a7781a );
 a7790a <=( A167  and  A168 );
 a7794a <=( (not A201)  and  A200 );
 a7795a <=( A199  and  a7794a );
 a7796a <=( a7795a  and  a7790a );
 a7799a <=( A235  and  (not A202) );
 a7803a <=( A269  and  (not A266) );
 a7804a <=( A265  and  a7803a );
 a7805a <=( a7804a  and  a7799a );
 a7808a <=( A167  and  A168 );
 a7812a <=( (not A201)  and  A200 );
 a7813a <=( A199  and  a7812a );
 a7814a <=( a7813a  and  a7808a );
 a7817a <=( A232  and  (not A202) );
 a7821a <=( A300  and  A299 );
 a7822a <=( A234  and  a7821a );
 a7823a <=( a7822a  and  a7817a );
 a7826a <=( A167  and  A168 );
 a7830a <=( (not A201)  and  A200 );
 a7831a <=( A199  and  a7830a );
 a7832a <=( a7831a  and  a7826a );
 a7835a <=( A232  and  (not A202) );
 a7839a <=( A300  and  A298 );
 a7840a <=( A234  and  a7839a );
 a7841a <=( a7840a  and  a7835a );
 a7844a <=( A167  and  A168 );
 a7848a <=( (not A201)  and  A200 );
 a7849a <=( A199  and  a7848a );
 a7850a <=( a7849a  and  a7844a );
 a7853a <=( A232  and  (not A202) );
 a7857a <=( A267  and  A265 );
 a7858a <=( A234  and  a7857a );
 a7859a <=( a7858a  and  a7853a );
 a7862a <=( A167  and  A168 );
 a7866a <=( (not A201)  and  A200 );
 a7867a <=( A199  and  a7866a );
 a7868a <=( a7867a  and  a7862a );
 a7871a <=( A232  and  (not A202) );
 a7875a <=( A267  and  A266 );
 a7876a <=( A234  and  a7875a );
 a7877a <=( a7876a  and  a7871a );
 a7880a <=( A167  and  A168 );
 a7884a <=( (not A201)  and  A200 );
 a7885a <=( A199  and  a7884a );
 a7886a <=( a7885a  and  a7880a );
 a7889a <=( A233  and  (not A202) );
 a7893a <=( A300  and  A299 );
 a7894a <=( A234  and  a7893a );
 a7895a <=( a7894a  and  a7889a );
 a7898a <=( A167  and  A168 );
 a7902a <=( (not A201)  and  A200 );
 a7903a <=( A199  and  a7902a );
 a7904a <=( a7903a  and  a7898a );
 a7907a <=( A233  and  (not A202) );
 a7911a <=( A300  and  A298 );
 a7912a <=( A234  and  a7911a );
 a7913a <=( a7912a  and  a7907a );
 a7916a <=( A167  and  A168 );
 a7920a <=( (not A201)  and  A200 );
 a7921a <=( A199  and  a7920a );
 a7922a <=( a7921a  and  a7916a );
 a7925a <=( A233  and  (not A202) );
 a7929a <=( A267  and  A265 );
 a7930a <=( A234  and  a7929a );
 a7931a <=( a7930a  and  a7925a );
 a7934a <=( A167  and  A168 );
 a7938a <=( (not A201)  and  A200 );
 a7939a <=( A199  and  a7938a );
 a7940a <=( a7939a  and  a7934a );
 a7943a <=( A233  and  (not A202) );
 a7947a <=( A267  and  A266 );
 a7948a <=( A234  and  a7947a );
 a7949a <=( a7948a  and  a7943a );
 a7952a <=( A167  and  A168 );
 a7956a <=( (not A201)  and  A200 );
 a7957a <=( A199  and  a7956a );
 a7958a <=( a7957a  and  a7952a );
 a7961a <=( (not A232)  and  (not A202) );
 a7965a <=( A301  and  A236 );
 a7966a <=( A233  and  a7965a );
 a7967a <=( a7966a  and  a7961a );
 a7970a <=( A167  and  A168 );
 a7974a <=( (not A201)  and  A200 );
 a7975a <=( A199  and  a7974a );
 a7976a <=( a7975a  and  a7970a );
 a7979a <=( (not A232)  and  (not A202) );
 a7983a <=( A268  and  A236 );
 a7984a <=( A233  and  a7983a );
 a7985a <=( a7984a  and  a7979a );
 a7988a <=( A167  and  A168 );
 a7992a <=( (not A201)  and  A200 );
 a7993a <=( A199  and  a7992a );
 a7994a <=( a7993a  and  a7988a );
 a7997a <=( A232  and  (not A202) );
 a8001a <=( A301  and  A236 );
 a8002a <=( (not A233)  and  a8001a );
 a8003a <=( a8002a  and  a7997a );
 a8006a <=( A167  and  A168 );
 a8010a <=( (not A201)  and  A200 );
 a8011a <=( A199  and  a8010a );
 a8012a <=( a8011a  and  a8006a );
 a8015a <=( A232  and  (not A202) );
 a8019a <=( A268  and  A236 );
 a8020a <=( (not A233)  and  a8019a );
 a8021a <=( a8020a  and  a8015a );
 a8024a <=( A167  and  A168 );
 a8028a <=( (not A202)  and  (not A200) );
 a8029a <=( (not A199)  and  a8028a );
 a8030a <=( a8029a  and  a8024a );
 a8033a <=( A234  and  A232 );
 a8037a <=( A302  and  (not A299) );
 a8038a <=( A298  and  a8037a );
 a8039a <=( a8038a  and  a8033a );
 a8042a <=( A167  and  A168 );
 a8046a <=( (not A202)  and  (not A200) );
 a8047a <=( (not A199)  and  a8046a );
 a8048a <=( a8047a  and  a8042a );
 a8051a <=( A234  and  A232 );
 a8055a <=( A302  and  A299 );
 a8056a <=( (not A298)  and  a8055a );
 a8057a <=( a8056a  and  a8051a );
 a8060a <=( A167  and  A168 );
 a8064a <=( (not A202)  and  (not A200) );
 a8065a <=( (not A199)  and  a8064a );
 a8066a <=( a8065a  and  a8060a );
 a8069a <=( A234  and  A232 );
 a8073a <=( A269  and  A266 );
 a8074a <=( (not A265)  and  a8073a );
 a8075a <=( a8074a  and  a8069a );
 a8078a <=( A167  and  A168 );
 a8082a <=( (not A202)  and  (not A200) );
 a8083a <=( (not A199)  and  a8082a );
 a8084a <=( a8083a  and  a8078a );
 a8087a <=( A234  and  A232 );
 a8091a <=( A269  and  (not A266) );
 a8092a <=( A265  and  a8091a );
 a8093a <=( a8092a  and  a8087a );
 a8096a <=( A167  and  A168 );
 a8100a <=( (not A202)  and  (not A200) );
 a8101a <=( (not A199)  and  a8100a );
 a8102a <=( a8101a  and  a8096a );
 a8105a <=( A234  and  A233 );
 a8109a <=( A302  and  (not A299) );
 a8110a <=( A298  and  a8109a );
 a8111a <=( a8110a  and  a8105a );
 a8114a <=( A167  and  A168 );
 a8118a <=( (not A202)  and  (not A200) );
 a8119a <=( (not A199)  and  a8118a );
 a8120a <=( a8119a  and  a8114a );
 a8123a <=( A234  and  A233 );
 a8127a <=( A302  and  A299 );
 a8128a <=( (not A298)  and  a8127a );
 a8129a <=( a8128a  and  a8123a );
 a8132a <=( A167  and  A168 );
 a8136a <=( (not A202)  and  (not A200) );
 a8137a <=( (not A199)  and  a8136a );
 a8138a <=( a8137a  and  a8132a );
 a8141a <=( A234  and  A233 );
 a8145a <=( A269  and  A266 );
 a8146a <=( (not A265)  and  a8145a );
 a8147a <=( a8146a  and  a8141a );
 a8150a <=( A167  and  A168 );
 a8154a <=( (not A202)  and  (not A200) );
 a8155a <=( (not A199)  and  a8154a );
 a8156a <=( a8155a  and  a8150a );
 a8159a <=( A234  and  A233 );
 a8163a <=( A269  and  (not A266) );
 a8164a <=( A265  and  a8163a );
 a8165a <=( a8164a  and  a8159a );
 a8168a <=( A167  and  A168 );
 a8172a <=( (not A202)  and  (not A200) );
 a8173a <=( (not A199)  and  a8172a );
 a8174a <=( a8173a  and  a8168a );
 a8177a <=( A233  and  (not A232) );
 a8181a <=( A300  and  A299 );
 a8182a <=( A236  and  a8181a );
 a8183a <=( a8182a  and  a8177a );
 a8186a <=( A167  and  A168 );
 a8190a <=( (not A202)  and  (not A200) );
 a8191a <=( (not A199)  and  a8190a );
 a8192a <=( a8191a  and  a8186a );
 a8195a <=( A233  and  (not A232) );
 a8199a <=( A300  and  A298 );
 a8200a <=( A236  and  a8199a );
 a8201a <=( a8200a  and  a8195a );
 a8204a <=( A167  and  A168 );
 a8208a <=( (not A202)  and  (not A200) );
 a8209a <=( (not A199)  and  a8208a );
 a8210a <=( a8209a  and  a8204a );
 a8213a <=( A233  and  (not A232) );
 a8217a <=( A267  and  A265 );
 a8218a <=( A236  and  a8217a );
 a8219a <=( a8218a  and  a8213a );
 a8222a <=( A167  and  A168 );
 a8226a <=( (not A202)  and  (not A200) );
 a8227a <=( (not A199)  and  a8226a );
 a8228a <=( a8227a  and  a8222a );
 a8231a <=( A233  and  (not A232) );
 a8235a <=( A267  and  A266 );
 a8236a <=( A236  and  a8235a );
 a8237a <=( a8236a  and  a8231a );
 a8240a <=( A167  and  A168 );
 a8244a <=( (not A202)  and  (not A200) );
 a8245a <=( (not A199)  and  a8244a );
 a8246a <=( a8245a  and  a8240a );
 a8249a <=( (not A233)  and  A232 );
 a8253a <=( A300  and  A299 );
 a8254a <=( A236  and  a8253a );
 a8255a <=( a8254a  and  a8249a );
 a8258a <=( A167  and  A168 );
 a8262a <=( (not A202)  and  (not A200) );
 a8263a <=( (not A199)  and  a8262a );
 a8264a <=( a8263a  and  a8258a );
 a8267a <=( (not A233)  and  A232 );
 a8271a <=( A300  and  A298 );
 a8272a <=( A236  and  a8271a );
 a8273a <=( a8272a  and  a8267a );
 a8276a <=( A167  and  A168 );
 a8280a <=( (not A202)  and  (not A200) );
 a8281a <=( (not A199)  and  a8280a );
 a8282a <=( a8281a  and  a8276a );
 a8285a <=( (not A233)  and  A232 );
 a8289a <=( A267  and  A265 );
 a8290a <=( A236  and  a8289a );
 a8291a <=( a8290a  and  a8285a );
 a8294a <=( A167  and  A168 );
 a8298a <=( (not A202)  and  (not A200) );
 a8299a <=( (not A199)  and  a8298a );
 a8300a <=( a8299a  and  a8294a );
 a8303a <=( (not A233)  and  A232 );
 a8307a <=( A267  and  A266 );
 a8308a <=( A236  and  a8307a );
 a8309a <=( a8308a  and  a8303a );
 a8312a <=( A167  and  A170 );
 a8316a <=( (not A202)  and  (not A201) );
 a8317a <=( (not A166)  and  a8316a );
 a8318a <=( a8317a  and  a8312a );
 a8321a <=( A235  and  (not A203) );
 a8325a <=( A302  and  (not A299) );
 a8326a <=( A298  and  a8325a );
 a8327a <=( a8326a  and  a8321a );
 a8330a <=( A167  and  A170 );
 a8334a <=( (not A202)  and  (not A201) );
 a8335a <=( (not A166)  and  a8334a );
 a8336a <=( a8335a  and  a8330a );
 a8339a <=( A235  and  (not A203) );
 a8343a <=( A302  and  A299 );
 a8344a <=( (not A298)  and  a8343a );
 a8345a <=( a8344a  and  a8339a );
 a8348a <=( A167  and  A170 );
 a8352a <=( (not A202)  and  (not A201) );
 a8353a <=( (not A166)  and  a8352a );
 a8354a <=( a8353a  and  a8348a );
 a8357a <=( A235  and  (not A203) );
 a8361a <=( A269  and  A266 );
 a8362a <=( (not A265)  and  a8361a );
 a8363a <=( a8362a  and  a8357a );
 a8366a <=( A167  and  A170 );
 a8370a <=( (not A202)  and  (not A201) );
 a8371a <=( (not A166)  and  a8370a );
 a8372a <=( a8371a  and  a8366a );
 a8375a <=( A235  and  (not A203) );
 a8379a <=( A269  and  (not A266) );
 a8380a <=( A265  and  a8379a );
 a8381a <=( a8380a  and  a8375a );
 a8384a <=( A167  and  A170 );
 a8388a <=( (not A202)  and  (not A201) );
 a8389a <=( (not A166)  and  a8388a );
 a8390a <=( a8389a  and  a8384a );
 a8393a <=( A232  and  (not A203) );
 a8397a <=( A300  and  A299 );
 a8398a <=( A234  and  a8397a );
 a8399a <=( a8398a  and  a8393a );
 a8402a <=( A167  and  A170 );
 a8406a <=( (not A202)  and  (not A201) );
 a8407a <=( (not A166)  and  a8406a );
 a8408a <=( a8407a  and  a8402a );
 a8411a <=( A232  and  (not A203) );
 a8415a <=( A300  and  A298 );
 a8416a <=( A234  and  a8415a );
 a8417a <=( a8416a  and  a8411a );
 a8420a <=( A167  and  A170 );
 a8424a <=( (not A202)  and  (not A201) );
 a8425a <=( (not A166)  and  a8424a );
 a8426a <=( a8425a  and  a8420a );
 a8429a <=( A232  and  (not A203) );
 a8433a <=( A267  and  A265 );
 a8434a <=( A234  and  a8433a );
 a8435a <=( a8434a  and  a8429a );
 a8438a <=( A167  and  A170 );
 a8442a <=( (not A202)  and  (not A201) );
 a8443a <=( (not A166)  and  a8442a );
 a8444a <=( a8443a  and  a8438a );
 a8447a <=( A232  and  (not A203) );
 a8451a <=( A267  and  A266 );
 a8452a <=( A234  and  a8451a );
 a8453a <=( a8452a  and  a8447a );
 a8456a <=( A167  and  A170 );
 a8460a <=( (not A202)  and  (not A201) );
 a8461a <=( (not A166)  and  a8460a );
 a8462a <=( a8461a  and  a8456a );
 a8465a <=( A233  and  (not A203) );
 a8469a <=( A300  and  A299 );
 a8470a <=( A234  and  a8469a );
 a8471a <=( a8470a  and  a8465a );
 a8474a <=( A167  and  A170 );
 a8478a <=( (not A202)  and  (not A201) );
 a8479a <=( (not A166)  and  a8478a );
 a8480a <=( a8479a  and  a8474a );
 a8483a <=( A233  and  (not A203) );
 a8487a <=( A300  and  A298 );
 a8488a <=( A234  and  a8487a );
 a8489a <=( a8488a  and  a8483a );
 a8492a <=( A167  and  A170 );
 a8496a <=( (not A202)  and  (not A201) );
 a8497a <=( (not A166)  and  a8496a );
 a8498a <=( a8497a  and  a8492a );
 a8501a <=( A233  and  (not A203) );
 a8505a <=( A267  and  A265 );
 a8506a <=( A234  and  a8505a );
 a8507a <=( a8506a  and  a8501a );
 a8510a <=( A167  and  A170 );
 a8514a <=( (not A202)  and  (not A201) );
 a8515a <=( (not A166)  and  a8514a );
 a8516a <=( a8515a  and  a8510a );
 a8519a <=( A233  and  (not A203) );
 a8523a <=( A267  and  A266 );
 a8524a <=( A234  and  a8523a );
 a8525a <=( a8524a  and  a8519a );
 a8528a <=( A167  and  A170 );
 a8532a <=( (not A202)  and  (not A201) );
 a8533a <=( (not A166)  and  a8532a );
 a8534a <=( a8533a  and  a8528a );
 a8537a <=( (not A232)  and  (not A203) );
 a8541a <=( A301  and  A236 );
 a8542a <=( A233  and  a8541a );
 a8543a <=( a8542a  and  a8537a );
 a8546a <=( A167  and  A170 );
 a8550a <=( (not A202)  and  (not A201) );
 a8551a <=( (not A166)  and  a8550a );
 a8552a <=( a8551a  and  a8546a );
 a8555a <=( (not A232)  and  (not A203) );
 a8559a <=( A268  and  A236 );
 a8560a <=( A233  and  a8559a );
 a8561a <=( a8560a  and  a8555a );
 a8564a <=( A167  and  A170 );
 a8568a <=( (not A202)  and  (not A201) );
 a8569a <=( (not A166)  and  a8568a );
 a8570a <=( a8569a  and  a8564a );
 a8573a <=( A232  and  (not A203) );
 a8577a <=( A301  and  A236 );
 a8578a <=( (not A233)  and  a8577a );
 a8579a <=( a8578a  and  a8573a );
 a8582a <=( A167  and  A170 );
 a8586a <=( (not A202)  and  (not A201) );
 a8587a <=( (not A166)  and  a8586a );
 a8588a <=( a8587a  and  a8582a );
 a8591a <=( A232  and  (not A203) );
 a8595a <=( A268  and  A236 );
 a8596a <=( (not A233)  and  a8595a );
 a8597a <=( a8596a  and  a8591a );
 a8600a <=( A167  and  A170 );
 a8604a <=( A200  and  A199 );
 a8605a <=( (not A166)  and  a8604a );
 a8606a <=( a8605a  and  a8600a );
 a8609a <=( (not A202)  and  (not A201) );
 a8613a <=( A300  and  A299 );
 a8614a <=( A235  and  a8613a );
 a8615a <=( a8614a  and  a8609a );
 a8618a <=( A167  and  A170 );
 a8622a <=( A200  and  A199 );
 a8623a <=( (not A166)  and  a8622a );
 a8624a <=( a8623a  and  a8618a );
 a8627a <=( (not A202)  and  (not A201) );
 a8631a <=( A300  and  A298 );
 a8632a <=( A235  and  a8631a );
 a8633a <=( a8632a  and  a8627a );
 a8636a <=( A167  and  A170 );
 a8640a <=( A200  and  A199 );
 a8641a <=( (not A166)  and  a8640a );
 a8642a <=( a8641a  and  a8636a );
 a8645a <=( (not A202)  and  (not A201) );
 a8649a <=( A267  and  A265 );
 a8650a <=( A235  and  a8649a );
 a8651a <=( a8650a  and  a8645a );
 a8654a <=( A167  and  A170 );
 a8658a <=( A200  and  A199 );
 a8659a <=( (not A166)  and  a8658a );
 a8660a <=( a8659a  and  a8654a );
 a8663a <=( (not A202)  and  (not A201) );
 a8667a <=( A267  and  A266 );
 a8668a <=( A235  and  a8667a );
 a8669a <=( a8668a  and  a8663a );
 a8672a <=( A167  and  A170 );
 a8676a <=( A200  and  A199 );
 a8677a <=( (not A166)  and  a8676a );
 a8678a <=( a8677a  and  a8672a );
 a8681a <=( (not A202)  and  (not A201) );
 a8685a <=( A301  and  A234 );
 a8686a <=( A232  and  a8685a );
 a8687a <=( a8686a  and  a8681a );
 a8690a <=( A167  and  A170 );
 a8694a <=( A200  and  A199 );
 a8695a <=( (not A166)  and  a8694a );
 a8696a <=( a8695a  and  a8690a );
 a8699a <=( (not A202)  and  (not A201) );
 a8703a <=( A268  and  A234 );
 a8704a <=( A232  and  a8703a );
 a8705a <=( a8704a  and  a8699a );
 a8708a <=( A167  and  A170 );
 a8712a <=( A200  and  A199 );
 a8713a <=( (not A166)  and  a8712a );
 a8714a <=( a8713a  and  a8708a );
 a8717a <=( (not A202)  and  (not A201) );
 a8721a <=( A301  and  A234 );
 a8722a <=( A233  and  a8721a );
 a8723a <=( a8722a  and  a8717a );
 a8726a <=( A167  and  A170 );
 a8730a <=( A200  and  A199 );
 a8731a <=( (not A166)  and  a8730a );
 a8732a <=( a8731a  and  a8726a );
 a8735a <=( (not A202)  and  (not A201) );
 a8739a <=( A268  and  A234 );
 a8740a <=( A233  and  a8739a );
 a8741a <=( a8740a  and  a8735a );
 a8744a <=( A167  and  A170 );
 a8748a <=( (not A200)  and  (not A199) );
 a8749a <=( (not A166)  and  a8748a );
 a8750a <=( a8749a  and  a8744a );
 a8753a <=( A235  and  (not A202) );
 a8757a <=( A302  and  (not A299) );
 a8758a <=( A298  and  a8757a );
 a8759a <=( a8758a  and  a8753a );
 a8762a <=( A167  and  A170 );
 a8766a <=( (not A200)  and  (not A199) );
 a8767a <=( (not A166)  and  a8766a );
 a8768a <=( a8767a  and  a8762a );
 a8771a <=( A235  and  (not A202) );
 a8775a <=( A302  and  A299 );
 a8776a <=( (not A298)  and  a8775a );
 a8777a <=( a8776a  and  a8771a );
 a8780a <=( A167  and  A170 );
 a8784a <=( (not A200)  and  (not A199) );
 a8785a <=( (not A166)  and  a8784a );
 a8786a <=( a8785a  and  a8780a );
 a8789a <=( A235  and  (not A202) );
 a8793a <=( A269  and  A266 );
 a8794a <=( (not A265)  and  a8793a );
 a8795a <=( a8794a  and  a8789a );
 a8798a <=( A167  and  A170 );
 a8802a <=( (not A200)  and  (not A199) );
 a8803a <=( (not A166)  and  a8802a );
 a8804a <=( a8803a  and  a8798a );
 a8807a <=( A235  and  (not A202) );
 a8811a <=( A269  and  (not A266) );
 a8812a <=( A265  and  a8811a );
 a8813a <=( a8812a  and  a8807a );
 a8816a <=( A167  and  A170 );
 a8820a <=( (not A200)  and  (not A199) );
 a8821a <=( (not A166)  and  a8820a );
 a8822a <=( a8821a  and  a8816a );
 a8825a <=( A232  and  (not A202) );
 a8829a <=( A300  and  A299 );
 a8830a <=( A234  and  a8829a );
 a8831a <=( a8830a  and  a8825a );
 a8834a <=( A167  and  A170 );
 a8838a <=( (not A200)  and  (not A199) );
 a8839a <=( (not A166)  and  a8838a );
 a8840a <=( a8839a  and  a8834a );
 a8843a <=( A232  and  (not A202) );
 a8847a <=( A300  and  A298 );
 a8848a <=( A234  and  a8847a );
 a8849a <=( a8848a  and  a8843a );
 a8852a <=( A167  and  A170 );
 a8856a <=( (not A200)  and  (not A199) );
 a8857a <=( (not A166)  and  a8856a );
 a8858a <=( a8857a  and  a8852a );
 a8861a <=( A232  and  (not A202) );
 a8865a <=( A267  and  A265 );
 a8866a <=( A234  and  a8865a );
 a8867a <=( a8866a  and  a8861a );
 a8870a <=( A167  and  A170 );
 a8874a <=( (not A200)  and  (not A199) );
 a8875a <=( (not A166)  and  a8874a );
 a8876a <=( a8875a  and  a8870a );
 a8879a <=( A232  and  (not A202) );
 a8883a <=( A267  and  A266 );
 a8884a <=( A234  and  a8883a );
 a8885a <=( a8884a  and  a8879a );
 a8888a <=( A167  and  A170 );
 a8892a <=( (not A200)  and  (not A199) );
 a8893a <=( (not A166)  and  a8892a );
 a8894a <=( a8893a  and  a8888a );
 a8897a <=( A233  and  (not A202) );
 a8901a <=( A300  and  A299 );
 a8902a <=( A234  and  a8901a );
 a8903a <=( a8902a  and  a8897a );
 a8906a <=( A167  and  A170 );
 a8910a <=( (not A200)  and  (not A199) );
 a8911a <=( (not A166)  and  a8910a );
 a8912a <=( a8911a  and  a8906a );
 a8915a <=( A233  and  (not A202) );
 a8919a <=( A300  and  A298 );
 a8920a <=( A234  and  a8919a );
 a8921a <=( a8920a  and  a8915a );
 a8924a <=( A167  and  A170 );
 a8928a <=( (not A200)  and  (not A199) );
 a8929a <=( (not A166)  and  a8928a );
 a8930a <=( a8929a  and  a8924a );
 a8933a <=( A233  and  (not A202) );
 a8937a <=( A267  and  A265 );
 a8938a <=( A234  and  a8937a );
 a8939a <=( a8938a  and  a8933a );
 a8942a <=( A167  and  A170 );
 a8946a <=( (not A200)  and  (not A199) );
 a8947a <=( (not A166)  and  a8946a );
 a8948a <=( a8947a  and  a8942a );
 a8951a <=( A233  and  (not A202) );
 a8955a <=( A267  and  A266 );
 a8956a <=( A234  and  a8955a );
 a8957a <=( a8956a  and  a8951a );
 a8960a <=( A167  and  A170 );
 a8964a <=( (not A200)  and  (not A199) );
 a8965a <=( (not A166)  and  a8964a );
 a8966a <=( a8965a  and  a8960a );
 a8969a <=( (not A232)  and  (not A202) );
 a8973a <=( A301  and  A236 );
 a8974a <=( A233  and  a8973a );
 a8975a <=( a8974a  and  a8969a );
 a8978a <=( A167  and  A170 );
 a8982a <=( (not A200)  and  (not A199) );
 a8983a <=( (not A166)  and  a8982a );
 a8984a <=( a8983a  and  a8978a );
 a8987a <=( (not A232)  and  (not A202) );
 a8991a <=( A268  and  A236 );
 a8992a <=( A233  and  a8991a );
 a8993a <=( a8992a  and  a8987a );
 a8996a <=( A167  and  A170 );
 a9000a <=( (not A200)  and  (not A199) );
 a9001a <=( (not A166)  and  a9000a );
 a9002a <=( a9001a  and  a8996a );
 a9005a <=( A232  and  (not A202) );
 a9009a <=( A301  and  A236 );
 a9010a <=( (not A233)  and  a9009a );
 a9011a <=( a9010a  and  a9005a );
 a9014a <=( A167  and  A170 );
 a9018a <=( (not A200)  and  (not A199) );
 a9019a <=( (not A166)  and  a9018a );
 a9020a <=( a9019a  and  a9014a );
 a9023a <=( A232  and  (not A202) );
 a9027a <=( A268  and  A236 );
 a9028a <=( (not A233)  and  a9027a );
 a9029a <=( a9028a  and  a9023a );
 a9032a <=( (not A167)  and  A170 );
 a9036a <=( (not A202)  and  (not A201) );
 a9037a <=( A166  and  a9036a );
 a9038a <=( a9037a  and  a9032a );
 a9041a <=( A235  and  (not A203) );
 a9045a <=( A302  and  (not A299) );
 a9046a <=( A298  and  a9045a );
 a9047a <=( a9046a  and  a9041a );
 a9050a <=( (not A167)  and  A170 );
 a9054a <=( (not A202)  and  (not A201) );
 a9055a <=( A166  and  a9054a );
 a9056a <=( a9055a  and  a9050a );
 a9059a <=( A235  and  (not A203) );
 a9063a <=( A302  and  A299 );
 a9064a <=( (not A298)  and  a9063a );
 a9065a <=( a9064a  and  a9059a );
 a9068a <=( (not A167)  and  A170 );
 a9072a <=( (not A202)  and  (not A201) );
 a9073a <=( A166  and  a9072a );
 a9074a <=( a9073a  and  a9068a );
 a9077a <=( A235  and  (not A203) );
 a9081a <=( A269  and  A266 );
 a9082a <=( (not A265)  and  a9081a );
 a9083a <=( a9082a  and  a9077a );
 a9086a <=( (not A167)  and  A170 );
 a9090a <=( (not A202)  and  (not A201) );
 a9091a <=( A166  and  a9090a );
 a9092a <=( a9091a  and  a9086a );
 a9095a <=( A235  and  (not A203) );
 a9099a <=( A269  and  (not A266) );
 a9100a <=( A265  and  a9099a );
 a9101a <=( a9100a  and  a9095a );
 a9104a <=( (not A167)  and  A170 );
 a9108a <=( (not A202)  and  (not A201) );
 a9109a <=( A166  and  a9108a );
 a9110a <=( a9109a  and  a9104a );
 a9113a <=( A232  and  (not A203) );
 a9117a <=( A300  and  A299 );
 a9118a <=( A234  and  a9117a );
 a9119a <=( a9118a  and  a9113a );
 a9122a <=( (not A167)  and  A170 );
 a9126a <=( (not A202)  and  (not A201) );
 a9127a <=( A166  and  a9126a );
 a9128a <=( a9127a  and  a9122a );
 a9131a <=( A232  and  (not A203) );
 a9135a <=( A300  and  A298 );
 a9136a <=( A234  and  a9135a );
 a9137a <=( a9136a  and  a9131a );
 a9140a <=( (not A167)  and  A170 );
 a9144a <=( (not A202)  and  (not A201) );
 a9145a <=( A166  and  a9144a );
 a9146a <=( a9145a  and  a9140a );
 a9149a <=( A232  and  (not A203) );
 a9153a <=( A267  and  A265 );
 a9154a <=( A234  and  a9153a );
 a9155a <=( a9154a  and  a9149a );
 a9158a <=( (not A167)  and  A170 );
 a9162a <=( (not A202)  and  (not A201) );
 a9163a <=( A166  and  a9162a );
 a9164a <=( a9163a  and  a9158a );
 a9167a <=( A232  and  (not A203) );
 a9171a <=( A267  and  A266 );
 a9172a <=( A234  and  a9171a );
 a9173a <=( a9172a  and  a9167a );
 a9176a <=( (not A167)  and  A170 );
 a9180a <=( (not A202)  and  (not A201) );
 a9181a <=( A166  and  a9180a );
 a9182a <=( a9181a  and  a9176a );
 a9185a <=( A233  and  (not A203) );
 a9189a <=( A300  and  A299 );
 a9190a <=( A234  and  a9189a );
 a9191a <=( a9190a  and  a9185a );
 a9194a <=( (not A167)  and  A170 );
 a9198a <=( (not A202)  and  (not A201) );
 a9199a <=( A166  and  a9198a );
 a9200a <=( a9199a  and  a9194a );
 a9203a <=( A233  and  (not A203) );
 a9207a <=( A300  and  A298 );
 a9208a <=( A234  and  a9207a );
 a9209a <=( a9208a  and  a9203a );
 a9212a <=( (not A167)  and  A170 );
 a9216a <=( (not A202)  and  (not A201) );
 a9217a <=( A166  and  a9216a );
 a9218a <=( a9217a  and  a9212a );
 a9221a <=( A233  and  (not A203) );
 a9225a <=( A267  and  A265 );
 a9226a <=( A234  and  a9225a );
 a9227a <=( a9226a  and  a9221a );
 a9230a <=( (not A167)  and  A170 );
 a9234a <=( (not A202)  and  (not A201) );
 a9235a <=( A166  and  a9234a );
 a9236a <=( a9235a  and  a9230a );
 a9239a <=( A233  and  (not A203) );
 a9243a <=( A267  and  A266 );
 a9244a <=( A234  and  a9243a );
 a9245a <=( a9244a  and  a9239a );
 a9248a <=( (not A167)  and  A170 );
 a9252a <=( (not A202)  and  (not A201) );
 a9253a <=( A166  and  a9252a );
 a9254a <=( a9253a  and  a9248a );
 a9257a <=( (not A232)  and  (not A203) );
 a9261a <=( A301  and  A236 );
 a9262a <=( A233  and  a9261a );
 a9263a <=( a9262a  and  a9257a );
 a9266a <=( (not A167)  and  A170 );
 a9270a <=( (not A202)  and  (not A201) );
 a9271a <=( A166  and  a9270a );
 a9272a <=( a9271a  and  a9266a );
 a9275a <=( (not A232)  and  (not A203) );
 a9279a <=( A268  and  A236 );
 a9280a <=( A233  and  a9279a );
 a9281a <=( a9280a  and  a9275a );
 a9284a <=( (not A167)  and  A170 );
 a9288a <=( (not A202)  and  (not A201) );
 a9289a <=( A166  and  a9288a );
 a9290a <=( a9289a  and  a9284a );
 a9293a <=( A232  and  (not A203) );
 a9297a <=( A301  and  A236 );
 a9298a <=( (not A233)  and  a9297a );
 a9299a <=( a9298a  and  a9293a );
 a9302a <=( (not A167)  and  A170 );
 a9306a <=( (not A202)  and  (not A201) );
 a9307a <=( A166  and  a9306a );
 a9308a <=( a9307a  and  a9302a );
 a9311a <=( A232  and  (not A203) );
 a9315a <=( A268  and  A236 );
 a9316a <=( (not A233)  and  a9315a );
 a9317a <=( a9316a  and  a9311a );
 a9320a <=( (not A167)  and  A170 );
 a9324a <=( A200  and  A199 );
 a9325a <=( A166  and  a9324a );
 a9326a <=( a9325a  and  a9320a );
 a9329a <=( (not A202)  and  (not A201) );
 a9333a <=( A300  and  A299 );
 a9334a <=( A235  and  a9333a );
 a9335a <=( a9334a  and  a9329a );
 a9338a <=( (not A167)  and  A170 );
 a9342a <=( A200  and  A199 );
 a9343a <=( A166  and  a9342a );
 a9344a <=( a9343a  and  a9338a );
 a9347a <=( (not A202)  and  (not A201) );
 a9351a <=( A300  and  A298 );
 a9352a <=( A235  and  a9351a );
 a9353a <=( a9352a  and  a9347a );
 a9356a <=( (not A167)  and  A170 );
 a9360a <=( A200  and  A199 );
 a9361a <=( A166  and  a9360a );
 a9362a <=( a9361a  and  a9356a );
 a9365a <=( (not A202)  and  (not A201) );
 a9369a <=( A267  and  A265 );
 a9370a <=( A235  and  a9369a );
 a9371a <=( a9370a  and  a9365a );
 a9374a <=( (not A167)  and  A170 );
 a9378a <=( A200  and  A199 );
 a9379a <=( A166  and  a9378a );
 a9380a <=( a9379a  and  a9374a );
 a9383a <=( (not A202)  and  (not A201) );
 a9387a <=( A267  and  A266 );
 a9388a <=( A235  and  a9387a );
 a9389a <=( a9388a  and  a9383a );
 a9392a <=( (not A167)  and  A170 );
 a9396a <=( A200  and  A199 );
 a9397a <=( A166  and  a9396a );
 a9398a <=( a9397a  and  a9392a );
 a9401a <=( (not A202)  and  (not A201) );
 a9405a <=( A301  and  A234 );
 a9406a <=( A232  and  a9405a );
 a9407a <=( a9406a  and  a9401a );
 a9410a <=( (not A167)  and  A170 );
 a9414a <=( A200  and  A199 );
 a9415a <=( A166  and  a9414a );
 a9416a <=( a9415a  and  a9410a );
 a9419a <=( (not A202)  and  (not A201) );
 a9423a <=( A268  and  A234 );
 a9424a <=( A232  and  a9423a );
 a9425a <=( a9424a  and  a9419a );
 a9428a <=( (not A167)  and  A170 );
 a9432a <=( A200  and  A199 );
 a9433a <=( A166  and  a9432a );
 a9434a <=( a9433a  and  a9428a );
 a9437a <=( (not A202)  and  (not A201) );
 a9441a <=( A301  and  A234 );
 a9442a <=( A233  and  a9441a );
 a9443a <=( a9442a  and  a9437a );
 a9446a <=( (not A167)  and  A170 );
 a9450a <=( A200  and  A199 );
 a9451a <=( A166  and  a9450a );
 a9452a <=( a9451a  and  a9446a );
 a9455a <=( (not A202)  and  (not A201) );
 a9459a <=( A268  and  A234 );
 a9460a <=( A233  and  a9459a );
 a9461a <=( a9460a  and  a9455a );
 a9464a <=( (not A167)  and  A170 );
 a9468a <=( (not A200)  and  (not A199) );
 a9469a <=( A166  and  a9468a );
 a9470a <=( a9469a  and  a9464a );
 a9473a <=( A235  and  (not A202) );
 a9477a <=( A302  and  (not A299) );
 a9478a <=( A298  and  a9477a );
 a9479a <=( a9478a  and  a9473a );
 a9482a <=( (not A167)  and  A170 );
 a9486a <=( (not A200)  and  (not A199) );
 a9487a <=( A166  and  a9486a );
 a9488a <=( a9487a  and  a9482a );
 a9491a <=( A235  and  (not A202) );
 a9495a <=( A302  and  A299 );
 a9496a <=( (not A298)  and  a9495a );
 a9497a <=( a9496a  and  a9491a );
 a9500a <=( (not A167)  and  A170 );
 a9504a <=( (not A200)  and  (not A199) );
 a9505a <=( A166  and  a9504a );
 a9506a <=( a9505a  and  a9500a );
 a9509a <=( A235  and  (not A202) );
 a9513a <=( A269  and  A266 );
 a9514a <=( (not A265)  and  a9513a );
 a9515a <=( a9514a  and  a9509a );
 a9518a <=( (not A167)  and  A170 );
 a9522a <=( (not A200)  and  (not A199) );
 a9523a <=( A166  and  a9522a );
 a9524a <=( a9523a  and  a9518a );
 a9527a <=( A235  and  (not A202) );
 a9531a <=( A269  and  (not A266) );
 a9532a <=( A265  and  a9531a );
 a9533a <=( a9532a  and  a9527a );
 a9536a <=( (not A167)  and  A170 );
 a9540a <=( (not A200)  and  (not A199) );
 a9541a <=( A166  and  a9540a );
 a9542a <=( a9541a  and  a9536a );
 a9545a <=( A232  and  (not A202) );
 a9549a <=( A300  and  A299 );
 a9550a <=( A234  and  a9549a );
 a9551a <=( a9550a  and  a9545a );
 a9554a <=( (not A167)  and  A170 );
 a9558a <=( (not A200)  and  (not A199) );
 a9559a <=( A166  and  a9558a );
 a9560a <=( a9559a  and  a9554a );
 a9563a <=( A232  and  (not A202) );
 a9567a <=( A300  and  A298 );
 a9568a <=( A234  and  a9567a );
 a9569a <=( a9568a  and  a9563a );
 a9572a <=( (not A167)  and  A170 );
 a9576a <=( (not A200)  and  (not A199) );
 a9577a <=( A166  and  a9576a );
 a9578a <=( a9577a  and  a9572a );
 a9581a <=( A232  and  (not A202) );
 a9585a <=( A267  and  A265 );
 a9586a <=( A234  and  a9585a );
 a9587a <=( a9586a  and  a9581a );
 a9590a <=( (not A167)  and  A170 );
 a9594a <=( (not A200)  and  (not A199) );
 a9595a <=( A166  and  a9594a );
 a9596a <=( a9595a  and  a9590a );
 a9599a <=( A232  and  (not A202) );
 a9603a <=( A267  and  A266 );
 a9604a <=( A234  and  a9603a );
 a9605a <=( a9604a  and  a9599a );
 a9608a <=( (not A167)  and  A170 );
 a9612a <=( (not A200)  and  (not A199) );
 a9613a <=( A166  and  a9612a );
 a9614a <=( a9613a  and  a9608a );
 a9617a <=( A233  and  (not A202) );
 a9621a <=( A300  and  A299 );
 a9622a <=( A234  and  a9621a );
 a9623a <=( a9622a  and  a9617a );
 a9626a <=( (not A167)  and  A170 );
 a9630a <=( (not A200)  and  (not A199) );
 a9631a <=( A166  and  a9630a );
 a9632a <=( a9631a  and  a9626a );
 a9635a <=( A233  and  (not A202) );
 a9639a <=( A300  and  A298 );
 a9640a <=( A234  and  a9639a );
 a9641a <=( a9640a  and  a9635a );
 a9644a <=( (not A167)  and  A170 );
 a9648a <=( (not A200)  and  (not A199) );
 a9649a <=( A166  and  a9648a );
 a9650a <=( a9649a  and  a9644a );
 a9653a <=( A233  and  (not A202) );
 a9657a <=( A267  and  A265 );
 a9658a <=( A234  and  a9657a );
 a9659a <=( a9658a  and  a9653a );
 a9662a <=( (not A167)  and  A170 );
 a9666a <=( (not A200)  and  (not A199) );
 a9667a <=( A166  and  a9666a );
 a9668a <=( a9667a  and  a9662a );
 a9671a <=( A233  and  (not A202) );
 a9675a <=( A267  and  A266 );
 a9676a <=( A234  and  a9675a );
 a9677a <=( a9676a  and  a9671a );
 a9680a <=( (not A167)  and  A170 );
 a9684a <=( (not A200)  and  (not A199) );
 a9685a <=( A166  and  a9684a );
 a9686a <=( a9685a  and  a9680a );
 a9689a <=( (not A232)  and  (not A202) );
 a9693a <=( A301  and  A236 );
 a9694a <=( A233  and  a9693a );
 a9695a <=( a9694a  and  a9689a );
 a9698a <=( (not A167)  and  A170 );
 a9702a <=( (not A200)  and  (not A199) );
 a9703a <=( A166  and  a9702a );
 a9704a <=( a9703a  and  a9698a );
 a9707a <=( (not A232)  and  (not A202) );
 a9711a <=( A268  and  A236 );
 a9712a <=( A233  and  a9711a );
 a9713a <=( a9712a  and  a9707a );
 a9716a <=( (not A167)  and  A170 );
 a9720a <=( (not A200)  and  (not A199) );
 a9721a <=( A166  and  a9720a );
 a9722a <=( a9721a  and  a9716a );
 a9725a <=( A232  and  (not A202) );
 a9729a <=( A301  and  A236 );
 a9730a <=( (not A233)  and  a9729a );
 a9731a <=( a9730a  and  a9725a );
 a9734a <=( (not A167)  and  A170 );
 a9738a <=( (not A200)  and  (not A199) );
 a9739a <=( A166  and  a9738a );
 a9740a <=( a9739a  and  a9734a );
 a9743a <=( A232  and  (not A202) );
 a9747a <=( A268  and  A236 );
 a9748a <=( (not A233)  and  a9747a );
 a9749a <=( a9748a  and  a9743a );
 a9752a <=( (not A201)  and  A169 );
 a9756a <=( (not A232)  and  (not A203) );
 a9757a <=( (not A202)  and  a9756a );
 a9758a <=( a9757a  and  a9752a );
 a9761a <=( A236  and  A233 );
 a9765a <=( A302  and  (not A299) );
 a9766a <=( A298  and  a9765a );
 a9767a <=( a9766a  and  a9761a );
 a9770a <=( (not A201)  and  A169 );
 a9774a <=( (not A232)  and  (not A203) );
 a9775a <=( (not A202)  and  a9774a );
 a9776a <=( a9775a  and  a9770a );
 a9779a <=( A236  and  A233 );
 a9783a <=( A302  and  A299 );
 a9784a <=( (not A298)  and  a9783a );
 a9785a <=( a9784a  and  a9779a );
 a9788a <=( (not A201)  and  A169 );
 a9792a <=( (not A232)  and  (not A203) );
 a9793a <=( (not A202)  and  a9792a );
 a9794a <=( a9793a  and  a9788a );
 a9797a <=( A236  and  A233 );
 a9801a <=( A269  and  A266 );
 a9802a <=( (not A265)  and  a9801a );
 a9803a <=( a9802a  and  a9797a );
 a9806a <=( (not A201)  and  A169 );
 a9810a <=( (not A232)  and  (not A203) );
 a9811a <=( (not A202)  and  a9810a );
 a9812a <=( a9811a  and  a9806a );
 a9815a <=( A236  and  A233 );
 a9819a <=( A269  and  (not A266) );
 a9820a <=( A265  and  a9819a );
 a9821a <=( a9820a  and  a9815a );
 a9824a <=( (not A201)  and  A169 );
 a9828a <=( A232  and  (not A203) );
 a9829a <=( (not A202)  and  a9828a );
 a9830a <=( a9829a  and  a9824a );
 a9833a <=( A236  and  (not A233) );
 a9837a <=( A302  and  (not A299) );
 a9838a <=( A298  and  a9837a );
 a9839a <=( a9838a  and  a9833a );
 a9842a <=( (not A201)  and  A169 );
 a9846a <=( A232  and  (not A203) );
 a9847a <=( (not A202)  and  a9846a );
 a9848a <=( a9847a  and  a9842a );
 a9851a <=( A236  and  (not A233) );
 a9855a <=( A302  and  A299 );
 a9856a <=( (not A298)  and  a9855a );
 a9857a <=( a9856a  and  a9851a );
 a9860a <=( (not A201)  and  A169 );
 a9864a <=( A232  and  (not A203) );
 a9865a <=( (not A202)  and  a9864a );
 a9866a <=( a9865a  and  a9860a );
 a9869a <=( A236  and  (not A233) );
 a9873a <=( A269  and  A266 );
 a9874a <=( (not A265)  and  a9873a );
 a9875a <=( a9874a  and  a9869a );
 a9878a <=( (not A201)  and  A169 );
 a9882a <=( A232  and  (not A203) );
 a9883a <=( (not A202)  and  a9882a );
 a9884a <=( a9883a  and  a9878a );
 a9887a <=( A236  and  (not A233) );
 a9891a <=( A269  and  (not A266) );
 a9892a <=( A265  and  a9891a );
 a9893a <=( a9892a  and  a9887a );
 a9896a <=( A199  and  A169 );
 a9900a <=( (not A202)  and  (not A201) );
 a9901a <=( A200  and  a9900a );
 a9902a <=( a9901a  and  a9896a );
 a9905a <=( A234  and  A232 );
 a9909a <=( A302  and  (not A299) );
 a9910a <=( A298  and  a9909a );
 a9911a <=( a9910a  and  a9905a );
 a9914a <=( A199  and  A169 );
 a9918a <=( (not A202)  and  (not A201) );
 a9919a <=( A200  and  a9918a );
 a9920a <=( a9919a  and  a9914a );
 a9923a <=( A234  and  A232 );
 a9927a <=( A302  and  A299 );
 a9928a <=( (not A298)  and  a9927a );
 a9929a <=( a9928a  and  a9923a );
 a9932a <=( A199  and  A169 );
 a9936a <=( (not A202)  and  (not A201) );
 a9937a <=( A200  and  a9936a );
 a9938a <=( a9937a  and  a9932a );
 a9941a <=( A234  and  A232 );
 a9945a <=( A269  and  A266 );
 a9946a <=( (not A265)  and  a9945a );
 a9947a <=( a9946a  and  a9941a );
 a9950a <=( A199  and  A169 );
 a9954a <=( (not A202)  and  (not A201) );
 a9955a <=( A200  and  a9954a );
 a9956a <=( a9955a  and  a9950a );
 a9959a <=( A234  and  A232 );
 a9963a <=( A269  and  (not A266) );
 a9964a <=( A265  and  a9963a );
 a9965a <=( a9964a  and  a9959a );
 a9968a <=( A199  and  A169 );
 a9972a <=( (not A202)  and  (not A201) );
 a9973a <=( A200  and  a9972a );
 a9974a <=( a9973a  and  a9968a );
 a9977a <=( A234  and  A233 );
 a9981a <=( A302  and  (not A299) );
 a9982a <=( A298  and  a9981a );
 a9983a <=( a9982a  and  a9977a );
 a9986a <=( A199  and  A169 );
 a9990a <=( (not A202)  and  (not A201) );
 a9991a <=( A200  and  a9990a );
 a9992a <=( a9991a  and  a9986a );
 a9995a <=( A234  and  A233 );
 a9999a <=( A302  and  A299 );
 a10000a <=( (not A298)  and  a9999a );
 a10001a <=( a10000a  and  a9995a );
 a10004a <=( A199  and  A169 );
 a10008a <=( (not A202)  and  (not A201) );
 a10009a <=( A200  and  a10008a );
 a10010a <=( a10009a  and  a10004a );
 a10013a <=( A234  and  A233 );
 a10017a <=( A269  and  A266 );
 a10018a <=( (not A265)  and  a10017a );
 a10019a <=( a10018a  and  a10013a );
 a10022a <=( A199  and  A169 );
 a10026a <=( (not A202)  and  (not A201) );
 a10027a <=( A200  and  a10026a );
 a10028a <=( a10027a  and  a10022a );
 a10031a <=( A234  and  A233 );
 a10035a <=( A269  and  (not A266) );
 a10036a <=( A265  and  a10035a );
 a10037a <=( a10036a  and  a10031a );
 a10040a <=( A199  and  A169 );
 a10044a <=( (not A202)  and  (not A201) );
 a10045a <=( A200  and  a10044a );
 a10046a <=( a10045a  and  a10040a );
 a10049a <=( A233  and  (not A232) );
 a10053a <=( A300  and  A299 );
 a10054a <=( A236  and  a10053a );
 a10055a <=( a10054a  and  a10049a );
 a10058a <=( A199  and  A169 );
 a10062a <=( (not A202)  and  (not A201) );
 a10063a <=( A200  and  a10062a );
 a10064a <=( a10063a  and  a10058a );
 a10067a <=( A233  and  (not A232) );
 a10071a <=( A300  and  A298 );
 a10072a <=( A236  and  a10071a );
 a10073a <=( a10072a  and  a10067a );
 a10076a <=( A199  and  A169 );
 a10080a <=( (not A202)  and  (not A201) );
 a10081a <=( A200  and  a10080a );
 a10082a <=( a10081a  and  a10076a );
 a10085a <=( A233  and  (not A232) );
 a10089a <=( A267  and  A265 );
 a10090a <=( A236  and  a10089a );
 a10091a <=( a10090a  and  a10085a );
 a10094a <=( A199  and  A169 );
 a10098a <=( (not A202)  and  (not A201) );
 a10099a <=( A200  and  a10098a );
 a10100a <=( a10099a  and  a10094a );
 a10103a <=( A233  and  (not A232) );
 a10107a <=( A267  and  A266 );
 a10108a <=( A236  and  a10107a );
 a10109a <=( a10108a  and  a10103a );
 a10112a <=( A199  and  A169 );
 a10116a <=( (not A202)  and  (not A201) );
 a10117a <=( A200  and  a10116a );
 a10118a <=( a10117a  and  a10112a );
 a10121a <=( (not A233)  and  A232 );
 a10125a <=( A300  and  A299 );
 a10126a <=( A236  and  a10125a );
 a10127a <=( a10126a  and  a10121a );
 a10130a <=( A199  and  A169 );
 a10134a <=( (not A202)  and  (not A201) );
 a10135a <=( A200  and  a10134a );
 a10136a <=( a10135a  and  a10130a );
 a10139a <=( (not A233)  and  A232 );
 a10143a <=( A300  and  A298 );
 a10144a <=( A236  and  a10143a );
 a10145a <=( a10144a  and  a10139a );
 a10148a <=( A199  and  A169 );
 a10152a <=( (not A202)  and  (not A201) );
 a10153a <=( A200  and  a10152a );
 a10154a <=( a10153a  and  a10148a );
 a10157a <=( (not A233)  and  A232 );
 a10161a <=( A267  and  A265 );
 a10162a <=( A236  and  a10161a );
 a10163a <=( a10162a  and  a10157a );
 a10166a <=( A199  and  A169 );
 a10170a <=( (not A202)  and  (not A201) );
 a10171a <=( A200  and  a10170a );
 a10172a <=( a10171a  and  a10166a );
 a10175a <=( (not A233)  and  A232 );
 a10179a <=( A267  and  A266 );
 a10180a <=( A236  and  a10179a );
 a10181a <=( a10180a  and  a10175a );
 a10184a <=( (not A199)  and  A169 );
 a10188a <=( (not A232)  and  (not A202) );
 a10189a <=( (not A200)  and  a10188a );
 a10190a <=( a10189a  and  a10184a );
 a10193a <=( A236  and  A233 );
 a10197a <=( A302  and  (not A299) );
 a10198a <=( A298  and  a10197a );
 a10199a <=( a10198a  and  a10193a );
 a10202a <=( (not A199)  and  A169 );
 a10206a <=( (not A232)  and  (not A202) );
 a10207a <=( (not A200)  and  a10206a );
 a10208a <=( a10207a  and  a10202a );
 a10211a <=( A236  and  A233 );
 a10215a <=( A302  and  A299 );
 a10216a <=( (not A298)  and  a10215a );
 a10217a <=( a10216a  and  a10211a );
 a10220a <=( (not A199)  and  A169 );
 a10224a <=( (not A232)  and  (not A202) );
 a10225a <=( (not A200)  and  a10224a );
 a10226a <=( a10225a  and  a10220a );
 a10229a <=( A236  and  A233 );
 a10233a <=( A269  and  A266 );
 a10234a <=( (not A265)  and  a10233a );
 a10235a <=( a10234a  and  a10229a );
 a10238a <=( (not A199)  and  A169 );
 a10242a <=( (not A232)  and  (not A202) );
 a10243a <=( (not A200)  and  a10242a );
 a10244a <=( a10243a  and  a10238a );
 a10247a <=( A236  and  A233 );
 a10251a <=( A269  and  (not A266) );
 a10252a <=( A265  and  a10251a );
 a10253a <=( a10252a  and  a10247a );
 a10256a <=( (not A199)  and  A169 );
 a10260a <=( A232  and  (not A202) );
 a10261a <=( (not A200)  and  a10260a );
 a10262a <=( a10261a  and  a10256a );
 a10265a <=( A236  and  (not A233) );
 a10269a <=( A302  and  (not A299) );
 a10270a <=( A298  and  a10269a );
 a10271a <=( a10270a  and  a10265a );
 a10274a <=( (not A199)  and  A169 );
 a10278a <=( A232  and  (not A202) );
 a10279a <=( (not A200)  and  a10278a );
 a10280a <=( a10279a  and  a10274a );
 a10283a <=( A236  and  (not A233) );
 a10287a <=( A302  and  A299 );
 a10288a <=( (not A298)  and  a10287a );
 a10289a <=( a10288a  and  a10283a );
 a10292a <=( (not A199)  and  A169 );
 a10296a <=( A232  and  (not A202) );
 a10297a <=( (not A200)  and  a10296a );
 a10298a <=( a10297a  and  a10292a );
 a10301a <=( A236  and  (not A233) );
 a10305a <=( A269  and  A266 );
 a10306a <=( (not A265)  and  a10305a );
 a10307a <=( a10306a  and  a10301a );
 a10310a <=( (not A199)  and  A169 );
 a10314a <=( A232  and  (not A202) );
 a10315a <=( (not A200)  and  a10314a );
 a10316a <=( a10315a  and  a10310a );
 a10319a <=( A236  and  (not A233) );
 a10323a <=( A269  and  (not A266) );
 a10324a <=( A265  and  a10323a );
 a10325a <=( a10324a  and  a10319a );
 a10328a <=( A166  and  A168 );
 a10332a <=( (not A203)  and  (not A202) );
 a10333a <=( (not A201)  and  a10332a );
 a10334a <=( a10333a  and  a10328a );
 a10338a <=( A236  and  A233 );
 a10339a <=( (not A232)  and  a10338a );
 a10343a <=( A302  and  (not A299) );
 a10344a <=( A298  and  a10343a );
 a10345a <=( a10344a  and  a10339a );
 a10348a <=( A166  and  A168 );
 a10352a <=( (not A203)  and  (not A202) );
 a10353a <=( (not A201)  and  a10352a );
 a10354a <=( a10353a  and  a10348a );
 a10358a <=( A236  and  A233 );
 a10359a <=( (not A232)  and  a10358a );
 a10363a <=( A302  and  A299 );
 a10364a <=( (not A298)  and  a10363a );
 a10365a <=( a10364a  and  a10359a );
 a10368a <=( A166  and  A168 );
 a10372a <=( (not A203)  and  (not A202) );
 a10373a <=( (not A201)  and  a10372a );
 a10374a <=( a10373a  and  a10368a );
 a10378a <=( A236  and  A233 );
 a10379a <=( (not A232)  and  a10378a );
 a10383a <=( A269  and  A266 );
 a10384a <=( (not A265)  and  a10383a );
 a10385a <=( a10384a  and  a10379a );
 a10388a <=( A166  and  A168 );
 a10392a <=( (not A203)  and  (not A202) );
 a10393a <=( (not A201)  and  a10392a );
 a10394a <=( a10393a  and  a10388a );
 a10398a <=( A236  and  A233 );
 a10399a <=( (not A232)  and  a10398a );
 a10403a <=( A269  and  (not A266) );
 a10404a <=( A265  and  a10403a );
 a10405a <=( a10404a  and  a10399a );
 a10408a <=( A166  and  A168 );
 a10412a <=( (not A203)  and  (not A202) );
 a10413a <=( (not A201)  and  a10412a );
 a10414a <=( a10413a  and  a10408a );
 a10418a <=( A236  and  (not A233) );
 a10419a <=( A232  and  a10418a );
 a10423a <=( A302  and  (not A299) );
 a10424a <=( A298  and  a10423a );
 a10425a <=( a10424a  and  a10419a );
 a10428a <=( A166  and  A168 );
 a10432a <=( (not A203)  and  (not A202) );
 a10433a <=( (not A201)  and  a10432a );
 a10434a <=( a10433a  and  a10428a );
 a10438a <=( A236  and  (not A233) );
 a10439a <=( A232  and  a10438a );
 a10443a <=( A302  and  A299 );
 a10444a <=( (not A298)  and  a10443a );
 a10445a <=( a10444a  and  a10439a );
 a10448a <=( A166  and  A168 );
 a10452a <=( (not A203)  and  (not A202) );
 a10453a <=( (not A201)  and  a10452a );
 a10454a <=( a10453a  and  a10448a );
 a10458a <=( A236  and  (not A233) );
 a10459a <=( A232  and  a10458a );
 a10463a <=( A269  and  A266 );
 a10464a <=( (not A265)  and  a10463a );
 a10465a <=( a10464a  and  a10459a );
 a10468a <=( A166  and  A168 );
 a10472a <=( (not A203)  and  (not A202) );
 a10473a <=( (not A201)  and  a10472a );
 a10474a <=( a10473a  and  a10468a );
 a10478a <=( A236  and  (not A233) );
 a10479a <=( A232  and  a10478a );
 a10483a <=( A269  and  (not A266) );
 a10484a <=( A265  and  a10483a );
 a10485a <=( a10484a  and  a10479a );
 a10488a <=( A166  and  A168 );
 a10492a <=( (not A201)  and  A200 );
 a10493a <=( A199  and  a10492a );
 a10494a <=( a10493a  and  a10488a );
 a10498a <=( A234  and  A232 );
 a10499a <=( (not A202)  and  a10498a );
 a10503a <=( A302  and  (not A299) );
 a10504a <=( A298  and  a10503a );
 a10505a <=( a10504a  and  a10499a );
 a10508a <=( A166  and  A168 );
 a10512a <=( (not A201)  and  A200 );
 a10513a <=( A199  and  a10512a );
 a10514a <=( a10513a  and  a10508a );
 a10518a <=( A234  and  A232 );
 a10519a <=( (not A202)  and  a10518a );
 a10523a <=( A302  and  A299 );
 a10524a <=( (not A298)  and  a10523a );
 a10525a <=( a10524a  and  a10519a );
 a10528a <=( A166  and  A168 );
 a10532a <=( (not A201)  and  A200 );
 a10533a <=( A199  and  a10532a );
 a10534a <=( a10533a  and  a10528a );
 a10538a <=( A234  and  A232 );
 a10539a <=( (not A202)  and  a10538a );
 a10543a <=( A269  and  A266 );
 a10544a <=( (not A265)  and  a10543a );
 a10545a <=( a10544a  and  a10539a );
 a10548a <=( A166  and  A168 );
 a10552a <=( (not A201)  and  A200 );
 a10553a <=( A199  and  a10552a );
 a10554a <=( a10553a  and  a10548a );
 a10558a <=( A234  and  A232 );
 a10559a <=( (not A202)  and  a10558a );
 a10563a <=( A269  and  (not A266) );
 a10564a <=( A265  and  a10563a );
 a10565a <=( a10564a  and  a10559a );
 a10568a <=( A166  and  A168 );
 a10572a <=( (not A201)  and  A200 );
 a10573a <=( A199  and  a10572a );
 a10574a <=( a10573a  and  a10568a );
 a10578a <=( A234  and  A233 );
 a10579a <=( (not A202)  and  a10578a );
 a10583a <=( A302  and  (not A299) );
 a10584a <=( A298  and  a10583a );
 a10585a <=( a10584a  and  a10579a );
 a10588a <=( A166  and  A168 );
 a10592a <=( (not A201)  and  A200 );
 a10593a <=( A199  and  a10592a );
 a10594a <=( a10593a  and  a10588a );
 a10598a <=( A234  and  A233 );
 a10599a <=( (not A202)  and  a10598a );
 a10603a <=( A302  and  A299 );
 a10604a <=( (not A298)  and  a10603a );
 a10605a <=( a10604a  and  a10599a );
 a10608a <=( A166  and  A168 );
 a10612a <=( (not A201)  and  A200 );
 a10613a <=( A199  and  a10612a );
 a10614a <=( a10613a  and  a10608a );
 a10618a <=( A234  and  A233 );
 a10619a <=( (not A202)  and  a10618a );
 a10623a <=( A269  and  A266 );
 a10624a <=( (not A265)  and  a10623a );
 a10625a <=( a10624a  and  a10619a );
 a10628a <=( A166  and  A168 );
 a10632a <=( (not A201)  and  A200 );
 a10633a <=( A199  and  a10632a );
 a10634a <=( a10633a  and  a10628a );
 a10638a <=( A234  and  A233 );
 a10639a <=( (not A202)  and  a10638a );
 a10643a <=( A269  and  (not A266) );
 a10644a <=( A265  and  a10643a );
 a10645a <=( a10644a  and  a10639a );
 a10648a <=( A166  and  A168 );
 a10652a <=( (not A201)  and  A200 );
 a10653a <=( A199  and  a10652a );
 a10654a <=( a10653a  and  a10648a );
 a10658a <=( A233  and  (not A232) );
 a10659a <=( (not A202)  and  a10658a );
 a10663a <=( A300  and  A299 );
 a10664a <=( A236  and  a10663a );
 a10665a <=( a10664a  and  a10659a );
 a10668a <=( A166  and  A168 );
 a10672a <=( (not A201)  and  A200 );
 a10673a <=( A199  and  a10672a );
 a10674a <=( a10673a  and  a10668a );
 a10678a <=( A233  and  (not A232) );
 a10679a <=( (not A202)  and  a10678a );
 a10683a <=( A300  and  A298 );
 a10684a <=( A236  and  a10683a );
 a10685a <=( a10684a  and  a10679a );
 a10688a <=( A166  and  A168 );
 a10692a <=( (not A201)  and  A200 );
 a10693a <=( A199  and  a10692a );
 a10694a <=( a10693a  and  a10688a );
 a10698a <=( A233  and  (not A232) );
 a10699a <=( (not A202)  and  a10698a );
 a10703a <=( A267  and  A265 );
 a10704a <=( A236  and  a10703a );
 a10705a <=( a10704a  and  a10699a );
 a10708a <=( A166  and  A168 );
 a10712a <=( (not A201)  and  A200 );
 a10713a <=( A199  and  a10712a );
 a10714a <=( a10713a  and  a10708a );
 a10718a <=( A233  and  (not A232) );
 a10719a <=( (not A202)  and  a10718a );
 a10723a <=( A267  and  A266 );
 a10724a <=( A236  and  a10723a );
 a10725a <=( a10724a  and  a10719a );
 a10728a <=( A166  and  A168 );
 a10732a <=( (not A201)  and  A200 );
 a10733a <=( A199  and  a10732a );
 a10734a <=( a10733a  and  a10728a );
 a10738a <=( (not A233)  and  A232 );
 a10739a <=( (not A202)  and  a10738a );
 a10743a <=( A300  and  A299 );
 a10744a <=( A236  and  a10743a );
 a10745a <=( a10744a  and  a10739a );
 a10748a <=( A166  and  A168 );
 a10752a <=( (not A201)  and  A200 );
 a10753a <=( A199  and  a10752a );
 a10754a <=( a10753a  and  a10748a );
 a10758a <=( (not A233)  and  A232 );
 a10759a <=( (not A202)  and  a10758a );
 a10763a <=( A300  and  A298 );
 a10764a <=( A236  and  a10763a );
 a10765a <=( a10764a  and  a10759a );
 a10768a <=( A166  and  A168 );
 a10772a <=( (not A201)  and  A200 );
 a10773a <=( A199  and  a10772a );
 a10774a <=( a10773a  and  a10768a );
 a10778a <=( (not A233)  and  A232 );
 a10779a <=( (not A202)  and  a10778a );
 a10783a <=( A267  and  A265 );
 a10784a <=( A236  and  a10783a );
 a10785a <=( a10784a  and  a10779a );
 a10788a <=( A166  and  A168 );
 a10792a <=( (not A201)  and  A200 );
 a10793a <=( A199  and  a10792a );
 a10794a <=( a10793a  and  a10788a );
 a10798a <=( (not A233)  and  A232 );
 a10799a <=( (not A202)  and  a10798a );
 a10803a <=( A267  and  A266 );
 a10804a <=( A236  and  a10803a );
 a10805a <=( a10804a  and  a10799a );
 a10808a <=( A166  and  A168 );
 a10812a <=( (not A202)  and  (not A200) );
 a10813a <=( (not A199)  and  a10812a );
 a10814a <=( a10813a  and  a10808a );
 a10818a <=( A236  and  A233 );
 a10819a <=( (not A232)  and  a10818a );
 a10823a <=( A302  and  (not A299) );
 a10824a <=( A298  and  a10823a );
 a10825a <=( a10824a  and  a10819a );
 a10828a <=( A166  and  A168 );
 a10832a <=( (not A202)  and  (not A200) );
 a10833a <=( (not A199)  and  a10832a );
 a10834a <=( a10833a  and  a10828a );
 a10838a <=( A236  and  A233 );
 a10839a <=( (not A232)  and  a10838a );
 a10843a <=( A302  and  A299 );
 a10844a <=( (not A298)  and  a10843a );
 a10845a <=( a10844a  and  a10839a );
 a10848a <=( A166  and  A168 );
 a10852a <=( (not A202)  and  (not A200) );
 a10853a <=( (not A199)  and  a10852a );
 a10854a <=( a10853a  and  a10848a );
 a10858a <=( A236  and  A233 );
 a10859a <=( (not A232)  and  a10858a );
 a10863a <=( A269  and  A266 );
 a10864a <=( (not A265)  and  a10863a );
 a10865a <=( a10864a  and  a10859a );
 a10868a <=( A166  and  A168 );
 a10872a <=( (not A202)  and  (not A200) );
 a10873a <=( (not A199)  and  a10872a );
 a10874a <=( a10873a  and  a10868a );
 a10878a <=( A236  and  A233 );
 a10879a <=( (not A232)  and  a10878a );
 a10883a <=( A269  and  (not A266) );
 a10884a <=( A265  and  a10883a );
 a10885a <=( a10884a  and  a10879a );
 a10888a <=( A166  and  A168 );
 a10892a <=( (not A202)  and  (not A200) );
 a10893a <=( (not A199)  and  a10892a );
 a10894a <=( a10893a  and  a10888a );
 a10898a <=( A236  and  (not A233) );
 a10899a <=( A232  and  a10898a );
 a10903a <=( A302  and  (not A299) );
 a10904a <=( A298  and  a10903a );
 a10905a <=( a10904a  and  a10899a );
 a10908a <=( A166  and  A168 );
 a10912a <=( (not A202)  and  (not A200) );
 a10913a <=( (not A199)  and  a10912a );
 a10914a <=( a10913a  and  a10908a );
 a10918a <=( A236  and  (not A233) );
 a10919a <=( A232  and  a10918a );
 a10923a <=( A302  and  A299 );
 a10924a <=( (not A298)  and  a10923a );
 a10925a <=( a10924a  and  a10919a );
 a10928a <=( A166  and  A168 );
 a10932a <=( (not A202)  and  (not A200) );
 a10933a <=( (not A199)  and  a10932a );
 a10934a <=( a10933a  and  a10928a );
 a10938a <=( A236  and  (not A233) );
 a10939a <=( A232  and  a10938a );
 a10943a <=( A269  and  A266 );
 a10944a <=( (not A265)  and  a10943a );
 a10945a <=( a10944a  and  a10939a );
 a10948a <=( A166  and  A168 );
 a10952a <=( (not A202)  and  (not A200) );
 a10953a <=( (not A199)  and  a10952a );
 a10954a <=( a10953a  and  a10948a );
 a10958a <=( A236  and  (not A233) );
 a10959a <=( A232  and  a10958a );
 a10963a <=( A269  and  (not A266) );
 a10964a <=( A265  and  a10963a );
 a10965a <=( a10964a  and  a10959a );
 a10968a <=( A167  and  A168 );
 a10972a <=( (not A203)  and  (not A202) );
 a10973a <=( (not A201)  and  a10972a );
 a10974a <=( a10973a  and  a10968a );
 a10978a <=( A236  and  A233 );
 a10979a <=( (not A232)  and  a10978a );
 a10983a <=( A302  and  (not A299) );
 a10984a <=( A298  and  a10983a );
 a10985a <=( a10984a  and  a10979a );
 a10988a <=( A167  and  A168 );
 a10992a <=( (not A203)  and  (not A202) );
 a10993a <=( (not A201)  and  a10992a );
 a10994a <=( a10993a  and  a10988a );
 a10998a <=( A236  and  A233 );
 a10999a <=( (not A232)  and  a10998a );
 a11003a <=( A302  and  A299 );
 a11004a <=( (not A298)  and  a11003a );
 a11005a <=( a11004a  and  a10999a );
 a11008a <=( A167  and  A168 );
 a11012a <=( (not A203)  and  (not A202) );
 a11013a <=( (not A201)  and  a11012a );
 a11014a <=( a11013a  and  a11008a );
 a11018a <=( A236  and  A233 );
 a11019a <=( (not A232)  and  a11018a );
 a11023a <=( A269  and  A266 );
 a11024a <=( (not A265)  and  a11023a );
 a11025a <=( a11024a  and  a11019a );
 a11028a <=( A167  and  A168 );
 a11032a <=( (not A203)  and  (not A202) );
 a11033a <=( (not A201)  and  a11032a );
 a11034a <=( a11033a  and  a11028a );
 a11038a <=( A236  and  A233 );
 a11039a <=( (not A232)  and  a11038a );
 a11043a <=( A269  and  (not A266) );
 a11044a <=( A265  and  a11043a );
 a11045a <=( a11044a  and  a11039a );
 a11048a <=( A167  and  A168 );
 a11052a <=( (not A203)  and  (not A202) );
 a11053a <=( (not A201)  and  a11052a );
 a11054a <=( a11053a  and  a11048a );
 a11058a <=( A236  and  (not A233) );
 a11059a <=( A232  and  a11058a );
 a11063a <=( A302  and  (not A299) );
 a11064a <=( A298  and  a11063a );
 a11065a <=( a11064a  and  a11059a );
 a11068a <=( A167  and  A168 );
 a11072a <=( (not A203)  and  (not A202) );
 a11073a <=( (not A201)  and  a11072a );
 a11074a <=( a11073a  and  a11068a );
 a11078a <=( A236  and  (not A233) );
 a11079a <=( A232  and  a11078a );
 a11083a <=( A302  and  A299 );
 a11084a <=( (not A298)  and  a11083a );
 a11085a <=( a11084a  and  a11079a );
 a11088a <=( A167  and  A168 );
 a11092a <=( (not A203)  and  (not A202) );
 a11093a <=( (not A201)  and  a11092a );
 a11094a <=( a11093a  and  a11088a );
 a11098a <=( A236  and  (not A233) );
 a11099a <=( A232  and  a11098a );
 a11103a <=( A269  and  A266 );
 a11104a <=( (not A265)  and  a11103a );
 a11105a <=( a11104a  and  a11099a );
 a11108a <=( A167  and  A168 );
 a11112a <=( (not A203)  and  (not A202) );
 a11113a <=( (not A201)  and  a11112a );
 a11114a <=( a11113a  and  a11108a );
 a11118a <=( A236  and  (not A233) );
 a11119a <=( A232  and  a11118a );
 a11123a <=( A269  and  (not A266) );
 a11124a <=( A265  and  a11123a );
 a11125a <=( a11124a  and  a11119a );
 a11128a <=( A167  and  A168 );
 a11132a <=( (not A201)  and  A200 );
 a11133a <=( A199  and  a11132a );
 a11134a <=( a11133a  and  a11128a );
 a11138a <=( A234  and  A232 );
 a11139a <=( (not A202)  and  a11138a );
 a11143a <=( A302  and  (not A299) );
 a11144a <=( A298  and  a11143a );
 a11145a <=( a11144a  and  a11139a );
 a11148a <=( A167  and  A168 );
 a11152a <=( (not A201)  and  A200 );
 a11153a <=( A199  and  a11152a );
 a11154a <=( a11153a  and  a11148a );
 a11158a <=( A234  and  A232 );
 a11159a <=( (not A202)  and  a11158a );
 a11163a <=( A302  and  A299 );
 a11164a <=( (not A298)  and  a11163a );
 a11165a <=( a11164a  and  a11159a );
 a11168a <=( A167  and  A168 );
 a11172a <=( (not A201)  and  A200 );
 a11173a <=( A199  and  a11172a );
 a11174a <=( a11173a  and  a11168a );
 a11178a <=( A234  and  A232 );
 a11179a <=( (not A202)  and  a11178a );
 a11183a <=( A269  and  A266 );
 a11184a <=( (not A265)  and  a11183a );
 a11185a <=( a11184a  and  a11179a );
 a11188a <=( A167  and  A168 );
 a11192a <=( (not A201)  and  A200 );
 a11193a <=( A199  and  a11192a );
 a11194a <=( a11193a  and  a11188a );
 a11198a <=( A234  and  A232 );
 a11199a <=( (not A202)  and  a11198a );
 a11203a <=( A269  and  (not A266) );
 a11204a <=( A265  and  a11203a );
 a11205a <=( a11204a  and  a11199a );
 a11208a <=( A167  and  A168 );
 a11212a <=( (not A201)  and  A200 );
 a11213a <=( A199  and  a11212a );
 a11214a <=( a11213a  and  a11208a );
 a11218a <=( A234  and  A233 );
 a11219a <=( (not A202)  and  a11218a );
 a11223a <=( A302  and  (not A299) );
 a11224a <=( A298  and  a11223a );
 a11225a <=( a11224a  and  a11219a );
 a11228a <=( A167  and  A168 );
 a11232a <=( (not A201)  and  A200 );
 a11233a <=( A199  and  a11232a );
 a11234a <=( a11233a  and  a11228a );
 a11238a <=( A234  and  A233 );
 a11239a <=( (not A202)  and  a11238a );
 a11243a <=( A302  and  A299 );
 a11244a <=( (not A298)  and  a11243a );
 a11245a <=( a11244a  and  a11239a );
 a11248a <=( A167  and  A168 );
 a11252a <=( (not A201)  and  A200 );
 a11253a <=( A199  and  a11252a );
 a11254a <=( a11253a  and  a11248a );
 a11258a <=( A234  and  A233 );
 a11259a <=( (not A202)  and  a11258a );
 a11263a <=( A269  and  A266 );
 a11264a <=( (not A265)  and  a11263a );
 a11265a <=( a11264a  and  a11259a );
 a11268a <=( A167  and  A168 );
 a11272a <=( (not A201)  and  A200 );
 a11273a <=( A199  and  a11272a );
 a11274a <=( a11273a  and  a11268a );
 a11278a <=( A234  and  A233 );
 a11279a <=( (not A202)  and  a11278a );
 a11283a <=( A269  and  (not A266) );
 a11284a <=( A265  and  a11283a );
 a11285a <=( a11284a  and  a11279a );
 a11288a <=( A167  and  A168 );
 a11292a <=( (not A201)  and  A200 );
 a11293a <=( A199  and  a11292a );
 a11294a <=( a11293a  and  a11288a );
 a11298a <=( A233  and  (not A232) );
 a11299a <=( (not A202)  and  a11298a );
 a11303a <=( A300  and  A299 );
 a11304a <=( A236  and  a11303a );
 a11305a <=( a11304a  and  a11299a );
 a11308a <=( A167  and  A168 );
 a11312a <=( (not A201)  and  A200 );
 a11313a <=( A199  and  a11312a );
 a11314a <=( a11313a  and  a11308a );
 a11318a <=( A233  and  (not A232) );
 a11319a <=( (not A202)  and  a11318a );
 a11323a <=( A300  and  A298 );
 a11324a <=( A236  and  a11323a );
 a11325a <=( a11324a  and  a11319a );
 a11328a <=( A167  and  A168 );
 a11332a <=( (not A201)  and  A200 );
 a11333a <=( A199  and  a11332a );
 a11334a <=( a11333a  and  a11328a );
 a11338a <=( A233  and  (not A232) );
 a11339a <=( (not A202)  and  a11338a );
 a11343a <=( A267  and  A265 );
 a11344a <=( A236  and  a11343a );
 a11345a <=( a11344a  and  a11339a );
 a11348a <=( A167  and  A168 );
 a11352a <=( (not A201)  and  A200 );
 a11353a <=( A199  and  a11352a );
 a11354a <=( a11353a  and  a11348a );
 a11358a <=( A233  and  (not A232) );
 a11359a <=( (not A202)  and  a11358a );
 a11363a <=( A267  and  A266 );
 a11364a <=( A236  and  a11363a );
 a11365a <=( a11364a  and  a11359a );
 a11368a <=( A167  and  A168 );
 a11372a <=( (not A201)  and  A200 );
 a11373a <=( A199  and  a11372a );
 a11374a <=( a11373a  and  a11368a );
 a11378a <=( (not A233)  and  A232 );
 a11379a <=( (not A202)  and  a11378a );
 a11383a <=( A300  and  A299 );
 a11384a <=( A236  and  a11383a );
 a11385a <=( a11384a  and  a11379a );
 a11388a <=( A167  and  A168 );
 a11392a <=( (not A201)  and  A200 );
 a11393a <=( A199  and  a11392a );
 a11394a <=( a11393a  and  a11388a );
 a11398a <=( (not A233)  and  A232 );
 a11399a <=( (not A202)  and  a11398a );
 a11403a <=( A300  and  A298 );
 a11404a <=( A236  and  a11403a );
 a11405a <=( a11404a  and  a11399a );
 a11408a <=( A167  and  A168 );
 a11412a <=( (not A201)  and  A200 );
 a11413a <=( A199  and  a11412a );
 a11414a <=( a11413a  and  a11408a );
 a11418a <=( (not A233)  and  A232 );
 a11419a <=( (not A202)  and  a11418a );
 a11423a <=( A267  and  A265 );
 a11424a <=( A236  and  a11423a );
 a11425a <=( a11424a  and  a11419a );
 a11428a <=( A167  and  A168 );
 a11432a <=( (not A201)  and  A200 );
 a11433a <=( A199  and  a11432a );
 a11434a <=( a11433a  and  a11428a );
 a11438a <=( (not A233)  and  A232 );
 a11439a <=( (not A202)  and  a11438a );
 a11443a <=( A267  and  A266 );
 a11444a <=( A236  and  a11443a );
 a11445a <=( a11444a  and  a11439a );
 a11448a <=( A167  and  A168 );
 a11452a <=( (not A202)  and  (not A200) );
 a11453a <=( (not A199)  and  a11452a );
 a11454a <=( a11453a  and  a11448a );
 a11458a <=( A236  and  A233 );
 a11459a <=( (not A232)  and  a11458a );
 a11463a <=( A302  and  (not A299) );
 a11464a <=( A298  and  a11463a );
 a11465a <=( a11464a  and  a11459a );
 a11468a <=( A167  and  A168 );
 a11472a <=( (not A202)  and  (not A200) );
 a11473a <=( (not A199)  and  a11472a );
 a11474a <=( a11473a  and  a11468a );
 a11478a <=( A236  and  A233 );
 a11479a <=( (not A232)  and  a11478a );
 a11483a <=( A302  and  A299 );
 a11484a <=( (not A298)  and  a11483a );
 a11485a <=( a11484a  and  a11479a );
 a11488a <=( A167  and  A168 );
 a11492a <=( (not A202)  and  (not A200) );
 a11493a <=( (not A199)  and  a11492a );
 a11494a <=( a11493a  and  a11488a );
 a11498a <=( A236  and  A233 );
 a11499a <=( (not A232)  and  a11498a );
 a11503a <=( A269  and  A266 );
 a11504a <=( (not A265)  and  a11503a );
 a11505a <=( a11504a  and  a11499a );
 a11508a <=( A167  and  A168 );
 a11512a <=( (not A202)  and  (not A200) );
 a11513a <=( (not A199)  and  a11512a );
 a11514a <=( a11513a  and  a11508a );
 a11518a <=( A236  and  A233 );
 a11519a <=( (not A232)  and  a11518a );
 a11523a <=( A269  and  (not A266) );
 a11524a <=( A265  and  a11523a );
 a11525a <=( a11524a  and  a11519a );
 a11528a <=( A167  and  A168 );
 a11532a <=( (not A202)  and  (not A200) );
 a11533a <=( (not A199)  and  a11532a );
 a11534a <=( a11533a  and  a11528a );
 a11538a <=( A236  and  (not A233) );
 a11539a <=( A232  and  a11538a );
 a11543a <=( A302  and  (not A299) );
 a11544a <=( A298  and  a11543a );
 a11545a <=( a11544a  and  a11539a );
 a11548a <=( A167  and  A168 );
 a11552a <=( (not A202)  and  (not A200) );
 a11553a <=( (not A199)  and  a11552a );
 a11554a <=( a11553a  and  a11548a );
 a11558a <=( A236  and  (not A233) );
 a11559a <=( A232  and  a11558a );
 a11563a <=( A302  and  A299 );
 a11564a <=( (not A298)  and  a11563a );
 a11565a <=( a11564a  and  a11559a );
 a11568a <=( A167  and  A168 );
 a11572a <=( (not A202)  and  (not A200) );
 a11573a <=( (not A199)  and  a11572a );
 a11574a <=( a11573a  and  a11568a );
 a11578a <=( A236  and  (not A233) );
 a11579a <=( A232  and  a11578a );
 a11583a <=( A269  and  A266 );
 a11584a <=( (not A265)  and  a11583a );
 a11585a <=( a11584a  and  a11579a );
 a11588a <=( A167  and  A168 );
 a11592a <=( (not A202)  and  (not A200) );
 a11593a <=( (not A199)  and  a11592a );
 a11594a <=( a11593a  and  a11588a );
 a11598a <=( A236  and  (not A233) );
 a11599a <=( A232  and  a11598a );
 a11603a <=( A269  and  (not A266) );
 a11604a <=( A265  and  a11603a );
 a11605a <=( a11604a  and  a11599a );
 a11608a <=( A167  and  A170 );
 a11612a <=( (not A202)  and  (not A201) );
 a11613a <=( (not A166)  and  a11612a );
 a11614a <=( a11613a  and  a11608a );
 a11618a <=( A234  and  A232 );
 a11619a <=( (not A203)  and  a11618a );
 a11623a <=( A302  and  (not A299) );
 a11624a <=( A298  and  a11623a );
 a11625a <=( a11624a  and  a11619a );
 a11628a <=( A167  and  A170 );
 a11632a <=( (not A202)  and  (not A201) );
 a11633a <=( (not A166)  and  a11632a );
 a11634a <=( a11633a  and  a11628a );
 a11638a <=( A234  and  A232 );
 a11639a <=( (not A203)  and  a11638a );
 a11643a <=( A302  and  A299 );
 a11644a <=( (not A298)  and  a11643a );
 a11645a <=( a11644a  and  a11639a );
 a11648a <=( A167  and  A170 );
 a11652a <=( (not A202)  and  (not A201) );
 a11653a <=( (not A166)  and  a11652a );
 a11654a <=( a11653a  and  a11648a );
 a11658a <=( A234  and  A232 );
 a11659a <=( (not A203)  and  a11658a );
 a11663a <=( A269  and  A266 );
 a11664a <=( (not A265)  and  a11663a );
 a11665a <=( a11664a  and  a11659a );
 a11668a <=( A167  and  A170 );
 a11672a <=( (not A202)  and  (not A201) );
 a11673a <=( (not A166)  and  a11672a );
 a11674a <=( a11673a  and  a11668a );
 a11678a <=( A234  and  A232 );
 a11679a <=( (not A203)  and  a11678a );
 a11683a <=( A269  and  (not A266) );
 a11684a <=( A265  and  a11683a );
 a11685a <=( a11684a  and  a11679a );
 a11688a <=( A167  and  A170 );
 a11692a <=( (not A202)  and  (not A201) );
 a11693a <=( (not A166)  and  a11692a );
 a11694a <=( a11693a  and  a11688a );
 a11698a <=( A234  and  A233 );
 a11699a <=( (not A203)  and  a11698a );
 a11703a <=( A302  and  (not A299) );
 a11704a <=( A298  and  a11703a );
 a11705a <=( a11704a  and  a11699a );
 a11708a <=( A167  and  A170 );
 a11712a <=( (not A202)  and  (not A201) );
 a11713a <=( (not A166)  and  a11712a );
 a11714a <=( a11713a  and  a11708a );
 a11718a <=( A234  and  A233 );
 a11719a <=( (not A203)  and  a11718a );
 a11723a <=( A302  and  A299 );
 a11724a <=( (not A298)  and  a11723a );
 a11725a <=( a11724a  and  a11719a );
 a11728a <=( A167  and  A170 );
 a11732a <=( (not A202)  and  (not A201) );
 a11733a <=( (not A166)  and  a11732a );
 a11734a <=( a11733a  and  a11728a );
 a11738a <=( A234  and  A233 );
 a11739a <=( (not A203)  and  a11738a );
 a11743a <=( A269  and  A266 );
 a11744a <=( (not A265)  and  a11743a );
 a11745a <=( a11744a  and  a11739a );
 a11748a <=( A167  and  A170 );
 a11752a <=( (not A202)  and  (not A201) );
 a11753a <=( (not A166)  and  a11752a );
 a11754a <=( a11753a  and  a11748a );
 a11758a <=( A234  and  A233 );
 a11759a <=( (not A203)  and  a11758a );
 a11763a <=( A269  and  (not A266) );
 a11764a <=( A265  and  a11763a );
 a11765a <=( a11764a  and  a11759a );
 a11768a <=( A167  and  A170 );
 a11772a <=( (not A202)  and  (not A201) );
 a11773a <=( (not A166)  and  a11772a );
 a11774a <=( a11773a  and  a11768a );
 a11778a <=( A233  and  (not A232) );
 a11779a <=( (not A203)  and  a11778a );
 a11783a <=( A300  and  A299 );
 a11784a <=( A236  and  a11783a );
 a11785a <=( a11784a  and  a11779a );
 a11788a <=( A167  and  A170 );
 a11792a <=( (not A202)  and  (not A201) );
 a11793a <=( (not A166)  and  a11792a );
 a11794a <=( a11793a  and  a11788a );
 a11798a <=( A233  and  (not A232) );
 a11799a <=( (not A203)  and  a11798a );
 a11803a <=( A300  and  A298 );
 a11804a <=( A236  and  a11803a );
 a11805a <=( a11804a  and  a11799a );
 a11808a <=( A167  and  A170 );
 a11812a <=( (not A202)  and  (not A201) );
 a11813a <=( (not A166)  and  a11812a );
 a11814a <=( a11813a  and  a11808a );
 a11818a <=( A233  and  (not A232) );
 a11819a <=( (not A203)  and  a11818a );
 a11823a <=( A267  and  A265 );
 a11824a <=( A236  and  a11823a );
 a11825a <=( a11824a  and  a11819a );
 a11828a <=( A167  and  A170 );
 a11832a <=( (not A202)  and  (not A201) );
 a11833a <=( (not A166)  and  a11832a );
 a11834a <=( a11833a  and  a11828a );
 a11838a <=( A233  and  (not A232) );
 a11839a <=( (not A203)  and  a11838a );
 a11843a <=( A267  and  A266 );
 a11844a <=( A236  and  a11843a );
 a11845a <=( a11844a  and  a11839a );
 a11848a <=( A167  and  A170 );
 a11852a <=( (not A202)  and  (not A201) );
 a11853a <=( (not A166)  and  a11852a );
 a11854a <=( a11853a  and  a11848a );
 a11858a <=( (not A233)  and  A232 );
 a11859a <=( (not A203)  and  a11858a );
 a11863a <=( A300  and  A299 );
 a11864a <=( A236  and  a11863a );
 a11865a <=( a11864a  and  a11859a );
 a11868a <=( A167  and  A170 );
 a11872a <=( (not A202)  and  (not A201) );
 a11873a <=( (not A166)  and  a11872a );
 a11874a <=( a11873a  and  a11868a );
 a11878a <=( (not A233)  and  A232 );
 a11879a <=( (not A203)  and  a11878a );
 a11883a <=( A300  and  A298 );
 a11884a <=( A236  and  a11883a );
 a11885a <=( a11884a  and  a11879a );
 a11888a <=( A167  and  A170 );
 a11892a <=( (not A202)  and  (not A201) );
 a11893a <=( (not A166)  and  a11892a );
 a11894a <=( a11893a  and  a11888a );
 a11898a <=( (not A233)  and  A232 );
 a11899a <=( (not A203)  and  a11898a );
 a11903a <=( A267  and  A265 );
 a11904a <=( A236  and  a11903a );
 a11905a <=( a11904a  and  a11899a );
 a11908a <=( A167  and  A170 );
 a11912a <=( (not A202)  and  (not A201) );
 a11913a <=( (not A166)  and  a11912a );
 a11914a <=( a11913a  and  a11908a );
 a11918a <=( (not A233)  and  A232 );
 a11919a <=( (not A203)  and  a11918a );
 a11923a <=( A267  and  A266 );
 a11924a <=( A236  and  a11923a );
 a11925a <=( a11924a  and  a11919a );
 a11928a <=( A167  and  A170 );
 a11932a <=( A200  and  A199 );
 a11933a <=( (not A166)  and  a11932a );
 a11934a <=( a11933a  and  a11928a );
 a11938a <=( A235  and  (not A202) );
 a11939a <=( (not A201)  and  a11938a );
 a11943a <=( A302  and  (not A299) );
 a11944a <=( A298  and  a11943a );
 a11945a <=( a11944a  and  a11939a );
 a11948a <=( A167  and  A170 );
 a11952a <=( A200  and  A199 );
 a11953a <=( (not A166)  and  a11952a );
 a11954a <=( a11953a  and  a11948a );
 a11958a <=( A235  and  (not A202) );
 a11959a <=( (not A201)  and  a11958a );
 a11963a <=( A302  and  A299 );
 a11964a <=( (not A298)  and  a11963a );
 a11965a <=( a11964a  and  a11959a );
 a11968a <=( A167  and  A170 );
 a11972a <=( A200  and  A199 );
 a11973a <=( (not A166)  and  a11972a );
 a11974a <=( a11973a  and  a11968a );
 a11978a <=( A235  and  (not A202) );
 a11979a <=( (not A201)  and  a11978a );
 a11983a <=( A269  and  A266 );
 a11984a <=( (not A265)  and  a11983a );
 a11985a <=( a11984a  and  a11979a );
 a11988a <=( A167  and  A170 );
 a11992a <=( A200  and  A199 );
 a11993a <=( (not A166)  and  a11992a );
 a11994a <=( a11993a  and  a11988a );
 a11998a <=( A235  and  (not A202) );
 a11999a <=( (not A201)  and  a11998a );
 a12003a <=( A269  and  (not A266) );
 a12004a <=( A265  and  a12003a );
 a12005a <=( a12004a  and  a11999a );
 a12008a <=( A167  and  A170 );
 a12012a <=( A200  and  A199 );
 a12013a <=( (not A166)  and  a12012a );
 a12014a <=( a12013a  and  a12008a );
 a12018a <=( A232  and  (not A202) );
 a12019a <=( (not A201)  and  a12018a );
 a12023a <=( A300  and  A299 );
 a12024a <=( A234  and  a12023a );
 a12025a <=( a12024a  and  a12019a );
 a12028a <=( A167  and  A170 );
 a12032a <=( A200  and  A199 );
 a12033a <=( (not A166)  and  a12032a );
 a12034a <=( a12033a  and  a12028a );
 a12038a <=( A232  and  (not A202) );
 a12039a <=( (not A201)  and  a12038a );
 a12043a <=( A300  and  A298 );
 a12044a <=( A234  and  a12043a );
 a12045a <=( a12044a  and  a12039a );
 a12048a <=( A167  and  A170 );
 a12052a <=( A200  and  A199 );
 a12053a <=( (not A166)  and  a12052a );
 a12054a <=( a12053a  and  a12048a );
 a12058a <=( A232  and  (not A202) );
 a12059a <=( (not A201)  and  a12058a );
 a12063a <=( A267  and  A265 );
 a12064a <=( A234  and  a12063a );
 a12065a <=( a12064a  and  a12059a );
 a12068a <=( A167  and  A170 );
 a12072a <=( A200  and  A199 );
 a12073a <=( (not A166)  and  a12072a );
 a12074a <=( a12073a  and  a12068a );
 a12078a <=( A232  and  (not A202) );
 a12079a <=( (not A201)  and  a12078a );
 a12083a <=( A267  and  A266 );
 a12084a <=( A234  and  a12083a );
 a12085a <=( a12084a  and  a12079a );
 a12088a <=( A167  and  A170 );
 a12092a <=( A200  and  A199 );
 a12093a <=( (not A166)  and  a12092a );
 a12094a <=( a12093a  and  a12088a );
 a12098a <=( A233  and  (not A202) );
 a12099a <=( (not A201)  and  a12098a );
 a12103a <=( A300  and  A299 );
 a12104a <=( A234  and  a12103a );
 a12105a <=( a12104a  and  a12099a );
 a12108a <=( A167  and  A170 );
 a12112a <=( A200  and  A199 );
 a12113a <=( (not A166)  and  a12112a );
 a12114a <=( a12113a  and  a12108a );
 a12118a <=( A233  and  (not A202) );
 a12119a <=( (not A201)  and  a12118a );
 a12123a <=( A300  and  A298 );
 a12124a <=( A234  and  a12123a );
 a12125a <=( a12124a  and  a12119a );
 a12128a <=( A167  and  A170 );
 a12132a <=( A200  and  A199 );
 a12133a <=( (not A166)  and  a12132a );
 a12134a <=( a12133a  and  a12128a );
 a12138a <=( A233  and  (not A202) );
 a12139a <=( (not A201)  and  a12138a );
 a12143a <=( A267  and  A265 );
 a12144a <=( A234  and  a12143a );
 a12145a <=( a12144a  and  a12139a );
 a12148a <=( A167  and  A170 );
 a12152a <=( A200  and  A199 );
 a12153a <=( (not A166)  and  a12152a );
 a12154a <=( a12153a  and  a12148a );
 a12158a <=( A233  and  (not A202) );
 a12159a <=( (not A201)  and  a12158a );
 a12163a <=( A267  and  A266 );
 a12164a <=( A234  and  a12163a );
 a12165a <=( a12164a  and  a12159a );
 a12168a <=( A167  and  A170 );
 a12172a <=( A200  and  A199 );
 a12173a <=( (not A166)  and  a12172a );
 a12174a <=( a12173a  and  a12168a );
 a12178a <=( (not A232)  and  (not A202) );
 a12179a <=( (not A201)  and  a12178a );
 a12183a <=( A301  and  A236 );
 a12184a <=( A233  and  a12183a );
 a12185a <=( a12184a  and  a12179a );
 a12188a <=( A167  and  A170 );
 a12192a <=( A200  and  A199 );
 a12193a <=( (not A166)  and  a12192a );
 a12194a <=( a12193a  and  a12188a );
 a12198a <=( (not A232)  and  (not A202) );
 a12199a <=( (not A201)  and  a12198a );
 a12203a <=( A268  and  A236 );
 a12204a <=( A233  and  a12203a );
 a12205a <=( a12204a  and  a12199a );
 a12208a <=( A167  and  A170 );
 a12212a <=( A200  and  A199 );
 a12213a <=( (not A166)  and  a12212a );
 a12214a <=( a12213a  and  a12208a );
 a12218a <=( A232  and  (not A202) );
 a12219a <=( (not A201)  and  a12218a );
 a12223a <=( A301  and  A236 );
 a12224a <=( (not A233)  and  a12223a );
 a12225a <=( a12224a  and  a12219a );
 a12228a <=( A167  and  A170 );
 a12232a <=( A200  and  A199 );
 a12233a <=( (not A166)  and  a12232a );
 a12234a <=( a12233a  and  a12228a );
 a12238a <=( A232  and  (not A202) );
 a12239a <=( (not A201)  and  a12238a );
 a12243a <=( A268  and  A236 );
 a12244a <=( (not A233)  and  a12243a );
 a12245a <=( a12244a  and  a12239a );
 a12248a <=( A167  and  A170 );
 a12252a <=( (not A200)  and  (not A199) );
 a12253a <=( (not A166)  and  a12252a );
 a12254a <=( a12253a  and  a12248a );
 a12258a <=( A234  and  A232 );
 a12259a <=( (not A202)  and  a12258a );
 a12263a <=( A302  and  (not A299) );
 a12264a <=( A298  and  a12263a );
 a12265a <=( a12264a  and  a12259a );
 a12268a <=( A167  and  A170 );
 a12272a <=( (not A200)  and  (not A199) );
 a12273a <=( (not A166)  and  a12272a );
 a12274a <=( a12273a  and  a12268a );
 a12278a <=( A234  and  A232 );
 a12279a <=( (not A202)  and  a12278a );
 a12283a <=( A302  and  A299 );
 a12284a <=( (not A298)  and  a12283a );
 a12285a <=( a12284a  and  a12279a );
 a12288a <=( A167  and  A170 );
 a12292a <=( (not A200)  and  (not A199) );
 a12293a <=( (not A166)  and  a12292a );
 a12294a <=( a12293a  and  a12288a );
 a12298a <=( A234  and  A232 );
 a12299a <=( (not A202)  and  a12298a );
 a12303a <=( A269  and  A266 );
 a12304a <=( (not A265)  and  a12303a );
 a12305a <=( a12304a  and  a12299a );
 a12308a <=( A167  and  A170 );
 a12312a <=( (not A200)  and  (not A199) );
 a12313a <=( (not A166)  and  a12312a );
 a12314a <=( a12313a  and  a12308a );
 a12318a <=( A234  and  A232 );
 a12319a <=( (not A202)  and  a12318a );
 a12323a <=( A269  and  (not A266) );
 a12324a <=( A265  and  a12323a );
 a12325a <=( a12324a  and  a12319a );
 a12328a <=( A167  and  A170 );
 a12332a <=( (not A200)  and  (not A199) );
 a12333a <=( (not A166)  and  a12332a );
 a12334a <=( a12333a  and  a12328a );
 a12338a <=( A234  and  A233 );
 a12339a <=( (not A202)  and  a12338a );
 a12343a <=( A302  and  (not A299) );
 a12344a <=( A298  and  a12343a );
 a12345a <=( a12344a  and  a12339a );
 a12348a <=( A167  and  A170 );
 a12352a <=( (not A200)  and  (not A199) );
 a12353a <=( (not A166)  and  a12352a );
 a12354a <=( a12353a  and  a12348a );
 a12358a <=( A234  and  A233 );
 a12359a <=( (not A202)  and  a12358a );
 a12363a <=( A302  and  A299 );
 a12364a <=( (not A298)  and  a12363a );
 a12365a <=( a12364a  and  a12359a );
 a12368a <=( A167  and  A170 );
 a12372a <=( (not A200)  and  (not A199) );
 a12373a <=( (not A166)  and  a12372a );
 a12374a <=( a12373a  and  a12368a );
 a12378a <=( A234  and  A233 );
 a12379a <=( (not A202)  and  a12378a );
 a12383a <=( A269  and  A266 );
 a12384a <=( (not A265)  and  a12383a );
 a12385a <=( a12384a  and  a12379a );
 a12388a <=( A167  and  A170 );
 a12392a <=( (not A200)  and  (not A199) );
 a12393a <=( (not A166)  and  a12392a );
 a12394a <=( a12393a  and  a12388a );
 a12398a <=( A234  and  A233 );
 a12399a <=( (not A202)  and  a12398a );
 a12403a <=( A269  and  (not A266) );
 a12404a <=( A265  and  a12403a );
 a12405a <=( a12404a  and  a12399a );
 a12408a <=( A167  and  A170 );
 a12412a <=( (not A200)  and  (not A199) );
 a12413a <=( (not A166)  and  a12412a );
 a12414a <=( a12413a  and  a12408a );
 a12418a <=( A233  and  (not A232) );
 a12419a <=( (not A202)  and  a12418a );
 a12423a <=( A300  and  A299 );
 a12424a <=( A236  and  a12423a );
 a12425a <=( a12424a  and  a12419a );
 a12428a <=( A167  and  A170 );
 a12432a <=( (not A200)  and  (not A199) );
 a12433a <=( (not A166)  and  a12432a );
 a12434a <=( a12433a  and  a12428a );
 a12438a <=( A233  and  (not A232) );
 a12439a <=( (not A202)  and  a12438a );
 a12443a <=( A300  and  A298 );
 a12444a <=( A236  and  a12443a );
 a12445a <=( a12444a  and  a12439a );
 a12448a <=( A167  and  A170 );
 a12452a <=( (not A200)  and  (not A199) );
 a12453a <=( (not A166)  and  a12452a );
 a12454a <=( a12453a  and  a12448a );
 a12458a <=( A233  and  (not A232) );
 a12459a <=( (not A202)  and  a12458a );
 a12463a <=( A267  and  A265 );
 a12464a <=( A236  and  a12463a );
 a12465a <=( a12464a  and  a12459a );
 a12468a <=( A167  and  A170 );
 a12472a <=( (not A200)  and  (not A199) );
 a12473a <=( (not A166)  and  a12472a );
 a12474a <=( a12473a  and  a12468a );
 a12478a <=( A233  and  (not A232) );
 a12479a <=( (not A202)  and  a12478a );
 a12483a <=( A267  and  A266 );
 a12484a <=( A236  and  a12483a );
 a12485a <=( a12484a  and  a12479a );
 a12488a <=( A167  and  A170 );
 a12492a <=( (not A200)  and  (not A199) );
 a12493a <=( (not A166)  and  a12492a );
 a12494a <=( a12493a  and  a12488a );
 a12498a <=( (not A233)  and  A232 );
 a12499a <=( (not A202)  and  a12498a );
 a12503a <=( A300  and  A299 );
 a12504a <=( A236  and  a12503a );
 a12505a <=( a12504a  and  a12499a );
 a12508a <=( A167  and  A170 );
 a12512a <=( (not A200)  and  (not A199) );
 a12513a <=( (not A166)  and  a12512a );
 a12514a <=( a12513a  and  a12508a );
 a12518a <=( (not A233)  and  A232 );
 a12519a <=( (not A202)  and  a12518a );
 a12523a <=( A300  and  A298 );
 a12524a <=( A236  and  a12523a );
 a12525a <=( a12524a  and  a12519a );
 a12528a <=( A167  and  A170 );
 a12532a <=( (not A200)  and  (not A199) );
 a12533a <=( (not A166)  and  a12532a );
 a12534a <=( a12533a  and  a12528a );
 a12538a <=( (not A233)  and  A232 );
 a12539a <=( (not A202)  and  a12538a );
 a12543a <=( A267  and  A265 );
 a12544a <=( A236  and  a12543a );
 a12545a <=( a12544a  and  a12539a );
 a12548a <=( A167  and  A170 );
 a12552a <=( (not A200)  and  (not A199) );
 a12553a <=( (not A166)  and  a12552a );
 a12554a <=( a12553a  and  a12548a );
 a12558a <=( (not A233)  and  A232 );
 a12559a <=( (not A202)  and  a12558a );
 a12563a <=( A267  and  A266 );
 a12564a <=( A236  and  a12563a );
 a12565a <=( a12564a  and  a12559a );
 a12568a <=( (not A167)  and  A170 );
 a12572a <=( (not A202)  and  (not A201) );
 a12573a <=( A166  and  a12572a );
 a12574a <=( a12573a  and  a12568a );
 a12578a <=( A234  and  A232 );
 a12579a <=( (not A203)  and  a12578a );
 a12583a <=( A302  and  (not A299) );
 a12584a <=( A298  and  a12583a );
 a12585a <=( a12584a  and  a12579a );
 a12588a <=( (not A167)  and  A170 );
 a12592a <=( (not A202)  and  (not A201) );
 a12593a <=( A166  and  a12592a );
 a12594a <=( a12593a  and  a12588a );
 a12598a <=( A234  and  A232 );
 a12599a <=( (not A203)  and  a12598a );
 a12603a <=( A302  and  A299 );
 a12604a <=( (not A298)  and  a12603a );
 a12605a <=( a12604a  and  a12599a );
 a12608a <=( (not A167)  and  A170 );
 a12612a <=( (not A202)  and  (not A201) );
 a12613a <=( A166  and  a12612a );
 a12614a <=( a12613a  and  a12608a );
 a12618a <=( A234  and  A232 );
 a12619a <=( (not A203)  and  a12618a );
 a12623a <=( A269  and  A266 );
 a12624a <=( (not A265)  and  a12623a );
 a12625a <=( a12624a  and  a12619a );
 a12628a <=( (not A167)  and  A170 );
 a12632a <=( (not A202)  and  (not A201) );
 a12633a <=( A166  and  a12632a );
 a12634a <=( a12633a  and  a12628a );
 a12638a <=( A234  and  A232 );
 a12639a <=( (not A203)  and  a12638a );
 a12643a <=( A269  and  (not A266) );
 a12644a <=( A265  and  a12643a );
 a12645a <=( a12644a  and  a12639a );
 a12648a <=( (not A167)  and  A170 );
 a12652a <=( (not A202)  and  (not A201) );
 a12653a <=( A166  and  a12652a );
 a12654a <=( a12653a  and  a12648a );
 a12658a <=( A234  and  A233 );
 a12659a <=( (not A203)  and  a12658a );
 a12663a <=( A302  and  (not A299) );
 a12664a <=( A298  and  a12663a );
 a12665a <=( a12664a  and  a12659a );
 a12668a <=( (not A167)  and  A170 );
 a12672a <=( (not A202)  and  (not A201) );
 a12673a <=( A166  and  a12672a );
 a12674a <=( a12673a  and  a12668a );
 a12678a <=( A234  and  A233 );
 a12679a <=( (not A203)  and  a12678a );
 a12683a <=( A302  and  A299 );
 a12684a <=( (not A298)  and  a12683a );
 a12685a <=( a12684a  and  a12679a );
 a12688a <=( (not A167)  and  A170 );
 a12692a <=( (not A202)  and  (not A201) );
 a12693a <=( A166  and  a12692a );
 a12694a <=( a12693a  and  a12688a );
 a12698a <=( A234  and  A233 );
 a12699a <=( (not A203)  and  a12698a );
 a12703a <=( A269  and  A266 );
 a12704a <=( (not A265)  and  a12703a );
 a12705a <=( a12704a  and  a12699a );
 a12708a <=( (not A167)  and  A170 );
 a12712a <=( (not A202)  and  (not A201) );
 a12713a <=( A166  and  a12712a );
 a12714a <=( a12713a  and  a12708a );
 a12718a <=( A234  and  A233 );
 a12719a <=( (not A203)  and  a12718a );
 a12723a <=( A269  and  (not A266) );
 a12724a <=( A265  and  a12723a );
 a12725a <=( a12724a  and  a12719a );
 a12728a <=( (not A167)  and  A170 );
 a12732a <=( (not A202)  and  (not A201) );
 a12733a <=( A166  and  a12732a );
 a12734a <=( a12733a  and  a12728a );
 a12738a <=( A233  and  (not A232) );
 a12739a <=( (not A203)  and  a12738a );
 a12743a <=( A300  and  A299 );
 a12744a <=( A236  and  a12743a );
 a12745a <=( a12744a  and  a12739a );
 a12748a <=( (not A167)  and  A170 );
 a12752a <=( (not A202)  and  (not A201) );
 a12753a <=( A166  and  a12752a );
 a12754a <=( a12753a  and  a12748a );
 a12758a <=( A233  and  (not A232) );
 a12759a <=( (not A203)  and  a12758a );
 a12763a <=( A300  and  A298 );
 a12764a <=( A236  and  a12763a );
 a12765a <=( a12764a  and  a12759a );
 a12768a <=( (not A167)  and  A170 );
 a12772a <=( (not A202)  and  (not A201) );
 a12773a <=( A166  and  a12772a );
 a12774a <=( a12773a  and  a12768a );
 a12778a <=( A233  and  (not A232) );
 a12779a <=( (not A203)  and  a12778a );
 a12783a <=( A267  and  A265 );
 a12784a <=( A236  and  a12783a );
 a12785a <=( a12784a  and  a12779a );
 a12788a <=( (not A167)  and  A170 );
 a12792a <=( (not A202)  and  (not A201) );
 a12793a <=( A166  and  a12792a );
 a12794a <=( a12793a  and  a12788a );
 a12798a <=( A233  and  (not A232) );
 a12799a <=( (not A203)  and  a12798a );
 a12803a <=( A267  and  A266 );
 a12804a <=( A236  and  a12803a );
 a12805a <=( a12804a  and  a12799a );
 a12808a <=( (not A167)  and  A170 );
 a12812a <=( (not A202)  and  (not A201) );
 a12813a <=( A166  and  a12812a );
 a12814a <=( a12813a  and  a12808a );
 a12818a <=( (not A233)  and  A232 );
 a12819a <=( (not A203)  and  a12818a );
 a12823a <=( A300  and  A299 );
 a12824a <=( A236  and  a12823a );
 a12825a <=( a12824a  and  a12819a );
 a12828a <=( (not A167)  and  A170 );
 a12832a <=( (not A202)  and  (not A201) );
 a12833a <=( A166  and  a12832a );
 a12834a <=( a12833a  and  a12828a );
 a12838a <=( (not A233)  and  A232 );
 a12839a <=( (not A203)  and  a12838a );
 a12843a <=( A300  and  A298 );
 a12844a <=( A236  and  a12843a );
 a12845a <=( a12844a  and  a12839a );
 a12848a <=( (not A167)  and  A170 );
 a12852a <=( (not A202)  and  (not A201) );
 a12853a <=( A166  and  a12852a );
 a12854a <=( a12853a  and  a12848a );
 a12858a <=( (not A233)  and  A232 );
 a12859a <=( (not A203)  and  a12858a );
 a12863a <=( A267  and  A265 );
 a12864a <=( A236  and  a12863a );
 a12865a <=( a12864a  and  a12859a );
 a12868a <=( (not A167)  and  A170 );
 a12872a <=( (not A202)  and  (not A201) );
 a12873a <=( A166  and  a12872a );
 a12874a <=( a12873a  and  a12868a );
 a12878a <=( (not A233)  and  A232 );
 a12879a <=( (not A203)  and  a12878a );
 a12883a <=( A267  and  A266 );
 a12884a <=( A236  and  a12883a );
 a12885a <=( a12884a  and  a12879a );
 a12888a <=( (not A167)  and  A170 );
 a12892a <=( A200  and  A199 );
 a12893a <=( A166  and  a12892a );
 a12894a <=( a12893a  and  a12888a );
 a12898a <=( A235  and  (not A202) );
 a12899a <=( (not A201)  and  a12898a );
 a12903a <=( A302  and  (not A299) );
 a12904a <=( A298  and  a12903a );
 a12905a <=( a12904a  and  a12899a );
 a12908a <=( (not A167)  and  A170 );
 a12912a <=( A200  and  A199 );
 a12913a <=( A166  and  a12912a );
 a12914a <=( a12913a  and  a12908a );
 a12918a <=( A235  and  (not A202) );
 a12919a <=( (not A201)  and  a12918a );
 a12923a <=( A302  and  A299 );
 a12924a <=( (not A298)  and  a12923a );
 a12925a <=( a12924a  and  a12919a );
 a12928a <=( (not A167)  and  A170 );
 a12932a <=( A200  and  A199 );
 a12933a <=( A166  and  a12932a );
 a12934a <=( a12933a  and  a12928a );
 a12938a <=( A235  and  (not A202) );
 a12939a <=( (not A201)  and  a12938a );
 a12943a <=( A269  and  A266 );
 a12944a <=( (not A265)  and  a12943a );
 a12945a <=( a12944a  and  a12939a );
 a12948a <=( (not A167)  and  A170 );
 a12952a <=( A200  and  A199 );
 a12953a <=( A166  and  a12952a );
 a12954a <=( a12953a  and  a12948a );
 a12958a <=( A235  and  (not A202) );
 a12959a <=( (not A201)  and  a12958a );
 a12963a <=( A269  and  (not A266) );
 a12964a <=( A265  and  a12963a );
 a12965a <=( a12964a  and  a12959a );
 a12968a <=( (not A167)  and  A170 );
 a12972a <=( A200  and  A199 );
 a12973a <=( A166  and  a12972a );
 a12974a <=( a12973a  and  a12968a );
 a12978a <=( A232  and  (not A202) );
 a12979a <=( (not A201)  and  a12978a );
 a12983a <=( A300  and  A299 );
 a12984a <=( A234  and  a12983a );
 a12985a <=( a12984a  and  a12979a );
 a12988a <=( (not A167)  and  A170 );
 a12992a <=( A200  and  A199 );
 a12993a <=( A166  and  a12992a );
 a12994a <=( a12993a  and  a12988a );
 a12998a <=( A232  and  (not A202) );
 a12999a <=( (not A201)  and  a12998a );
 a13003a <=( A300  and  A298 );
 a13004a <=( A234  and  a13003a );
 a13005a <=( a13004a  and  a12999a );
 a13008a <=( (not A167)  and  A170 );
 a13012a <=( A200  and  A199 );
 a13013a <=( A166  and  a13012a );
 a13014a <=( a13013a  and  a13008a );
 a13018a <=( A232  and  (not A202) );
 a13019a <=( (not A201)  and  a13018a );
 a13023a <=( A267  and  A265 );
 a13024a <=( A234  and  a13023a );
 a13025a <=( a13024a  and  a13019a );
 a13028a <=( (not A167)  and  A170 );
 a13032a <=( A200  and  A199 );
 a13033a <=( A166  and  a13032a );
 a13034a <=( a13033a  and  a13028a );
 a13038a <=( A232  and  (not A202) );
 a13039a <=( (not A201)  and  a13038a );
 a13043a <=( A267  and  A266 );
 a13044a <=( A234  and  a13043a );
 a13045a <=( a13044a  and  a13039a );
 a13048a <=( (not A167)  and  A170 );
 a13052a <=( A200  and  A199 );
 a13053a <=( A166  and  a13052a );
 a13054a <=( a13053a  and  a13048a );
 a13058a <=( A233  and  (not A202) );
 a13059a <=( (not A201)  and  a13058a );
 a13063a <=( A300  and  A299 );
 a13064a <=( A234  and  a13063a );
 a13065a <=( a13064a  and  a13059a );
 a13068a <=( (not A167)  and  A170 );
 a13072a <=( A200  and  A199 );
 a13073a <=( A166  and  a13072a );
 a13074a <=( a13073a  and  a13068a );
 a13078a <=( A233  and  (not A202) );
 a13079a <=( (not A201)  and  a13078a );
 a13083a <=( A300  and  A298 );
 a13084a <=( A234  and  a13083a );
 a13085a <=( a13084a  and  a13079a );
 a13088a <=( (not A167)  and  A170 );
 a13092a <=( A200  and  A199 );
 a13093a <=( A166  and  a13092a );
 a13094a <=( a13093a  and  a13088a );
 a13098a <=( A233  and  (not A202) );
 a13099a <=( (not A201)  and  a13098a );
 a13103a <=( A267  and  A265 );
 a13104a <=( A234  and  a13103a );
 a13105a <=( a13104a  and  a13099a );
 a13108a <=( (not A167)  and  A170 );
 a13112a <=( A200  and  A199 );
 a13113a <=( A166  and  a13112a );
 a13114a <=( a13113a  and  a13108a );
 a13118a <=( A233  and  (not A202) );
 a13119a <=( (not A201)  and  a13118a );
 a13123a <=( A267  and  A266 );
 a13124a <=( A234  and  a13123a );
 a13125a <=( a13124a  and  a13119a );
 a13128a <=( (not A167)  and  A170 );
 a13132a <=( A200  and  A199 );
 a13133a <=( A166  and  a13132a );
 a13134a <=( a13133a  and  a13128a );
 a13138a <=( (not A232)  and  (not A202) );
 a13139a <=( (not A201)  and  a13138a );
 a13143a <=( A301  and  A236 );
 a13144a <=( A233  and  a13143a );
 a13145a <=( a13144a  and  a13139a );
 a13148a <=( (not A167)  and  A170 );
 a13152a <=( A200  and  A199 );
 a13153a <=( A166  and  a13152a );
 a13154a <=( a13153a  and  a13148a );
 a13158a <=( (not A232)  and  (not A202) );
 a13159a <=( (not A201)  and  a13158a );
 a13163a <=( A268  and  A236 );
 a13164a <=( A233  and  a13163a );
 a13165a <=( a13164a  and  a13159a );
 a13168a <=( (not A167)  and  A170 );
 a13172a <=( A200  and  A199 );
 a13173a <=( A166  and  a13172a );
 a13174a <=( a13173a  and  a13168a );
 a13178a <=( A232  and  (not A202) );
 a13179a <=( (not A201)  and  a13178a );
 a13183a <=( A301  and  A236 );
 a13184a <=( (not A233)  and  a13183a );
 a13185a <=( a13184a  and  a13179a );
 a13188a <=( (not A167)  and  A170 );
 a13192a <=( A200  and  A199 );
 a13193a <=( A166  and  a13192a );
 a13194a <=( a13193a  and  a13188a );
 a13198a <=( A232  and  (not A202) );
 a13199a <=( (not A201)  and  a13198a );
 a13203a <=( A268  and  A236 );
 a13204a <=( (not A233)  and  a13203a );
 a13205a <=( a13204a  and  a13199a );
 a13208a <=( (not A167)  and  A170 );
 a13212a <=( (not A200)  and  (not A199) );
 a13213a <=( A166  and  a13212a );
 a13214a <=( a13213a  and  a13208a );
 a13218a <=( A234  and  A232 );
 a13219a <=( (not A202)  and  a13218a );
 a13223a <=( A302  and  (not A299) );
 a13224a <=( A298  and  a13223a );
 a13225a <=( a13224a  and  a13219a );
 a13228a <=( (not A167)  and  A170 );
 a13232a <=( (not A200)  and  (not A199) );
 a13233a <=( A166  and  a13232a );
 a13234a <=( a13233a  and  a13228a );
 a13238a <=( A234  and  A232 );
 a13239a <=( (not A202)  and  a13238a );
 a13243a <=( A302  and  A299 );
 a13244a <=( (not A298)  and  a13243a );
 a13245a <=( a13244a  and  a13239a );
 a13248a <=( (not A167)  and  A170 );
 a13252a <=( (not A200)  and  (not A199) );
 a13253a <=( A166  and  a13252a );
 a13254a <=( a13253a  and  a13248a );
 a13258a <=( A234  and  A232 );
 a13259a <=( (not A202)  and  a13258a );
 a13263a <=( A269  and  A266 );
 a13264a <=( (not A265)  and  a13263a );
 a13265a <=( a13264a  and  a13259a );
 a13268a <=( (not A167)  and  A170 );
 a13272a <=( (not A200)  and  (not A199) );
 a13273a <=( A166  and  a13272a );
 a13274a <=( a13273a  and  a13268a );
 a13278a <=( A234  and  A232 );
 a13279a <=( (not A202)  and  a13278a );
 a13283a <=( A269  and  (not A266) );
 a13284a <=( A265  and  a13283a );
 a13285a <=( a13284a  and  a13279a );
 a13288a <=( (not A167)  and  A170 );
 a13292a <=( (not A200)  and  (not A199) );
 a13293a <=( A166  and  a13292a );
 a13294a <=( a13293a  and  a13288a );
 a13298a <=( A234  and  A233 );
 a13299a <=( (not A202)  and  a13298a );
 a13303a <=( A302  and  (not A299) );
 a13304a <=( A298  and  a13303a );
 a13305a <=( a13304a  and  a13299a );
 a13308a <=( (not A167)  and  A170 );
 a13312a <=( (not A200)  and  (not A199) );
 a13313a <=( A166  and  a13312a );
 a13314a <=( a13313a  and  a13308a );
 a13318a <=( A234  and  A233 );
 a13319a <=( (not A202)  and  a13318a );
 a13323a <=( A302  and  A299 );
 a13324a <=( (not A298)  and  a13323a );
 a13325a <=( a13324a  and  a13319a );
 a13328a <=( (not A167)  and  A170 );
 a13332a <=( (not A200)  and  (not A199) );
 a13333a <=( A166  and  a13332a );
 a13334a <=( a13333a  and  a13328a );
 a13338a <=( A234  and  A233 );
 a13339a <=( (not A202)  and  a13338a );
 a13343a <=( A269  and  A266 );
 a13344a <=( (not A265)  and  a13343a );
 a13345a <=( a13344a  and  a13339a );
 a13348a <=( (not A167)  and  A170 );
 a13352a <=( (not A200)  and  (not A199) );
 a13353a <=( A166  and  a13352a );
 a13354a <=( a13353a  and  a13348a );
 a13358a <=( A234  and  A233 );
 a13359a <=( (not A202)  and  a13358a );
 a13363a <=( A269  and  (not A266) );
 a13364a <=( A265  and  a13363a );
 a13365a <=( a13364a  and  a13359a );
 a13368a <=( (not A167)  and  A170 );
 a13372a <=( (not A200)  and  (not A199) );
 a13373a <=( A166  and  a13372a );
 a13374a <=( a13373a  and  a13368a );
 a13378a <=( A233  and  (not A232) );
 a13379a <=( (not A202)  and  a13378a );
 a13383a <=( A300  and  A299 );
 a13384a <=( A236  and  a13383a );
 a13385a <=( a13384a  and  a13379a );
 a13388a <=( (not A167)  and  A170 );
 a13392a <=( (not A200)  and  (not A199) );
 a13393a <=( A166  and  a13392a );
 a13394a <=( a13393a  and  a13388a );
 a13398a <=( A233  and  (not A232) );
 a13399a <=( (not A202)  and  a13398a );
 a13403a <=( A300  and  A298 );
 a13404a <=( A236  and  a13403a );
 a13405a <=( a13404a  and  a13399a );
 a13408a <=( (not A167)  and  A170 );
 a13412a <=( (not A200)  and  (not A199) );
 a13413a <=( A166  and  a13412a );
 a13414a <=( a13413a  and  a13408a );
 a13418a <=( A233  and  (not A232) );
 a13419a <=( (not A202)  and  a13418a );
 a13423a <=( A267  and  A265 );
 a13424a <=( A236  and  a13423a );
 a13425a <=( a13424a  and  a13419a );
 a13428a <=( (not A167)  and  A170 );
 a13432a <=( (not A200)  and  (not A199) );
 a13433a <=( A166  and  a13432a );
 a13434a <=( a13433a  and  a13428a );
 a13438a <=( A233  and  (not A232) );
 a13439a <=( (not A202)  and  a13438a );
 a13443a <=( A267  and  A266 );
 a13444a <=( A236  and  a13443a );
 a13445a <=( a13444a  and  a13439a );
 a13448a <=( (not A167)  and  A170 );
 a13452a <=( (not A200)  and  (not A199) );
 a13453a <=( A166  and  a13452a );
 a13454a <=( a13453a  and  a13448a );
 a13458a <=( (not A233)  and  A232 );
 a13459a <=( (not A202)  and  a13458a );
 a13463a <=( A300  and  A299 );
 a13464a <=( A236  and  a13463a );
 a13465a <=( a13464a  and  a13459a );
 a13468a <=( (not A167)  and  A170 );
 a13472a <=( (not A200)  and  (not A199) );
 a13473a <=( A166  and  a13472a );
 a13474a <=( a13473a  and  a13468a );
 a13478a <=( (not A233)  and  A232 );
 a13479a <=( (not A202)  and  a13478a );
 a13483a <=( A300  and  A298 );
 a13484a <=( A236  and  a13483a );
 a13485a <=( a13484a  and  a13479a );
 a13488a <=( (not A167)  and  A170 );
 a13492a <=( (not A200)  and  (not A199) );
 a13493a <=( A166  and  a13492a );
 a13494a <=( a13493a  and  a13488a );
 a13498a <=( (not A233)  and  A232 );
 a13499a <=( (not A202)  and  a13498a );
 a13503a <=( A267  and  A265 );
 a13504a <=( A236  and  a13503a );
 a13505a <=( a13504a  and  a13499a );
 a13508a <=( (not A167)  and  A170 );
 a13512a <=( (not A200)  and  (not A199) );
 a13513a <=( A166  and  a13512a );
 a13514a <=( a13513a  and  a13508a );
 a13518a <=( (not A233)  and  A232 );
 a13519a <=( (not A202)  and  a13518a );
 a13523a <=( A267  and  A266 );
 a13524a <=( A236  and  a13523a );
 a13525a <=( a13524a  and  a13519a );
 a13528a <=( A199  and  A169 );
 a13532a <=( (not A202)  and  (not A201) );
 a13533a <=( A200  and  a13532a );
 a13534a <=( a13533a  and  a13528a );
 a13538a <=( A236  and  A233 );
 a13539a <=( (not A232)  and  a13538a );
 a13543a <=( A302  and  (not A299) );
 a13544a <=( A298  and  a13543a );
 a13545a <=( a13544a  and  a13539a );
 a13548a <=( A199  and  A169 );
 a13552a <=( (not A202)  and  (not A201) );
 a13553a <=( A200  and  a13552a );
 a13554a <=( a13553a  and  a13548a );
 a13558a <=( A236  and  A233 );
 a13559a <=( (not A232)  and  a13558a );
 a13563a <=( A302  and  A299 );
 a13564a <=( (not A298)  and  a13563a );
 a13565a <=( a13564a  and  a13559a );
 a13568a <=( A199  and  A169 );
 a13572a <=( (not A202)  and  (not A201) );
 a13573a <=( A200  and  a13572a );
 a13574a <=( a13573a  and  a13568a );
 a13578a <=( A236  and  A233 );
 a13579a <=( (not A232)  and  a13578a );
 a13583a <=( A269  and  A266 );
 a13584a <=( (not A265)  and  a13583a );
 a13585a <=( a13584a  and  a13579a );
 a13588a <=( A199  and  A169 );
 a13592a <=( (not A202)  and  (not A201) );
 a13593a <=( A200  and  a13592a );
 a13594a <=( a13593a  and  a13588a );
 a13598a <=( A236  and  A233 );
 a13599a <=( (not A232)  and  a13598a );
 a13603a <=( A269  and  (not A266) );
 a13604a <=( A265  and  a13603a );
 a13605a <=( a13604a  and  a13599a );
 a13608a <=( A199  and  A169 );
 a13612a <=( (not A202)  and  (not A201) );
 a13613a <=( A200  and  a13612a );
 a13614a <=( a13613a  and  a13608a );
 a13618a <=( A236  and  (not A233) );
 a13619a <=( A232  and  a13618a );
 a13623a <=( A302  and  (not A299) );
 a13624a <=( A298  and  a13623a );
 a13625a <=( a13624a  and  a13619a );
 a13628a <=( A199  and  A169 );
 a13632a <=( (not A202)  and  (not A201) );
 a13633a <=( A200  and  a13632a );
 a13634a <=( a13633a  and  a13628a );
 a13638a <=( A236  and  (not A233) );
 a13639a <=( A232  and  a13638a );
 a13643a <=( A302  and  A299 );
 a13644a <=( (not A298)  and  a13643a );
 a13645a <=( a13644a  and  a13639a );
 a13648a <=( A199  and  A169 );
 a13652a <=( (not A202)  and  (not A201) );
 a13653a <=( A200  and  a13652a );
 a13654a <=( a13653a  and  a13648a );
 a13658a <=( A236  and  (not A233) );
 a13659a <=( A232  and  a13658a );
 a13663a <=( A269  and  A266 );
 a13664a <=( (not A265)  and  a13663a );
 a13665a <=( a13664a  and  a13659a );
 a13668a <=( A199  and  A169 );
 a13672a <=( (not A202)  and  (not A201) );
 a13673a <=( A200  and  a13672a );
 a13674a <=( a13673a  and  a13668a );
 a13678a <=( A236  and  (not A233) );
 a13679a <=( A232  and  a13678a );
 a13683a <=( A269  and  (not A266) );
 a13684a <=( A265  and  a13683a );
 a13685a <=( a13684a  and  a13679a );
 a13689a <=( A199  and  A166 );
 a13690a <=( A168  and  a13689a );
 a13694a <=( (not A202)  and  (not A201) );
 a13695a <=( A200  and  a13694a );
 a13696a <=( a13695a  and  a13690a );
 a13700a <=( A236  and  A233 );
 a13701a <=( (not A232)  and  a13700a );
 a13705a <=( A302  and  (not A299) );
 a13706a <=( A298  and  a13705a );
 a13707a <=( a13706a  and  a13701a );
 a13711a <=( A199  and  A166 );
 a13712a <=( A168  and  a13711a );
 a13716a <=( (not A202)  and  (not A201) );
 a13717a <=( A200  and  a13716a );
 a13718a <=( a13717a  and  a13712a );
 a13722a <=( A236  and  A233 );
 a13723a <=( (not A232)  and  a13722a );
 a13727a <=( A302  and  A299 );
 a13728a <=( (not A298)  and  a13727a );
 a13729a <=( a13728a  and  a13723a );
 a13733a <=( A199  and  A166 );
 a13734a <=( A168  and  a13733a );
 a13738a <=( (not A202)  and  (not A201) );
 a13739a <=( A200  and  a13738a );
 a13740a <=( a13739a  and  a13734a );
 a13744a <=( A236  and  A233 );
 a13745a <=( (not A232)  and  a13744a );
 a13749a <=( A269  and  A266 );
 a13750a <=( (not A265)  and  a13749a );
 a13751a <=( a13750a  and  a13745a );
 a13755a <=( A199  and  A166 );
 a13756a <=( A168  and  a13755a );
 a13760a <=( (not A202)  and  (not A201) );
 a13761a <=( A200  and  a13760a );
 a13762a <=( a13761a  and  a13756a );
 a13766a <=( A236  and  A233 );
 a13767a <=( (not A232)  and  a13766a );
 a13771a <=( A269  and  (not A266) );
 a13772a <=( A265  and  a13771a );
 a13773a <=( a13772a  and  a13767a );
 a13777a <=( A199  and  A166 );
 a13778a <=( A168  and  a13777a );
 a13782a <=( (not A202)  and  (not A201) );
 a13783a <=( A200  and  a13782a );
 a13784a <=( a13783a  and  a13778a );
 a13788a <=( A236  and  (not A233) );
 a13789a <=( A232  and  a13788a );
 a13793a <=( A302  and  (not A299) );
 a13794a <=( A298  and  a13793a );
 a13795a <=( a13794a  and  a13789a );
 a13799a <=( A199  and  A166 );
 a13800a <=( A168  and  a13799a );
 a13804a <=( (not A202)  and  (not A201) );
 a13805a <=( A200  and  a13804a );
 a13806a <=( a13805a  and  a13800a );
 a13810a <=( A236  and  (not A233) );
 a13811a <=( A232  and  a13810a );
 a13815a <=( A302  and  A299 );
 a13816a <=( (not A298)  and  a13815a );
 a13817a <=( a13816a  and  a13811a );
 a13821a <=( A199  and  A166 );
 a13822a <=( A168  and  a13821a );
 a13826a <=( (not A202)  and  (not A201) );
 a13827a <=( A200  and  a13826a );
 a13828a <=( a13827a  and  a13822a );
 a13832a <=( A236  and  (not A233) );
 a13833a <=( A232  and  a13832a );
 a13837a <=( A269  and  A266 );
 a13838a <=( (not A265)  and  a13837a );
 a13839a <=( a13838a  and  a13833a );
 a13843a <=( A199  and  A166 );
 a13844a <=( A168  and  a13843a );
 a13848a <=( (not A202)  and  (not A201) );
 a13849a <=( A200  and  a13848a );
 a13850a <=( a13849a  and  a13844a );
 a13854a <=( A236  and  (not A233) );
 a13855a <=( A232  and  a13854a );
 a13859a <=( A269  and  (not A266) );
 a13860a <=( A265  and  a13859a );
 a13861a <=( a13860a  and  a13855a );
 a13865a <=( A199  and  A167 );
 a13866a <=( A168  and  a13865a );
 a13870a <=( (not A202)  and  (not A201) );
 a13871a <=( A200  and  a13870a );
 a13872a <=( a13871a  and  a13866a );
 a13876a <=( A236  and  A233 );
 a13877a <=( (not A232)  and  a13876a );
 a13881a <=( A302  and  (not A299) );
 a13882a <=( A298  and  a13881a );
 a13883a <=( a13882a  and  a13877a );
 a13887a <=( A199  and  A167 );
 a13888a <=( A168  and  a13887a );
 a13892a <=( (not A202)  and  (not A201) );
 a13893a <=( A200  and  a13892a );
 a13894a <=( a13893a  and  a13888a );
 a13898a <=( A236  and  A233 );
 a13899a <=( (not A232)  and  a13898a );
 a13903a <=( A302  and  A299 );
 a13904a <=( (not A298)  and  a13903a );
 a13905a <=( a13904a  and  a13899a );
 a13909a <=( A199  and  A167 );
 a13910a <=( A168  and  a13909a );
 a13914a <=( (not A202)  and  (not A201) );
 a13915a <=( A200  and  a13914a );
 a13916a <=( a13915a  and  a13910a );
 a13920a <=( A236  and  A233 );
 a13921a <=( (not A232)  and  a13920a );
 a13925a <=( A269  and  A266 );
 a13926a <=( (not A265)  and  a13925a );
 a13927a <=( a13926a  and  a13921a );
 a13931a <=( A199  and  A167 );
 a13932a <=( A168  and  a13931a );
 a13936a <=( (not A202)  and  (not A201) );
 a13937a <=( A200  and  a13936a );
 a13938a <=( a13937a  and  a13932a );
 a13942a <=( A236  and  A233 );
 a13943a <=( (not A232)  and  a13942a );
 a13947a <=( A269  and  (not A266) );
 a13948a <=( A265  and  a13947a );
 a13949a <=( a13948a  and  a13943a );
 a13953a <=( A199  and  A167 );
 a13954a <=( A168  and  a13953a );
 a13958a <=( (not A202)  and  (not A201) );
 a13959a <=( A200  and  a13958a );
 a13960a <=( a13959a  and  a13954a );
 a13964a <=( A236  and  (not A233) );
 a13965a <=( A232  and  a13964a );
 a13969a <=( A302  and  (not A299) );
 a13970a <=( A298  and  a13969a );
 a13971a <=( a13970a  and  a13965a );
 a13975a <=( A199  and  A167 );
 a13976a <=( A168  and  a13975a );
 a13980a <=( (not A202)  and  (not A201) );
 a13981a <=( A200  and  a13980a );
 a13982a <=( a13981a  and  a13976a );
 a13986a <=( A236  and  (not A233) );
 a13987a <=( A232  and  a13986a );
 a13991a <=( A302  and  A299 );
 a13992a <=( (not A298)  and  a13991a );
 a13993a <=( a13992a  and  a13987a );
 a13997a <=( A199  and  A167 );
 a13998a <=( A168  and  a13997a );
 a14002a <=( (not A202)  and  (not A201) );
 a14003a <=( A200  and  a14002a );
 a14004a <=( a14003a  and  a13998a );
 a14008a <=( A236  and  (not A233) );
 a14009a <=( A232  and  a14008a );
 a14013a <=( A269  and  A266 );
 a14014a <=( (not A265)  and  a14013a );
 a14015a <=( a14014a  and  a14009a );
 a14019a <=( A199  and  A167 );
 a14020a <=( A168  and  a14019a );
 a14024a <=( (not A202)  and  (not A201) );
 a14025a <=( A200  and  a14024a );
 a14026a <=( a14025a  and  a14020a );
 a14030a <=( A236  and  (not A233) );
 a14031a <=( A232  and  a14030a );
 a14035a <=( A269  and  (not A266) );
 a14036a <=( A265  and  a14035a );
 a14037a <=( a14036a  and  a14031a );
 a14041a <=( (not A166)  and  A167 );
 a14042a <=( A170  and  a14041a );
 a14046a <=( (not A203)  and  (not A202) );
 a14047a <=( (not A201)  and  a14046a );
 a14048a <=( a14047a  and  a14042a );
 a14052a <=( A236  and  A233 );
 a14053a <=( (not A232)  and  a14052a );
 a14057a <=( A302  and  (not A299) );
 a14058a <=( A298  and  a14057a );
 a14059a <=( a14058a  and  a14053a );
 a14063a <=( (not A166)  and  A167 );
 a14064a <=( A170  and  a14063a );
 a14068a <=( (not A203)  and  (not A202) );
 a14069a <=( (not A201)  and  a14068a );
 a14070a <=( a14069a  and  a14064a );
 a14074a <=( A236  and  A233 );
 a14075a <=( (not A232)  and  a14074a );
 a14079a <=( A302  and  A299 );
 a14080a <=( (not A298)  and  a14079a );
 a14081a <=( a14080a  and  a14075a );
 a14085a <=( (not A166)  and  A167 );
 a14086a <=( A170  and  a14085a );
 a14090a <=( (not A203)  and  (not A202) );
 a14091a <=( (not A201)  and  a14090a );
 a14092a <=( a14091a  and  a14086a );
 a14096a <=( A236  and  A233 );
 a14097a <=( (not A232)  and  a14096a );
 a14101a <=( A269  and  A266 );
 a14102a <=( (not A265)  and  a14101a );
 a14103a <=( a14102a  and  a14097a );
 a14107a <=( (not A166)  and  A167 );
 a14108a <=( A170  and  a14107a );
 a14112a <=( (not A203)  and  (not A202) );
 a14113a <=( (not A201)  and  a14112a );
 a14114a <=( a14113a  and  a14108a );
 a14118a <=( A236  and  A233 );
 a14119a <=( (not A232)  and  a14118a );
 a14123a <=( A269  and  (not A266) );
 a14124a <=( A265  and  a14123a );
 a14125a <=( a14124a  and  a14119a );
 a14129a <=( (not A166)  and  A167 );
 a14130a <=( A170  and  a14129a );
 a14134a <=( (not A203)  and  (not A202) );
 a14135a <=( (not A201)  and  a14134a );
 a14136a <=( a14135a  and  a14130a );
 a14140a <=( A236  and  (not A233) );
 a14141a <=( A232  and  a14140a );
 a14145a <=( A302  and  (not A299) );
 a14146a <=( A298  and  a14145a );
 a14147a <=( a14146a  and  a14141a );
 a14151a <=( (not A166)  and  A167 );
 a14152a <=( A170  and  a14151a );
 a14156a <=( (not A203)  and  (not A202) );
 a14157a <=( (not A201)  and  a14156a );
 a14158a <=( a14157a  and  a14152a );
 a14162a <=( A236  and  (not A233) );
 a14163a <=( A232  and  a14162a );
 a14167a <=( A302  and  A299 );
 a14168a <=( (not A298)  and  a14167a );
 a14169a <=( a14168a  and  a14163a );
 a14173a <=( (not A166)  and  A167 );
 a14174a <=( A170  and  a14173a );
 a14178a <=( (not A203)  and  (not A202) );
 a14179a <=( (not A201)  and  a14178a );
 a14180a <=( a14179a  and  a14174a );
 a14184a <=( A236  and  (not A233) );
 a14185a <=( A232  and  a14184a );
 a14189a <=( A269  and  A266 );
 a14190a <=( (not A265)  and  a14189a );
 a14191a <=( a14190a  and  a14185a );
 a14195a <=( (not A166)  and  A167 );
 a14196a <=( A170  and  a14195a );
 a14200a <=( (not A203)  and  (not A202) );
 a14201a <=( (not A201)  and  a14200a );
 a14202a <=( a14201a  and  a14196a );
 a14206a <=( A236  and  (not A233) );
 a14207a <=( A232  and  a14206a );
 a14211a <=( A269  and  (not A266) );
 a14212a <=( A265  and  a14211a );
 a14213a <=( a14212a  and  a14207a );
 a14217a <=( (not A166)  and  A167 );
 a14218a <=( A170  and  a14217a );
 a14222a <=( (not A201)  and  A200 );
 a14223a <=( A199  and  a14222a );
 a14224a <=( a14223a  and  a14218a );
 a14228a <=( A234  and  A232 );
 a14229a <=( (not A202)  and  a14228a );
 a14233a <=( A302  and  (not A299) );
 a14234a <=( A298  and  a14233a );
 a14235a <=( a14234a  and  a14229a );
 a14239a <=( (not A166)  and  A167 );
 a14240a <=( A170  and  a14239a );
 a14244a <=( (not A201)  and  A200 );
 a14245a <=( A199  and  a14244a );
 a14246a <=( a14245a  and  a14240a );
 a14250a <=( A234  and  A232 );
 a14251a <=( (not A202)  and  a14250a );
 a14255a <=( A302  and  A299 );
 a14256a <=( (not A298)  and  a14255a );
 a14257a <=( a14256a  and  a14251a );
 a14261a <=( (not A166)  and  A167 );
 a14262a <=( A170  and  a14261a );
 a14266a <=( (not A201)  and  A200 );
 a14267a <=( A199  and  a14266a );
 a14268a <=( a14267a  and  a14262a );
 a14272a <=( A234  and  A232 );
 a14273a <=( (not A202)  and  a14272a );
 a14277a <=( A269  and  A266 );
 a14278a <=( (not A265)  and  a14277a );
 a14279a <=( a14278a  and  a14273a );
 a14283a <=( (not A166)  and  A167 );
 a14284a <=( A170  and  a14283a );
 a14288a <=( (not A201)  and  A200 );
 a14289a <=( A199  and  a14288a );
 a14290a <=( a14289a  and  a14284a );
 a14294a <=( A234  and  A232 );
 a14295a <=( (not A202)  and  a14294a );
 a14299a <=( A269  and  (not A266) );
 a14300a <=( A265  and  a14299a );
 a14301a <=( a14300a  and  a14295a );
 a14305a <=( (not A166)  and  A167 );
 a14306a <=( A170  and  a14305a );
 a14310a <=( (not A201)  and  A200 );
 a14311a <=( A199  and  a14310a );
 a14312a <=( a14311a  and  a14306a );
 a14316a <=( A234  and  A233 );
 a14317a <=( (not A202)  and  a14316a );
 a14321a <=( A302  and  (not A299) );
 a14322a <=( A298  and  a14321a );
 a14323a <=( a14322a  and  a14317a );
 a14327a <=( (not A166)  and  A167 );
 a14328a <=( A170  and  a14327a );
 a14332a <=( (not A201)  and  A200 );
 a14333a <=( A199  and  a14332a );
 a14334a <=( a14333a  and  a14328a );
 a14338a <=( A234  and  A233 );
 a14339a <=( (not A202)  and  a14338a );
 a14343a <=( A302  and  A299 );
 a14344a <=( (not A298)  and  a14343a );
 a14345a <=( a14344a  and  a14339a );
 a14349a <=( (not A166)  and  A167 );
 a14350a <=( A170  and  a14349a );
 a14354a <=( (not A201)  and  A200 );
 a14355a <=( A199  and  a14354a );
 a14356a <=( a14355a  and  a14350a );
 a14360a <=( A234  and  A233 );
 a14361a <=( (not A202)  and  a14360a );
 a14365a <=( A269  and  A266 );
 a14366a <=( (not A265)  and  a14365a );
 a14367a <=( a14366a  and  a14361a );
 a14371a <=( (not A166)  and  A167 );
 a14372a <=( A170  and  a14371a );
 a14376a <=( (not A201)  and  A200 );
 a14377a <=( A199  and  a14376a );
 a14378a <=( a14377a  and  a14372a );
 a14382a <=( A234  and  A233 );
 a14383a <=( (not A202)  and  a14382a );
 a14387a <=( A269  and  (not A266) );
 a14388a <=( A265  and  a14387a );
 a14389a <=( a14388a  and  a14383a );
 a14393a <=( (not A166)  and  A167 );
 a14394a <=( A170  and  a14393a );
 a14398a <=( (not A201)  and  A200 );
 a14399a <=( A199  and  a14398a );
 a14400a <=( a14399a  and  a14394a );
 a14404a <=( A233  and  (not A232) );
 a14405a <=( (not A202)  and  a14404a );
 a14409a <=( A300  and  A299 );
 a14410a <=( A236  and  a14409a );
 a14411a <=( a14410a  and  a14405a );
 a14415a <=( (not A166)  and  A167 );
 a14416a <=( A170  and  a14415a );
 a14420a <=( (not A201)  and  A200 );
 a14421a <=( A199  and  a14420a );
 a14422a <=( a14421a  and  a14416a );
 a14426a <=( A233  and  (not A232) );
 a14427a <=( (not A202)  and  a14426a );
 a14431a <=( A300  and  A298 );
 a14432a <=( A236  and  a14431a );
 a14433a <=( a14432a  and  a14427a );
 a14437a <=( (not A166)  and  A167 );
 a14438a <=( A170  and  a14437a );
 a14442a <=( (not A201)  and  A200 );
 a14443a <=( A199  and  a14442a );
 a14444a <=( a14443a  and  a14438a );
 a14448a <=( A233  and  (not A232) );
 a14449a <=( (not A202)  and  a14448a );
 a14453a <=( A267  and  A265 );
 a14454a <=( A236  and  a14453a );
 a14455a <=( a14454a  and  a14449a );
 a14459a <=( (not A166)  and  A167 );
 a14460a <=( A170  and  a14459a );
 a14464a <=( (not A201)  and  A200 );
 a14465a <=( A199  and  a14464a );
 a14466a <=( a14465a  and  a14460a );
 a14470a <=( A233  and  (not A232) );
 a14471a <=( (not A202)  and  a14470a );
 a14475a <=( A267  and  A266 );
 a14476a <=( A236  and  a14475a );
 a14477a <=( a14476a  and  a14471a );
 a14481a <=( (not A166)  and  A167 );
 a14482a <=( A170  and  a14481a );
 a14486a <=( (not A201)  and  A200 );
 a14487a <=( A199  and  a14486a );
 a14488a <=( a14487a  and  a14482a );
 a14492a <=( (not A233)  and  A232 );
 a14493a <=( (not A202)  and  a14492a );
 a14497a <=( A300  and  A299 );
 a14498a <=( A236  and  a14497a );
 a14499a <=( a14498a  and  a14493a );
 a14503a <=( (not A166)  and  A167 );
 a14504a <=( A170  and  a14503a );
 a14508a <=( (not A201)  and  A200 );
 a14509a <=( A199  and  a14508a );
 a14510a <=( a14509a  and  a14504a );
 a14514a <=( (not A233)  and  A232 );
 a14515a <=( (not A202)  and  a14514a );
 a14519a <=( A300  and  A298 );
 a14520a <=( A236  and  a14519a );
 a14521a <=( a14520a  and  a14515a );
 a14525a <=( (not A166)  and  A167 );
 a14526a <=( A170  and  a14525a );
 a14530a <=( (not A201)  and  A200 );
 a14531a <=( A199  and  a14530a );
 a14532a <=( a14531a  and  a14526a );
 a14536a <=( (not A233)  and  A232 );
 a14537a <=( (not A202)  and  a14536a );
 a14541a <=( A267  and  A265 );
 a14542a <=( A236  and  a14541a );
 a14543a <=( a14542a  and  a14537a );
 a14547a <=( (not A166)  and  A167 );
 a14548a <=( A170  and  a14547a );
 a14552a <=( (not A201)  and  A200 );
 a14553a <=( A199  and  a14552a );
 a14554a <=( a14553a  and  a14548a );
 a14558a <=( (not A233)  and  A232 );
 a14559a <=( (not A202)  and  a14558a );
 a14563a <=( A267  and  A266 );
 a14564a <=( A236  and  a14563a );
 a14565a <=( a14564a  and  a14559a );
 a14569a <=( (not A166)  and  A167 );
 a14570a <=( A170  and  a14569a );
 a14574a <=( (not A202)  and  (not A200) );
 a14575a <=( (not A199)  and  a14574a );
 a14576a <=( a14575a  and  a14570a );
 a14580a <=( A236  and  A233 );
 a14581a <=( (not A232)  and  a14580a );
 a14585a <=( A302  and  (not A299) );
 a14586a <=( A298  and  a14585a );
 a14587a <=( a14586a  and  a14581a );
 a14591a <=( (not A166)  and  A167 );
 a14592a <=( A170  and  a14591a );
 a14596a <=( (not A202)  and  (not A200) );
 a14597a <=( (not A199)  and  a14596a );
 a14598a <=( a14597a  and  a14592a );
 a14602a <=( A236  and  A233 );
 a14603a <=( (not A232)  and  a14602a );
 a14607a <=( A302  and  A299 );
 a14608a <=( (not A298)  and  a14607a );
 a14609a <=( a14608a  and  a14603a );
 a14613a <=( (not A166)  and  A167 );
 a14614a <=( A170  and  a14613a );
 a14618a <=( (not A202)  and  (not A200) );
 a14619a <=( (not A199)  and  a14618a );
 a14620a <=( a14619a  and  a14614a );
 a14624a <=( A236  and  A233 );
 a14625a <=( (not A232)  and  a14624a );
 a14629a <=( A269  and  A266 );
 a14630a <=( (not A265)  and  a14629a );
 a14631a <=( a14630a  and  a14625a );
 a14635a <=( (not A166)  and  A167 );
 a14636a <=( A170  and  a14635a );
 a14640a <=( (not A202)  and  (not A200) );
 a14641a <=( (not A199)  and  a14640a );
 a14642a <=( a14641a  and  a14636a );
 a14646a <=( A236  and  A233 );
 a14647a <=( (not A232)  and  a14646a );
 a14651a <=( A269  and  (not A266) );
 a14652a <=( A265  and  a14651a );
 a14653a <=( a14652a  and  a14647a );
 a14657a <=( (not A166)  and  A167 );
 a14658a <=( A170  and  a14657a );
 a14662a <=( (not A202)  and  (not A200) );
 a14663a <=( (not A199)  and  a14662a );
 a14664a <=( a14663a  and  a14658a );
 a14668a <=( A236  and  (not A233) );
 a14669a <=( A232  and  a14668a );
 a14673a <=( A302  and  (not A299) );
 a14674a <=( A298  and  a14673a );
 a14675a <=( a14674a  and  a14669a );
 a14679a <=( (not A166)  and  A167 );
 a14680a <=( A170  and  a14679a );
 a14684a <=( (not A202)  and  (not A200) );
 a14685a <=( (not A199)  and  a14684a );
 a14686a <=( a14685a  and  a14680a );
 a14690a <=( A236  and  (not A233) );
 a14691a <=( A232  and  a14690a );
 a14695a <=( A302  and  A299 );
 a14696a <=( (not A298)  and  a14695a );
 a14697a <=( a14696a  and  a14691a );
 a14701a <=( (not A166)  and  A167 );
 a14702a <=( A170  and  a14701a );
 a14706a <=( (not A202)  and  (not A200) );
 a14707a <=( (not A199)  and  a14706a );
 a14708a <=( a14707a  and  a14702a );
 a14712a <=( A236  and  (not A233) );
 a14713a <=( A232  and  a14712a );
 a14717a <=( A269  and  A266 );
 a14718a <=( (not A265)  and  a14717a );
 a14719a <=( a14718a  and  a14713a );
 a14723a <=( (not A166)  and  A167 );
 a14724a <=( A170  and  a14723a );
 a14728a <=( (not A202)  and  (not A200) );
 a14729a <=( (not A199)  and  a14728a );
 a14730a <=( a14729a  and  a14724a );
 a14734a <=( A236  and  (not A233) );
 a14735a <=( A232  and  a14734a );
 a14739a <=( A269  and  (not A266) );
 a14740a <=( A265  and  a14739a );
 a14741a <=( a14740a  and  a14735a );
 a14745a <=( A166  and  (not A167) );
 a14746a <=( A170  and  a14745a );
 a14750a <=( (not A203)  and  (not A202) );
 a14751a <=( (not A201)  and  a14750a );
 a14752a <=( a14751a  and  a14746a );
 a14756a <=( A236  and  A233 );
 a14757a <=( (not A232)  and  a14756a );
 a14761a <=( A302  and  (not A299) );
 a14762a <=( A298  and  a14761a );
 a14763a <=( a14762a  and  a14757a );
 a14767a <=( A166  and  (not A167) );
 a14768a <=( A170  and  a14767a );
 a14772a <=( (not A203)  and  (not A202) );
 a14773a <=( (not A201)  and  a14772a );
 a14774a <=( a14773a  and  a14768a );
 a14778a <=( A236  and  A233 );
 a14779a <=( (not A232)  and  a14778a );
 a14783a <=( A302  and  A299 );
 a14784a <=( (not A298)  and  a14783a );
 a14785a <=( a14784a  and  a14779a );
 a14789a <=( A166  and  (not A167) );
 a14790a <=( A170  and  a14789a );
 a14794a <=( (not A203)  and  (not A202) );
 a14795a <=( (not A201)  and  a14794a );
 a14796a <=( a14795a  and  a14790a );
 a14800a <=( A236  and  A233 );
 a14801a <=( (not A232)  and  a14800a );
 a14805a <=( A269  and  A266 );
 a14806a <=( (not A265)  and  a14805a );
 a14807a <=( a14806a  and  a14801a );
 a14811a <=( A166  and  (not A167) );
 a14812a <=( A170  and  a14811a );
 a14816a <=( (not A203)  and  (not A202) );
 a14817a <=( (not A201)  and  a14816a );
 a14818a <=( a14817a  and  a14812a );
 a14822a <=( A236  and  A233 );
 a14823a <=( (not A232)  and  a14822a );
 a14827a <=( A269  and  (not A266) );
 a14828a <=( A265  and  a14827a );
 a14829a <=( a14828a  and  a14823a );
 a14833a <=( A166  and  (not A167) );
 a14834a <=( A170  and  a14833a );
 a14838a <=( (not A203)  and  (not A202) );
 a14839a <=( (not A201)  and  a14838a );
 a14840a <=( a14839a  and  a14834a );
 a14844a <=( A236  and  (not A233) );
 a14845a <=( A232  and  a14844a );
 a14849a <=( A302  and  (not A299) );
 a14850a <=( A298  and  a14849a );
 a14851a <=( a14850a  and  a14845a );
 a14855a <=( A166  and  (not A167) );
 a14856a <=( A170  and  a14855a );
 a14860a <=( (not A203)  and  (not A202) );
 a14861a <=( (not A201)  and  a14860a );
 a14862a <=( a14861a  and  a14856a );
 a14866a <=( A236  and  (not A233) );
 a14867a <=( A232  and  a14866a );
 a14871a <=( A302  and  A299 );
 a14872a <=( (not A298)  and  a14871a );
 a14873a <=( a14872a  and  a14867a );
 a14877a <=( A166  and  (not A167) );
 a14878a <=( A170  and  a14877a );
 a14882a <=( (not A203)  and  (not A202) );
 a14883a <=( (not A201)  and  a14882a );
 a14884a <=( a14883a  and  a14878a );
 a14888a <=( A236  and  (not A233) );
 a14889a <=( A232  and  a14888a );
 a14893a <=( A269  and  A266 );
 a14894a <=( (not A265)  and  a14893a );
 a14895a <=( a14894a  and  a14889a );
 a14899a <=( A166  and  (not A167) );
 a14900a <=( A170  and  a14899a );
 a14904a <=( (not A203)  and  (not A202) );
 a14905a <=( (not A201)  and  a14904a );
 a14906a <=( a14905a  and  a14900a );
 a14910a <=( A236  and  (not A233) );
 a14911a <=( A232  and  a14910a );
 a14915a <=( A269  and  (not A266) );
 a14916a <=( A265  and  a14915a );
 a14917a <=( a14916a  and  a14911a );
 a14921a <=( A166  and  (not A167) );
 a14922a <=( A170  and  a14921a );
 a14926a <=( (not A201)  and  A200 );
 a14927a <=( A199  and  a14926a );
 a14928a <=( a14927a  and  a14922a );
 a14932a <=( A234  and  A232 );
 a14933a <=( (not A202)  and  a14932a );
 a14937a <=( A302  and  (not A299) );
 a14938a <=( A298  and  a14937a );
 a14939a <=( a14938a  and  a14933a );
 a14943a <=( A166  and  (not A167) );
 a14944a <=( A170  and  a14943a );
 a14948a <=( (not A201)  and  A200 );
 a14949a <=( A199  and  a14948a );
 a14950a <=( a14949a  and  a14944a );
 a14954a <=( A234  and  A232 );
 a14955a <=( (not A202)  and  a14954a );
 a14959a <=( A302  and  A299 );
 a14960a <=( (not A298)  and  a14959a );
 a14961a <=( a14960a  and  a14955a );
 a14965a <=( A166  and  (not A167) );
 a14966a <=( A170  and  a14965a );
 a14970a <=( (not A201)  and  A200 );
 a14971a <=( A199  and  a14970a );
 a14972a <=( a14971a  and  a14966a );
 a14976a <=( A234  and  A232 );
 a14977a <=( (not A202)  and  a14976a );
 a14981a <=( A269  and  A266 );
 a14982a <=( (not A265)  and  a14981a );
 a14983a <=( a14982a  and  a14977a );
 a14987a <=( A166  and  (not A167) );
 a14988a <=( A170  and  a14987a );
 a14992a <=( (not A201)  and  A200 );
 a14993a <=( A199  and  a14992a );
 a14994a <=( a14993a  and  a14988a );
 a14998a <=( A234  and  A232 );
 a14999a <=( (not A202)  and  a14998a );
 a15003a <=( A269  and  (not A266) );
 a15004a <=( A265  and  a15003a );
 a15005a <=( a15004a  and  a14999a );
 a15009a <=( A166  and  (not A167) );
 a15010a <=( A170  and  a15009a );
 a15014a <=( (not A201)  and  A200 );
 a15015a <=( A199  and  a15014a );
 a15016a <=( a15015a  and  a15010a );
 a15020a <=( A234  and  A233 );
 a15021a <=( (not A202)  and  a15020a );
 a15025a <=( A302  and  (not A299) );
 a15026a <=( A298  and  a15025a );
 a15027a <=( a15026a  and  a15021a );
 a15031a <=( A166  and  (not A167) );
 a15032a <=( A170  and  a15031a );
 a15036a <=( (not A201)  and  A200 );
 a15037a <=( A199  and  a15036a );
 a15038a <=( a15037a  and  a15032a );
 a15042a <=( A234  and  A233 );
 a15043a <=( (not A202)  and  a15042a );
 a15047a <=( A302  and  A299 );
 a15048a <=( (not A298)  and  a15047a );
 a15049a <=( a15048a  and  a15043a );
 a15053a <=( A166  and  (not A167) );
 a15054a <=( A170  and  a15053a );
 a15058a <=( (not A201)  and  A200 );
 a15059a <=( A199  and  a15058a );
 a15060a <=( a15059a  and  a15054a );
 a15064a <=( A234  and  A233 );
 a15065a <=( (not A202)  and  a15064a );
 a15069a <=( A269  and  A266 );
 a15070a <=( (not A265)  and  a15069a );
 a15071a <=( a15070a  and  a15065a );
 a15075a <=( A166  and  (not A167) );
 a15076a <=( A170  and  a15075a );
 a15080a <=( (not A201)  and  A200 );
 a15081a <=( A199  and  a15080a );
 a15082a <=( a15081a  and  a15076a );
 a15086a <=( A234  and  A233 );
 a15087a <=( (not A202)  and  a15086a );
 a15091a <=( A269  and  (not A266) );
 a15092a <=( A265  and  a15091a );
 a15093a <=( a15092a  and  a15087a );
 a15097a <=( A166  and  (not A167) );
 a15098a <=( A170  and  a15097a );
 a15102a <=( (not A201)  and  A200 );
 a15103a <=( A199  and  a15102a );
 a15104a <=( a15103a  and  a15098a );
 a15108a <=( A233  and  (not A232) );
 a15109a <=( (not A202)  and  a15108a );
 a15113a <=( A300  and  A299 );
 a15114a <=( A236  and  a15113a );
 a15115a <=( a15114a  and  a15109a );
 a15119a <=( A166  and  (not A167) );
 a15120a <=( A170  and  a15119a );
 a15124a <=( (not A201)  and  A200 );
 a15125a <=( A199  and  a15124a );
 a15126a <=( a15125a  and  a15120a );
 a15130a <=( A233  and  (not A232) );
 a15131a <=( (not A202)  and  a15130a );
 a15135a <=( A300  and  A298 );
 a15136a <=( A236  and  a15135a );
 a15137a <=( a15136a  and  a15131a );
 a15141a <=( A166  and  (not A167) );
 a15142a <=( A170  and  a15141a );
 a15146a <=( (not A201)  and  A200 );
 a15147a <=( A199  and  a15146a );
 a15148a <=( a15147a  and  a15142a );
 a15152a <=( A233  and  (not A232) );
 a15153a <=( (not A202)  and  a15152a );
 a15157a <=( A267  and  A265 );
 a15158a <=( A236  and  a15157a );
 a15159a <=( a15158a  and  a15153a );
 a15163a <=( A166  and  (not A167) );
 a15164a <=( A170  and  a15163a );
 a15168a <=( (not A201)  and  A200 );
 a15169a <=( A199  and  a15168a );
 a15170a <=( a15169a  and  a15164a );
 a15174a <=( A233  and  (not A232) );
 a15175a <=( (not A202)  and  a15174a );
 a15179a <=( A267  and  A266 );
 a15180a <=( A236  and  a15179a );
 a15181a <=( a15180a  and  a15175a );
 a15185a <=( A166  and  (not A167) );
 a15186a <=( A170  and  a15185a );
 a15190a <=( (not A201)  and  A200 );
 a15191a <=( A199  and  a15190a );
 a15192a <=( a15191a  and  a15186a );
 a15196a <=( (not A233)  and  A232 );
 a15197a <=( (not A202)  and  a15196a );
 a15201a <=( A300  and  A299 );
 a15202a <=( A236  and  a15201a );
 a15203a <=( a15202a  and  a15197a );
 a15207a <=( A166  and  (not A167) );
 a15208a <=( A170  and  a15207a );
 a15212a <=( (not A201)  and  A200 );
 a15213a <=( A199  and  a15212a );
 a15214a <=( a15213a  and  a15208a );
 a15218a <=( (not A233)  and  A232 );
 a15219a <=( (not A202)  and  a15218a );
 a15223a <=( A300  and  A298 );
 a15224a <=( A236  and  a15223a );
 a15225a <=( a15224a  and  a15219a );
 a15229a <=( A166  and  (not A167) );
 a15230a <=( A170  and  a15229a );
 a15234a <=( (not A201)  and  A200 );
 a15235a <=( A199  and  a15234a );
 a15236a <=( a15235a  and  a15230a );
 a15240a <=( (not A233)  and  A232 );
 a15241a <=( (not A202)  and  a15240a );
 a15245a <=( A267  and  A265 );
 a15246a <=( A236  and  a15245a );
 a15247a <=( a15246a  and  a15241a );
 a15251a <=( A166  and  (not A167) );
 a15252a <=( A170  and  a15251a );
 a15256a <=( (not A201)  and  A200 );
 a15257a <=( A199  and  a15256a );
 a15258a <=( a15257a  and  a15252a );
 a15262a <=( (not A233)  and  A232 );
 a15263a <=( (not A202)  and  a15262a );
 a15267a <=( A267  and  A266 );
 a15268a <=( A236  and  a15267a );
 a15269a <=( a15268a  and  a15263a );
 a15273a <=( A166  and  (not A167) );
 a15274a <=( A170  and  a15273a );
 a15278a <=( (not A202)  and  (not A200) );
 a15279a <=( (not A199)  and  a15278a );
 a15280a <=( a15279a  and  a15274a );
 a15284a <=( A236  and  A233 );
 a15285a <=( (not A232)  and  a15284a );
 a15289a <=( A302  and  (not A299) );
 a15290a <=( A298  and  a15289a );
 a15291a <=( a15290a  and  a15285a );
 a15295a <=( A166  and  (not A167) );
 a15296a <=( A170  and  a15295a );
 a15300a <=( (not A202)  and  (not A200) );
 a15301a <=( (not A199)  and  a15300a );
 a15302a <=( a15301a  and  a15296a );
 a15306a <=( A236  and  A233 );
 a15307a <=( (not A232)  and  a15306a );
 a15311a <=( A302  and  A299 );
 a15312a <=( (not A298)  and  a15311a );
 a15313a <=( a15312a  and  a15307a );
 a15317a <=( A166  and  (not A167) );
 a15318a <=( A170  and  a15317a );
 a15322a <=( (not A202)  and  (not A200) );
 a15323a <=( (not A199)  and  a15322a );
 a15324a <=( a15323a  and  a15318a );
 a15328a <=( A236  and  A233 );
 a15329a <=( (not A232)  and  a15328a );
 a15333a <=( A269  and  A266 );
 a15334a <=( (not A265)  and  a15333a );
 a15335a <=( a15334a  and  a15329a );
 a15339a <=( A166  and  (not A167) );
 a15340a <=( A170  and  a15339a );
 a15344a <=( (not A202)  and  (not A200) );
 a15345a <=( (not A199)  and  a15344a );
 a15346a <=( a15345a  and  a15340a );
 a15350a <=( A236  and  A233 );
 a15351a <=( (not A232)  and  a15350a );
 a15355a <=( A269  and  (not A266) );
 a15356a <=( A265  and  a15355a );
 a15357a <=( a15356a  and  a15351a );
 a15361a <=( A166  and  (not A167) );
 a15362a <=( A170  and  a15361a );
 a15366a <=( (not A202)  and  (not A200) );
 a15367a <=( (not A199)  and  a15366a );
 a15368a <=( a15367a  and  a15362a );
 a15372a <=( A236  and  (not A233) );
 a15373a <=( A232  and  a15372a );
 a15377a <=( A302  and  (not A299) );
 a15378a <=( A298  and  a15377a );
 a15379a <=( a15378a  and  a15373a );
 a15383a <=( A166  and  (not A167) );
 a15384a <=( A170  and  a15383a );
 a15388a <=( (not A202)  and  (not A200) );
 a15389a <=( (not A199)  and  a15388a );
 a15390a <=( a15389a  and  a15384a );
 a15394a <=( A236  and  (not A233) );
 a15395a <=( A232  and  a15394a );
 a15399a <=( A302  and  A299 );
 a15400a <=( (not A298)  and  a15399a );
 a15401a <=( a15400a  and  a15395a );
 a15405a <=( A166  and  (not A167) );
 a15406a <=( A170  and  a15405a );
 a15410a <=( (not A202)  and  (not A200) );
 a15411a <=( (not A199)  and  a15410a );
 a15412a <=( a15411a  and  a15406a );
 a15416a <=( A236  and  (not A233) );
 a15417a <=( A232  and  a15416a );
 a15421a <=( A269  and  A266 );
 a15422a <=( (not A265)  and  a15421a );
 a15423a <=( a15422a  and  a15417a );
 a15427a <=( A166  and  (not A167) );
 a15428a <=( A170  and  a15427a );
 a15432a <=( (not A202)  and  (not A200) );
 a15433a <=( (not A199)  and  a15432a );
 a15434a <=( a15433a  and  a15428a );
 a15438a <=( A236  and  (not A233) );
 a15439a <=( A232  and  a15438a );
 a15443a <=( A269  and  (not A266) );
 a15444a <=( A265  and  a15443a );
 a15445a <=( a15444a  and  a15439a );
 a15449a <=( (not A166)  and  A167 );
 a15450a <=( A170  and  a15449a );
 a15454a <=( (not A201)  and  A200 );
 a15455a <=( A199  and  a15454a );
 a15456a <=( a15455a  and  a15450a );
 a15460a <=( A233  and  (not A232) );
 a15461a <=( (not A202)  and  a15460a );
 a15464a <=( A298  and  A236 );
 a15467a <=( A302  and  (not A299) );
 a15468a <=( a15467a  and  a15464a );
 a15469a <=( a15468a  and  a15461a );
 a15473a <=( (not A166)  and  A167 );
 a15474a <=( A170  and  a15473a );
 a15478a <=( (not A201)  and  A200 );
 a15479a <=( A199  and  a15478a );
 a15480a <=( a15479a  and  a15474a );
 a15484a <=( A233  and  (not A232) );
 a15485a <=( (not A202)  and  a15484a );
 a15488a <=( (not A298)  and  A236 );
 a15491a <=( A302  and  A299 );
 a15492a <=( a15491a  and  a15488a );
 a15493a <=( a15492a  and  a15485a );
 a15497a <=( (not A166)  and  A167 );
 a15498a <=( A170  and  a15497a );
 a15502a <=( (not A201)  and  A200 );
 a15503a <=( A199  and  a15502a );
 a15504a <=( a15503a  and  a15498a );
 a15508a <=( A233  and  (not A232) );
 a15509a <=( (not A202)  and  a15508a );
 a15512a <=( (not A265)  and  A236 );
 a15515a <=( A269  and  A266 );
 a15516a <=( a15515a  and  a15512a );
 a15517a <=( a15516a  and  a15509a );
 a15521a <=( (not A166)  and  A167 );
 a15522a <=( A170  and  a15521a );
 a15526a <=( (not A201)  and  A200 );
 a15527a <=( A199  and  a15526a );
 a15528a <=( a15527a  and  a15522a );
 a15532a <=( A233  and  (not A232) );
 a15533a <=( (not A202)  and  a15532a );
 a15536a <=( A265  and  A236 );
 a15539a <=( A269  and  (not A266) );
 a15540a <=( a15539a  and  a15536a );
 a15541a <=( a15540a  and  a15533a );
 a15545a <=( (not A166)  and  A167 );
 a15546a <=( A170  and  a15545a );
 a15550a <=( (not A201)  and  A200 );
 a15551a <=( A199  and  a15550a );
 a15552a <=( a15551a  and  a15546a );
 a15556a <=( (not A233)  and  A232 );
 a15557a <=( (not A202)  and  a15556a );
 a15560a <=( A298  and  A236 );
 a15563a <=( A302  and  (not A299) );
 a15564a <=( a15563a  and  a15560a );
 a15565a <=( a15564a  and  a15557a );
 a15569a <=( (not A166)  and  A167 );
 a15570a <=( A170  and  a15569a );
 a15574a <=( (not A201)  and  A200 );
 a15575a <=( A199  and  a15574a );
 a15576a <=( a15575a  and  a15570a );
 a15580a <=( (not A233)  and  A232 );
 a15581a <=( (not A202)  and  a15580a );
 a15584a <=( (not A298)  and  A236 );
 a15587a <=( A302  and  A299 );
 a15588a <=( a15587a  and  a15584a );
 a15589a <=( a15588a  and  a15581a );
 a15593a <=( (not A166)  and  A167 );
 a15594a <=( A170  and  a15593a );
 a15598a <=( (not A201)  and  A200 );
 a15599a <=( A199  and  a15598a );
 a15600a <=( a15599a  and  a15594a );
 a15604a <=( (not A233)  and  A232 );
 a15605a <=( (not A202)  and  a15604a );
 a15608a <=( (not A265)  and  A236 );
 a15611a <=( A269  and  A266 );
 a15612a <=( a15611a  and  a15608a );
 a15613a <=( a15612a  and  a15605a );
 a15617a <=( (not A166)  and  A167 );
 a15618a <=( A170  and  a15617a );
 a15622a <=( (not A201)  and  A200 );
 a15623a <=( A199  and  a15622a );
 a15624a <=( a15623a  and  a15618a );
 a15628a <=( (not A233)  and  A232 );
 a15629a <=( (not A202)  and  a15628a );
 a15632a <=( A265  and  A236 );
 a15635a <=( A269  and  (not A266) );
 a15636a <=( a15635a  and  a15632a );
 a15637a <=( a15636a  and  a15629a );
 a15641a <=( A166  and  (not A167) );
 a15642a <=( A170  and  a15641a );
 a15646a <=( (not A201)  and  A200 );
 a15647a <=( A199  and  a15646a );
 a15648a <=( a15647a  and  a15642a );
 a15652a <=( A233  and  (not A232) );
 a15653a <=( (not A202)  and  a15652a );
 a15656a <=( A298  and  A236 );
 a15659a <=( A302  and  (not A299) );
 a15660a <=( a15659a  and  a15656a );
 a15661a <=( a15660a  and  a15653a );
 a15665a <=( A166  and  (not A167) );
 a15666a <=( A170  and  a15665a );
 a15670a <=( (not A201)  and  A200 );
 a15671a <=( A199  and  a15670a );
 a15672a <=( a15671a  and  a15666a );
 a15676a <=( A233  and  (not A232) );
 a15677a <=( (not A202)  and  a15676a );
 a15680a <=( (not A298)  and  A236 );
 a15683a <=( A302  and  A299 );
 a15684a <=( a15683a  and  a15680a );
 a15685a <=( a15684a  and  a15677a );
 a15689a <=( A166  and  (not A167) );
 a15690a <=( A170  and  a15689a );
 a15694a <=( (not A201)  and  A200 );
 a15695a <=( A199  and  a15694a );
 a15696a <=( a15695a  and  a15690a );
 a15700a <=( A233  and  (not A232) );
 a15701a <=( (not A202)  and  a15700a );
 a15704a <=( (not A265)  and  A236 );
 a15707a <=( A269  and  A266 );
 a15708a <=( a15707a  and  a15704a );
 a15709a <=( a15708a  and  a15701a );
 a15713a <=( A166  and  (not A167) );
 a15714a <=( A170  and  a15713a );
 a15718a <=( (not A201)  and  A200 );
 a15719a <=( A199  and  a15718a );
 a15720a <=( a15719a  and  a15714a );
 a15724a <=( A233  and  (not A232) );
 a15725a <=( (not A202)  and  a15724a );
 a15728a <=( A265  and  A236 );
 a15731a <=( A269  and  (not A266) );
 a15732a <=( a15731a  and  a15728a );
 a15733a <=( a15732a  and  a15725a );
 a15737a <=( A166  and  (not A167) );
 a15738a <=( A170  and  a15737a );
 a15742a <=( (not A201)  and  A200 );
 a15743a <=( A199  and  a15742a );
 a15744a <=( a15743a  and  a15738a );
 a15748a <=( (not A233)  and  A232 );
 a15749a <=( (not A202)  and  a15748a );
 a15752a <=( A298  and  A236 );
 a15755a <=( A302  and  (not A299) );
 a15756a <=( a15755a  and  a15752a );
 a15757a <=( a15756a  and  a15749a );
 a15761a <=( A166  and  (not A167) );
 a15762a <=( A170  and  a15761a );
 a15766a <=( (not A201)  and  A200 );
 a15767a <=( A199  and  a15766a );
 a15768a <=( a15767a  and  a15762a );
 a15772a <=( (not A233)  and  A232 );
 a15773a <=( (not A202)  and  a15772a );
 a15776a <=( (not A298)  and  A236 );
 a15779a <=( A302  and  A299 );
 a15780a <=( a15779a  and  a15776a );
 a15781a <=( a15780a  and  a15773a );
 a15785a <=( A166  and  (not A167) );
 a15786a <=( A170  and  a15785a );
 a15790a <=( (not A201)  and  A200 );
 a15791a <=( A199  and  a15790a );
 a15792a <=( a15791a  and  a15786a );
 a15796a <=( (not A233)  and  A232 );
 a15797a <=( (not A202)  and  a15796a );
 a15800a <=( (not A265)  and  A236 );
 a15803a <=( A269  and  A266 );
 a15804a <=( a15803a  and  a15800a );
 a15805a <=( a15804a  and  a15797a );
 a15809a <=( A166  and  (not A167) );
 a15810a <=( A170  and  a15809a );
 a15814a <=( (not A201)  and  A200 );
 a15815a <=( A199  and  a15814a );
 a15816a <=( a15815a  and  a15810a );
 a15820a <=( (not A233)  and  A232 );
 a15821a <=( (not A202)  and  a15820a );
 a15824a <=( A265  and  A236 );
 a15827a <=( A269  and  (not A266) );
 a15828a <=( a15827a  and  a15824a );
 a15829a <=( a15828a  and  a15821a );


end x25_12x_behav;
