Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_10x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A105: buffer std_logic
);
end x25_10x;

architecture x25_10x_behav of x25_10x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1753a,a1754a,a1755a,a1756a,a1757a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1765a,a1766a,a1767a,a1768a,a1769a,a1770a,a1771a,a1772a,a1773a,a1774a,a1775a,a1776a,a1777a,a1778a,a1779a,a1780a,a1781a,a1782a,a1783a,a1784a,a1785a,a1786a,a1787a,a1788a,a1789a,a1790a,a1791a,a1792a,a1793a,a1794a,a1795a,a1796a,a1797a,a1798a,a1799a,a1800a,a1801a,a1802a,a1803a,a1804a,a1805a,a1806a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1816a,a1817a,a1818a,a1819a,a1820a,a1821a,a1822a,a1823a,a1824a,a1825a,a1826a,a1827a,a1828a,a1829a,a1830a,a1831a,a1832a,a1833a,a1834a,a1835a,a1836a,a1837a,a1838a,a1839a,a1840a,a1841a,a1842a,a1843a,a1844a,a1845a,a1846a,a1847a,a1848a,a1849a,a1850a,a1851a,a1852a,a1853a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1860a,a1861a,a1862a,a1863a,a1864a,a1865a,a1866a,a1867a,a1868a,a1869a,a1870a,a1871a,a1872a,a1873a,a1874a,a1875a,a1876a,a1877a,a1878a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1890a,a1891a,a1892a,a1893a,a1894a,a1895a,a1896a,a1897a,a1898a,a1899a,a1900a,a1901a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1910a,a1911a,a1912a,a1913a,a1914a,a1915a,a1916a,a1917a,a1918a,a1919a,a1920a,a1921a,a1922a,a1923a,a1924a,a1925a,a1926a,a1927a,a1928a,a1929a,a1930a,a1931a,a1932a,a1933a,a1934a,a1935a,a1936a,a1937a,a1938a,a1939a,a1940a,a1941a,a1942a,a1943a,a1944a,a1945a,a1946a,a1947a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1956a,a1957a,a1958a,a1959a,a1960a,a1961a,a1962a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1970a,a1971a,a1972a,a1973a,a1974a,a1975a,a1976a,a1977a,a1978a,a1979a,a1980a,a1981a,a1982a,a1983a,a1984a,a1985a,a1986a,a1987a,a1988a,a1989a,a1990a,a1991a,a1992a,a1993a,a1994a,a1995a,a1996a,a1997a,a1998a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2005a,a2006a,a2007a,a2008a,a2009a,a2010a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2025a,a2026a,a2027a,a2028a,a2029a,a2030a,a2031a,a2032a,a2033a,a2034a,a2035a,a2036a,a2037a,a2038a,a2039a,a2040a,a2041a,a2042a,a2043a,a2044a,a2045a,a2046a,a2047a,a2048a,a2049a,a2050a,a2051a,a2052a,a2053a,a2054a,a2055a,a2056a,a2057a,a2058a,a2059a,a2060a,a2061a,a2062a,a2063a,a2064a,a2065a,a2066a,a2067a,a2068a,a2069a,a2070a,a2071a,a2072a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2079a,a2080a,a2081a,a2082a,a2083a,a2084a,a2085a,a2086a,a2087a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2101a,a2102a,a2103a,a2104a,a2105a,a2106a,a2107a,a2108a,a2109a,a2110a,a2111a,a2112a,a2113a,a2114a,a2115a,a2116a,a2117a,a2118a,a2119a,a2120a,a2121a,a2122a,a2123a,a2124a,a2125a,a2126a,a2127a,a2128a,a2129a,a2130a,a2131a,a2132a,a2133a,a2134a,a2135a,a2136a,a2137a,a2138a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2145a,a2146a,a2147a,a2148a,a2149a,a2150a,a2151a,a2152a,a2153a,a2154a,a2155a,a2156a,a2157a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2164a,a2165a,a2166a,a2167a,a2168a,a2169a,a2170a,a2171a,a2172a,a2173a,a2174a,a2175a,a2176a,a2177a,a2178a,a2179a,a2180a,a2181a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2190a,a2191a,a2192a,a2193a,a2194a,a2195a,a2196a,a2197a,a2198a,a2199a,a2200a,a2201a,a2202a,a2203a,a2204a,a2205a,a2206a,a2207a,a2208a,a2209a,a2210a,a2211a,a2212a,a2213a,a2214a,a2215a,a2216a,a2217a,a2218a,a2219a,a2220a,a2221a,a2222a,a2223a,a2224a,a2225a,a2226a,a2227a,a2228a,a2229a,a2230a,a2231a,a2232a,a2233a,a2234a,a2235a,a2236a,a2237a,a2238a,a2239a,a2240a,a2241a,a2242a,a2243a,a2244a,a2245a,a2246a,a2247a,a2248a,a2249a,a2250a,a2251a,a2252a,a2253a,a2254a,a2255a,a2256a,a2257a,a2258a,a2259a,a2260a,a2261a,a2262a,a2263a,a2264a,a2265a,a2266a,a2267a,a2268a,a2269a,a2270a,a2271a,a2272a,a2273a,a2274a,a2275a,a2276a,a2277a,a2278a,a2279a,a2280a,a2281a,a2282a,a2283a,a2284a,a2285a,a2286a,a2287a,a2288a,a2289a,a2290a,a2291a,a2292a,a2293a,a2294a,a2295a,a2296a,a2297a,a2298a,a2299a,a2300a,a2301a,a2302a,a2303a,a2304a,a2305a,a2306a,a2307a,a2308a,a2309a,a2310a,a2311a,a2312a,a2313a,a2314a,a2315a,a2316a,a2317a,a2318a,a2319a,a2320a,a2321a,a2322a,a2323a,a2324a,a2325a,a2326a,a2327a,a2328a,a2329a,a2330a,a2331a,a2332a,a2333a,a2334a,a2335a,a2336a,a2337a,a2338a,a2339a,a2340a,a2341a,a2342a,a2343a,a2344a,a2345a,a2346a,a2347a,a2348a,a2349a,a2350a,a2351a,a2352a,a2353a,a2354a,a2355a,a2356a,a2357a,a2358a,a2359a,a2360a,a2361a,a2362a,a2363a,a2364a,a2365a,a2366a,a2367a,a2368a,a2369a,a2370a,a2371a,a2372a,a2373a,a2374a,a2375a,a2376a,a2377a,a2378a,a2379a,a2380a,a2381a,a2382a,a2383a,a2384a,a2385a,a2386a,a2387a,a2388a,a2389a,a2390a,a2391a,a2392a,a2393a,a2394a,a2395a,a2396a,a2397a,a2398a,a2399a,a2400a,a2401a,a2402a,a2403a,a2404a,a2405a,a2406a,a2407a,a2408a,a2409a,a2410a,a2411a,a2412a,a2413a,a2414a,a2415a,a2416a,a2417a,a2418a,a2419a,a2420a,a2421a,a2422a,a2423a,a2424a,a2425a,a2426a,a2427a,a2428a,a2429a,a2430a,a2431a,a2432a,a2433a,a2434a,a2435a,a2436a,a2437a,a2438a,a2439a,a2440a,a2441a,a2442a,a2443a,a2444a,a2445a,a2446a,a2447a,a2448a,a2449a,a2450a,a2451a,a2452a,a2453a,a2454a,a2455a,a2456a,a2457a,a2458a,a2459a,a2460a,a2461a,a2462a,a2463a,a2464a,a2465a,a2466a,a2467a,a2468a,a2469a,a2470a,a2471a,a2472a,a2473a,a2474a,a2475a,a2476a,a2477a,a2478a,a2479a,a2480a,a2481a,a2482a,a2483a,a2484a,a2485a,a2486a,a2487a,a2488a,a2489a,a2490a,a2491a,a2492a,a2493a,a2494a,a2495a,a2496a,a2497a,a2498a,a2499a,a2500a,a2501a,a2502a,a2503a,a2504a,a2505a,a2506a,a2507a,a2508a,a2509a,a2510a,a2511a,a2512a,a2513a,a2514a,a2515a,a2516a,a2517a,a2518a,a2519a,a2520a,a2521a,a2522a,a2523a,a2524a,a2525a,a2526a,a2527a,a2528a,a2529a,a2530a,a2531a,a2532a,a2533a,a2534a,a2535a,a2536a,a2537a,a2538a,a2539a,a2540a,a2541a,a2542a,a2543a,a2544a,a2545a,a2546a,a2547a,a2548a,a2549a,a2550a,a2551a,a2552a,a2553a,a2554a,a2555a,a2556a,a2557a,a2558a,a2559a,a2560a,a2561a,a2562a,a2563a,a2564a,a2565a,a2566a,a2567a,a2568a,a2569a,a2570a,a2571a,a2572a,a2573a,a2574a,a2575a,a2576a,a2577a,a2578a,a2579a,a2580a,a2581a,a2582a,a2583a,a2584a,a2585a,a2586a,a2587a,a2588a,a2589a,a2590a,a2591a,a2592a,a2593a,a2594a,a2595a,a2596a,a2597a,a2598a,a2599a,a2600a,a2601a,a2602a,a2603a,a2604a,a2605a,a2606a,a2607a,a2608a,a2609a,a2610a,a2611a,a2612a,a2613a,a2614a,a2615a,a2616a,a2617a,a2618a,a2619a,a2620a,a2621a,a2622a,a2623a,a2624a,a2625a,a2626a,a2627a,a2628a,a2629a,a2630a,a2631a,a2632a,a2633a,a2634a,a2635a,a2636a,a2637a,a2638a,a2639a,a2640a,a2641a,a2642a,a2643a,a2644a,a2645a,a2646a,a2647a,a2648a,a2649a,a2650a,a2651a,a2652a,a2653a,a2654a,a2655a,a2656a,a2657a,a2658a,a2659a,a2660a,a2661a,a2662a,a2663a,a2664a,a2665a,a2666a,a2667a,a2668a,a2669a,a2670a,a2671a,a2672a,a2673a,a2674a,a2675a,a2676a,a2677a,a2678a,a2679a,a2680a,a2681a,a2682a,a2683a,a2684a,a2685a,a2686a,a2687a,a2688a,a2689a,a2690a,a2691a,a2692a,a2693a,a2694a,a2695a,a2696a,a2697a,a2698a,a2699a,a2700a,a2701a,a2702a,a2703a,a2704a,a2705a,a2706a,a2707a,a2708a,a2709a,a2710a,a2711a,a2712a,a2713a,a2714a,a2715a,a2716a,a2717a,a2718a,a2719a,a2720a,a2721a,a2722a,a2723a,a2724a,a2725a,a2726a,a2727a,a2728a,a2729a,a2730a,a2731a,a2732a,a2733a,a2734a,a2735a,a2736a,a2737a,a2738a,a2739a,a2740a,a2741a,a2742a,a2743a,a2744a,a2745a,a2746a,a2747a,a2748a,a2749a,a2750a,a2751a,a2752a,a2753a,a2754a,a2755a,a2756a,a2757a,a2758a,a2759a,a2760a,a2761a,a2762a,a2763a,a2764a,a2765a,a2766a,a2767a,a2768a,a2769a,a2770a,a2771a,a2772a,a2773a,a2774a,a2775a,a2776a,a2777a,a2778a,a2779a,a2780a,a2781a,a2782a,a2783a,a2784a,a2785a,a2786a,a2787a,a2788a,a2789a,a2790a,a2791a,a2792a,a2793a,a2794a,a2795a,a2796a,a2797a,a2798a,a2799a,a2800a,a2801a,a2802a,a2803a,a2804a,a2805a,a2806a,a2807a,a2808a,a2809a,a2810a,a2811a,a2812a,a2813a,a2814a,a2815a,a2816a,a2817a,a2818a,a2819a,a2820a,a2821a,a2822a,a2823a,a2824a,a2825a,a2826a,a2827a,a2828a,a2829a,a2830a,a2831a,a2832a,a2833a,a2834a,a2835a,a2836a,a2837a,a2838a,a2839a,a2840a,a2841a,a2842a,a2843a,a2844a,a2845a,a2846a,a2847a,a2848a,a2849a,a2850a,a2851a,a2852a,a2853a,a2854a,a2855a,a2856a,a2857a,a2858a,a2859a,a2860a,a2861a,a2862a,a2863a,a2864a,a2865a,a2866a,a2867a,a2868a,a2869a,a2870a,a2871a,a2872a,a2873a,a2874a,a2875a,a2876a,a2877a,a2878a,a2879a,a2880a,a2881a,a2882a,a2883a,a2884a,a2885a,a2886a,a2887a,a2888a,a2889a,a2890a,a2891a,a2892a,a2893a,a2894a,a2895a,a2896a,a2897a,a2898a,a2899a,a2900a,a2901a,a2902a,a2903a,a2904a,a2905a,a2906a,a2907a,a2908a,a2909a,a2910a,a2911a,a2912a,a2913a,a2914a,a2915a,a2916a,a2917a,a2918a,a2919a,a2920a,a2921a,a2922a,a2923a,a2924a,a2925a,a2926a,a2927a,a2928a,a2929a,a2930a,a2931a,a2932a,a2933a,a2934a,a2935a,a2936a,a2937a,a2938a,a2939a,a2940a,a2941a,a2942a,a2943a,a2944a,a2945a,a2946a,a2947a,a2948a,a2949a,a2950a,a2951a,a2952a,a2953a,a2954a,a2955a,a2956a,a2957a,a2958a,a2959a,a2960a,a2961a,a2962a,a2963a,a2964a,a2965a,a2966a,a2967a,a2968a,a2969a,a2970a,a2971a,a2972a,a2973a,a2974a,a2975a,a2976a,a2977a,a2978a,a2979a,a2980a,a2981a,a2982a,a2983a,a2984a,a2985a,a2986a,a2987a,a2988a,a2989a,a2990a,a2991a,a2992a,a2993a,a2994a,a2995a,a2996a,a2997a,a2998a,a2999a,a3000a,a3001a,a3002a,a3003a,a3004a,a3005a,a3006a,a3007a,a3008a,a3009a,a3010a,a3011a,a3012a,a3013a,a3014a,a3015a,a3016a,a3017a,a3018a,a3019a,a3020a,a3021a,a3022a,a3023a,a3024a,a3025a,a3026a,a3027a,a3028a,a3029a,a3030a,a3031a,a3032a,a3033a,a3034a,a3035a,a3036a,a3037a,a3038a,a3039a,a3040a,a3041a,a3042a,a3043a,a3044a,a3045a,a3046a,a3047a,a3048a,a3049a,a3050a,a3051a,a3052a,a3053a,a3054a,a3055a,a3056a,a3057a,a3058a,a3059a,a3060a,a3061a,a3062a,a3063a,a3064a,a3065a,a3066a,a3067a,a3068a,a3069a,a3070a,a3071a,a3072a,a3073a,a3074a,a3075a,a3076a,a3077a,a3078a,a3079a,a3080a,a3081a,a3082a,a3083a,a3084a,a3085a,a3086a,a3087a,a3088a,a3089a,a3090a,a3091a,a3092a,a3093a,a3094a,a3095a,a3096a,a3097a,a3098a,a3099a,a3100a,a3101a,a3102a,a3103a,a3104a,a3105a,a3106a,a3107a,a3108a,a3109a,a3110a,a3111a,a3112a,a3113a,a3114a,a3115a,a3116a,a3117a,a3118a,a3119a,a3120a,a3121a,a3122a,a3123a,a3124a,a3125a,a3126a,a3127a,a3128a,a3129a,a3130a,a3131a,a3132a,a3133a,a3134a,a3135a,a3136a,a3137a,a3138a,a3139a,a3140a,a3141a,a3142a,a3143a,a3144a,a3145a,a3146a,a3147a,a3148a,a3149a,a3150a,a3151a,a3152a,a3153a,a3154a,a3155a,a3156a,a3157a,a3158a,a3159a,a3160a,a3161a,a3162a,a3163a,a3164a,a3165a,a3166a,a3167a,a3168a,a3169a,a3170a,a3171a,a3172a,a3173a,a3174a,a3178a,a3179a,a3183a,a3184a,a3185a,a3189a,a3190a,a3194a,a3195a,a3196a,a3197a,a3201a,a3202a,a3206a,a3207a,a3208a,a3212a,a3213a,a3217a,a3218a,a3219a,a3220a,a3221a,a3225a,a3226a,a3230a,a3231a,a3232a,a3236a,a3237a,a3241a,a3242a,a3243a,a3244a,a3248a,a3249a,a3253a,a3254a,a3255a,a3259a,a3260a,a3263a,a3266a,a3267a,a3268a,a3269a,a3270a,a3271a,a3275a,a3276a,a3280a,a3281a,a3282a,a3286a,a3287a,a3291a,a3292a,a3293a,a3294a,a3298a,a3299a,a3303a,a3304a,a3305a,a3309a,a3310a,a3313a,a3316a,a3317a,a3318a,a3319a,a3320a,a3324a,a3325a,a3329a,a3330a,a3331a,a3335a,a3336a,a3340a,a3341a,a3342a,a3343a,a3347a,a3348a,a3352a,a3353a,a3354a,a3358a,a3359a,a3362a,a3365a,a3366a,a3367a,a3368a,a3369a,a3370a,a3371a,a3375a,a3376a,a3380a,a3381a,a3382a,a3386a,a3387a,a3391a,a3392a,a3393a,a3394a,a3398a,a3399a,a3403a,a3404a,a3405a,a3409a,a3410a,a3414a,a3415a,a3416a,a3417a,a3418a,a3422a,a3423a,a3427a,a3428a,a3429a,a3433a,a3434a,a3438a,a3439a,a3440a,a3441a,a3445a,a3446a,a3450a,a3451a,a3452a,a3456a,a3457a,a3460a,a3463a,a3464a,a3465a,a3466a,a3467a,a3468a,a3472a,a3473a,a3477a,a3478a,a3479a,a3483a,a3484a,a3488a,a3489a,a3490a,a3491a,a3495a,a3496a,a3500a,a3501a,a3502a,a3506a,a3507a,a3510a,a3513a,a3514a,a3515a,a3516a,a3517a,a3521a,a3522a,a3526a,a3527a,a3528a,a3532a,a3533a,a3537a,a3538a,a3539a,a3540a,a3544a,a3545a,a3549a,a3550a,a3551a,a3555a,a3556a,a3559a,a3562a,a3563a,a3564a,a3565a,a3566a,a3567a,a3568a,a3569a,a3573a,a3574a,a3578a,a3579a,a3580a,a3584a,a3585a,a3589a,a3590a,a3591a,a3592a,a3596a,a3597a,a3601a,a3602a,a3603a,a3607a,a3608a,a3612a,a3613a,a3614a,a3615a,a3616a,a3620a,a3621a,a3625a,a3626a,a3627a,a3631a,a3632a,a3636a,a3637a,a3638a,a3639a,a3643a,a3644a,a3648a,a3649a,a3650a,a3654a,a3655a,a3658a,a3661a,a3662a,a3663a,a3664a,a3665a,a3666a,a3670a,a3671a,a3675a,a3676a,a3677a,a3681a,a3682a,a3686a,a3687a,a3688a,a3689a,a3693a,a3694a,a3698a,a3699a,a3700a,a3704a,a3705a,a3708a,a3711a,a3712a,a3713a,a3714a,a3715a,a3719a,a3720a,a3724a,a3725a,a3726a,a3730a,a3731a,a3735a,a3736a,a3737a,a3738a,a3742a,a3743a,a3747a,a3748a,a3749a,a3753a,a3754a,a3757a,a3760a,a3761a,a3762a,a3763a,a3764a,a3765a,a3766a,a3770a,a3771a,a3775a,a3776a,a3777a,a3781a,a3782a,a3786a,a3787a,a3788a,a3789a,a3793a,a3794a,a3798a,a3799a,a3800a,a3804a,a3805a,a3809a,a3810a,a3811a,a3812a,a3813a,a3817a,a3818a,a3822a,a3823a,a3824a,a3828a,a3829a,a3833a,a3834a,a3835a,a3836a,a3840a,a3841a,a3845a,a3846a,a3847a,a3851a,a3852a,a3855a,a3858a,a3859a,a3860a,a3861a,a3862a,a3863a,a3867a,a3868a,a3872a,a3873a,a3874a,a3878a,a3879a,a3883a,a3884a,a3885a,a3886a,a3890a,a3891a,a3895a,a3896a,a3897a,a3901a,a3902a,a3905a,a3908a,a3909a,a3910a,a3911a,a3912a,a3916a,a3917a,a3921a,a3922a,a3923a,a3927a,a3928a,a3932a,a3933a,a3934a,a3935a,a3939a,a3940a,a3944a,a3945a,a3946a,a3950a,a3951a,a3954a,a3957a,a3958a,a3959a,a3960a,a3961a,a3962a,a3963a,a3964a,a3965a,a3969a,a3970a,a3974a,a3975a,a3976a,a3980a,a3981a,a3985a,a3986a,a3987a,a3988a,a3992a,a3993a,a3997a,a3998a,a3999a,a4003a,a4004a,a4008a,a4009a,a4010a,a4011a,a4012a,a4016a,a4017a,a4021a,a4022a,a4023a,a4027a,a4028a,a4032a,a4033a,a4034a,a4035a,a4039a,a4040a,a4044a,a4045a,a4046a,a4050a,a4051a,a4054a,a4057a,a4058a,a4059a,a4060a,a4061a,a4062a,a4066a,a4067a,a4071a,a4072a,a4073a,a4077a,a4078a,a4082a,a4083a,a4084a,a4085a,a4089a,a4090a,a4094a,a4095a,a4096a,a4100a,a4101a,a4104a,a4107a,a4108a,a4109a,a4110a,a4111a,a4115a,a4116a,a4120a,a4121a,a4122a,a4126a,a4127a,a4131a,a4132a,a4133a,a4134a,a4138a,a4139a,a4143a,a4144a,a4145a,a4149a,a4150a,a4153a,a4156a,a4157a,a4158a,a4159a,a4160a,a4161a,a4162a,a4166a,a4167a,a4171a,a4172a,a4173a,a4177a,a4178a,a4182a,a4183a,a4184a,a4185a,a4189a,a4190a,a4194a,a4195a,a4196a,a4200a,a4201a,a4205a,a4206a,a4207a,a4208a,a4209a,a4213a,a4214a,a4218a,a4219a,a4220a,a4224a,a4225a,a4229a,a4230a,a4231a,a4232a,a4236a,a4237a,a4241a,a4242a,a4243a,a4247a,a4248a,a4251a,a4254a,a4255a,a4256a,a4257a,a4258a,a4259a,a4263a,a4264a,a4268a,a4269a,a4270a,a4274a,a4275a,a4279a,a4280a,a4281a,a4282a,a4286a,a4287a,a4291a,a4292a,a4293a,a4297a,a4298a,a4301a,a4304a,a4305a,a4306a,a4307a,a4308a,a4312a,a4313a,a4317a,a4318a,a4319a,a4323a,a4324a,a4328a,a4329a,a4330a,a4331a,a4335a,a4336a,a4340a,a4341a,a4342a,a4346a,a4347a,a4350a,a4353a,a4354a,a4355a,a4356a,a4357a,a4358a,a4359a,a4360a,a4364a,a4365a,a4369a,a4370a,a4371a,a4375a,a4376a,a4380a,a4381a,a4382a,a4383a,a4387a,a4388a,a4392a,a4393a,a4394a,a4398a,a4399a,a4403a,a4404a,a4405a,a4406a,a4407a,a4411a,a4412a,a4416a,a4417a,a4418a,a4422a,a4423a,a4427a,a4428a,a4429a,a4430a,a4434a,a4435a,a4439a,a4440a,a4441a,a4445a,a4446a,a4449a,a4452a,a4453a,a4454a,a4455a,a4456a,a4457a,a4461a,a4462a,a4466a,a4467a,a4468a,a4472a,a4473a,a4477a,a4478a,a4479a,a4480a,a4484a,a4485a,a4489a,a4490a,a4491a,a4495a,a4496a,a4499a,a4502a,a4503a,a4504a,a4505a,a4506a,a4510a,a4511a,a4515a,a4516a,a4517a,a4521a,a4522a,a4526a,a4527a,a4528a,a4529a,a4533a,a4534a,a4538a,a4539a,a4540a,a4544a,a4545a,a4548a,a4551a,a4552a,a4553a,a4554a,a4555a,a4556a,a4557a,a4561a,a4562a,a4566a,a4567a,a4568a,a4572a,a4573a,a4577a,a4578a,a4579a,a4580a,a4584a,a4585a,a4589a,a4590a,a4591a,a4595a,a4596a,a4599a,a4602a,a4603a,a4604a,a4605a,a4606a,a4610a,a4611a,a4615a,a4616a,a4617a,a4621a,a4622a,a4626a,a4627a,a4628a,a4629a,a4633a,a4634a,a4638a,a4639a,a4640a,a4644a,a4645a,a4648a,a4651a,a4652a,a4653a,a4654a,a4655a,a4656a,a4660a,a4661a,a4665a,a4666a,a4667a,a4671a,a4672a,a4676a,a4677a,a4678a,a4679a,a4683a,a4684a,a4688a,a4689a,a4690a,a4694a,a4695a,a4698a,a4701a,a4702a,a4703a,a4704a,a4705a,a4709a,a4710a,a4714a,a4715a,a4716a,a4720a,a4721a,a4725a,a4726a,a4727a,a4728a,a4732a,a4733a,a4737a,a4738a,a4739a,a4743a,a4744a,a4747a,a4750a,a4751a,a4752a,a4753a,a4754a,a4755a,a4756a,a4757a,a4758a,a4759a,a4763a,a4764a,a4768a,a4769a,a4770a,a4774a,a4775a,a4779a,a4780a,a4781a,a4782a,a4786a,a4787a,a4791a,a4792a,a4793a,a4797a,a4798a,a4802a,a4803a,a4804a,a4805a,a4806a,a4810a,a4811a,a4815a,a4816a,a4817a,a4821a,a4822a,a4826a,a4827a,a4828a,a4829a,a4833a,a4834a,a4838a,a4839a,a4840a,a4844a,a4845a,a4848a,a4851a,a4852a,a4853a,a4854a,a4855a,a4856a,a4860a,a4861a,a4865a,a4866a,a4867a,a4871a,a4872a,a4876a,a4877a,a4878a,a4879a,a4883a,a4884a,a4888a,a4889a,a4890a,a4894a,a4895a,a4898a,a4901a,a4902a,a4903a,a4904a,a4905a,a4909a,a4910a,a4914a,a4915a,a4916a,a4920a,a4921a,a4925a,a4926a,a4927a,a4928a,a4932a,a4933a,a4937a,a4938a,a4939a,a4943a,a4944a,a4947a,a4950a,a4951a,a4952a,a4953a,a4954a,a4955a,a4956a,a4960a,a4961a,a4965a,a4966a,a4967a,a4971a,a4972a,a4976a,a4977a,a4978a,a4979a,a4983a,a4984a,a4988a,a4989a,a4990a,a4994a,a4995a,a4999a,a5000a,a5001a,a5002a,a5003a,a5007a,a5008a,a5012a,a5013a,a5014a,a5018a,a5019a,a5023a,a5024a,a5025a,a5026a,a5030a,a5031a,a5035a,a5036a,a5037a,a5041a,a5042a,a5045a,a5048a,a5049a,a5050a,a5051a,a5052a,a5053a,a5057a,a5058a,a5062a,a5063a,a5064a,a5068a,a5069a,a5073a,a5074a,a5075a,a5076a,a5080a,a5081a,a5085a,a5086a,a5087a,a5091a,a5092a,a5095a,a5098a,a5099a,a5100a,a5101a,a5102a,a5106a,a5107a,a5111a,a5112a,a5113a,a5117a,a5118a,a5122a,a5123a,a5124a,a5125a,a5129a,a5130a,a5134a,a5135a,a5136a,a5140a,a5141a,a5144a,a5147a,a5148a,a5149a,a5150a,a5151a,a5152a,a5153a,a5154a,a5158a,a5159a,a5163a,a5164a,a5165a,a5169a,a5170a,a5174a,a5175a,a5176a,a5177a,a5181a,a5182a,a5186a,a5187a,a5188a,a5192a,a5193a,a5197a,a5198a,a5199a,a5200a,a5201a,a5205a,a5206a,a5210a,a5211a,a5212a,a5216a,a5217a,a5221a,a5222a,a5223a,a5224a,a5228a,a5229a,a5233a,a5234a,a5235a,a5239a,a5240a,a5243a,a5246a,a5247a,a5248a,a5249a,a5250a,a5251a,a5255a,a5256a,a5260a,a5261a,a5262a,a5266a,a5267a,a5271a,a5272a,a5273a,a5274a,a5278a,a5279a,a5283a,a5284a,a5285a,a5289a,a5290a,a5293a,a5296a,a5297a,a5298a,a5299a,a5300a,a5304a,a5305a,a5309a,a5310a,a5311a,a5315a,a5316a,a5320a,a5321a,a5322a,a5323a,a5327a,a5328a,a5332a,a5333a,a5334a,a5338a,a5339a,a5342a,a5345a,a5346a,a5347a,a5348a,a5349a,a5350a,a5351a,a5355a,a5356a,a5360a,a5361a,a5362a,a5366a,a5367a,a5371a,a5372a,a5373a,a5374a,a5378a,a5379a,a5383a,a5384a,a5385a,a5389a,a5390a,a5393a,a5396a,a5397a,a5398a,a5399a,a5400a,a5404a,a5405a,a5409a,a5410a,a5411a,a5415a,a5416a,a5420a,a5421a,a5422a,a5423a,a5427a,a5428a,a5432a,a5433a,a5434a,a5438a,a5439a,a5442a,a5445a,a5446a,a5447a,a5448a,a5449a,a5450a,a5454a,a5455a,a5459a,a5460a,a5461a,a5465a,a5466a,a5470a,a5471a,a5472a,a5473a,a5477a,a5478a,a5482a,a5483a,a5484a,a5488a,a5489a,a5492a,a5495a,a5496a,a5497a,a5498a,a5499a,a5503a,a5504a,a5508a,a5509a,a5510a,a5514a,a5515a,a5519a,a5520a,a5521a,a5522a,a5526a,a5527a,a5531a,a5532a,a5533a,a5537a,a5538a,a5541a,a5544a,a5545a,a5546a,a5547a,a5548a,a5549a,a5550a,a5551a,a5552a,a5556a,a5557a,a5561a,a5562a,a5563a,a5567a,a5568a,a5572a,a5573a,a5574a,a5575a,a5579a,a5580a,a5584a,a5585a,a5586a,a5590a,a5591a,a5595a,a5596a,a5597a,a5598a,a5599a,a5603a,a5604a,a5608a,a5609a,a5610a,a5614a,a5615a,a5619a,a5620a,a5621a,a5622a,a5626a,a5627a,a5631a,a5632a,a5633a,a5637a,a5638a,a5641a,a5644a,a5645a,a5646a,a5647a,a5648a,a5649a,a5653a,a5654a,a5658a,a5659a,a5660a,a5664a,a5665a,a5669a,a5670a,a5671a,a5672a,a5676a,a5677a,a5681a,a5682a,a5683a,a5687a,a5688a,a5691a,a5694a,a5695a,a5696a,a5697a,a5698a,a5702a,a5703a,a5707a,a5708a,a5709a,a5713a,a5714a,a5718a,a5719a,a5720a,a5721a,a5725a,a5726a,a5730a,a5731a,a5732a,a5736a,a5737a,a5740a,a5743a,a5744a,a5745a,a5746a,a5747a,a5748a,a5749a,a5753a,a5754a,a5758a,a5759a,a5760a,a5764a,a5765a,a5769a,a5770a,a5771a,a5772a,a5776a,a5777a,a5781a,a5782a,a5783a,a5787a,a5788a,a5792a,a5793a,a5794a,a5795a,a5796a,a5800a,a5801a,a5805a,a5806a,a5807a,a5811a,a5812a,a5816a,a5817a,a5818a,a5819a,a5823a,a5824a,a5828a,a5829a,a5830a,a5834a,a5835a,a5838a,a5841a,a5842a,a5843a,a5844a,a5845a,a5846a,a5850a,a5851a,a5855a,a5856a,a5857a,a5861a,a5862a,a5866a,a5867a,a5868a,a5869a,a5873a,a5874a,a5878a,a5879a,a5880a,a5884a,a5885a,a5888a,a5891a,a5892a,a5893a,a5894a,a5895a,a5899a,a5900a,a5904a,a5905a,a5906a,a5910a,a5911a,a5915a,a5916a,a5917a,a5918a,a5922a,a5923a,a5927a,a5928a,a5929a,a5933a,a5934a,a5937a,a5940a,a5941a,a5942a,a5943a,a5944a,a5945a,a5946a,a5947a,a5951a,a5952a,a5956a,a5957a,a5958a,a5962a,a5963a,a5967a,a5968a,a5969a,a5970a,a5974a,a5975a,a5979a,a5980a,a5981a,a5985a,a5986a,a5990a,a5991a,a5992a,a5993a,a5994a,a5998a,a5999a,a6003a,a6004a,a6005a,a6009a,a6010a,a6014a,a6015a,a6016a,a6017a,a6021a,a6022a,a6026a,a6027a,a6028a,a6032a,a6033a,a6036a,a6039a,a6040a,a6041a,a6042a,a6043a,a6044a,a6048a,a6049a,a6053a,a6054a,a6055a,a6059a,a6060a,a6064a,a6065a,a6066a,a6067a,a6071a,a6072a,a6076a,a6077a,a6078a,a6082a,a6083a,a6086a,a6089a,a6090a,a6091a,a6092a,a6093a,a6097a,a6098a,a6102a,a6103a,a6104a,a6108a,a6109a,a6113a,a6114a,a6115a,a6116a,a6120a,a6121a,a6125a,a6126a,a6127a,a6131a,a6132a,a6135a,a6138a,a6139a,a6140a,a6141a,a6142a,a6143a,a6144a,a6148a,a6149a,a6153a,a6154a,a6155a,a6159a,a6160a,a6164a,a6165a,a6166a,a6167a,a6171a,a6172a,a6176a,a6177a,a6178a,a6182a,a6183a,a6186a,a6189a,a6190a,a6191a,a6192a,a6193a,a6197a,a6198a,a6202a,a6203a,a6204a,a6208a,a6209a,a6213a,a6214a,a6215a,a6216a,a6220a,a6221a,a6225a,a6226a,a6227a,a6231a,a6232a,a6235a,a6238a,a6239a,a6240a,a6241a,a6242a,a6243a,a6247a,a6248a,a6252a,a6253a,a6254a,a6258a,a6259a,a6263a,a6264a,a6265a,a6266a,a6270a,a6271a,a6275a,a6276a,a6277a,a6281a,a6282a,a6285a,a6288a,a6289a,a6290a,a6291a,a6292a,a6296a,a6297a,a6301a,a6302a,a6303a,a6307a,a6308a,a6312a,a6313a,a6314a,a6315a,a6319a,a6320a,a6324a,a6325a,a6326a,a6330a,a6331a,a6334a,a6337a,a6338a,a6339a,a6340a,a6341a,a6342a,a6343a,a6344a,a6345a,a6346a,a6347a,a6351a,a6352a,a6356a,a6357a,a6358a,a6362a,a6363a,a6367a,a6368a,a6369a,a6370a,a6374a,a6375a,a6379a,a6380a,a6381a,a6385a,a6386a,a6390a,a6391a,a6392a,a6393a,a6394a,a6398a,a6399a,a6403a,a6404a,a6405a,a6409a,a6410a,a6414a,a6415a,a6416a,a6417a,a6421a,a6422a,a6426a,a6427a,a6428a,a6432a,a6433a,a6436a,a6439a,a6440a,a6441a,a6442a,a6443a,a6444a,a6448a,a6449a,a6453a,a6454a,a6455a,a6459a,a6460a,a6464a,a6465a,a6466a,a6467a,a6471a,a6472a,a6476a,a6477a,a6478a,a6482a,a6483a,a6486a,a6489a,a6490a,a6491a,a6492a,a6493a,a6497a,a6498a,a6502a,a6503a,a6504a,a6508a,a6509a,a6513a,a6514a,a6515a,a6516a,a6520a,a6521a,a6525a,a6526a,a6527a,a6531a,a6532a,a6535a,a6538a,a6539a,a6540a,a6541a,a6542a,a6543a,a6544a,a6548a,a6549a,a6553a,a6554a,a6555a,a6559a,a6560a,a6564a,a6565a,a6566a,a6567a,a6571a,a6572a,a6576a,a6577a,a6578a,a6582a,a6583a,a6587a,a6588a,a6589a,a6590a,a6591a,a6595a,a6596a,a6600a,a6601a,a6602a,a6606a,a6607a,a6611a,a6612a,a6613a,a6614a,a6618a,a6619a,a6623a,a6624a,a6625a,a6629a,a6630a,a6633a,a6636a,a6637a,a6638a,a6639a,a6640a,a6641a,a6645a,a6646a,a6650a,a6651a,a6652a,a6656a,a6657a,a6661a,a6662a,a6663a,a6664a,a6668a,a6669a,a6673a,a6674a,a6675a,a6679a,a6680a,a6683a,a6686a,a6687a,a6688a,a6689a,a6690a,a6694a,a6695a,a6699a,a6700a,a6701a,a6705a,a6706a,a6710a,a6711a,a6712a,a6713a,a6717a,a6718a,a6722a,a6723a,a6724a,a6728a,a6729a,a6732a,a6735a,a6736a,a6737a,a6738a,a6739a,a6740a,a6741a,a6742a,a6746a,a6747a,a6751a,a6752a,a6753a,a6757a,a6758a,a6762a,a6763a,a6764a,a6765a,a6769a,a6770a,a6774a,a6775a,a6776a,a6780a,a6781a,a6785a,a6786a,a6787a,a6788a,a6789a,a6793a,a6794a,a6798a,a6799a,a6800a,a6804a,a6805a,a6809a,a6810a,a6811a,a6812a,a6816a,a6817a,a6821a,a6822a,a6823a,a6827a,a6828a,a6831a,a6834a,a6835a,a6836a,a6837a,a6838a,a6839a,a6843a,a6844a,a6848a,a6849a,a6850a,a6854a,a6855a,a6859a,a6860a,a6861a,a6862a,a6866a,a6867a,a6871a,a6872a,a6873a,a6877a,a6878a,a6881a,a6884a,a6885a,a6886a,a6887a,a6888a,a6892a,a6893a,a6897a,a6898a,a6899a,a6903a,a6904a,a6908a,a6909a,a6910a,a6911a,a6915a,a6916a,a6920a,a6921a,a6922a,a6926a,a6927a,a6930a,a6933a,a6934a,a6935a,a6936a,a6937a,a6938a,a6939a,a6943a,a6944a,a6948a,a6949a,a6950a,a6954a,a6955a,a6959a,a6960a,a6961a,a6962a,a6966a,a6967a,a6971a,a6972a,a6973a,a6977a,a6978a,a6982a,a6983a,a6984a,a6985a,a6986a,a6990a,a6991a,a6995a,a6996a,a6997a,a7001a,a7002a,a7006a,a7007a,a7008a,a7009a,a7013a,a7014a,a7018a,a7019a,a7020a,a7024a,a7025a,a7028a,a7031a,a7032a,a7033a,a7034a,a7035a,a7036a,a7040a,a7041a,a7045a,a7046a,a7047a,a7051a,a7052a,a7056a,a7057a,a7058a,a7059a,a7063a,a7064a,a7068a,a7069a,a7070a,a7074a,a7075a,a7078a,a7081a,a7082a,a7083a,a7084a,a7085a,a7089a,a7090a,a7094a,a7095a,a7096a,a7100a,a7101a,a7105a,a7106a,a7107a,a7108a,a7112a,a7113a,a7117a,a7118a,a7119a,a7123a,a7124a,a7127a,a7130a,a7131a,a7132a,a7133a,a7134a,a7135a,a7136a,a7137a,a7138a,a7142a,a7143a,a7147a,a7148a,a7149a,a7153a,a7154a,a7158a,a7159a,a7160a,a7161a,a7165a,a7166a,a7170a,a7171a,a7172a,a7176a,a7177a,a7181a,a7182a,a7183a,a7184a,a7185a,a7189a,a7190a,a7194a,a7195a,a7196a,a7200a,a7201a,a7205a,a7206a,a7207a,a7208a,a7212a,a7213a,a7217a,a7218a,a7219a,a7223a,a7224a,a7227a,a7230a,a7231a,a7232a,a7233a,a7234a,a7235a,a7239a,a7240a,a7244a,a7245a,a7246a,a7250a,a7251a,a7255a,a7256a,a7257a,a7258a,a7262a,a7263a,a7267a,a7268a,a7269a,a7273a,a7274a,a7277a,a7280a,a7281a,a7282a,a7283a,a7284a,a7288a,a7289a,a7293a,a7294a,a7295a,a7299a,a7300a,a7304a,a7305a,a7306a,a7307a,a7311a,a7312a,a7316a,a7317a,a7318a,a7322a,a7323a,a7326a,a7329a,a7330a,a7331a,a7332a,a7333a,a7334a,a7335a,a7339a,a7340a,a7344a,a7345a,a7346a,a7350a,a7351a,a7355a,a7356a,a7357a,a7358a,a7362a,a7363a,a7367a,a7368a,a7369a,a7373a,a7374a,a7378a,a7379a,a7380a,a7381a,a7382a,a7386a,a7387a,a7391a,a7392a,a7393a,a7397a,a7398a,a7402a,a7403a,a7404a,a7405a,a7409a,a7410a,a7414a,a7415a,a7416a,a7420a,a7421a,a7424a,a7427a,a7428a,a7429a,a7430a,a7431a,a7432a,a7436a,a7437a,a7441a,a7442a,a7443a,a7447a,a7448a,a7452a,a7453a,a7454a,a7455a,a7459a,a7460a,a7464a,a7465a,a7466a,a7470a,a7471a,a7474a,a7477a,a7478a,a7479a,a7480a,a7481a,a7485a,a7486a,a7490a,a7491a,a7492a,a7496a,a7497a,a7501a,a7502a,a7503a,a7504a,a7508a,a7509a,a7513a,a7514a,a7515a,a7519a,a7520a,a7523a,a7526a,a7527a,a7528a,a7529a,a7530a,a7531a,a7532a,a7533a,a7537a,a7538a,a7542a,a7543a,a7544a,a7548a,a7549a,a7553a,a7554a,a7555a,a7556a,a7560a,a7561a,a7565a,a7566a,a7567a,a7571a,a7572a,a7576a,a7577a,a7578a,a7579a,a7580a,a7584a,a7585a,a7589a,a7590a,a7591a,a7595a,a7596a,a7600a,a7601a,a7602a,a7603a,a7607a,a7608a,a7612a,a7613a,a7614a,a7618a,a7619a,a7622a,a7625a,a7626a,a7627a,a7628a,a7629a,a7630a,a7634a,a7635a,a7639a,a7640a,a7641a,a7645a,a7646a,a7650a,a7651a,a7652a,a7653a,a7657a,a7658a,a7662a,a7663a,a7664a,a7668a,a7669a,a7672a,a7675a,a7676a,a7677a,a7678a,a7679a,a7683a,a7684a,a7688a,a7689a,a7690a,a7694a,a7695a,a7699a,a7700a,a7701a,a7702a,a7706a,a7707a,a7711a,a7712a,a7713a,a7717a,a7718a,a7721a,a7724a,a7725a,a7726a,a7727a,a7728a,a7729a,a7730a,a7734a,a7735a,a7739a,a7740a,a7741a,a7745a,a7746a,a7750a,a7751a,a7752a,a7753a,a7757a,a7758a,a7762a,a7763a,a7764a,a7768a,a7769a,a7772a,a7775a,a7776a,a7777a,a7778a,a7779a,a7783a,a7784a,a7788a,a7789a,a7790a,a7794a,a7795a,a7799a,a7800a,a7801a,a7802a,a7806a,a7807a,a7811a,a7812a,a7813a,a7817a,a7818a,a7821a,a7824a,a7825a,a7826a,a7827a,a7828a,a7829a,a7833a,a7834a,a7838a,a7839a,a7840a,a7844a,a7845a,a7849a,a7850a,a7851a,a7852a,a7856a,a7857a,a7861a,a7862a,a7863a,a7867a,a7868a,a7871a,a7874a,a7875a,a7876a,a7877a,a7878a,a7882a,a7883a,a7887a,a7888a,a7889a,a7893a,a7894a,a7898a,a7899a,a7900a,a7901a,a7905a,a7906a,a7910a,a7911a,a7912a,a7916a,a7917a,a7920a,a7923a,a7924a,a7925a,a7926a,a7927a,a7928a,a7929a,a7930a,a7931a,a7932a,a7936a,a7937a,a7941a,a7942a,a7943a,a7947a,a7948a,a7952a,a7953a,a7954a,a7955a,a7959a,a7960a,a7964a,a7965a,a7966a,a7970a,a7971a,a7975a,a7976a,a7977a,a7978a,a7979a,a7983a,a7984a,a7988a,a7989a,a7990a,a7994a,a7995a,a7999a,a8000a,a8001a,a8002a,a8006a,a8007a,a8011a,a8012a,a8013a,a8017a,a8018a,a8021a,a8024a,a8025a,a8026a,a8027a,a8028a,a8029a,a8033a,a8034a,a8038a,a8039a,a8040a,a8044a,a8045a,a8049a,a8050a,a8051a,a8052a,a8056a,a8057a,a8061a,a8062a,a8063a,a8067a,a8068a,a8071a,a8074a,a8075a,a8076a,a8077a,a8078a,a8082a,a8083a,a8087a,a8088a,a8089a,a8093a,a8094a,a8098a,a8099a,a8100a,a8101a,a8105a,a8106a,a8110a,a8111a,a8112a,a8116a,a8117a,a8120a,a8123a,a8124a,a8125a,a8126a,a8127a,a8128a,a8129a,a8133a,a8134a,a8138a,a8139a,a8140a,a8144a,a8145a,a8149a,a8150a,a8151a,a8152a,a8156a,a8157a,a8161a,a8162a,a8163a,a8167a,a8168a,a8172a,a8173a,a8174a,a8175a,a8176a,a8180a,a8181a,a8185a,a8186a,a8187a,a8191a,a8192a,a8196a,a8197a,a8198a,a8199a,a8203a,a8204a,a8208a,a8209a,a8210a,a8214a,a8215a,a8218a,a8221a,a8222a,a8223a,a8224a,a8225a,a8226a,a8230a,a8231a,a8235a,a8236a,a8237a,a8241a,a8242a,a8246a,a8247a,a8248a,a8249a,a8253a,a8254a,a8258a,a8259a,a8260a,a8264a,a8265a,a8268a,a8271a,a8272a,a8273a,a8274a,a8275a,a8279a,a8280a,a8284a,a8285a,a8286a,a8290a,a8291a,a8295a,a8296a,a8297a,a8298a,a8302a,a8303a,a8307a,a8308a,a8309a,a8313a,a8314a,a8317a,a8320a,a8321a,a8322a,a8323a,a8324a,a8325a,a8326a,a8327a,a8331a,a8332a,a8336a,a8337a,a8338a,a8342a,a8343a,a8347a,a8348a,a8349a,a8350a,a8354a,a8355a,a8359a,a8360a,a8361a,a8365a,a8366a,a8370a,a8371a,a8372a,a8373a,a8374a,a8378a,a8379a,a8383a,a8384a,a8385a,a8389a,a8390a,a8394a,a8395a,a8396a,a8397a,a8401a,a8402a,a8406a,a8407a,a8408a,a8412a,a8413a,a8416a,a8419a,a8420a,a8421a,a8422a,a8423a,a8424a,a8428a,a8429a,a8433a,a8434a,a8435a,a8439a,a8440a,a8444a,a8445a,a8446a,a8447a,a8451a,a8452a,a8456a,a8457a,a8458a,a8462a,a8463a,a8466a,a8469a,a8470a,a8471a,a8472a,a8473a,a8477a,a8478a,a8482a,a8483a,a8484a,a8488a,a8489a,a8493a,a8494a,a8495a,a8496a,a8500a,a8501a,a8505a,a8506a,a8507a,a8511a,a8512a,a8515a,a8518a,a8519a,a8520a,a8521a,a8522a,a8523a,a8524a,a8528a,a8529a,a8533a,a8534a,a8535a,a8539a,a8540a,a8544a,a8545a,a8546a,a8547a,a8551a,a8552a,a8556a,a8557a,a8558a,a8562a,a8563a,a8566a,a8569a,a8570a,a8571a,a8572a,a8573a,a8577a,a8578a,a8582a,a8583a,a8584a,a8588a,a8589a,a8593a,a8594a,a8595a,a8596a,a8600a,a8601a,a8605a,a8606a,a8607a,a8611a,a8612a,a8615a,a8618a,a8619a,a8620a,a8621a,a8622a,a8623a,a8627a,a8628a,a8632a,a8633a,a8634a,a8638a,a8639a,a8643a,a8644a,a8645a,a8646a,a8650a,a8651a,a8655a,a8656a,a8657a,a8661a,a8662a,a8665a,a8668a,a8669a,a8670a,a8671a,a8672a,a8676a,a8677a,a8681a,a8682a,a8683a,a8687a,a8688a,a8692a,a8693a,a8694a,a8695a,a8699a,a8700a,a8704a,a8705a,a8706a,a8710a,a8711a,a8714a,a8717a,a8718a,a8719a,a8720a,a8721a,a8722a,a8723a,a8724a,a8725a,a8729a,a8730a,a8734a,a8735a,a8736a,a8740a,a8741a,a8745a,a8746a,a8747a,a8748a,a8752a,a8753a,a8757a,a8758a,a8759a,a8763a,a8764a,a8768a,a8769a,a8770a,a8771a,a8772a,a8776a,a8777a,a8781a,a8782a,a8783a,a8787a,a8788a,a8792a,a8793a,a8794a,a8795a,a8799a,a8800a,a8804a,a8805a,a8806a,a8810a,a8811a,a8814a,a8817a,a8818a,a8819a,a8820a,a8821a,a8822a,a8826a,a8827a,a8831a,a8832a,a8833a,a8837a,a8838a,a8842a,a8843a,a8844a,a8845a,a8849a,a8850a,a8854a,a8855a,a8856a,a8860a,a8861a,a8864a,a8867a,a8868a,a8869a,a8870a,a8871a,a8875a,a8876a,a8880a,a8881a,a8882a,a8886a,a8887a,a8891a,a8892a,a8893a,a8894a,a8898a,a8899a,a8903a,a8904a,a8905a,a8909a,a8910a,a8913a,a8916a,a8917a,a8918a,a8919a,a8920a,a8921a,a8922a,a8926a,a8927a,a8931a,a8932a,a8933a,a8937a,a8938a,a8942a,a8943a,a8944a,a8945a,a8949a,a8950a,a8954a,a8955a,a8956a,a8960a,a8961a,a8965a,a8966a,a8967a,a8968a,a8969a,a8973a,a8974a,a8978a,a8979a,a8980a,a8984a,a8985a,a8989a,a8990a,a8991a,a8992a,a8996a,a8997a,a9001a,a9002a,a9003a,a9007a,a9008a,a9011a,a9014a,a9015a,a9016a,a9017a,a9018a,a9019a,a9023a,a9024a,a9028a,a9029a,a9030a,a9034a,a9035a,a9039a,a9040a,a9041a,a9042a,a9046a,a9047a,a9051a,a9052a,a9053a,a9057a,a9058a,a9061a,a9064a,a9065a,a9066a,a9067a,a9068a,a9072a,a9073a,a9077a,a9078a,a9079a,a9083a,a9084a,a9088a,a9089a,a9090a,a9091a,a9095a,a9096a,a9100a,a9101a,a9102a,a9106a,a9107a,a9110a,a9113a,a9114a,a9115a,a9116a,a9117a,a9118a,a9119a,a9120a,a9124a,a9125a,a9129a,a9130a,a9131a,a9135a,a9136a,a9140a,a9141a,a9142a,a9143a,a9147a,a9148a,a9152a,a9153a,a9154a,a9158a,a9159a,a9163a,a9164a,a9165a,a9166a,a9167a,a9171a,a9172a,a9176a,a9177a,a9178a,a9182a,a9183a,a9187a,a9188a,a9189a,a9190a,a9194a,a9195a,a9199a,a9200a,a9201a,a9205a,a9206a,a9209a,a9212a,a9213a,a9214a,a9215a,a9216a,a9217a,a9221a,a9222a,a9226a,a9227a,a9228a,a9232a,a9233a,a9237a,a9238a,a9239a,a9240a,a9244a,a9245a,a9249a,a9250a,a9251a,a9255a,a9256a,a9259a,a9262a,a9263a,a9264a,a9265a,a9266a,a9270a,a9271a,a9275a,a9276a,a9277a,a9281a,a9282a,a9286a,a9287a,a9288a,a9289a,a9293a,a9294a,a9298a,a9299a,a9300a,a9304a,a9305a,a9308a,a9311a,a9312a,a9313a,a9314a,a9315a,a9316a,a9317a,a9321a,a9322a,a9326a,a9327a,a9328a,a9332a,a9333a,a9337a,a9338a,a9339a,a9340a,a9344a,a9345a,a9349a,a9350a,a9351a,a9355a,a9356a,a9359a,a9362a,a9363a,a9364a,a9365a,a9366a,a9370a,a9371a,a9375a,a9376a,a9377a,a9381a,a9382a,a9386a,a9387a,a9388a,a9389a,a9393a,a9394a,a9398a,a9399a,a9400a,a9404a,a9405a,a9408a,a9411a,a9412a,a9413a,a9414a,a9415a,a9416a,a9420a,a9421a,a9425a,a9426a,a9427a,a9431a,a9432a,a9436a,a9437a,a9438a,a9439a,a9443a,a9444a,a9448a,a9449a,a9450a,a9454a,a9455a,a9458a,a9461a,a9462a,a9463a,a9464a,a9465a,a9469a,a9470a,a9474a,a9475a,a9476a,a9480a,a9481a,a9485a,a9486a,a9487a,a9488a,a9492a,a9493a,a9497a,a9498a,a9499a,a9503a,a9504a,a9507a,a9510a,a9511a,a9512a,a9513a,a9514a,a9515a,a9516a,a9517a,a9518a,a9519a,a9520a,a9523a,a9526a,a9527a,a9530a,a9533a,a9534a,a9537a,a9540a,a9541a,a9544a,a9547a,a9548a,a9551a,a9554a,a9555a,a9558a,a9561a,a9562a,a9565a,a9568a,a9569a,a9572a,a9575a,a9576a,a9579a,a9582a,a9583a,a9586a,a9589a,a9590a,a9593a,a9596a,a9597a,a9600a,a9603a,a9604a,a9607a,a9610a,a9611a,a9614a,a9617a,a9618a,a9621a,a9624a,a9625a,a9628a,a9631a,a9632a,a9635a,a9638a,a9639a,a9642a,a9645a,a9646a,a9649a,a9652a,a9653a,a9656a,a9659a,a9660a,a9663a,a9666a,a9667a,a9670a,a9673a,a9674a,a9677a,a9680a,a9681a,a9684a,a9687a,a9688a,a9691a,a9694a,a9695a,a9698a,a9701a,a9702a,a9705a,a9708a,a9709a,a9712a,a9715a,a9716a,a9719a,a9722a,a9723a,a9726a,a9729a,a9730a,a9733a,a9736a,a9737a,a9740a,a9743a,a9744a,a9747a,a9750a,a9751a,a9754a,a9757a,a9758a,a9761a,a9764a,a9765a,a9768a,a9771a,a9772a,a9775a,a9778a,a9779a,a9782a,a9785a,a9786a,a9789a,a9792a,a9793a,a9796a,a9799a,a9800a,a9803a,a9806a,a9807a,a9810a,a9813a,a9814a,a9817a,a9820a,a9821a,a9824a,a9827a,a9828a,a9831a,a9834a,a9835a,a9838a,a9841a,a9842a,a9845a,a9848a,a9849a,a9852a,a9855a,a9856a,a9859a,a9862a,a9863a,a9866a,a9870a,a9871a,a9872a,a9875a,a9878a,a9879a,a9882a,a9886a,a9887a,a9888a,a9891a,a9894a,a9895a,a9898a,a9902a,a9903a,a9904a,a9907a,a9910a,a9911a,a9914a,a9918a,a9919a,a9920a,a9923a,a9926a,a9927a,a9930a,a9934a,a9935a,a9936a,a9939a,a9942a,a9943a,a9946a,a9950a,a9951a,a9952a,a9955a,a9958a,a9959a,a9962a,a9966a,a9967a,a9968a,a9971a,a9974a,a9975a,a9978a,a9982a,a9983a,a9984a,a9987a,a9990a,a9991a,a9994a,a9998a,a9999a,a10000a,a10003a,a10006a,a10007a,a10010a,a10014a,a10015a,a10016a,a10019a,a10022a,a10023a,a10026a,a10030a,a10031a,a10032a,a10035a,a10038a,a10039a,a10042a,a10046a,a10047a,a10048a,a10051a,a10054a,a10055a,a10058a,a10062a,a10063a,a10064a,a10067a,a10070a,a10071a,a10074a,a10078a,a10079a,a10080a,a10083a,a10086a,a10087a,a10090a,a10094a,a10095a,a10096a,a10099a,a10102a,a10103a,a10106a,a10110a,a10111a,a10112a,a10115a,a10118a,a10119a,a10122a,a10126a,a10127a,a10128a,a10131a,a10134a,a10135a,a10138a,a10142a,a10143a,a10144a,a10147a,a10150a,a10151a,a10154a,a10158a,a10159a,a10160a,a10163a,a10166a,a10167a,a10170a,a10174a,a10175a,a10176a,a10179a,a10182a,a10183a,a10186a,a10190a,a10191a,a10192a,a10195a,a10198a,a10199a,a10202a,a10206a,a10207a,a10208a,a10211a,a10215a,a10216a,a10217a,a10220a,a10224a,a10225a,a10226a,a10229a,a10233a,a10234a,a10235a,a10238a,a10242a,a10243a,a10244a,a10247a,a10251a,a10252a,a10253a,a10256a,a10260a,a10261a,a10262a,a10265a,a10269a,a10270a,a10271a,a10274a,a10278a,a10279a,a10280a,a10283a,a10287a,a10288a,a10289a,a10292a,a10296a,a10297a,a10298a,a10301a,a10305a,a10306a,a10307a,a10310a,a10314a,a10315a,a10316a,a10319a,a10323a,a10324a,a10325a,a10328a,a10332a,a10333a,a10334a,a10337a,a10341a,a10342a,a10343a,a10346a,a10350a,a10351a,a10352a,a10355a,a10359a,a10360a,a10361a,a10364a,a10368a,a10369a,a10370a,a10373a,a10377a,a10378a,a10379a,a10382a,a10386a,a10387a,a10388a,a10391a,a10395a,a10396a,a10397a,a10400a,a10404a,a10405a,a10406a,a10409a,a10413a,a10414a,a10415a,a10418a,a10422a,a10423a,a10424a,a10427a,a10431a,a10432a,a10433a,a10436a,a10440a,a10441a,a10442a,a10445a,a10449a,a10450a,a10451a,a10454a,a10458a,a10459a,a10460a,a10463a,a10467a,a10468a,a10469a,a10472a,a10476a,a10477a,a10478a,a10481a,a10485a,a10486a,a10487a,a10490a,a10494a,a10495a,a10496a,a10499a,a10503a,a10504a,a10505a,a10508a,a10512a,a10513a,a10514a,a10517a,a10521a,a10522a,a10523a,a10526a,a10530a,a10531a,a10532a,a10535a,a10539a,a10540a,a10541a,a10544a,a10548a,a10549a,a10550a,a10553a,a10557a,a10558a,a10559a,a10562a,a10566a,a10567a,a10568a,a10571a,a10575a,a10576a,a10577a,a10580a,a10584a,a10585a,a10586a,a10589a,a10593a,a10594a,a10595a,a10598a,a10602a,a10603a,a10604a,a10607a,a10611a,a10612a,a10613a,a10616a,a10620a,a10621a,a10622a,a10625a,a10629a,a10630a,a10631a,a10634a,a10638a,a10639a,a10640a,a10643a,a10647a,a10648a,a10649a,a10652a,a10656a,a10657a,a10658a,a10661a,a10665a,a10666a,a10667a,a10670a,a10674a,a10675a,a10676a,a10679a,a10683a,a10684a,a10685a,a10688a,a10692a,a10693a,a10694a,a10697a,a10701a,a10702a,a10703a,a10706a,a10710a,a10711a,a10712a,a10715a,a10719a,a10720a,a10721a,a10724a,a10728a,a10729a,a10730a,a10733a,a10737a,a10738a,a10739a,a10742a,a10746a,a10747a,a10748a,a10751a,a10755a,a10756a,a10757a,a10760a,a10764a,a10765a,a10766a,a10769a,a10773a,a10774a,a10775a,a10778a,a10782a,a10783a,a10784a,a10787a,a10791a,a10792a,a10793a,a10796a,a10800a,a10801a,a10802a,a10805a,a10809a,a10810a,a10811a,a10814a,a10818a,a10819a,a10820a,a10823a,a10827a,a10828a,a10829a,a10832a,a10836a,a10837a,a10838a,a10841a,a10845a,a10846a,a10847a,a10850a,a10854a,a10855a,a10856a,a10859a,a10863a,a10864a,a10865a,a10868a,a10872a,a10873a,a10874a,a10877a,a10881a,a10882a,a10883a,a10886a,a10890a,a10891a,a10892a,a10895a,a10899a,a10900a,a10901a,a10904a,a10908a,a10909a,a10910a,a10913a,a10917a,a10918a,a10919a,a10922a,a10926a,a10927a,a10928a,a10931a,a10935a,a10936a,a10937a,a10940a,a10944a,a10945a,a10946a,a10949a,a10953a,a10954a,a10955a,a10958a,a10962a,a10963a,a10964a,a10967a,a10971a,a10972a,a10973a,a10976a,a10980a,a10981a,a10982a,a10985a,a10989a,a10990a,a10991a,a10994a,a10998a,a10999a,a11000a,a11003a,a11007a,a11008a,a11009a,a11012a,a11016a,a11017a,a11018a,a11021a,a11025a,a11026a,a11027a,a11030a,a11034a,a11035a,a11036a,a11039a,a11043a,a11044a,a11045a,a11048a,a11052a,a11053a,a11054a,a11057a,a11061a,a11062a,a11063a,a11066a,a11070a,a11071a,a11072a,a11075a,a11079a,a11080a,a11081a,a11084a,a11088a,a11089a,a11090a,a11093a,a11097a,a11098a,a11099a,a11102a,a11106a,a11107a,a11108a,a11111a,a11115a,a11116a,a11117a,a11120a,a11124a,a11125a,a11126a,a11129a,a11133a,a11134a,a11135a,a11138a,a11142a,a11143a,a11144a,a11147a,a11151a,a11152a,a11153a,a11156a,a11160a,a11161a,a11162a,a11165a,a11169a,a11170a,a11171a,a11174a,a11178a,a11179a,a11180a,a11183a,a11187a,a11188a,a11189a,a11192a,a11196a,a11197a,a11198a,a11201a,a11205a,a11206a,a11207a,a11210a,a11214a,a11215a,a11216a,a11219a,a11223a,a11224a,a11225a,a11228a,a11232a,a11233a,a11234a,a11237a,a11241a,a11242a,a11243a,a11246a,a11250a,a11251a,a11252a,a11255a,a11259a,a11260a,a11261a,a11264a,a11268a,a11269a,a11270a,a11273a,a11277a,a11278a,a11279a,a11282a,a11286a,a11287a,a11288a,a11291a,a11295a,a11296a,a11297a,a11300a,a11304a,a11305a,a11306a,a11309a,a11313a,a11314a,a11315a,a11318a,a11322a,a11323a,a11324a,a11327a,a11331a,a11332a,a11333a,a11336a,a11340a,a11341a,a11342a,a11345a,a11349a,a11350a,a11351a,a11354a,a11358a,a11359a,a11360a,a11363a,a11367a,a11368a,a11369a,a11372a,a11376a,a11377a,a11378a,a11381a,a11385a,a11386a,a11387a,a11390a,a11394a,a11395a,a11396a,a11399a,a11403a,a11404a,a11405a,a11408a,a11412a,a11413a,a11414a,a11417a,a11421a,a11422a,a11423a,a11426a,a11430a,a11431a,a11432a,a11435a,a11439a,a11440a,a11441a,a11444a,a11448a,a11449a,a11450a,a11453a,a11457a,a11458a,a11459a,a11462a,a11466a,a11467a,a11468a,a11471a,a11475a,a11476a,a11477a,a11480a,a11484a,a11485a,a11486a,a11489a,a11493a,a11494a,a11495a,a11498a,a11502a,a11503a,a11504a,a11507a,a11511a,a11512a,a11513a,a11516a,a11520a,a11521a,a11522a,a11525a,a11529a,a11530a,a11531a,a11534a,a11538a,a11539a,a11540a,a11543a,a11547a,a11548a,a11549a,a11552a,a11556a,a11557a,a11558a,a11561a,a11565a,a11566a,a11567a,a11570a,a11574a,a11575a,a11576a,a11579a,a11583a,a11584a,a11585a,a11588a,a11592a,a11593a,a11594a,a11597a,a11601a,a11602a,a11603a,a11606a,a11610a,a11611a,a11612a,a11615a,a11619a,a11620a,a11621a,a11624a,a11628a,a11629a,a11630a,a11633a,a11637a,a11638a,a11639a,a11642a,a11646a,a11647a,a11648a,a11651a,a11655a,a11656a,a11657a,a11660a,a11664a,a11665a,a11666a,a11669a,a11673a,a11674a,a11675a,a11678a,a11682a,a11683a,a11684a,a11687a,a11691a,a11692a,a11693a,a11696a,a11700a,a11701a,a11702a,a11705a,a11709a,a11710a,a11711a,a11714a,a11718a,a11719a,a11720a,a11723a,a11727a,a11728a,a11729a,a11732a,a11736a,a11737a,a11738a,a11741a,a11745a,a11746a,a11747a,a11750a,a11754a,a11755a,a11756a,a11759a,a11763a,a11764a,a11765a,a11768a,a11772a,a11773a,a11774a,a11777a,a11781a,a11782a,a11783a,a11786a,a11790a,a11791a,a11792a,a11795a,a11799a,a11800a,a11801a,a11804a,a11808a,a11809a,a11810a,a11813a,a11817a,a11818a,a11819a,a11822a,a11826a,a11827a,a11828a,a11831a,a11835a,a11836a,a11837a,a11840a,a11844a,a11845a,a11846a,a11849a,a11853a,a11854a,a11855a,a11858a,a11862a,a11863a,a11864a,a11867a,a11871a,a11872a,a11873a,a11876a,a11880a,a11881a,a11882a,a11885a,a11889a,a11890a,a11891a,a11894a,a11898a,a11899a,a11900a,a11903a,a11907a,a11908a,a11909a,a11912a,a11916a,a11917a,a11918a,a11921a,a11925a,a11926a,a11927a,a11930a,a11934a,a11935a,a11936a,a11939a,a11943a,a11944a,a11945a,a11948a,a11952a,a11953a,a11954a,a11957a,a11961a,a11962a,a11963a,a11966a,a11970a,a11971a,a11972a,a11975a,a11979a,a11980a,a11981a,a11984a,a11988a,a11989a,a11990a,a11993a,a11997a,a11998a,a11999a,a12002a,a12006a,a12007a,a12008a,a12011a,a12015a,a12016a,a12017a,a12020a,a12024a,a12025a,a12026a,a12029a,a12033a,a12034a,a12035a,a12038a,a12042a,a12043a,a12044a,a12047a,a12051a,a12052a,a12053a,a12056a,a12060a,a12061a,a12062a,a12065a,a12069a,a12070a,a12071a,a12074a,a12078a,a12079a,a12080a,a12083a,a12087a,a12088a,a12089a,a12092a,a12096a,a12097a,a12098a,a12101a,a12105a,a12106a,a12107a,a12110a,a12114a,a12115a,a12116a,a12119a,a12123a,a12124a,a12125a,a12128a,a12132a,a12133a,a12134a,a12137a,a12141a,a12142a,a12143a,a12146a,a12150a,a12151a,a12152a,a12155a,a12159a,a12160a,a12161a,a12164a,a12168a,a12169a,a12170a,a12173a,a12177a,a12178a,a12179a,a12182a,a12186a,a12187a,a12188a,a12191a,a12195a,a12196a,a12197a,a12200a,a12204a,a12205a,a12206a,a12209a,a12213a,a12214a,a12215a,a12218a,a12222a,a12223a,a12224a,a12227a,a12231a,a12232a,a12233a,a12236a,a12240a,a12241a,a12242a,a12245a,a12249a,a12250a,a12251a,a12254a,a12258a,a12259a,a12260a,a12263a,a12267a,a12268a,a12269a,a12272a,a12276a,a12277a,a12278a,a12281a,a12285a,a12286a,a12287a,a12290a,a12294a,a12295a,a12296a,a12299a,a12303a,a12304a,a12305a,a12308a,a12312a,a12313a,a12314a,a12317a,a12321a,a12322a,a12323a,a12326a,a12330a,a12331a,a12332a,a12335a,a12339a,a12340a,a12341a,a12344a,a12348a,a12349a,a12350a,a12353a,a12357a,a12358a,a12359a,a12362a,a12366a,a12367a,a12368a,a12371a,a12375a,a12376a,a12377a,a12380a,a12384a,a12385a,a12386a,a12389a,a12393a,a12394a,a12395a,a12398a,a12402a,a12403a,a12404a,a12407a,a12411a,a12412a,a12413a,a12416a,a12420a,a12421a,a12422a,a12425a,a12429a,a12430a,a12431a,a12434a,a12438a,a12439a,a12440a,a12443a,a12447a,a12448a,a12449a,a12452a,a12456a,a12457a,a12458a,a12461a,a12465a,a12466a,a12467a,a12470a,a12474a,a12475a,a12476a,a12479a,a12483a,a12484a,a12485a,a12488a,a12492a,a12493a,a12494a,a12497a,a12501a,a12502a,a12503a,a12506a,a12510a,a12511a,a12512a,a12515a,a12519a,a12520a,a12521a,a12524a,a12528a,a12529a,a12530a,a12533a,a12537a,a12538a,a12539a,a12542a,a12546a,a12547a,a12548a,a12551a,a12555a,a12556a,a12557a,a12560a,a12564a,a12565a,a12566a,a12569a,a12573a,a12574a,a12575a,a12578a,a12582a,a12583a,a12584a,a12587a,a12591a,a12592a,a12593a,a12596a,a12600a,a12601a,a12602a,a12605a,a12609a,a12610a,a12611a,a12614a,a12618a,a12619a,a12620a,a12623a,a12627a,a12628a,a12629a,a12632a,a12636a,a12637a,a12638a,a12641a,a12645a,a12646a,a12647a,a12650a,a12654a,a12655a,a12656a,a12659a,a12663a,a12664a,a12665a,a12668a,a12672a,a12673a,a12674a,a12677a,a12681a,a12682a,a12683a,a12686a,a12690a,a12691a,a12692a,a12695a,a12699a,a12700a,a12701a,a12704a,a12708a,a12709a,a12710a,a12713a,a12717a,a12718a,a12719a,a12722a,a12726a,a12727a,a12728a,a12731a,a12735a,a12736a,a12737a,a12740a,a12744a,a12745a,a12746a,a12749a,a12753a,a12754a,a12755a,a12758a,a12762a,a12763a,a12764a,a12767a,a12771a,a12772a,a12773a,a12776a,a12780a,a12781a,a12782a,a12785a,a12789a,a12790a,a12791a,a12794a,a12798a,a12799a,a12800a,a12803a,a12807a,a12808a,a12809a,a12812a,a12816a,a12817a,a12818a,a12821a,a12825a,a12826a,a12827a,a12830a,a12834a,a12835a,a12836a,a12839a,a12843a,a12844a,a12845a,a12848a,a12852a,a12853a,a12854a,a12857a,a12861a,a12862a,a12863a,a12866a,a12870a,a12871a,a12872a,a12875a,a12879a,a12880a,a12881a,a12884a,a12888a,a12889a,a12890a,a12893a,a12897a,a12898a,a12899a,a12902a,a12906a,a12907a,a12908a,a12911a,a12915a,a12916a,a12917a,a12920a,a12924a,a12925a,a12926a,a12929a,a12933a,a12934a,a12935a,a12938a,a12942a,a12943a,a12944a,a12947a,a12951a,a12952a,a12953a,a12956a,a12960a,a12961a,a12962a,a12965a,a12969a,a12970a,a12971a,a12974a,a12978a,a12979a,a12980a,a12983a,a12987a,a12988a,a12989a,a12992a,a12996a,a12997a,a12998a,a13001a,a13005a,a13006a,a13007a,a13010a,a13014a,a13015a,a13016a,a13019a,a13023a,a13024a,a13025a,a13028a,a13032a,a13033a,a13034a,a13037a,a13041a,a13042a,a13043a,a13046a,a13050a,a13051a,a13052a,a13055a,a13059a,a13060a,a13061a,a13064a,a13068a,a13069a,a13070a,a13073a,a13077a,a13078a,a13079a,a13082a,a13086a,a13087a,a13088a,a13091a,a13095a,a13096a,a13097a,a13100a,a13104a,a13105a,a13106a,a13109a,a13113a,a13114a,a13115a,a13118a,a13122a,a13123a,a13124a,a13127a,a13131a,a13132a,a13133a,a13136a,a13140a,a13141a,a13142a,a13145a,a13149a,a13150a,a13151a,a13154a,a13158a,a13159a,a13160a,a13163a,a13167a,a13168a,a13169a,a13172a,a13176a,a13177a,a13178a,a13181a,a13185a,a13186a,a13187a,a13190a,a13194a,a13195a,a13196a,a13199a,a13203a,a13204a,a13205a,a13208a,a13212a,a13213a,a13214a,a13217a,a13221a,a13222a,a13223a,a13226a,a13230a,a13231a,a13232a,a13235a,a13239a,a13240a,a13241a,a13244a,a13248a,a13249a,a13250a,a13253a,a13257a,a13258a,a13259a,a13262a,a13266a,a13267a,a13268a,a13271a,a13275a,a13276a,a13277a,a13280a,a13284a,a13285a,a13286a,a13289a,a13293a,a13294a,a13295a,a13298a,a13302a,a13303a,a13304a,a13307a,a13311a,a13312a,a13313a,a13316a,a13320a,a13321a,a13322a,a13325a,a13329a,a13330a,a13331a,a13334a,a13338a,a13339a,a13340a,a13343a,a13347a,a13348a,a13349a,a13352a,a13356a,a13357a,a13358a,a13361a,a13365a,a13366a,a13367a,a13370a,a13374a,a13375a,a13376a,a13379a,a13383a,a13384a,a13385a,a13388a,a13392a,a13393a,a13394a,a13397a,a13401a,a13402a,a13403a,a13406a,a13410a,a13411a,a13412a,a13415a,a13419a,a13420a,a13421a,a13424a,a13428a,a13429a,a13430a,a13433a,a13437a,a13438a,a13439a,a13442a,a13446a,a13447a,a13448a,a13451a,a13455a,a13456a,a13457a,a13460a,a13464a,a13465a,a13466a,a13469a,a13473a,a13474a,a13475a,a13478a,a13482a,a13483a,a13484a,a13487a,a13491a,a13492a,a13493a,a13496a,a13500a,a13501a,a13502a,a13505a,a13509a,a13510a,a13511a,a13514a,a13518a,a13519a,a13520a,a13523a,a13527a,a13528a,a13529a,a13532a,a13536a,a13537a,a13538a,a13541a,a13545a,a13546a,a13547a,a13550a,a13554a,a13555a,a13556a,a13559a,a13563a,a13564a,a13565a,a13568a,a13572a,a13573a,a13574a,a13577a,a13581a,a13582a,a13583a,a13586a,a13590a,a13591a,a13592a,a13595a,a13599a,a13600a,a13601a,a13604a,a13608a,a13609a,a13610a,a13613a,a13617a,a13618a,a13619a,a13622a,a13626a,a13627a,a13628a,a13631a,a13635a,a13636a,a13637a,a13641a,a13642a,a13646a,a13647a,a13648a,a13651a,a13655a,a13656a,a13657a,a13661a,a13662a,a13666a,a13667a,a13668a,a13671a,a13675a,a13676a,a13677a,a13681a,a13682a,a13686a,a13687a,a13688a,a13691a,a13695a,a13696a,a13697a,a13701a,a13702a,a13706a,a13707a,a13708a,a13711a,a13715a,a13716a,a13717a,a13721a,a13722a,a13726a,a13727a,a13728a,a13731a,a13735a,a13736a,a13737a,a13741a,a13742a,a13746a,a13747a,a13748a,a13751a,a13755a,a13756a,a13757a,a13761a,a13762a,a13766a,a13767a,a13768a,a13771a,a13775a,a13776a,a13777a,a13781a,a13782a,a13786a,a13787a,a13788a,a13791a,a13795a,a13796a,a13797a,a13801a,a13802a,a13806a,a13807a,a13808a,a13811a,a13815a,a13816a,a13817a,a13821a,a13822a,a13826a,a13827a,a13828a,a13831a,a13835a,a13836a,a13837a,a13841a,a13842a,a13846a,a13847a,a13848a,a13851a,a13855a,a13856a,a13857a,a13861a,a13862a,a13866a,a13867a,a13868a,a13871a,a13875a,a13876a,a13877a,a13881a,a13882a,a13886a,a13887a,a13888a,a13891a,a13895a,a13896a,a13897a,a13901a,a13902a,a13906a,a13907a,a13908a,a13911a,a13915a,a13916a,a13917a,a13921a,a13922a,a13926a,a13927a,a13928a,a13931a,a13935a,a13936a,a13937a,a13941a,a13942a,a13946a,a13947a,a13948a,a13951a,a13955a,a13956a,a13957a,a13961a,a13962a,a13966a,a13967a,a13968a,a13971a,a13975a,a13976a,a13977a,a13981a,a13982a,a13986a,a13987a,a13988a,a13991a,a13995a,a13996a,a13997a,a14001a,a14002a,a14006a,a14007a,a14008a,a14011a,a14015a,a14016a,a14017a,a14021a,a14022a,a14026a,a14027a,a14028a,a14031a,a14035a,a14036a,a14037a,a14041a,a14042a,a14046a,a14047a,a14048a,a14051a,a14055a,a14056a,a14057a,a14061a,a14062a,a14066a,a14067a,a14068a,a14071a,a14075a,a14076a,a14077a,a14081a,a14082a,a14086a,a14087a,a14088a,a14091a,a14095a,a14096a,a14097a,a14101a,a14102a,a14106a,a14107a,a14108a,a14111a,a14115a,a14116a,a14117a,a14121a,a14122a,a14126a,a14127a,a14128a,a14131a,a14135a,a14136a,a14137a,a14141a,a14142a,a14146a,a14147a,a14148a,a14151a,a14155a,a14156a,a14157a,a14161a,a14162a,a14166a,a14167a,a14168a,a14171a,a14175a,a14176a,a14177a,a14181a,a14182a,a14186a,a14187a,a14188a,a14191a,a14195a,a14196a,a14197a,a14201a,a14202a,a14206a,a14207a,a14208a,a14211a,a14215a,a14216a,a14217a,a14221a,a14222a,a14226a,a14227a,a14228a,a14231a,a14235a,a14236a,a14237a,a14241a,a14242a,a14246a,a14247a,a14248a,a14251a,a14255a,a14256a,a14257a,a14261a,a14262a,a14266a,a14267a,a14268a,a14271a,a14275a,a14276a,a14277a,a14281a,a14282a,a14286a,a14287a,a14288a,a14291a,a14295a,a14296a,a14297a,a14301a,a14302a,a14306a,a14307a,a14308a,a14311a,a14315a,a14316a,a14317a,a14321a,a14322a,a14326a,a14327a,a14328a,a14331a,a14335a,a14336a,a14337a,a14341a,a14342a,a14346a,a14347a,a14348a,a14351a,a14355a,a14356a,a14357a,a14361a,a14362a,a14366a,a14367a,a14368a,a14371a,a14375a,a14376a,a14377a,a14381a,a14382a,a14386a,a14387a,a14388a,a14391a,a14395a,a14396a,a14397a,a14401a,a14402a,a14406a,a14407a,a14408a,a14411a,a14415a,a14416a,a14417a,a14421a,a14422a,a14426a,a14427a,a14428a,a14431a,a14435a,a14436a,a14437a,a14441a,a14442a,a14446a,a14447a,a14448a,a14451a,a14455a,a14456a,a14457a,a14461a,a14462a,a14466a,a14467a,a14468a,a14471a,a14475a,a14476a,a14477a,a14481a,a14482a,a14486a,a14487a,a14488a,a14491a,a14495a,a14496a,a14497a,a14501a,a14502a,a14506a,a14507a,a14508a,a14511a,a14515a,a14516a,a14517a,a14521a,a14522a,a14526a,a14527a,a14528a,a14531a,a14535a,a14536a,a14537a,a14541a,a14542a,a14546a,a14547a,a14548a,a14551a,a14555a,a14556a,a14557a,a14561a,a14562a,a14566a,a14567a,a14568a,a14571a,a14575a,a14576a,a14577a,a14581a,a14582a,a14586a,a14587a,a14588a,a14591a,a14595a,a14596a,a14597a,a14601a,a14602a,a14606a,a14607a,a14608a,a14611a,a14615a,a14616a,a14617a,a14621a,a14622a,a14626a,a14627a,a14628a,a14631a,a14635a,a14636a,a14637a,a14641a,a14642a,a14646a,a14647a,a14648a,a14651a,a14655a,a14656a,a14657a,a14661a,a14662a,a14666a,a14667a,a14668a,a14671a,a14675a,a14676a,a14677a,a14681a,a14682a,a14686a,a14687a,a14688a,a14691a,a14695a,a14696a,a14697a,a14701a,a14702a,a14706a,a14707a,a14708a,a14711a,a14715a,a14716a,a14717a,a14721a,a14722a,a14726a,a14727a,a14728a,a14731a,a14735a,a14736a,a14737a,a14741a,a14742a,a14746a,a14747a,a14748a,a14751a,a14755a,a14756a,a14757a,a14761a,a14762a,a14766a,a14767a,a14768a,a14771a,a14775a,a14776a,a14777a,a14781a,a14782a,a14786a,a14787a,a14788a,a14791a,a14795a,a14796a,a14797a,a14801a,a14802a,a14806a,a14807a,a14808a,a14811a,a14815a,a14816a,a14817a,a14821a,a14822a,a14826a,a14827a,a14828a,a14831a,a14835a,a14836a,a14837a,a14841a,a14842a,a14846a,a14847a,a14848a,a14851a,a14855a,a14856a,a14857a,a14861a,a14862a,a14866a,a14867a,a14868a,a14871a,a14875a,a14876a,a14877a,a14881a,a14882a,a14886a,a14887a,a14888a,a14891a,a14895a,a14896a,a14897a,a14901a,a14902a,a14906a,a14907a,a14908a,a14911a,a14915a,a14916a,a14917a,a14921a,a14922a,a14926a,a14927a,a14928a,a14931a,a14935a,a14936a,a14937a,a14941a,a14942a,a14946a,a14947a,a14948a,a14951a,a14955a,a14956a,a14957a,a14961a,a14962a,a14966a,a14967a,a14968a,a14971a,a14975a,a14976a,a14977a,a14981a,a14982a,a14986a,a14987a,a14988a,a14991a,a14995a,a14996a,a14997a,a15001a,a15002a,a15006a,a15007a,a15008a,a15011a,a15015a,a15016a,a15017a,a15021a,a15022a,a15026a,a15027a,a15028a,a15031a,a15035a,a15036a,a15037a,a15041a,a15042a,a15046a,a15047a,a15048a,a15051a,a15055a,a15056a,a15057a,a15061a,a15062a,a15066a,a15067a,a15068a,a15071a,a15075a,a15076a,a15077a,a15081a,a15082a,a15086a,a15087a,a15088a,a15091a,a15095a,a15096a,a15097a,a15101a,a15102a,a15106a,a15107a,a15108a,a15111a,a15115a,a15116a,a15117a,a15121a,a15122a,a15126a,a15127a,a15128a,a15131a,a15135a,a15136a,a15137a,a15141a,a15142a,a15146a,a15147a,a15148a,a15151a,a15155a,a15156a,a15157a,a15161a,a15162a,a15166a,a15167a,a15168a,a15171a,a15175a,a15176a,a15177a,a15181a,a15182a,a15186a,a15187a,a15188a,a15191a,a15195a,a15196a,a15197a,a15201a,a15202a,a15206a,a15207a,a15208a,a15211a,a15215a,a15216a,a15217a,a15221a,a15222a,a15226a,a15227a,a15228a,a15231a,a15235a,a15236a,a15237a,a15241a,a15242a,a15246a,a15247a,a15248a,a15251a,a15255a,a15256a,a15257a,a15261a,a15262a,a15266a,a15267a,a15268a,a15271a,a15275a,a15276a,a15277a,a15281a,a15282a,a15286a,a15287a,a15288a,a15291a,a15295a,a15296a,a15297a,a15301a,a15302a,a15306a,a15307a,a15308a,a15311a,a15315a,a15316a,a15317a,a15321a,a15322a,a15326a,a15327a,a15328a,a15331a,a15335a,a15336a,a15337a,a15341a,a15342a,a15346a,a15347a,a15348a,a15351a,a15355a,a15356a,a15357a,a15361a,a15362a,a15366a,a15367a,a15368a,a15371a,a15375a,a15376a,a15377a,a15381a,a15382a,a15386a,a15387a,a15388a,a15391a,a15395a,a15396a,a15397a,a15401a,a15402a,a15406a,a15407a,a15408a,a15411a,a15415a,a15416a,a15417a,a15421a,a15422a,a15426a,a15427a,a15428a,a15431a,a15435a,a15436a,a15437a,a15441a,a15442a,a15446a,a15447a,a15448a,a15451a,a15455a,a15456a,a15457a,a15461a,a15462a,a15466a,a15467a,a15468a,a15471a,a15475a,a15476a,a15477a,a15481a,a15482a,a15486a,a15487a,a15488a,a15491a,a15495a,a15496a,a15497a,a15501a,a15502a,a15506a,a15507a,a15508a,a15511a,a15515a,a15516a,a15517a,a15521a,a15522a,a15526a,a15527a,a15528a,a15531a,a15535a,a15536a,a15537a,a15541a,a15542a,a15546a,a15547a,a15548a,a15551a,a15555a,a15556a,a15557a,a15561a,a15562a,a15566a,a15567a,a15568a,a15571a,a15575a,a15576a,a15577a,a15581a,a15582a,a15586a,a15587a,a15588a,a15591a,a15595a,a15596a,a15597a,a15601a,a15602a,a15606a,a15607a,a15608a,a15611a,a15615a,a15616a,a15617a,a15621a,a15622a,a15626a,a15627a,a15628a,a15631a,a15635a,a15636a,a15637a,a15641a,a15642a,a15646a,a15647a,a15648a,a15651a,a15655a,a15656a,a15657a,a15661a,a15662a,a15666a,a15667a,a15668a,a15671a,a15675a,a15676a,a15677a,a15681a,a15682a,a15686a,a15687a,a15688a,a15691a,a15695a,a15696a,a15697a,a15701a,a15702a,a15706a,a15707a,a15708a,a15711a,a15715a,a15716a,a15717a,a15721a,a15722a,a15726a,a15727a,a15728a,a15731a,a15735a,a15736a,a15737a,a15741a,a15742a,a15746a,a15747a,a15748a,a15751a,a15755a,a15756a,a15757a,a15761a,a15762a,a15766a,a15767a,a15768a,a15771a,a15775a,a15776a,a15777a,a15781a,a15782a,a15786a,a15787a,a15788a,a15791a,a15795a,a15796a,a15797a,a15801a,a15802a,a15806a,a15807a,a15808a,a15811a,a15815a,a15816a,a15817a,a15821a,a15822a,a15826a,a15827a,a15828a,a15831a,a15835a,a15836a,a15837a,a15841a,a15842a,a15846a,a15847a,a15848a,a15851a,a15855a,a15856a,a15857a,a15861a,a15862a,a15866a,a15867a,a15868a,a15871a,a15875a,a15876a,a15877a,a15881a,a15882a,a15886a,a15887a,a15888a,a15891a,a15895a,a15896a,a15897a,a15901a,a15902a,a15906a,a15907a,a15908a,a15911a,a15915a,a15916a,a15917a,a15921a,a15922a,a15926a,a15927a,a15928a,a15931a,a15935a,a15936a,a15937a,a15941a,a15942a,a15946a,a15947a,a15948a,a15951a,a15955a,a15956a,a15957a,a15961a,a15962a,a15966a,a15967a,a15968a,a15971a,a15975a,a15976a,a15977a,a15981a,a15982a,a15986a,a15987a,a15988a,a15991a,a15995a,a15996a,a15997a,a16001a,a16002a,a16006a,a16007a,a16008a,a16011a,a16015a,a16016a,a16017a,a16021a,a16022a,a16026a,a16027a,a16028a,a16031a,a16035a,a16036a,a16037a,a16041a,a16042a,a16046a,a16047a,a16048a,a16051a,a16055a,a16056a,a16057a,a16061a,a16062a,a16066a,a16067a,a16068a,a16071a,a16075a,a16076a,a16077a,a16081a,a16082a,a16086a,a16087a,a16088a,a16091a,a16095a,a16096a,a16097a,a16101a,a16102a,a16106a,a16107a,a16108a,a16111a,a16115a,a16116a,a16117a,a16121a,a16122a,a16126a,a16127a,a16128a,a16131a,a16135a,a16136a,a16137a,a16141a,a16142a,a16146a,a16147a,a16148a,a16151a,a16155a,a16156a,a16157a,a16161a,a16162a,a16166a,a16167a,a16168a,a16171a,a16175a,a16176a,a16177a,a16181a,a16182a,a16186a,a16187a,a16188a,a16191a,a16195a,a16196a,a16197a,a16201a,a16202a,a16206a,a16207a,a16208a,a16211a,a16215a,a16216a,a16217a,a16221a,a16222a,a16226a,a16227a,a16228a,a16231a,a16235a,a16236a,a16237a,a16241a,a16242a,a16246a,a16247a,a16248a,a16251a,a16255a,a16256a,a16257a,a16261a,a16262a,a16266a,a16267a,a16268a,a16271a,a16275a,a16276a,a16277a,a16281a,a16282a,a16286a,a16287a,a16288a,a16291a,a16295a,a16296a,a16297a,a16301a,a16302a,a16306a,a16307a,a16308a,a16311a,a16315a,a16316a,a16317a,a16321a,a16322a,a16326a,a16327a,a16328a,a16331a,a16335a,a16336a,a16337a,a16341a,a16342a,a16346a,a16347a,a16348a,a16351a,a16355a,a16356a,a16357a,a16361a,a16362a,a16366a,a16367a,a16368a,a16371a,a16375a,a16376a,a16377a,a16381a,a16382a,a16386a,a16387a,a16388a,a16391a,a16395a,a16396a,a16397a,a16401a,a16402a,a16406a,a16407a,a16408a,a16411a,a16415a,a16416a,a16417a,a16421a,a16422a,a16426a,a16427a,a16428a,a16431a,a16435a,a16436a,a16437a,a16441a,a16442a,a16446a,a16447a,a16448a,a16451a,a16455a,a16456a,a16457a,a16461a,a16462a,a16466a,a16467a,a16468a,a16471a,a16475a,a16476a,a16477a,a16481a,a16482a,a16486a,a16487a,a16488a,a16491a,a16495a,a16496a,a16497a,a16501a,a16502a,a16506a,a16507a,a16508a,a16511a,a16515a,a16516a,a16517a,a16521a,a16522a,a16526a,a16527a,a16528a,a16531a,a16535a,a16536a,a16537a,a16541a,a16542a,a16546a,a16547a,a16548a,a16551a,a16555a,a16556a,a16557a,a16561a,a16562a,a16566a,a16567a,a16568a,a16571a,a16575a,a16576a,a16577a,a16581a,a16582a,a16586a,a16587a,a16588a,a16591a,a16595a,a16596a,a16597a,a16601a,a16602a,a16606a,a16607a,a16608a,a16611a,a16615a,a16616a,a16617a,a16621a,a16622a,a16626a,a16627a,a16628a,a16631a,a16635a,a16636a,a16637a,a16641a,a16642a,a16646a,a16647a,a16648a,a16651a,a16655a,a16656a,a16657a,a16661a,a16662a,a16666a,a16667a,a16668a,a16671a,a16675a,a16676a,a16677a,a16681a,a16682a,a16686a,a16687a,a16688a,a16691a,a16695a,a16696a,a16697a,a16701a,a16702a,a16706a,a16707a,a16708a,a16711a,a16715a,a16716a,a16717a,a16721a,a16722a,a16726a,a16727a,a16728a,a16731a,a16735a,a16736a,a16737a,a16741a,a16742a,a16746a,a16747a,a16748a,a16751a,a16755a,a16756a,a16757a,a16761a,a16762a,a16766a,a16767a,a16768a,a16771a,a16775a,a16776a,a16777a,a16781a,a16782a,a16786a,a16787a,a16788a,a16791a,a16795a,a16796a,a16797a,a16801a,a16802a,a16806a,a16807a,a16808a,a16811a,a16815a,a16816a,a16817a,a16821a,a16822a,a16826a,a16827a,a16828a,a16831a,a16835a,a16836a,a16837a,a16841a,a16842a,a16846a,a16847a,a16848a,a16851a,a16855a,a16856a,a16857a,a16861a,a16862a,a16866a,a16867a,a16868a,a16871a,a16875a,a16876a,a16877a,a16881a,a16882a,a16886a,a16887a,a16888a,a16891a,a16895a,a16896a,a16897a,a16901a,a16902a,a16906a,a16907a,a16908a,a16911a,a16915a,a16916a,a16917a,a16921a,a16922a,a16926a,a16927a,a16928a,a16931a,a16935a,a16936a,a16937a,a16941a,a16942a,a16946a,a16947a,a16948a,a16951a,a16955a,a16956a,a16957a,a16961a,a16962a,a16966a,a16967a,a16968a,a16971a,a16975a,a16976a,a16977a,a16981a,a16982a,a16986a,a16987a,a16988a,a16991a,a16995a,a16996a,a16997a,a17001a,a17002a,a17006a,a17007a,a17008a,a17011a,a17015a,a17016a,a17017a,a17021a,a17022a,a17026a,a17027a,a17028a,a17031a,a17035a,a17036a,a17037a,a17041a,a17042a,a17046a,a17047a,a17048a,a17051a,a17055a,a17056a,a17057a,a17061a,a17062a,a17066a,a17067a,a17068a,a17071a,a17075a,a17076a,a17077a,a17081a,a17082a,a17086a,a17087a,a17088a,a17091a,a17095a,a17096a,a17097a,a17101a,a17102a,a17106a,a17107a,a17108a,a17111a,a17115a,a17116a,a17117a,a17121a,a17122a,a17126a,a17127a,a17128a,a17131a,a17135a,a17136a,a17137a,a17141a,a17142a,a17146a,a17147a,a17148a,a17151a,a17155a,a17156a,a17157a,a17161a,a17162a,a17166a,a17167a,a17168a,a17171a,a17175a,a17176a,a17177a,a17181a,a17182a,a17186a,a17187a,a17188a,a17191a,a17195a,a17196a,a17197a,a17201a,a17202a,a17206a,a17207a,a17208a,a17211a,a17215a,a17216a,a17217a,a17221a,a17222a,a17226a,a17227a,a17228a,a17231a,a17235a,a17236a,a17237a,a17241a,a17242a,a17246a,a17247a,a17248a,a17251a,a17255a,a17256a,a17257a,a17261a,a17262a,a17266a,a17267a,a17268a,a17271a,a17275a,a17276a,a17277a,a17281a,a17282a,a17286a,a17287a,a17288a,a17291a,a17295a,a17296a,a17297a,a17301a,a17302a,a17306a,a17307a,a17308a,a17311a,a17315a,a17316a,a17317a,a17321a,a17322a,a17326a,a17327a,a17328a,a17331a,a17335a,a17336a,a17337a,a17341a,a17342a,a17346a,a17347a,a17348a,a17351a,a17355a,a17356a,a17357a,a17361a,a17362a,a17366a,a17367a,a17368a,a17371a,a17375a,a17376a,a17377a,a17381a,a17382a,a17386a,a17387a,a17388a,a17391a,a17395a,a17396a,a17397a,a17401a,a17402a,a17406a,a17407a,a17408a,a17411a,a17415a,a17416a,a17417a,a17421a,a17422a,a17426a,a17427a,a17428a,a17432a,a17433a,a17437a,a17438a,a17439a,a17443a,a17444a,a17448a,a17449a,a17450a,a17454a,a17455a,a17459a,a17460a,a17461a,a17465a,a17466a,a17470a,a17471a,a17472a,a17476a,a17477a,a17481a,a17482a,a17483a,a17487a,a17488a,a17492a,a17493a,a17494a,a17498a,a17499a,a17503a,a17504a,a17505a,a17509a,a17510a,a17514a,a17515a,a17516a,a17520a,a17521a,a17525a,a17526a,a17527a,a17531a,a17532a,a17536a,a17537a,a17538a,a17542a,a17543a,a17547a,a17548a,a17549a,a17553a,a17554a,a17558a,a17559a,a17560a,a17564a,a17565a,a17569a,a17570a,a17571a,a17575a,a17576a,a17580a,a17581a,a17582a,a17586a,a17587a,a17591a,a17592a,a17593a,a17597a,a17598a,a17602a,a17603a,a17604a,a17608a,a17609a,a17613a,a17614a,a17615a,a17619a,a17620a,a17624a,a17625a,a17626a,a17630a,a17631a,a17635a,a17636a,a17637a,a17641a,a17642a,a17646a,a17647a,a17648a,a17652a,a17653a,a17657a,a17658a,a17659a,a17663a,a17664a,a17668a,a17669a,a17670a,a17674a,a17675a,a17679a,a17680a,a17681a,a17685a,a17686a,a17690a,a17691a,a17692a,a17696a,a17697a,a17701a,a17702a,a17703a,a17707a,a17708a,a17712a,a17713a,a17714a,a17718a,a17719a,a17723a,a17724a,a17725a,a17729a,a17730a,a17734a,a17735a,a17736a,a17740a,a17741a,a17745a,a17746a,a17747a,a17751a,a17752a,a17756a,a17757a,a17758a,a17762a,a17763a,a17767a,a17768a,a17769a,a17773a,a17774a,a17778a,a17779a,a17780a,a17784a,a17785a,a17789a,a17790a,a17791a,a17795a,a17796a,a17800a,a17801a,a17802a,a17806a,a17807a,a17811a,a17812a,a17813a,a17817a,a17818a,a17822a,a17823a,a17824a,a17828a,a17829a,a17833a,a17834a,a17835a,a17839a,a17840a,a17844a,a17845a,a17846a,a17850a,a17851a,a17855a,a17856a,a17857a,a17861a,a17862a,a17866a,a17867a,a17868a,a17872a,a17873a,a17877a,a17878a,a17879a,a17883a,a17884a,a17888a,a17889a,a17890a,a17894a,a17895a,a17899a,a17900a,a17901a,a17905a,a17906a,a17910a,a17911a,a17912a,a17916a,a17917a,a17921a,a17922a,a17923a,a17927a,a17928a,a17932a,a17933a,a17934a,a17938a,a17939a,a17943a,a17944a,a17945a,a17949a,a17950a,a17954a,a17955a,a17956a,a17960a,a17961a,a17965a,a17966a,a17967a,a17971a,a17972a,a17976a,a17977a,a17978a,a17982a,a17983a,a17987a,a17988a,a17989a,a17993a,a17994a,a17998a,a17999a,a18000a,a18004a,a18005a,a18009a,a18010a,a18011a,a18015a,a18016a,a18020a,a18021a,a18022a,a18026a,a18027a,a18031a,a18032a,a18033a,a18037a,a18038a,a18042a,a18043a,a18044a,a18048a,a18049a,a18053a,a18054a,a18055a,a18059a,a18060a,a18064a,a18065a,a18066a,a18070a,a18071a,a18075a,a18076a,a18077a,a18081a,a18082a,a18086a,a18087a,a18088a,a18092a,a18093a,a18097a,a18098a,a18099a,a18103a,a18104a,a18108a,a18109a,a18110a,a18114a,a18115a,a18119a,a18120a,a18121a,a18125a,a18126a,a18130a,a18131a,a18132a,a18136a,a18137a,a18141a,a18142a,a18143a,a18147a,a18148a,a18152a,a18153a,a18154a,a18158a,a18159a,a18163a,a18164a,a18165a,a18169a,a18170a,a18174a,a18175a,a18176a,a18180a,a18181a,a18185a,a18186a,a18187a,a18191a,a18192a,a18196a,a18197a,a18198a,a18202a,a18203a,a18207a,a18208a,a18209a,a18213a,a18214a,a18218a,a18219a,a18220a,a18224a,a18225a,a18229a,a18230a,a18231a,a18235a,a18236a,a18240a,a18241a,a18242a,a18246a,a18247a,a18251a,a18252a,a18253a,a18257a,a18258a,a18262a,a18263a,a18264a,a18268a,a18269a,a18273a,a18274a,a18275a,a18279a,a18280a,a18284a,a18285a,a18286a,a18290a,a18291a,a18295a,a18296a,a18297a,a18301a,a18302a,a18306a,a18307a,a18308a,a18312a,a18313a,a18317a,a18318a,a18319a,a18323a,a18324a,a18328a,a18329a,a18330a,a18334a,a18335a,a18339a,a18340a,a18341a,a18345a,a18346a,a18350a,a18351a,a18352a,a18356a,a18357a,a18361a,a18362a,a18363a,a18367a,a18368a,a18372a,a18373a,a18374a,a18378a,a18379a,a18383a,a18384a,a18385a,a18389a,a18390a,a18394a,a18395a,a18396a,a18400a,a18401a,a18405a,a18406a,a18407a,a18411a,a18412a,a18416a,a18417a,a18418a,a18422a,a18423a,a18427a,a18428a,a18429a,a18433a,a18434a,a18438a,a18439a,a18440a,a18444a,a18445a,a18449a,a18450a,a18451a,a18455a,a18456a,a18460a,a18461a,a18462a,a18466a,a18467a,a18471a,a18472a,a18473a,a18477a,a18478a,a18482a,a18483a,a18484a,a18488a,a18489a,a18493a,a18494a,a18495a,a18499a,a18500a,a18504a,a18505a,a18506a,a18510a,a18511a,a18515a,a18516a,a18517a,a18521a,a18522a,a18526a,a18527a,a18528a,a18532a,a18533a,a18537a,a18538a,a18539a,a18543a,a18544a,a18548a,a18549a,a18550a,a18554a,a18555a,a18559a,a18560a,a18561a,a18565a,a18566a,a18570a,a18571a,a18572a,a18576a,a18577a,a18581a,a18582a,a18583a,a18587a,a18588a,a18592a,a18593a,a18594a,a18598a,a18599a,a18603a,a18604a,a18605a,a18609a,a18610a,a18614a,a18615a,a18616a,a18620a,a18621a,a18625a,a18626a,a18627a,a18631a,a18632a,a18636a,a18637a,a18638a,a18642a,a18643a,a18647a,a18648a,a18649a,a18653a,a18654a,a18658a,a18659a,a18660a,a18664a,a18665a,a18669a,a18670a,a18671a,a18675a,a18676a,a18680a,a18681a,a18682a,a18686a,a18687a,a18691a,a18692a,a18693a,a18697a,a18698a,a18702a,a18703a,a18704a,a18708a,a18709a,a18713a,a18714a,a18715a,a18719a,a18720a,a18724a,a18725a,a18726a,a18730a,a18731a,a18735a,a18736a,a18737a,a18741a,a18742a,a18746a,a18747a,a18748a,a18752a,a18753a,a18757a,a18758a,a18759a,a18763a,a18764a,a18768a,a18769a,a18770a,a18774a,a18775a,a18779a,a18780a,a18781a,a18785a,a18786a,a18790a,a18791a,a18792a,a18796a,a18797a,a18801a,a18802a,a18803a,a18807a,a18808a,a18812a,a18813a,a18814a,a18818a,a18819a,a18823a,a18824a,a18825a,a18829a,a18830a,a18834a,a18835a,a18836a,a18840a,a18841a,a18845a,a18846a,a18847a,a18851a,a18852a,a18856a,a18857a,a18858a,a18862a,a18863a,a18867a,a18868a,a18869a,a18873a,a18874a,a18878a,a18879a,a18880a,a18884a,a18885a,a18889a,a18890a,a18891a,a18895a,a18896a,a18900a,a18901a,a18902a,a18906a,a18907a,a18911a,a18912a,a18913a,a18917a,a18918a,a18922a,a18923a,a18924a,a18928a,a18929a,a18933a,a18934a,a18935a,a18939a,a18940a,a18944a,a18945a,a18946a,a18950a,a18951a,a18955a,a18956a,a18957a,a18961a,a18962a,a18966a,a18967a,a18968a,a18972a,a18973a,a18977a,a18978a,a18979a,a18983a,a18984a,a18988a,a18989a,a18990a,a18994a,a18995a,a18999a,a19000a,a19001a,a19005a,a19006a,a19010a,a19011a,a19012a,a19016a,a19017a,a19021a,a19022a,a19023a,a19027a,a19028a,a19032a,a19033a,a19034a,a19038a,a19039a,a19043a,a19044a,a19045a,a19049a,a19050a,a19054a,a19055a,a19056a,a19060a,a19061a,a19065a,a19066a,a19067a,a19071a,a19072a,a19076a,a19077a,a19078a,a19082a,a19083a,a19087a,a19088a,a19089a,a19093a,a19094a,a19098a,a19099a,a19100a,a19104a,a19105a,a19109a,a19110a,a19111a,a19115a,a19116a,a19120a,a19121a,a19122a,a19126a,a19127a,a19131a,a19132a,a19133a,a19137a,a19138a,a19142a,a19143a,a19144a,a19148a,a19149a,a19153a,a19154a,a19155a,a19159a,a19160a,a19164a,a19165a,a19166a,a19170a,a19171a,a19175a,a19176a,a19177a,a19181a,a19182a,a19186a,a19187a,a19188a,a19192a,a19193a,a19197a,a19198a,a19199a,a19203a,a19204a,a19208a,a19209a,a19210a,a19214a,a19215a,a19219a,a19220a,a19221a,a19225a,a19226a,a19230a,a19231a,a19232a,a19236a,a19237a,a19241a,a19242a,a19243a,a19247a,a19248a,a19252a,a19253a,a19254a,a19258a,a19259a,a19263a,a19264a,a19265a,a19269a,a19270a,a19274a,a19275a,a19276a,a19280a,a19281a,a19285a,a19286a,a19287a,a19291a,a19292a,a19296a,a19297a,a19298a,a19302a,a19303a,a19307a,a19308a,a19309a,a19313a,a19314a,a19318a,a19319a,a19320a,a19324a,a19325a,a19329a,a19330a,a19331a,a19335a,a19336a,a19340a,a19341a,a19342a,a19346a,a19347a,a19351a,a19352a,a19353a,a19357a,a19358a,a19362a,a19363a,a19364a,a19368a,a19369a,a19373a,a19374a,a19375a,a19379a,a19380a,a19384a,a19385a,a19386a,a19390a,a19391a,a19395a,a19396a,a19397a,a19401a,a19402a,a19406a,a19407a,a19408a,a19412a,a19413a,a19417a,a19418a,a19419a,a19423a,a19424a,a19428a,a19429a,a19430a,a19434a,a19435a,a19439a,a19440a,a19441a,a19445a,a19446a,a19450a,a19451a,a19452a,a19456a,a19457a,a19461a,a19462a,a19463a,a19467a,a19468a,a19472a,a19473a,a19474a,a19478a,a19479a,a19483a,a19484a,a19485a,a19489a,a19490a,a19494a,a19495a,a19496a,a19500a,a19501a,a19505a,a19506a,a19507a,a19511a,a19512a,a19516a,a19517a,a19518a,a19522a,a19523a,a19527a,a19528a,a19529a,a19533a,a19534a,a19538a,a19539a,a19540a,a19544a,a19545a,a19549a,a19550a,a19551a,a19555a,a19556a,a19560a,a19561a,a19562a,a19566a,a19567a,a19571a,a19572a,a19573a,a19577a,a19578a,a19582a,a19583a,a19584a,a19588a,a19589a,a19593a,a19594a,a19595a,a19599a,a19600a,a19604a,a19605a,a19606a,a19610a,a19611a,a19615a,a19616a,a19617a,a19621a,a19622a,a19626a,a19627a,a19628a,a19632a,a19633a,a19637a,a19638a,a19639a,a19643a,a19644a,a19648a,a19649a,a19650a,a19654a,a19655a,a19659a,a19660a,a19661a,a19665a,a19666a,a19670a,a19671a,a19672a,a19676a,a19677a,a19681a,a19682a,a19683a,a19687a,a19688a,a19692a,a19693a,a19694a,a19698a,a19699a,a19703a,a19704a,a19705a,a19709a,a19710a,a19714a,a19715a,a19716a,a19720a,a19721a,a19725a,a19726a,a19727a,a19731a,a19732a,a19736a,a19737a,a19738a,a19742a,a19743a,a19747a,a19748a,a19749a,a19753a,a19754a,a19758a,a19759a,a19760a,a19764a,a19765a,a19769a,a19770a,a19771a,a19775a,a19776a,a19780a,a19781a,a19782a,a19786a,a19787a,a19791a,a19792a,a19793a,a19797a,a19798a,a19802a,a19803a,a19804a,a19808a,a19809a,a19813a,a19814a,a19815a,a19819a,a19820a,a19824a,a19825a,a19826a,a19830a,a19831a,a19835a,a19836a,a19837a,a19841a,a19842a,a19846a,a19847a,a19848a,a19852a,a19853a,a19857a,a19858a,a19859a,a19863a,a19864a,a19868a,a19869a,a19870a,a19874a,a19875a,a19879a,a19880a,a19881a,a19885a,a19886a,a19890a,a19891a,a19892a,a19896a,a19897a,a19901a,a19902a,a19903a,a19907a,a19908a,a19912a,a19913a,a19914a,a19918a,a19919a,a19923a,a19924a,a19925a,a19929a,a19930a,a19934a,a19935a,a19936a,a19940a,a19941a,a19945a,a19946a,a19947a,a19951a,a19952a,a19956a,a19957a,a19958a,a19962a,a19963a,a19967a,a19968a,a19969a,a19973a,a19974a,a19978a,a19979a,a19980a,a19984a,a19985a,a19989a,a19990a,a19991a,a19995a,a19996a,a20000a,a20001a,a20002a,a20006a,a20007a,a20011a,a20012a,a20013a,a20017a,a20018a,a20022a,a20023a,a20024a,a20028a,a20029a,a20033a,a20034a,a20035a,a20039a,a20040a,a20044a,a20045a,a20046a,a20050a,a20051a,a20055a,a20056a,a20057a,a20061a,a20062a,a20066a,a20067a,a20068a,a20072a,a20073a,a20077a,a20078a,a20079a,a20083a,a20084a,a20088a,a20089a,a20090a,a20094a,a20095a,a20099a,a20100a,a20101a,a20105a,a20106a,a20110a,a20111a,a20112a,a20116a,a20117a,a20121a,a20122a,a20123a,a20127a,a20128a,a20132a,a20133a,a20134a,a20138a,a20139a,a20143a,a20144a,a20145a,a20149a,a20150a,a20154a,a20155a,a20156a,a20160a,a20161a,a20165a,a20166a,a20167a,a20171a,a20172a,a20176a,a20177a,a20178a,a20182a,a20183a,a20187a,a20188a,a20189a,a20193a,a20194a,a20198a,a20199a,a20200a,a20204a,a20205a,a20209a,a20210a,a20211a,a20215a,a20216a,a20220a,a20221a,a20222a,a20226a,a20227a,a20231a,a20232a,a20233a,a20237a,a20238a,a20242a,a20243a,a20244a,a20248a,a20249a,a20253a,a20254a,a20255a,a20259a,a20260a,a20264a,a20265a,a20266a,a20270a,a20271a,a20275a,a20276a,a20277a,a20281a,a20282a,a20286a,a20287a,a20288a,a20292a,a20293a,a20297a,a20298a,a20299a,a20303a,a20304a,a20308a,a20309a,a20310a,a20314a,a20315a,a20319a,a20320a,a20321a,a20325a,a20326a,a20330a,a20331a,a20332a,a20336a,a20337a,a20341a,a20342a,a20343a,a20347a,a20348a,a20352a,a20353a,a20354a,a20358a,a20359a,a20363a,a20364a,a20365a,a20369a,a20370a,a20374a,a20375a,a20376a,a20380a,a20381a,a20385a,a20386a,a20387a,a20391a,a20392a,a20396a,a20397a,a20398a,a20402a,a20403a,a20407a,a20408a,a20409a,a20413a,a20414a,a20418a,a20419a,a20420a,a20424a,a20425a,a20429a,a20430a,a20431a,a20435a,a20436a,a20440a,a20441a,a20442a,a20446a,a20447a,a20451a,a20452a,a20453a,a20457a,a20458a,a20462a,a20463a,a20464a,a20468a,a20469a,a20473a,a20474a,a20475a,a20479a,a20480a,a20484a,a20485a,a20486a,a20490a,a20491a,a20495a,a20496a,a20497a,a20501a,a20502a,a20506a,a20507a,a20508a,a20512a,a20513a,a20517a,a20518a,a20519a,a20523a,a20524a,a20528a,a20529a,a20530a,a20534a,a20535a,a20539a,a20540a,a20541a,a20545a,a20546a,a20550a,a20551a,a20552a,a20556a,a20557a,a20561a,a20562a,a20563a,a20567a,a20568a,a20572a,a20573a,a20574a,a20578a,a20579a,a20583a,a20584a,a20585a,a20589a,a20590a,a20594a,a20595a,a20596a,a20600a,a20601a,a20605a,a20606a,a20607a,a20611a,a20612a,a20616a,a20617a,a20618a,a20622a,a20623a,a20627a,a20628a,a20629a,a20633a,a20634a,a20638a,a20639a,a20640a,a20644a,a20645a,a20649a,a20650a,a20651a,a20655a,a20656a,a20660a,a20661a,a20662a,a20666a,a20667a,a20671a,a20672a,a20673a,a20677a,a20678a,a20682a,a20683a,a20684a,a20688a,a20689a,a20693a,a20694a,a20695a,a20699a,a20700a,a20704a,a20705a,a20706a,a20710a,a20711a,a20715a,a20716a,a20717a,a20721a,a20722a,a20726a,a20727a,a20728a,a20732a,a20733a,a20737a,a20738a,a20739a,a20743a,a20744a,a20748a,a20749a,a20750a,a20754a,a20755a,a20759a,a20760a,a20761a,a20765a,a20766a,a20770a,a20771a,a20772a,a20776a,a20777a,a20781a,a20782a,a20783a,a20787a,a20788a,a20792a,a20793a,a20794a,a20798a,a20799a,a20803a,a20804a,a20805a,a20809a,a20810a,a20814a,a20815a,a20816a,a20820a,a20821a,a20825a,a20826a,a20827a,a20831a,a20832a,a20836a,a20837a,a20838a,a20842a,a20843a,a20847a,a20848a,a20849a,a20853a,a20854a,a20858a,a20859a,a20860a,a20864a,a20865a,a20869a,a20870a,a20871a,a20875a,a20876a,a20880a,a20881a,a20882a,a20886a,a20887a,a20891a,a20892a,a20893a,a20897a,a20898a,a20902a,a20903a,a20904a,a20908a,a20909a,a20913a,a20914a,a20915a,a20919a,a20920a,a20924a,a20925a,a20926a,a20930a,a20931a,a20935a,a20936a,a20937a,a20941a,a20942a,a20946a,a20947a,a20948a,a20952a,a20953a,a20957a,a20958a,a20959a,a20963a,a20964a,a20968a,a20969a,a20970a,a20974a,a20975a,a20979a,a20980a,a20981a,a20985a,a20986a,a20990a,a20991a,a20992a,a20996a,a20997a,a21001a,a21002a,a21003a,a21007a,a21008a,a21012a,a21013a,a21014a,a21018a,a21019a,a21023a,a21024a,a21025a,a21029a,a21030a,a21034a,a21035a,a21036a,a21040a,a21041a,a21045a,a21046a,a21047a,a21051a,a21052a,a21056a,a21057a,a21058a,a21062a,a21063a,a21067a,a21068a,a21069a,a21073a,a21074a,a21078a,a21079a,a21080a,a21084a,a21085a,a21089a,a21090a,a21091a,a21095a,a21096a,a21100a,a21101a,a21102a,a21106a,a21107a,a21111a,a21112a,a21113a,a21117a,a21118a,a21122a,a21123a,a21124a,a21128a,a21129a,a21133a,a21134a,a21135a,a21139a,a21140a,a21144a,a21145a,a21146a,a21150a,a21151a,a21155a,a21156a,a21157a,a21161a,a21162a,a21166a,a21167a,a21168a,a21172a,a21173a,a21177a,a21178a,a21179a,a21183a,a21184a,a21188a,a21189a,a21190a,a21194a,a21195a,a21199a,a21200a,a21201a,a21205a,a21206a,a21210a,a21211a,a21212a,a21216a,a21217a,a21221a,a21222a,a21223a,a21227a,a21228a,a21232a,a21233a,a21234a,a21238a,a21239a,a21243a,a21244a,a21245a,a21249a,a21250a,a21254a,a21255a,a21256a,a21260a,a21261a,a21265a,a21266a,a21267a,a21271a,a21272a,a21276a,a21277a,a21278a,a21282a,a21283a,a21287a,a21288a,a21289a,a21293a,a21294a,a21298a,a21299a,a21300a,a21304a,a21305a,a21309a,a21310a,a21311a,a21315a,a21316a,a21320a,a21321a,a21322a,a21326a,a21327a,a21331a,a21332a,a21333a,a21337a,a21338a,a21342a,a21343a,a21344a,a21348a,a21349a,a21353a,a21354a,a21355a,a21359a,a21360a,a21364a,a21365a,a21366a,a21370a,a21371a,a21375a,a21376a,a21377a,a21381a,a21382a,a21386a,a21387a,a21388a,a21392a,a21393a,a21397a,a21398a,a21399a,a21403a,a21404a,a21408a,a21409a,a21410a,a21414a,a21415a,a21419a,a21420a,a21421a,a21425a,a21426a,a21430a,a21431a,a21432a,a21436a,a21437a,a21441a,a21442a,a21443a,a21447a,a21448a,a21452a,a21453a,a21454a,a21458a,a21459a,a21463a,a21464a,a21465a,a21469a,a21470a,a21474a,a21475a,a21476a,a21480a,a21481a,a21485a,a21486a,a21487a,a21491a,a21492a,a21496a,a21497a,a21498a,a21502a,a21503a,a21507a,a21508a,a21509a,a21513a,a21514a,a21518a,a21519a,a21520a,a21524a,a21525a,a21529a,a21530a,a21531a,a21535a,a21536a,a21540a,a21541a,a21542a,a21546a,a21547a,a21551a,a21552a,a21553a,a21557a,a21558a,a21562a,a21563a,a21564a,a21568a,a21569a,a21573a,a21574a,a21575a,a21579a,a21580a,a21584a,a21585a,a21586a,a21590a,a21591a,a21595a,a21596a,a21597a,a21601a,a21602a,a21606a,a21607a,a21608a,a21612a,a21613a,a21617a,a21618a,a21619a,a21623a,a21624a,a21628a,a21629a,a21630a,a21634a,a21635a,a21639a,a21640a,a21641a,a21645a,a21646a,a21650a,a21651a,a21652a,a21656a,a21657a,a21661a,a21662a,a21663a,a21667a,a21668a,a21672a,a21673a,a21674a,a21678a,a21679a,a21683a,a21684a,a21685a,a21689a,a21690a,a21694a,a21695a,a21696a,a21700a,a21701a,a21705a,a21706a,a21707a,a21711a,a21712a,a21716a,a21717a,a21718a,a21722a,a21723a,a21727a,a21728a,a21729a,a21733a,a21734a,a21738a,a21739a,a21740a,a21744a,a21745a,a21749a,a21750a,a21751a,a21755a,a21756a,a21760a,a21761a,a21762a,a21766a,a21767a,a21771a,a21772a,a21773a,a21777a,a21778a,a21782a,a21783a,a21784a,a21788a,a21789a,a21793a,a21794a,a21795a,a21799a,a21800a,a21804a,a21805a,a21806a,a21810a,a21811a,a21815a,a21816a,a21817a,a21821a,a21822a,a21826a,a21827a,a21828a,a21832a,a21833a,a21837a,a21838a,a21839a,a21843a,a21844a,a21848a,a21849a,a21850a,a21854a,a21855a,a21859a,a21860a,a21861a,a21865a,a21866a,a21870a,a21871a,a21872a,a21876a,a21877a,a21881a,a21882a,a21883a,a21887a,a21888a,a21892a,a21893a,a21894a,a21898a,a21899a,a21903a,a21904a,a21905a,a21909a,a21910a,a21914a,a21915a,a21916a,a21920a,a21921a,a21925a,a21926a,a21927a,a21931a,a21932a,a21936a,a21937a,a21938a,a21942a,a21943a,a21947a,a21948a,a21949a,a21953a,a21954a,a21958a,a21959a,a21960a,a21964a,a21965a,a21969a,a21970a,a21971a,a21975a,a21976a,a21980a,a21981a,a21982a,a21986a,a21987a,a21991a,a21992a,a21993a,a21997a,a21998a,a22002a,a22003a,a22004a,a22008a,a22009a,a22013a,a22014a,a22015a,a22019a,a22020a,a22024a,a22025a,a22026a,a22030a,a22031a,a22035a,a22036a,a22037a,a22041a,a22042a,a22046a,a22047a,a22048a,a22052a,a22053a,a22057a,a22058a,a22059a,a22063a,a22064a,a22068a,a22069a,a22070a,a22074a,a22075a,a22079a,a22080a,a22081a,a22085a,a22086a,a22090a,a22091a,a22092a,a22096a,a22097a,a22101a,a22102a,a22103a,a22107a,a22108a,a22112a,a22113a,a22114a,a22118a,a22119a,a22123a,a22124a,a22125a,a22129a,a22130a,a22134a,a22135a,a22136a,a22140a,a22141a,a22145a,a22146a,a22147a,a22151a,a22152a,a22156a,a22157a,a22158a,a22162a,a22163a,a22167a,a22168a,a22169a,a22173a,a22174a,a22178a,a22179a,a22180a,a22184a,a22185a,a22189a,a22190a,a22191a,a22195a,a22196a,a22200a,a22201a,a22202a,a22206a,a22207a,a22211a,a22212a,a22213a,a22217a,a22218a,a22222a,a22223a,a22224a,a22228a,a22229a,a22233a,a22234a,a22235a,a22239a,a22240a,a22244a,a22245a,a22246a,a22250a,a22251a,a22255a,a22256a,a22257a,a22261a,a22262a,a22266a,a22267a,a22268a,a22272a,a22273a,a22277a,a22278a,a22279a,a22283a,a22284a,a22288a,a22289a,a22290a,a22294a,a22295a,a22299a,a22300a,a22301a,a22305a,a22306a,a22310a,a22311a,a22312a,a22316a,a22317a,a22321a,a22322a,a22323a,a22327a,a22328a,a22332a,a22333a,a22334a,a22338a,a22339a,a22343a,a22344a,a22345a,a22349a,a22350a,a22354a,a22355a,a22356a,a22360a,a22361a,a22365a,a22366a,a22367a,a22371a,a22372a,a22376a,a22377a,a22378a,a22382a,a22383a,a22387a,a22388a,a22389a,a22393a,a22394a,a22398a,a22399a,a22400a,a22404a,a22405a,a22409a,a22410a,a22411a,a22415a,a22416a,a22420a,a22421a,a22422a,a22426a,a22427a,a22431a,a22432a,a22433a,a22437a,a22438a,a22442a,a22443a,a22444a,a22448a,a22449a,a22453a,a22454a,a22455a,a22459a,a22460a,a22464a,a22465a,a22466a,a22470a,a22471a,a22475a,a22476a,a22477a,a22481a,a22482a,a22486a,a22487a,a22488a,a22492a,a22493a,a22497a,a22498a,a22499a,a22503a,a22504a,a22508a,a22509a,a22510a,a22514a,a22515a,a22519a,a22520a,a22521a,a22525a,a22526a,a22530a,a22531a,a22532a,a22536a,a22537a,a22541a,a22542a,a22543a,a22547a,a22548a,a22552a,a22553a,a22554a,a22558a,a22559a,a22563a,a22564a,a22565a,a22569a,a22570a,a22574a,a22575a,a22576a,a22580a,a22581a,a22585a,a22586a,a22587a,a22591a,a22592a,a22596a,a22597a,a22598a,a22602a,a22603a,a22607a,a22608a,a22609a,a22613a,a22614a,a22618a,a22619a,a22620a,a22624a,a22625a,a22629a,a22630a,a22631a,a22635a,a22636a,a22640a,a22641a,a22642a,a22646a,a22647a,a22651a,a22652a,a22653a,a22657a,a22658a,a22662a,a22663a,a22664a,a22668a,a22669a,a22673a,a22674a,a22675a,a22679a,a22680a,a22684a,a22685a,a22686a,a22690a,a22691a,a22695a,a22696a,a22697a,a22701a,a22702a,a22706a,a22707a,a22708a,a22712a,a22713a,a22717a,a22718a,a22719a,a22723a,a22724a,a22728a,a22729a,a22730a,a22734a,a22735a,a22739a,a22740a,a22741a,a22745a,a22746a,a22750a,a22751a,a22752a,a22756a,a22757a,a22761a,a22762a,a22763a,a22767a,a22768a,a22772a,a22773a,a22774a,a22778a,a22779a,a22783a,a22784a,a22785a,a22789a,a22790a,a22794a,a22795a,a22796a,a22800a,a22801a,a22805a,a22806a,a22807a,a22811a,a22812a,a22816a,a22817a,a22818a,a22822a,a22823a,a22827a,a22828a,a22829a,a22833a,a22834a,a22838a,a22839a,a22840a,a22844a,a22845a,a22849a,a22850a,a22851a,a22855a,a22856a,a22860a,a22861a,a22862a,a22866a,a22867a,a22871a,a22872a,a22873a,a22877a,a22878a,a22882a,a22883a,a22884a,a22888a,a22889a,a22893a,a22894a,a22895a,a22899a,a22900a,a22904a,a22905a,a22906a,a22910a,a22911a,a22915a,a22916a,a22917a,a22921a,a22922a,a22926a,a22927a,a22928a,a22932a,a22933a,a22937a,a22938a,a22939a,a22943a,a22944a,a22948a,a22949a,a22950a,a22954a,a22955a,a22959a,a22960a,a22961a,a22965a,a22966a,a22970a,a22971a,a22972a,a22976a,a22977a,a22981a,a22982a,a22983a,a22987a,a22988a,a22992a,a22993a,a22994a,a22998a,a22999a,a23003a,a23004a,a23005a,a23009a,a23010a,a23014a,a23015a,a23016a,a23020a,a23021a,a23025a,a23026a,a23027a,a23031a,a23032a,a23036a,a23037a,a23038a,a23042a,a23043a,a23047a,a23048a,a23049a,a23053a,a23054a,a23058a,a23059a,a23060a,a23064a,a23065a,a23069a,a23070a,a23071a,a23075a,a23076a,a23080a,a23081a,a23082a,a23086a,a23087a,a23091a,a23092a,a23093a,a23097a,a23098a,a23102a,a23103a,a23104a,a23108a,a23109a,a23113a,a23114a,a23115a,a23119a,a23120a,a23124a,a23125a,a23126a,a23130a,a23131a,a23135a,a23136a,a23137a,a23141a,a23142a,a23146a,a23147a,a23148a,a23152a,a23153a,a23157a,a23158a,a23159a,a23163a,a23164a,a23168a,a23169a,a23170a,a23174a,a23175a,a23179a,a23180a,a23181a,a23185a,a23186a,a23190a,a23191a,a23192a,a23196a,a23197a,a23201a,a23202a,a23203a,a23207a,a23208a,a23212a,a23213a,a23214a,a23218a,a23219a,a23223a,a23224a,a23225a,a23229a,a23230a,a23234a,a23235a,a23236a,a23240a,a23241a,a23245a,a23246a,a23247a,a23251a,a23252a,a23256a,a23257a,a23258a,a23262a,a23263a,a23267a,a23268a,a23269a,a23273a,a23274a,a23278a,a23279a,a23280a,a23284a,a23285a,a23289a,a23290a,a23291a,a23295a,a23296a,a23300a,a23301a,a23302a,a23306a,a23307a,a23311a,a23312a,a23313a,a23317a,a23318a,a23322a,a23323a,a23324a,a23328a,a23329a,a23333a,a23334a,a23335a,a23339a,a23340a,a23344a,a23345a,a23346a,a23350a,a23351a,a23355a,a23356a,a23357a,a23361a,a23362a,a23366a,a23367a,a23368a,a23372a,a23373a,a23377a,a23378a,a23379a,a23383a,a23384a,a23388a,a23389a,a23390a,a23394a,a23395a,a23399a,a23400a,a23401a,a23405a,a23406a,a23410a,a23411a,a23412a,a23416a,a23417a,a23421a,a23422a,a23423a,a23427a,a23428a,a23432a,a23433a,a23434a,a23438a,a23439a,a23443a,a23444a,a23445a,a23449a,a23450a,a23454a,a23455a,a23456a,a23460a,a23461a,a23465a,a23466a,a23467a,a23471a,a23472a,a23476a,a23477a,a23478a,a23482a,a23483a,a23487a,a23488a,a23489a,a23493a,a23494a,a23498a,a23499a,a23500a,a23504a,a23505a,a23509a,a23510a,a23511a,a23515a,a23516a,a23520a,a23521a,a23522a,a23526a,a23527a,a23531a,a23532a,a23533a,a23537a,a23538a,a23542a,a23543a,a23544a,a23548a,a23549a,a23553a,a23554a,a23555a,a23559a,a23560a,a23564a,a23565a,a23566a,a23570a,a23571a,a23575a,a23576a,a23577a,a23581a,a23582a,a23586a,a23587a,a23588a,a23592a,a23593a,a23597a,a23598a,a23599a,a23603a,a23604a,a23608a,a23609a,a23610a,a23614a,a23615a,a23619a,a23620a,a23621a,a23625a,a23626a,a23630a,a23631a,a23632a,a23636a,a23637a,a23641a,a23642a,a23643a,a23647a,a23648a,a23652a,a23653a,a23654a,a23658a,a23659a,a23663a,a23664a,a23665a,a23669a,a23670a,a23674a,a23675a,a23676a,a23680a,a23681a,a23685a,a23686a,a23687a,a23691a,a23692a,a23696a,a23697a,a23698a,a23702a,a23703a,a23707a,a23708a,a23709a,a23713a,a23714a,a23718a,a23719a,a23720a,a23724a,a23725a,a23729a,a23730a,a23731a,a23735a,a23736a,a23740a,a23741a,a23742a,a23746a,a23747a,a23751a,a23752a,a23753a,a23757a,a23758a,a23762a,a23763a,a23764a,a23768a,a23769a,a23773a,a23774a,a23775a,a23779a,a23780a,a23784a,a23785a,a23786a,a23790a,a23791a,a23795a,a23796a,a23797a,a23801a,a23802a,a23806a,a23807a,a23808a,a23812a,a23813a,a23817a,a23818a,a23819a,a23823a,a23824a,a23828a,a23829a,a23830a,a23834a,a23835a,a23839a,a23840a,a23841a,a23845a,a23846a,a23850a,a23851a,a23852a,a23856a,a23857a,a23861a,a23862a,a23863a,a23867a,a23868a,a23872a,a23873a,a23874a,a23878a,a23879a,a23883a,a23884a,a23885a,a23889a,a23890a,a23894a,a23895a,a23896a,a23900a,a23901a,a23905a,a23906a,a23907a,a23911a,a23912a,a23916a,a23917a,a23918a,a23922a,a23923a,a23927a,a23928a,a23929a,a23933a,a23934a,a23938a,a23939a,a23940a,a23944a,a23945a,a23949a,a23950a,a23951a,a23955a,a23956a,a23960a,a23961a,a23962a,a23966a,a23967a,a23971a,a23972a,a23973a,a23977a,a23978a,a23982a,a23983a,a23984a,a23988a,a23989a,a23993a,a23994a,a23995a,a23999a,a24000a,a24004a,a24005a,a24006a,a24010a,a24011a,a24015a,a24016a,a24017a,a24021a,a24022a,a24026a,a24027a,a24028a,a24032a,a24033a,a24037a,a24038a,a24039a,a24043a,a24044a,a24048a,a24049a,a24050a,a24054a,a24055a,a24059a,a24060a,a24061a,a24065a,a24066a,a24070a,a24071a,a24072a,a24076a,a24077a,a24081a,a24082a,a24083a,a24087a,a24088a,a24092a,a24093a,a24094a,a24098a,a24099a,a24103a,a24104a,a24105a,a24109a,a24110a,a24114a,a24115a,a24116a,a24120a,a24121a,a24125a,a24126a,a24127a,a24131a,a24132a,a24136a,a24137a,a24138a,a24142a,a24143a,a24147a,a24148a,a24149a,a24153a,a24154a,a24158a,a24159a,a24160a,a24164a,a24165a,a24169a,a24170a,a24171a,a24175a,a24176a,a24180a,a24181a,a24182a,a24186a,a24187a,a24191a,a24192a,a24193a,a24197a,a24198a,a24202a,a24203a,a24204a,a24208a,a24209a,a24213a,a24214a,a24215a,a24219a,a24220a,a24224a,a24225a,a24226a,a24230a,a24231a,a24235a,a24236a,a24237a,a24241a,a24242a,a24246a,a24247a,a24248a,a24252a,a24253a,a24257a,a24258a,a24259a,a24263a,a24264a,a24268a,a24269a,a24270a,a24274a,a24275a,a24279a,a24280a,a24281a,a24285a,a24286a,a24290a,a24291a,a24292a,a24296a,a24297a,a24301a,a24302a,a24303a,a24307a,a24308a,a24312a,a24313a,a24314a,a24318a,a24319a,a24323a,a24324a,a24325a,a24329a,a24330a,a24334a,a24335a,a24336a,a24340a,a24341a,a24345a,a24346a,a24347a,a24351a,a24352a,a24356a,a24357a,a24358a,a24362a,a24363a,a24367a,a24368a,a24369a,a24373a,a24374a,a24378a,a24379a,a24380a,a24384a,a24385a,a24389a,a24390a,a24391a,a24395a,a24396a,a24400a,a24401a,a24402a,a24406a,a24407a,a24411a,a24412a,a24413a,a24417a,a24418a,a24422a,a24423a,a24424a,a24428a,a24429a,a24433a,a24434a,a24435a,a24439a,a24440a,a24444a,a24445a,a24446a,a24450a,a24451a,a24455a,a24456a,a24457a,a24461a,a24462a,a24466a,a24467a,a24468a,a24472a,a24473a,a24477a,a24478a,a24479a,a24483a,a24484a,a24488a,a24489a,a24490a,a24494a,a24495a,a24499a,a24500a,a24501a,a24505a,a24506a,a24510a,a24511a,a24512a,a24516a,a24517a,a24521a,a24522a,a24523a,a24527a,a24528a,a24532a,a24533a,a24534a,a24538a,a24539a,a24543a,a24544a,a24545a,a24549a,a24550a,a24554a,a24555a,a24556a,a24560a,a24561a,a24565a,a24566a,a24567a,a24571a,a24572a,a24576a,a24577a,a24578a,a24582a,a24583a,a24587a,a24588a,a24589a,a24593a,a24594a,a24598a,a24599a,a24600a,a24604a,a24605a,a24609a,a24610a,a24611a,a24615a,a24616a,a24620a,a24621a,a24622a,a24626a,a24627a,a24631a,a24632a,a24633a,a24637a,a24638a,a24642a,a24643a,a24644a,a24648a,a24649a,a24653a,a24654a,a24655a,a24659a,a24660a,a24664a,a24665a,a24666a,a24670a,a24671a,a24675a,a24676a,a24677a,a24681a,a24682a,a24686a,a24687a,a24688a,a24692a,a24693a,a24697a,a24698a,a24699a,a24703a,a24704a,a24708a,a24709a,a24710a,a24714a,a24715a,a24719a,a24720a,a24721a,a24725a,a24726a,a24730a,a24731a,a24732a,a24736a,a24737a,a24741a,a24742a,a24743a,a24747a,a24748a,a24752a,a24753a,a24754a,a24758a,a24759a,a24763a,a24764a,a24765a,a24769a,a24770a,a24774a,a24775a,a24776a,a24780a,a24781a,a24785a,a24786a,a24787a,a24791a,a24792a,a24796a,a24797a,a24798a,a24802a,a24803a,a24807a,a24808a,a24809a,a24813a,a24814a,a24818a,a24819a,a24820a,a24824a,a24825a,a24829a,a24830a,a24831a,a24835a,a24836a,a24840a,a24841a,a24842a,a24846a,a24847a,a24851a,a24852a,a24853a,a24857a,a24858a,a24862a,a24863a,a24864a,a24868a,a24869a,a24873a,a24874a,a24875a,a24879a,a24880a,a24884a,a24885a,a24886a,a24890a,a24891a,a24895a,a24896a,a24897a,a24901a,a24902a,a24906a,a24907a,a24908a,a24912a,a24913a,a24917a,a24918a,a24919a,a24923a,a24924a,a24928a,a24929a,a24930a,a24934a,a24935a,a24939a,a24940a,a24941a,a24945a,a24946a,a24950a,a24951a,a24952a,a24956a,a24957a,a24961a,a24962a,a24963a,a24967a,a24968a,a24972a,a24973a,a24974a,a24978a,a24979a,a24983a,a24984a,a24985a,a24989a,a24990a,a24994a,a24995a,a24996a,a25000a,a25001a,a25005a,a25006a,a25007a,a25011a,a25012a,a25016a,a25017a,a25018a,a25022a,a25023a,a25027a,a25028a,a25029a,a25033a,a25034a,a25038a,a25039a,a25040a,a25044a,a25045a,a25049a,a25050a,a25051a,a25055a,a25056a,a25060a,a25061a,a25062a,a25066a,a25067a,a25071a,a25072a,a25073a,a25077a,a25078a,a25082a,a25083a,a25084a,a25088a,a25089a,a25093a,a25094a,a25095a,a25099a,a25100a,a25104a,a25105a,a25106a,a25110a,a25111a,a25115a,a25116a,a25117a,a25121a,a25122a,a25126a,a25127a,a25128a,a25132a,a25133a,a25137a,a25138a,a25139a,a25143a,a25144a,a25148a,a25149a,a25150a,a25154a,a25155a,a25159a,a25160a,a25161a,a25165a,a25166a,a25170a,a25171a,a25172a,a25176a,a25177a,a25181a,a25182a,a25183a,a25187a,a25188a,a25192a,a25193a,a25194a,a25198a,a25199a,a25203a,a25204a,a25205a,a25209a,a25210a,a25214a,a25215a,a25216a,a25220a,a25221a,a25225a,a25226a,a25227a,a25231a,a25232a,a25236a,a25237a,a25238a,a25242a,a25243a,a25247a,a25248a,a25249a,a25253a,a25254a,a25258a,a25259a,a25260a,a25264a,a25265a,a25269a,a25270a,a25271a,a25275a,a25276a,a25280a,a25281a,a25282a,a25286a,a25287a,a25291a,a25292a,a25293a,a25297a,a25298a,a25302a,a25303a,a25304a,a25308a,a25309a,a25313a,a25314a,a25315a,a25319a,a25320a,a25324a,a25325a,a25326a,a25330a,a25331a,a25335a,a25336a,a25337a,a25341a,a25342a,a25346a,a25347a,a25348a,a25352a,a25353a,a25357a,a25358a,a25359a,a25363a,a25364a,a25368a,a25369a,a25370a,a25374a,a25375a,a25379a,a25380a,a25381a,a25385a,a25386a,a25390a,a25391a,a25392a,a25396a,a25397a,a25401a,a25402a,a25403a,a25407a,a25408a,a25412a,a25413a,a25414a,a25418a,a25419a,a25423a,a25424a,a25425a,a25429a,a25430a,a25434a,a25435a,a25436a,a25440a,a25441a,a25445a,a25446a,a25447a,a25451a,a25452a,a25456a,a25457a,a25458a,a25462a,a25463a,a25467a,a25468a,a25469a,a25473a,a25474a,a25478a,a25479a,a25480a,a25484a,a25485a,a25489a,a25490a,a25491a,a25495a,a25496a,a25500a,a25501a,a25502a,a25506a,a25507a,a25511a,a25512a,a25513a,a25517a,a25518a,a25522a,a25523a,a25524a,a25528a,a25529a,a25533a,a25534a,a25535a,a25539a,a25540a,a25544a,a25545a,a25546a,a25550a,a25551a,a25555a,a25556a,a25557a,a25561a,a25562a,a25566a,a25567a,a25568a,a25572a,a25573a,a25577a,a25578a,a25579a,a25583a,a25584a,a25588a,a25589a,a25590a,a25594a,a25595a,a25599a,a25600a,a25601a,a25605a,a25606a,a25610a,a25611a,a25612a,a25616a,a25617a,a25621a,a25622a,a25623a,a25627a,a25628a,a25632a,a25633a,a25634a,a25638a,a25639a,a25643a,a25644a,a25645a,a25649a,a25650a,a25654a,a25655a,a25656a,a25660a,a25661a,a25665a,a25666a,a25667a,a25671a,a25672a,a25676a,a25677a,a25678a,a25682a,a25683a,a25687a,a25688a,a25689a,a25693a,a25694a,a25698a,a25699a,a25700a,a25704a,a25705a,a25709a,a25710a,a25711a,a25715a,a25716a,a25720a,a25721a,a25722a,a25726a,a25727a,a25731a,a25732a,a25733a,a25737a,a25738a,a25742a,a25743a,a25744a,a25748a,a25749a,a25753a,a25754a,a25755a,a25759a,a25760a,a25764a,a25765a,a25766a,a25770a,a25771a,a25775a,a25776a,a25777a,a25781a,a25782a,a25786a,a25787a,a25788a,a25792a,a25793a,a25797a,a25798a,a25799a,a25803a,a25804a,a25808a,a25809a,a25810a,a25814a,a25815a,a25819a,a25820a,a25821a,a25825a,a25826a,a25830a,a25831a,a25832a,a25836a,a25837a,a25841a,a25842a,a25843a,a25847a,a25848a,a25852a,a25853a,a25854a,a25858a,a25859a,a25863a,a25864a,a25865a,a25869a,a25870a,a25874a,a25875a,a25876a,a25880a,a25881a,a25885a,a25886a,a25887a,a25891a,a25892a,a25896a,a25897a,a25898a,a25902a,a25903a,a25907a,a25908a,a25909a,a25913a,a25914a,a25918a,a25919a,a25920a,a25924a,a25925a,a25929a,a25930a,a25931a,a25935a,a25936a,a25940a,a25941a,a25942a,a25946a,a25947a,a25951a,a25952a,a25953a,a25957a,a25958a,a25962a,a25963a,a25964a,a25968a,a25969a,a25973a,a25974a,a25975a,a25979a,a25980a,a25984a,a25985a,a25986a,a25990a,a25991a,a25995a,a25996a,a25997a,a26001a,a26002a,a26006a,a26007a,a26008a,a26012a,a26013a,a26017a,a26018a,a26019a,a26023a,a26024a,a26028a,a26029a,a26030a,a26034a,a26035a,a26039a,a26040a,a26041a,a26045a,a26046a,a26050a,a26051a,a26052a,a26056a,a26057a,a26061a,a26062a,a26063a,a26067a,a26068a,a26072a,a26073a,a26074a,a26078a,a26079a,a26083a,a26084a,a26085a,a26089a,a26090a,a26094a,a26095a,a26096a,a26100a,a26101a,a26105a,a26106a,a26107a,a26111a,a26112a,a26116a,a26117a,a26118a,a26122a,a26123a,a26127a,a26128a,a26129a,a26133a,a26134a,a26138a,a26139a,a26140a,a26144a,a26145a,a26149a,a26150a,a26151a,a26155a,a26156a,a26160a,a26161a,a26162a,a26166a,a26167a,a26171a,a26172a,a26173a,a26177a,a26178a,a26182a,a26183a,a26184a,a26188a,a26189a,a26193a,a26194a,a26195a,a26199a,a26200a,a26204a,a26205a,a26206a,a26210a,a26211a,a26215a,a26216a,a26217a,a26221a,a26222a,a26226a,a26227a,a26228a,a26232a,a26233a,a26237a,a26238a,a26239a,a26243a,a26244a,a26248a,a26249a,a26250a,a26254a,a26255a,a26259a,a26260a,a26261a,a26265a,a26266a,a26270a,a26271a,a26272a,a26276a,a26277a,a26281a,a26282a,a26283a,a26287a,a26288a,a26292a,a26293a,a26294a,a26298a,a26299a,a26303a,a26304a,a26305a,a26309a,a26310a,a26314a,a26315a,a26316a,a26320a,a26321a,a26325a,a26326a,a26327a,a26331a,a26332a,a26336a,a26337a,a26338a,a26342a,a26343a,a26347a,a26348a,a26349a,a26353a,a26354a,a26358a,a26359a,a26360a,a26364a,a26365a,a26369a,a26370a,a26371a,a26375a,a26376a,a26380a,a26381a,a26382a,a26386a,a26387a,a26391a,a26392a,a26393a,a26397a,a26398a,a26402a,a26403a,a26404a,a26408a,a26409a,a26413a,a26414a,a26415a,a26419a,a26420a,a26424a,a26425a,a26426a,a26430a,a26431a,a26435a,a26436a,a26437a,a26441a,a26442a,a26446a,a26447a,a26448a,a26452a,a26453a,a26457a,a26458a,a26459a,a26463a,a26464a,a26468a,a26469a,a26470a,a26474a,a26475a,a26479a,a26480a,a26481a,a26485a,a26486a,a26490a,a26491a,a26492a,a26496a,a26497a,a26501a,a26502a,a26503a,a26507a,a26508a,a26512a,a26513a,a26514a,a26518a,a26519a,a26523a,a26524a,a26525a,a26529a,a26530a,a26534a,a26535a,a26536a,a26540a,a26541a,a26545a,a26546a,a26547a,a26551a,a26552a,a26556a,a26557a,a26558a,a26562a,a26563a,a26567a,a26568a,a26569a,a26573a,a26574a,a26578a,a26579a,a26580a,a26584a,a26585a,a26589a,a26590a,a26591a,a26595a,a26596a,a26600a,a26601a,a26602a,a26606a,a26607a,a26611a,a26612a,a26613a,a26617a,a26618a,a26622a,a26623a,a26624a,a26628a,a26629a,a26633a,a26634a,a26635a,a26639a,a26640a,a26644a,a26645a,a26646a,a26650a,a26651a,a26655a,a26656a,a26657a,a26661a,a26662a,a26666a,a26667a,a26668a,a26672a,a26673a,a26677a,a26678a,a26679a,a26683a,a26684a,a26688a,a26689a,a26690a,a26694a,a26695a,a26699a,a26700a,a26701a,a26705a,a26706a,a26710a,a26711a,a26712a,a26716a,a26717a,a26721a,a26722a,a26723a,a26727a,a26728a,a26732a,a26733a,a26734a,a26738a,a26739a,a26743a,a26744a,a26745a,a26749a,a26750a,a26754a,a26755a,a26756a,a26760a,a26761a,a26765a,a26766a,a26767a,a26771a,a26772a,a26776a,a26777a,a26778a,a26782a,a26783a,a26787a,a26788a,a26789a,a26793a,a26794a,a26798a,a26799a,a26800a,a26804a,a26805a,a26809a,a26810a,a26811a,a26815a,a26816a,a26820a,a26821a,a26822a,a26826a,a26827a,a26831a,a26832a,a26833a,a26837a,a26838a,a26842a,a26843a,a26844a,a26848a,a26849a,a26853a,a26854a,a26855a,a26859a,a26860a,a26864a,a26865a,a26866a,a26870a,a26871a,a26875a,a26876a,a26877a,a26881a,a26882a,a26886a,a26887a,a26888a,a26892a,a26893a,a26897a,a26898a,a26899a,a26903a,a26904a,a26908a,a26909a,a26910a,a26914a,a26915a,a26919a,a26920a,a26921a,a26925a,a26926a,a26930a,a26931a,a26932a,a26936a,a26937a,a26941a,a26942a,a26943a,a26947a,a26948a,a26952a,a26953a,a26954a,a26958a,a26959a,a26963a,a26964a,a26965a,a26969a,a26970a,a26974a,a26975a,a26976a,a26980a,a26981a,a26985a,a26986a,a26987a,a26991a,a26992a,a26996a,a26997a,a26998a,a27002a,a27003a,a27007a,a27008a,a27009a,a27013a,a27014a,a27018a,a27019a,a27020a,a27024a,a27025a,a27029a,a27030a,a27031a,a27035a,a27036a,a27040a,a27041a,a27042a,a27046a,a27047a,a27051a,a27052a,a27053a,a27057a,a27058a,a27062a,a27063a,a27064a,a27068a,a27069a,a27073a,a27074a,a27075a,a27079a,a27080a,a27084a,a27085a,a27086a,a27090a,a27091a,a27095a,a27096a,a27097a,a27101a,a27102a,a27106a,a27107a,a27108a,a27112a,a27113a,a27117a,a27118a,a27119a,a27123a,a27124a,a27128a,a27129a,a27130a,a27134a,a27135a,a27139a,a27140a,a27141a,a27145a,a27146a,a27150a,a27151a,a27152a,a27156a,a27157a,a27161a,a27162a,a27163a,a27167a,a27168a,a27172a,a27173a,a27174a,a27178a,a27179a,a27183a,a27184a,a27185a,a27189a,a27190a,a27194a,a27195a,a27196a,a27200a,a27201a,a27205a,a27206a,a27207a,a27211a,a27212a,a27216a,a27217a,a27218a,a27222a,a27223a,a27227a,a27228a,a27229a,a27233a,a27234a,a27238a,a27239a,a27240a,a27244a,a27245a,a27249a,a27250a,a27251a,a27255a,a27256a,a27260a,a27261a,a27262a,a27266a,a27267a,a27271a,a27272a,a27273a,a27277a,a27278a,a27282a,a27283a,a27284a,a27288a,a27289a,a27293a,a27294a,a27295a,a27299a,a27300a,a27304a,a27305a,a27306a,a27310a,a27311a,a27315a,a27316a,a27317a,a27321a,a27322a,a27326a,a27327a,a27328a,a27332a,a27333a,a27337a,a27338a,a27339a,a27343a,a27344a,a27348a,a27349a,a27350a,a27354a,a27355a,a27359a,a27360a,a27361a,a27365a,a27366a,a27370a,a27371a,a27372a,a27376a,a27377a,a27381a,a27382a,a27383a,a27387a,a27388a,a27392a,a27393a,a27394a,a27398a,a27399a,a27403a,a27404a,a27405a,a27409a,a27410a,a27414a,a27415a,a27416a,a27420a,a27421a,a27425a,a27426a,a27427a,a27431a,a27432a,a27436a,a27437a,a27438a,a27442a,a27443a,a27447a,a27448a,a27449a,a27453a,a27454a,a27458a,a27459a,a27460a,a27464a,a27465a,a27469a,a27470a,a27471a,a27475a,a27476a,a27480a,a27481a,a27482a,a27486a,a27487a,a27491a,a27492a,a27493a,a27497a,a27498a,a27502a,a27503a,a27504a,a27508a,a27509a,a27513a,a27514a,a27515a,a27519a,a27520a,a27524a,a27525a,a27526a,a27530a,a27531a,a27535a,a27536a,a27537a,a27541a,a27542a,a27546a,a27547a,a27548a,a27552a,a27553a,a27557a,a27558a,a27559a,a27563a,a27564a,a27568a,a27569a,a27570a,a27574a,a27575a,a27579a,a27580a,a27581a,a27585a,a27586a,a27590a,a27591a,a27592a,a27596a,a27597a,a27601a,a27602a,a27603a,a27607a,a27608a,a27612a,a27613a,a27614a,a27618a,a27619a,a27623a,a27624a,a27625a,a27629a,a27630a,a27634a,a27635a,a27636a,a27640a,a27641a,a27645a,a27646a,a27647a,a27651a,a27652a,a27656a,a27657a,a27658a,a27662a,a27663a,a27667a,a27668a,a27669a,a27673a,a27674a,a27678a,a27679a,a27680a,a27684a,a27685a,a27689a,a27690a,a27691a,a27695a,a27696a,a27700a,a27701a,a27702a,a27706a,a27707a,a27711a,a27712a,a27713a,a27717a,a27718a,a27722a,a27723a,a27724a,a27728a,a27729a,a27733a,a27734a,a27735a,a27739a,a27740a,a27744a,a27745a,a27746a,a27750a,a27751a,a27755a,a27756a,a27757a,a27761a,a27762a,a27766a,a27767a,a27768a,a27772a,a27773a,a27777a,a27778a,a27779a,a27783a,a27784a,a27788a,a27789a,a27790a,a27794a,a27795a,a27799a,a27800a,a27801a,a27805a,a27806a,a27810a,a27811a,a27812a,a27816a,a27817a,a27821a,a27822a,a27823a,a27827a,a27828a,a27832a,a27833a,a27834a,a27838a,a27839a,a27843a,a27844a,a27845a,a27849a,a27850a,a27854a,a27855a,a27856a,a27860a,a27861a,a27865a,a27866a,a27867a,a27871a,a27872a,a27876a,a27877a,a27878a,a27882a,a27883a,a27887a,a27888a,a27889a,a27893a,a27894a,a27898a,a27899a,a27900a,a27904a,a27905a,a27909a,a27910a,a27911a,a27915a,a27916a,a27920a,a27921a,a27922a,a27926a,a27927a,a27931a,a27932a,a27933a,a27937a,a27938a,a27942a,a27943a,a27944a,a27948a,a27949a,a27953a,a27954a,a27955a,a27959a,a27960a,a27964a,a27965a,a27966a,a27970a,a27971a,a27975a,a27976a,a27977a,a27981a,a27982a,a27986a,a27987a,a27988a,a27992a,a27993a,a27997a,a27998a,a27999a,a28003a,a28004a,a28008a,a28009a,a28010a,a28014a,a28015a,a28019a,a28020a,a28021a,a28025a,a28026a,a28030a,a28031a,a28032a,a28036a,a28037a,a28041a,a28042a,a28043a,a28047a,a28048a,a28052a,a28053a,a28054a,a28058a,a28059a,a28063a,a28064a,a28065a,a28069a,a28070a,a28074a,a28075a,a28076a,a28080a,a28081a,a28085a,a28086a,a28087a,a28091a,a28092a,a28096a,a28097a,a28098a,a28102a,a28103a,a28107a,a28108a,a28109a,a28113a,a28114a,a28118a,a28119a,a28120a,a28124a,a28125a,a28129a,a28130a,a28131a,a28135a,a28136a,a28140a,a28141a,a28142a,a28146a,a28147a,a28151a,a28152a,a28153a,a28157a,a28158a,a28162a,a28163a,a28164a,a28168a,a28169a,a28173a,a28174a,a28175a,a28179a,a28180a,a28184a,a28185a,a28186a,a28190a,a28191a,a28195a,a28196a,a28197a,a28201a,a28202a,a28206a,a28207a,a28208a,a28212a,a28213a,a28217a,a28218a,a28219a,a28223a,a28224a,a28228a,a28229a,a28230a,a28234a,a28235a,a28239a,a28240a,a28241a,a28245a,a28246a,a28250a,a28251a,a28252a,a28256a,a28257a,a28261a,a28262a,a28263a,a28267a,a28268a,a28272a,a28273a,a28274a,a28278a,a28279a,a28283a,a28284a,a28285a,a28289a,a28290a,a28294a,a28295a,a28296a,a28300a,a28301a,a28305a,a28306a,a28307a,a28311a,a28312a,a28316a,a28317a,a28318a,a28322a,a28323a,a28327a,a28328a,a28329a,a28333a,a28334a,a28338a,a28339a,a28340a,a28344a,a28345a,a28349a,a28350a,a28351a,a28355a,a28356a,a28360a,a28361a,a28362a,a28366a,a28367a,a28371a,a28372a,a28373a,a28377a,a28378a,a28382a,a28383a,a28384a,a28388a,a28389a,a28393a,a28394a,a28395a,a28399a,a28400a,a28404a,a28405a,a28406a,a28410a,a28411a,a28415a,a28416a,a28417a,a28421a,a28422a,a28426a,a28427a,a28428a,a28432a,a28433a,a28437a,a28438a,a28439a,a28443a,a28444a,a28448a,a28449a,a28450a,a28454a,a28455a,a28459a,a28460a,a28461a,a28465a,a28466a,a28470a,a28471a,a28472a,a28476a,a28477a,a28481a,a28482a,a28483a,a28487a,a28488a,a28492a,a28493a,a28494a,a28498a,a28499a,a28503a,a28504a,a28505a,a28509a,a28510a,a28514a,a28515a,a28516a,a28520a,a28521a,a28525a,a28526a,a28527a,a28531a,a28532a,a28536a,a28537a,a28538a,a28542a,a28543a,a28547a,a28548a,a28549a,a28553a,a28554a,a28558a,a28559a,a28560a,a28564a,a28565a,a28569a,a28570a,a28571a,a28575a,a28576a,a28580a,a28581a,a28582a,a28586a,a28587a,a28591a,a28592a,a28593a,a28597a,a28598a,a28602a,a28603a,a28604a,a28608a,a28609a,a28613a,a28614a,a28615a,a28619a,a28620a,a28624a,a28625a,a28626a,a28630a,a28631a,a28635a,a28636a,a28637a,a28641a,a28642a,a28646a,a28647a,a28648a,a28652a,a28653a,a28657a,a28658a,a28659a,a28663a,a28664a,a28668a,a28669a,a28670a,a28674a,a28675a,a28679a,a28680a,a28681a,a28685a,a28686a,a28690a,a28691a,a28692a,a28696a,a28697a,a28701a,a28702a,a28703a,a28707a,a28708a,a28712a,a28713a,a28714a,a28718a,a28719a,a28723a,a28724a,a28725a,a28729a,a28730a,a28734a,a28735a,a28736a,a28740a,a28741a,a28745a,a28746a,a28747a,a28751a,a28752a,a28756a,a28757a,a28758a,a28762a,a28763a,a28767a,a28768a,a28769a,a28773a,a28774a,a28778a,a28779a,a28780a,a28784a,a28785a,a28789a,a28790a,a28791a,a28795a,a28796a,a28800a,a28801a,a28802a,a28806a,a28807a,a28811a,a28812a,a28813a,a28817a,a28818a,a28822a,a28823a,a28824a,a28828a,a28829a,a28833a,a28834a,a28835a,a28839a,a28840a,a28844a,a28845a,a28846a,a28850a,a28851a,a28855a,a28856a,a28857a,a28861a,a28862a,a28866a,a28867a,a28868a,a28872a,a28873a,a28877a,a28878a,a28879a,a28883a,a28884a,a28888a,a28889a,a28890a,a28894a,a28895a,a28899a,a28900a,a28901a,a28905a,a28906a,a28910a,a28911a,a28912a,a28916a,a28917a,a28921a,a28922a,a28923a,a28927a,a28928a,a28932a,a28933a,a28934a,a28938a,a28939a,a28943a,a28944a,a28945a,a28949a,a28950a,a28954a,a28955a,a28956a,a28960a,a28961a,a28965a,a28966a,a28967a,a28971a,a28972a,a28976a,a28977a,a28978a,a28982a,a28983a,a28987a,a28988a,a28989a,a28993a,a28994a,a28998a,a28999a,a29000a,a29004a,a29005a,a29009a,a29010a,a29011a,a29015a,a29016a,a29020a,a29021a,a29022a,a29026a,a29027a,a29031a,a29032a,a29033a,a29037a,a29038a,a29042a,a29043a,a29044a,a29048a,a29049a,a29053a,a29054a,a29055a,a29059a,a29060a,a29064a,a29065a,a29066a,a29070a,a29071a,a29075a,a29076a,a29077a,a29081a,a29082a,a29086a,a29087a,a29088a,a29092a,a29093a,a29097a,a29098a,a29099a,a29103a,a29104a,a29108a,a29109a,a29110a,a29114a,a29115a,a29119a,a29120a,a29121a,a29125a,a29126a,a29130a,a29131a,a29132a,a29136a,a29137a,a29141a,a29142a,a29143a,a29147a,a29148a,a29152a,a29153a,a29154a,a29158a,a29159a,a29163a,a29164a,a29165a,a29169a,a29170a,a29174a,a29175a,a29176a,a29180a,a29181a,a29185a,a29186a,a29187a,a29191a,a29192a,a29196a,a29197a,a29198a,a29202a,a29203a,a29207a,a29208a,a29209a,a29213a,a29214a,a29218a,a29219a,a29220a,a29224a,a29225a,a29229a,a29230a,a29231a,a29235a,a29236a,a29240a,a29241a,a29242a,a29246a,a29247a,a29251a,a29252a,a29253a,a29257a,a29258a,a29262a,a29263a,a29264a,a29268a,a29269a,a29273a,a29274a,a29275a,a29279a,a29280a,a29284a,a29285a,a29286a,a29290a,a29291a,a29295a,a29296a,a29297a,a29301a,a29302a,a29306a,a29307a,a29308a,a29312a,a29313a,a29317a,a29318a,a29319a,a29323a,a29324a,a29328a,a29329a,a29330a,a29334a,a29335a,a29339a,a29340a,a29341a,a29345a,a29346a,a29350a,a29351a,a29352a,a29356a,a29357a,a29361a,a29362a,a29363a,a29367a,a29368a,a29372a,a29373a,a29374a,a29378a,a29379a,a29383a,a29384a,a29385a,a29389a,a29390a,a29394a,a29395a,a29396a,a29400a,a29401a,a29405a,a29406a,a29407a,a29411a,a29412a,a29416a,a29417a,a29418a,a29422a,a29423a,a29427a,a29428a,a29429a,a29433a,a29434a,a29438a,a29439a,a29440a,a29444a,a29445a,a29449a,a29450a,a29451a,a29455a,a29456a,a29460a,a29461a,a29462a,a29466a,a29467a,a29471a,a29472a,a29473a,a29477a,a29478a,a29482a,a29483a,a29484a,a29488a,a29489a,a29493a,a29494a,a29495a,a29499a,a29500a,a29503a,a29506a,a29507a,a29508a,a29512a,a29513a,a29517a,a29518a,a29519a,a29523a,a29524a,a29527a,a29530a,a29531a,a29532a,a29536a,a29537a,a29541a,a29542a,a29543a,a29547a,a29548a,a29551a,a29554a,a29555a,a29556a,a29560a,a29561a,a29565a,a29566a,a29567a,a29571a,a29572a,a29575a,a29578a,a29579a,a29580a,a29584a,a29585a,a29589a,a29590a,a29591a,a29595a,a29596a,a29599a,a29602a,a29603a,a29604a,a29608a,a29609a,a29613a,a29614a,a29615a,a29619a,a29620a,a29623a,a29626a,a29627a,a29628a,a29632a,a29633a,a29637a,a29638a,a29639a,a29643a,a29644a,a29647a,a29650a,a29651a,a29652a,a29656a,a29657a,a29661a,a29662a,a29663a,a29667a,a29668a,a29671a,a29674a,a29675a,a29676a,a29680a,a29681a,a29685a,a29686a,a29687a,a29691a,a29692a,a29695a,a29698a,a29699a,a29700a,a29704a,a29705a,a29709a,a29710a,a29711a,a29715a,a29716a,a29719a,a29722a,a29723a,a29724a,a29728a,a29729a,a29733a,a29734a,a29735a,a29739a,a29740a,a29743a,a29746a,a29747a,a29748a,a29752a,a29753a,a29757a,a29758a,a29759a,a29763a,a29764a,a29767a,a29770a,a29771a,a29772a,a29776a,a29777a,a29781a,a29782a,a29783a,a29787a,a29788a,a29791a,a29794a,a29795a,a29796a,a29800a,a29801a,a29805a,a29806a,a29807a,a29811a,a29812a,a29815a,a29818a,a29819a,a29820a,a29824a,a29825a,a29829a,a29830a,a29831a,a29835a,a29836a,a29839a,a29842a,a29843a,a29844a,a29848a,a29849a,a29853a,a29854a,a29855a,a29859a,a29860a,a29863a,a29866a,a29867a,a29868a,a29872a,a29873a,a29877a,a29878a,a29879a,a29883a,a29884a,a29887a,a29890a,a29891a,a29892a,a29896a,a29897a,a29901a,a29902a,a29903a,a29907a,a29908a,a29911a,a29914a,a29915a,a29916a,a29920a,a29921a,a29925a,a29926a,a29927a,a29931a,a29932a,a29935a,a29938a,a29939a,a29940a,a29944a,a29945a,a29949a,a29950a,a29951a,a29955a,a29956a,a29959a,a29962a,a29963a,a29964a,a29968a,a29969a,a29973a,a29974a,a29975a,a29979a,a29980a,a29983a,a29986a,a29987a,a29988a,a29992a,a29993a,a29997a,a29998a,a29999a,a30003a,a30004a,a30007a,a30010a,a30011a,a30012a,a30016a,a30017a,a30021a,a30022a,a30023a,a30027a,a30028a,a30031a,a30034a,a30035a,a30036a,a30040a,a30041a,a30045a,a30046a,a30047a,a30051a,a30052a,a30055a,a30058a,a30059a,a30060a,a30064a,a30065a,a30069a,a30070a,a30071a,a30075a,a30076a,a30079a,a30082a,a30083a,a30084a,a30088a,a30089a,a30093a,a30094a,a30095a,a30099a,a30100a,a30103a,a30106a,a30107a,a30108a,a30112a,a30113a,a30117a,a30118a,a30119a,a30123a,a30124a,a30127a,a30130a,a30131a,a30132a,a30136a,a30137a,a30141a,a30142a,a30143a,a30147a,a30148a,a30151a,a30154a,a30155a,a30156a,a30160a,a30161a,a30165a,a30166a,a30167a,a30171a,a30172a,a30175a,a30178a,a30179a,a30180a,a30184a,a30185a,a30189a,a30190a,a30191a,a30195a,a30196a,a30199a,a30202a,a30203a,a30204a,a30208a,a30209a,a30213a,a30214a,a30215a,a30219a,a30220a,a30223a,a30226a,a30227a,a30228a,a30232a,a30233a,a30237a,a30238a,a30239a,a30243a,a30244a,a30247a,a30250a,a30251a,a30252a,a30256a,a30257a,a30261a,a30262a,a30263a,a30267a,a30268a,a30271a,a30274a,a30275a,a30276a,a30280a,a30281a,a30285a,a30286a,a30287a,a30291a,a30292a,a30295a,a30298a,a30299a,a30300a,a30304a,a30305a,a30309a,a30310a,a30311a,a30315a,a30316a,a30319a,a30322a,a30323a,a30324a,a30328a,a30329a,a30333a,a30334a,a30335a,a30339a,a30340a,a30343a,a30346a,a30347a,a30348a,a30352a,a30353a,a30357a,a30358a,a30359a,a30363a,a30364a,a30367a,a30370a,a30371a,a30372a,a30376a,a30377a,a30381a,a30382a,a30383a,a30387a,a30388a,a30391a,a30394a,a30395a,a30396a,a30400a,a30401a,a30405a,a30406a,a30407a,a30411a,a30412a,a30415a,a30418a,a30419a,a30420a,a30424a,a30425a,a30429a,a30430a,a30431a,a30435a,a30436a,a30439a,a30442a,a30443a,a30444a,a30448a,a30449a,a30453a,a30454a,a30455a,a30459a,a30460a,a30463a,a30466a,a30467a,a30468a,a30472a,a30473a,a30477a,a30478a,a30479a,a30483a,a30484a,a30487a,a30490a,a30491a,a30492a,a30496a,a30497a,a30501a,a30502a,a30503a,a30507a,a30508a,a30511a,a30514a,a30515a,a30516a,a30520a,a30521a,a30525a,a30526a,a30527a,a30531a,a30532a,a30535a,a30538a,a30539a,a30540a,a30544a,a30545a,a30549a,a30550a,a30551a,a30555a,a30556a,a30559a,a30562a,a30563a,a30564a,a30568a,a30569a,a30573a,a30574a,a30575a,a30579a,a30580a,a30583a,a30586a,a30587a,a30588a,a30592a,a30593a,a30597a,a30598a,a30599a,a30603a,a30604a,a30607a,a30610a,a30611a,a30612a,a30616a,a30617a,a30621a,a30622a,a30623a,a30627a,a30628a,a30631a,a30634a,a30635a,a30636a,a30640a,a30641a,a30645a,a30646a,a30647a,a30651a,a30652a,a30655a,a30658a,a30659a,a30660a,a30664a,a30665a,a30669a,a30670a,a30671a,a30675a,a30676a,a30679a,a30682a,a30683a,a30684a,a30688a,a30689a,a30693a,a30694a,a30695a,a30699a,a30700a,a30703a,a30706a,a30707a,a30708a,a30712a,a30713a,a30717a,a30718a,a30719a,a30723a,a30724a,a30727a,a30730a,a30731a,a30732a,a30736a,a30737a,a30741a,a30742a,a30743a,a30747a,a30748a,a30751a,a30754a,a30755a,a30756a,a30760a,a30761a,a30765a,a30766a,a30767a,a30771a,a30772a,a30775a,a30778a,a30779a,a30780a,a30784a,a30785a,a30789a,a30790a,a30791a,a30795a,a30796a,a30799a,a30802a,a30803a,a30804a,a30808a,a30809a,a30813a,a30814a,a30815a,a30819a,a30820a,a30823a,a30826a,a30827a,a30828a,a30832a,a30833a,a30837a,a30838a,a30839a,a30843a,a30844a,a30847a,a30850a,a30851a,a30852a,a30856a,a30857a,a30861a,a30862a,a30863a,a30867a,a30868a,a30871a,a30874a,a30875a,a30876a,a30880a,a30881a,a30885a,a30886a,a30887a,a30891a,a30892a,a30895a,a30898a,a30899a,a30900a,a30904a,a30905a,a30909a,a30910a,a30911a,a30915a,a30916a,a30919a,a30922a,a30923a,a30924a,a30928a,a30929a,a30933a,a30934a,a30935a,a30939a,a30940a,a30943a,a30946a,a30947a,a30948a,a30952a,a30953a,a30957a,a30958a,a30959a,a30963a,a30964a,a30967a,a30970a,a30971a,a30972a,a30976a,a30977a,a30981a,a30982a,a30983a,a30987a,a30988a,a30991a,a30994a,a30995a,a30996a,a31000a,a31001a,a31005a,a31006a,a31007a,a31011a,a31012a,a31015a,a31018a,a31019a,a31020a,a31024a,a31025a,a31029a,a31030a,a31031a,a31035a,a31036a,a31039a,a31042a,a31043a,a31044a,a31048a,a31049a,a31053a,a31054a,a31055a,a31059a,a31060a,a31063a,a31066a,a31067a,a31068a,a31072a,a31073a,a31077a,a31078a,a31079a,a31083a,a31084a,a31087a,a31090a,a31091a,a31092a,a31096a,a31097a,a31101a,a31102a,a31103a,a31107a,a31108a,a31111a,a31114a,a31115a,a31116a,a31120a,a31121a,a31125a,a31126a,a31127a,a31131a,a31132a,a31135a,a31138a,a31139a,a31140a,a31144a,a31145a,a31149a,a31150a,a31151a,a31155a,a31156a,a31159a,a31162a,a31163a,a31164a,a31168a,a31169a,a31173a,a31174a,a31175a,a31179a,a31180a,a31183a,a31186a,a31187a,a31188a,a31192a,a31193a,a31197a,a31198a,a31199a,a31203a,a31204a,a31207a,a31210a,a31211a,a31212a,a31216a,a31217a,a31221a,a31222a,a31223a,a31227a,a31228a,a31231a,a31234a,a31235a,a31236a,a31240a,a31241a,a31245a,a31246a,a31247a,a31251a,a31252a,a31255a,a31258a,a31259a,a31260a,a31264a,a31265a,a31269a,a31270a,a31271a,a31275a,a31276a,a31279a,a31282a,a31283a,a31284a,a31288a,a31289a,a31293a,a31294a,a31295a,a31299a,a31300a,a31303a,a31306a,a31307a,a31308a,a31312a,a31313a,a31317a,a31318a,a31319a,a31323a,a31324a,a31327a,a31330a,a31331a,a31332a,a31336a,a31337a,a31341a,a31342a,a31343a,a31347a,a31348a,a31351a,a31354a,a31355a,a31356a,a31360a,a31361a,a31365a,a31366a,a31367a,a31371a,a31372a,a31375a,a31378a,a31379a,a31380a,a31384a,a31385a,a31389a,a31390a,a31391a,a31395a,a31396a,a31399a,a31402a,a31403a,a31404a,a31408a,a31409a,a31413a,a31414a,a31415a,a31419a,a31420a,a31423a,a31426a,a31427a,a31428a,a31432a,a31433a,a31437a,a31438a,a31439a,a31443a,a31444a,a31447a,a31450a,a31451a,a31452a,a31456a,a31457a,a31461a,a31462a,a31463a,a31467a,a31468a,a31471a,a31474a,a31475a,a31476a,a31480a,a31481a,a31485a,a31486a,a31487a,a31491a,a31492a,a31495a,a31498a,a31499a,a31500a,a31504a,a31505a,a31509a,a31510a,a31511a,a31515a,a31516a,a31519a,a31522a,a31523a,a31524a,a31528a,a31529a,a31533a,a31534a,a31535a,a31539a,a31540a,a31543a,a31546a,a31547a,a31548a,a31552a,a31553a,a31557a,a31558a,a31559a,a31563a,a31564a,a31567a,a31570a,a31571a,a31572a,a31576a,a31577a,a31581a,a31582a,a31583a,a31587a,a31588a,a31591a,a31594a,a31595a,a31596a,a31600a,a31601a,a31605a,a31606a,a31607a,a31611a,a31612a,a31615a,a31618a,a31619a,a31620a,a31624a,a31625a,a31629a,a31630a,a31631a,a31635a,a31636a,a31639a,a31642a,a31643a,a31644a,a31648a,a31649a,a31653a,a31654a,a31655a,a31659a,a31660a,a31663a,a31666a,a31667a,a31668a,a31672a,a31673a,a31677a,a31678a,a31679a,a31683a,a31684a,a31687a,a31690a,a31691a,a31692a,a31696a,a31697a,a31701a,a31702a,a31703a,a31707a,a31708a,a31711a,a31714a,a31715a,a31716a,a31720a,a31721a,a31725a,a31726a,a31727a,a31731a,a31732a,a31735a,a31738a,a31739a,a31740a,a31744a,a31745a,a31749a,a31750a,a31751a,a31755a,a31756a,a31759a,a31762a,a31763a,a31764a,a31768a,a31769a,a31773a,a31774a,a31775a,a31779a,a31780a,a31783a,a31786a,a31787a,a31788a,a31792a,a31793a,a31797a,a31798a,a31799a,a31803a,a31804a,a31807a,a31810a,a31811a,a31812a,a31816a,a31817a,a31821a,a31822a,a31823a,a31827a,a31828a,a31831a,a31834a,a31835a,a31836a,a31840a,a31841a,a31845a,a31846a,a31847a,a31851a,a31852a,a31855a,a31858a,a31859a,a31860a,a31864a,a31865a,a31869a,a31870a,a31871a,a31875a,a31876a,a31879a,a31882a,a31883a,a31884a,a31888a,a31889a,a31893a,a31894a,a31895a,a31899a,a31900a,a31903a,a31906a,a31907a,a31908a,a31912a,a31913a,a31917a,a31918a,a31919a,a31923a,a31924a,a31927a,a31930a,a31931a,a31932a,a31936a,a31937a,a31941a,a31942a,a31943a,a31947a,a31948a,a31951a,a31954a,a31955a,a31956a,a31960a,a31961a,a31965a,a31966a,a31967a,a31971a,a31972a,a31975a,a31978a,a31979a,a31980a,a31984a,a31985a,a31989a,a31990a,a31991a,a31995a,a31996a,a31999a,a32002a,a32003a,a32004a,a32008a,a32009a,a32013a,a32014a,a32015a,a32019a,a32020a,a32023a,a32026a,a32027a,a32028a,a32032a,a32033a,a32037a,a32038a,a32039a,a32043a,a32044a,a32047a,a32050a,a32051a,a32052a,a32056a,a32057a,a32061a,a32062a,a32063a,a32067a,a32068a,a32071a,a32074a,a32075a,a32076a,a32080a,a32081a,a32085a,a32086a,a32087a,a32091a,a32092a,a32095a,a32098a,a32099a,a32100a,a32104a,a32105a,a32109a,a32110a,a32111a,a32115a,a32116a,a32119a,a32122a,a32123a,a32124a,a32128a,a32129a,a32133a,a32134a,a32135a,a32139a,a32140a,a32143a,a32146a,a32147a,a32148a,a32152a,a32153a,a32157a,a32158a,a32159a,a32163a,a32164a,a32167a,a32170a,a32171a,a32172a,a32176a,a32177a,a32181a,a32182a,a32183a,a32187a,a32188a,a32191a,a32194a,a32195a,a32196a,a32200a,a32201a,a32205a,a32206a,a32207a,a32211a,a32212a,a32215a,a32218a,a32219a,a32220a,a32224a,a32225a,a32229a,a32230a,a32231a,a32235a,a32236a,a32239a,a32242a,a32243a,a32244a,a32248a,a32249a,a32253a,a32254a,a32255a,a32259a,a32260a,a32263a,a32266a,a32267a,a32268a,a32272a,a32273a,a32277a,a32278a,a32279a,a32283a,a32284a,a32287a,a32290a,a32291a,a32292a,a32296a,a32297a,a32301a,a32302a,a32303a,a32307a,a32308a,a32311a,a32314a,a32315a,a32316a,a32320a,a32321a,a32325a,a32326a,a32327a,a32331a,a32332a,a32335a,a32338a,a32339a,a32340a,a32344a,a32345a,a32349a,a32350a,a32351a,a32355a,a32356a,a32359a,a32362a,a32363a,a32364a,a32368a,a32369a,a32373a,a32374a,a32375a,a32379a,a32380a,a32383a,a32386a,a32387a,a32388a,a32392a,a32393a,a32397a,a32398a,a32399a,a32403a,a32404a,a32407a,a32410a,a32411a,a32412a,a32416a,a32417a,a32421a,a32422a,a32423a,a32427a,a32428a,a32431a,a32434a,a32435a,a32436a,a32440a,a32441a,a32445a,a32446a,a32447a,a32451a,a32452a,a32455a,a32458a,a32459a,a32460a,a32464a,a32465a,a32469a,a32470a,a32471a,a32475a,a32476a,a32479a,a32482a,a32483a,a32484a,a32488a,a32489a,a32493a,a32494a,a32495a,a32499a,a32500a,a32503a,a32506a,a32507a,a32508a,a32512a,a32513a,a32517a,a32518a,a32519a,a32523a,a32524a,a32527a,a32530a,a32531a,a32532a,a32536a,a32537a,a32541a,a32542a,a32543a,a32547a,a32548a,a32551a,a32554a,a32555a,a32556a,a32560a,a32561a,a32565a,a32566a,a32567a,a32571a,a32572a,a32575a,a32578a,a32579a,a32580a,a32584a,a32585a,a32589a,a32590a,a32591a,a32595a,a32596a,a32599a,a32602a,a32603a,a32604a,a32608a,a32609a,a32613a,a32614a,a32615a,a32619a,a32620a,a32623a,a32626a,a32627a,a32628a,a32632a,a32633a,a32637a,a32638a,a32639a,a32643a,a32644a,a32647a,a32650a,a32651a,a32652a,a32656a,a32657a,a32661a,a32662a,a32663a,a32667a,a32668a,a32671a,a32674a,a32675a,a32676a,a32680a,a32681a,a32685a,a32686a,a32687a,a32691a,a32692a,a32695a,a32698a,a32699a,a32700a,a32704a,a32705a,a32709a,a32710a,a32711a,a32715a,a32716a,a32719a,a32722a,a32723a,a32724a,a32728a,a32729a,a32733a,a32734a,a32735a,a32739a,a32740a,a32743a,a32746a,a32747a,a32748a,a32752a,a32753a,a32757a,a32758a,a32759a,a32763a,a32764a,a32767a,a32770a,a32771a,a32772a,a32776a,a32777a,a32781a,a32782a,a32783a,a32787a,a32788a,a32791a,a32794a,a32795a,a32796a,a32800a,a32801a,a32805a,a32806a,a32807a,a32811a,a32812a,a32815a,a32818a,a32819a,a32820a,a32824a,a32825a,a32829a,a32830a,a32831a,a32835a,a32836a,a32839a,a32842a,a32843a,a32844a,a32848a,a32849a,a32853a,a32854a,a32855a,a32859a,a32860a,a32863a,a32866a,a32867a,a32868a,a32872a,a32873a,a32877a,a32878a,a32879a,a32883a,a32884a,a32887a,a32890a,a32891a,a32892a,a32896a,a32897a,a32901a,a32902a,a32903a,a32907a,a32908a,a32911a,a32914a,a32915a,a32916a,a32920a,a32921a,a32925a,a32926a,a32927a,a32931a,a32932a,a32935a,a32938a,a32939a,a32940a,a32944a,a32945a,a32949a,a32950a,a32951a,a32955a,a32956a,a32959a,a32962a,a32963a,a32964a,a32968a,a32969a,a32973a,a32974a,a32975a,a32979a,a32980a,a32983a,a32986a,a32987a,a32988a,a32992a,a32993a,a32997a,a32998a,a32999a,a33003a,a33004a,a33007a,a33010a,a33011a,a33012a,a33016a,a33017a,a33021a,a33022a,a33023a,a33027a,a33028a,a33031a,a33034a,a33035a,a33036a,a33040a,a33041a,a33045a,a33046a,a33047a,a33051a,a33052a,a33055a,a33058a,a33059a,a33060a,a33064a,a33065a,a33069a,a33070a,a33071a,a33075a,a33076a,a33079a,a33082a,a33083a,a33084a,a33088a,a33089a,a33093a,a33094a,a33095a,a33099a,a33100a,a33103a,a33106a,a33107a,a33108a,a33112a,a33113a,a33117a,a33118a,a33119a,a33123a,a33124a,a33127a,a33130a,a33131a,a33132a,a33136a,a33137a,a33141a,a33142a,a33143a,a33147a,a33148a,a33151a,a33154a,a33155a,a33156a,a33160a,a33161a,a33165a,a33166a,a33167a,a33171a,a33172a,a33175a,a33178a,a33179a,a33180a,a33184a,a33185a,a33189a,a33190a,a33191a,a33195a,a33196a,a33199a,a33202a,a33203a,a33204a,a33208a,a33209a,a33213a,a33214a,a33215a,a33219a,a33220a,a33223a,a33226a,a33227a,a33228a,a33232a,a33233a,a33237a,a33238a,a33239a,a33243a,a33244a,a33247a,a33250a,a33251a,a33252a,a33256a,a33257a,a33261a,a33262a,a33263a,a33267a,a33268a,a33271a,a33274a,a33275a,a33276a,a33280a,a33281a,a33285a,a33286a,a33287a,a33291a,a33292a,a33295a,a33298a,a33299a,a33300a,a33304a,a33305a,a33309a,a33310a,a33311a,a33315a,a33316a,a33319a,a33322a,a33323a,a33324a,a33328a,a33329a,a33333a,a33334a,a33335a,a33339a,a33340a,a33343a,a33346a,a33347a,a33348a,a33352a,a33353a,a33357a,a33358a,a33359a,a33363a,a33364a,a33367a,a33370a,a33371a,a33372a,a33376a,a33377a,a33381a,a33382a,a33383a,a33387a,a33388a,a33391a,a33394a,a33395a,a33396a,a33400a,a33401a,a33405a,a33406a,a33407a,a33411a,a33412a,a33415a,a33418a,a33419a,a33420a,a33424a,a33425a,a33429a,a33430a,a33431a,a33435a,a33436a,a33439a,a33442a,a33443a,a33444a,a33448a,a33449a,a33453a,a33454a,a33455a,a33459a,a33460a,a33463a,a33466a,a33467a,a33468a,a33472a,a33473a,a33477a,a33478a,a33479a,a33483a,a33484a,a33487a,a33490a,a33491a,a33492a,a33496a,a33497a,a33501a,a33502a,a33503a,a33507a,a33508a,a33511a,a33514a,a33515a,a33516a,a33520a,a33521a,a33525a,a33526a,a33527a,a33531a,a33532a,a33535a,a33538a,a33539a,a33540a,a33544a,a33545a,a33549a,a33550a,a33551a,a33555a,a33556a,a33559a,a33562a,a33563a,a33564a,a33568a,a33569a,a33573a,a33574a,a33575a,a33579a,a33580a,a33583a,a33586a,a33587a,a33588a,a33592a,a33593a,a33597a,a33598a,a33599a,a33603a,a33604a,a33607a,a33610a,a33611a,a33612a,a33616a,a33617a,a33621a,a33622a,a33623a,a33627a,a33628a,a33631a,a33634a,a33635a,a33636a,a33640a,a33641a,a33645a,a33646a,a33647a,a33651a,a33652a,a33655a,a33658a,a33659a,a33660a,a33664a,a33665a,a33669a,a33670a,a33671a,a33675a,a33676a,a33679a,a33682a,a33683a,a33684a,a33688a,a33689a,a33693a,a33694a,a33695a,a33699a,a33700a,a33703a,a33706a,a33707a,a33708a,a33712a,a33713a,a33717a,a33718a,a33719a,a33723a,a33724a,a33727a,a33730a,a33731a,a33732a,a33736a,a33737a,a33741a,a33742a,a33743a,a33747a,a33748a,a33751a,a33754a,a33755a,a33756a,a33760a,a33761a,a33765a,a33766a,a33767a,a33771a,a33772a,a33775a,a33778a,a33779a,a33780a,a33784a,a33785a,a33789a,a33790a,a33791a,a33795a,a33796a,a33799a,a33802a,a33803a,a33804a,a33808a,a33809a,a33813a,a33814a,a33815a,a33819a,a33820a,a33823a,a33826a,a33827a,a33828a,a33832a,a33833a,a33837a,a33838a,a33839a,a33843a,a33844a,a33847a,a33850a,a33851a,a33852a,a33856a,a33857a,a33861a,a33862a,a33863a,a33867a,a33868a,a33871a,a33874a,a33875a,a33876a,a33880a,a33881a,a33885a,a33886a,a33887a,a33891a,a33892a,a33895a,a33898a,a33899a,a33900a,a33904a,a33905a,a33909a,a33910a,a33911a,a33915a,a33916a,a33919a,a33922a,a33923a,a33924a,a33928a,a33929a,a33933a,a33934a,a33935a,a33939a,a33940a,a33943a,a33946a,a33947a,a33948a,a33952a,a33953a,a33957a,a33958a,a33959a,a33963a,a33964a,a33967a,a33970a,a33971a,a33972a,a33976a,a33977a,a33981a,a33982a,a33983a,a33987a,a33988a,a33991a,a33994a,a33995a,a33996a,a34000a,a34001a,a34005a,a34006a,a34007a,a34011a,a34012a,a34015a,a34018a,a34019a,a34020a,a34024a,a34025a,a34029a,a34030a,a34031a,a34035a,a34036a,a34039a,a34042a,a34043a,a34044a,a34048a,a34049a,a34053a,a34054a,a34055a,a34059a,a34060a,a34063a,a34066a,a34067a,a34068a,a34072a,a34073a,a34077a,a34078a,a34079a,a34083a,a34084a,a34087a,a34090a,a34091a,a34092a,a34096a,a34097a,a34101a,a34102a,a34103a,a34107a,a34108a,a34111a,a34114a,a34115a,a34116a,a34120a,a34121a,a34125a,a34126a,a34127a,a34131a,a34132a,a34135a,a34138a,a34139a,a34140a,a34144a,a34145a,a34149a,a34150a,a34151a,a34155a,a34156a,a34159a,a34162a,a34163a,a34164a,a34168a,a34169a,a34173a,a34174a,a34175a,a34179a,a34180a,a34183a,a34186a,a34187a,a34188a,a34192a,a34193a,a34197a,a34198a,a34199a,a34203a,a34204a,a34207a,a34210a,a34211a,a34212a,a34216a,a34217a,a34221a,a34222a,a34223a,a34227a,a34228a,a34231a,a34234a,a34235a,a34236a,a34240a,a34241a,a34245a,a34246a,a34247a,a34251a,a34252a,a34255a,a34258a,a34259a,a34260a,a34264a,a34265a,a34269a,a34270a,a34271a,a34275a,a34276a,a34279a,a34282a,a34283a,a34284a,a34288a,a34289a,a34293a,a34294a,a34295a,a34299a,a34300a,a34303a,a34306a,a34307a,a34308a,a34312a,a34313a,a34317a,a34318a,a34319a,a34323a,a34324a,a34327a,a34330a,a34331a,a34332a,a34336a,a34337a,a34341a,a34342a,a34343a,a34347a,a34348a,a34351a,a34354a,a34355a,a34356a,a34360a,a34361a,a34365a,a34366a,a34367a,a34371a,a34372a,a34375a,a34378a,a34379a,a34380a,a34384a,a34385a,a34389a,a34390a,a34391a,a34395a,a34396a,a34399a,a34402a,a34403a,a34404a,a34408a,a34409a,a34413a,a34414a,a34415a,a34419a,a34420a,a34423a,a34426a,a34427a,a34428a,a34432a,a34433a,a34437a,a34438a,a34439a,a34443a,a34444a,a34447a,a34450a,a34451a,a34452a,a34456a,a34457a,a34461a,a34462a,a34463a,a34467a,a34468a,a34471a,a34474a,a34475a,a34476a,a34480a,a34481a,a34485a,a34486a,a34487a,a34491a,a34492a,a34495a,a34498a,a34499a,a34500a,a34504a,a34505a,a34509a,a34510a,a34511a,a34515a,a34516a,a34519a,a34522a,a34523a,a34524a,a34528a,a34529a,a34533a,a34534a,a34535a,a34539a,a34540a,a34543a,a34546a,a34547a,a34548a,a34552a,a34553a,a34557a,a34558a,a34559a,a34563a,a34564a,a34567a,a34570a,a34571a,a34572a,a34576a,a34577a,a34581a,a34582a,a34583a,a34587a,a34588a,a34591a,a34594a,a34595a,a34596a,a34600a,a34601a,a34605a,a34606a,a34607a,a34611a,a34612a,a34615a,a34618a,a34619a,a34620a,a34624a,a34625a,a34629a,a34630a,a34631a,a34635a,a34636a,a34639a,a34642a,a34643a,a34644a,a34648a,a34649a,a34653a,a34654a,a34655a,a34659a,a34660a,a34663a,a34666a,a34667a,a34668a,a34672a,a34673a,a34677a,a34678a,a34679a,a34683a,a34684a,a34687a,a34690a,a34691a,a34692a,a34696a,a34697a,a34701a,a34702a,a34703a,a34707a,a34708a,a34711a,a34714a,a34715a,a34716a,a34720a,a34721a,a34725a,a34726a,a34727a,a34731a,a34732a,a34735a,a34738a,a34739a,a34740a,a34744a,a34745a,a34749a,a34750a,a34751a,a34755a,a34756a,a34759a,a34762a,a34763a,a34764a,a34768a,a34769a,a34773a,a34774a,a34775a,a34779a,a34780a,a34783a,a34786a,a34787a,a34788a,a34792a,a34793a,a34797a,a34798a,a34799a,a34803a,a34804a,a34807a,a34810a,a34811a,a34812a,a34816a,a34817a,a34821a,a34822a,a34823a,a34827a,a34828a,a34831a,a34834a,a34835a,a34836a,a34840a,a34841a,a34845a,a34846a,a34847a,a34851a,a34852a,a34855a,a34858a,a34859a,a34860a,a34864a,a34865a,a34869a,a34870a,a34871a,a34875a,a34876a,a34879a,a34882a,a34883a,a34884a,a34888a,a34889a,a34893a,a34894a,a34895a,a34899a,a34900a,a34903a,a34906a,a34907a,a34908a,a34912a,a34913a,a34917a,a34918a,a34919a,a34923a,a34924a,a34927a,a34930a,a34931a,a34932a,a34936a,a34937a,a34941a,a34942a,a34943a,a34947a,a34948a,a34951a,a34954a,a34955a,a34956a,a34960a,a34961a,a34965a,a34966a,a34967a,a34971a,a34972a,a34975a,a34978a,a34979a,a34980a,a34984a,a34985a,a34989a,a34990a,a34991a,a34995a,a34996a,a34999a,a35002a,a35003a,a35004a,a35008a,a35009a,a35013a,a35014a,a35015a,a35019a,a35020a,a35023a,a35026a,a35027a,a35028a,a35032a,a35033a,a35037a,a35038a,a35039a,a35043a,a35044a,a35047a,a35050a,a35051a,a35052a,a35056a,a35057a,a35061a,a35062a,a35063a,a35067a,a35068a,a35071a,a35074a,a35075a,a35076a,a35080a,a35081a,a35085a,a35086a,a35087a,a35091a,a35092a,a35095a,a35098a,a35099a,a35100a,a35104a,a35105a,a35109a,a35110a,a35111a,a35115a,a35116a,a35119a,a35122a,a35123a,a35124a,a35128a,a35129a,a35133a,a35134a,a35135a,a35139a,a35140a,a35143a,a35146a,a35147a,a35148a,a35152a,a35153a,a35157a,a35158a,a35159a,a35163a,a35164a,a35167a,a35170a,a35171a,a35172a,a35176a,a35177a,a35181a,a35182a,a35183a,a35187a,a35188a,a35191a,a35194a,a35195a,a35196a,a35200a,a35201a,a35205a,a35206a,a35207a,a35211a,a35212a,a35215a,a35218a,a35219a,a35220a,a35224a,a35225a,a35229a,a35230a,a35231a,a35235a,a35236a,a35239a,a35242a,a35243a,a35244a,a35248a,a35249a,a35253a,a35254a,a35255a,a35259a,a35260a,a35263a,a35266a,a35267a,a35268a,a35272a,a35273a,a35277a,a35278a,a35279a,a35283a,a35284a,a35287a,a35290a,a35291a,a35292a,a35296a,a35297a,a35301a,a35302a,a35303a,a35307a,a35308a,a35311a,a35314a,a35315a,a35316a,a35320a,a35321a,a35325a,a35326a,a35327a,a35331a,a35332a,a35335a,a35338a,a35339a,a35340a,a35344a,a35345a,a35349a,a35350a,a35351a,a35355a,a35356a,a35359a,a35362a,a35363a,a35364a,a35368a,a35369a,a35373a,a35374a,a35375a,a35379a,a35380a,a35383a,a35386a,a35387a,a35388a,a35392a,a35393a,a35397a,a35398a,a35399a,a35403a,a35404a,a35407a,a35410a,a35411a,a35412a,a35416a,a35417a,a35421a,a35422a,a35423a,a35427a,a35428a,a35431a,a35434a,a35435a,a35436a,a35440a,a35441a,a35445a,a35446a,a35447a,a35451a,a35452a,a35455a,a35458a,a35459a,a35460a,a35464a,a35465a,a35469a,a35470a,a35471a,a35475a,a35476a,a35479a,a35482a,a35483a,a35484a,a35488a,a35489a,a35493a,a35494a,a35495a,a35499a,a35500a,a35503a,a35506a,a35507a,a35508a,a35512a,a35513a,a35517a,a35518a,a35519a,a35523a,a35524a,a35527a,a35530a,a35531a,a35532a,a35536a,a35537a,a35541a,a35542a,a35543a,a35547a,a35548a,a35551a,a35554a,a35555a,a35556a,a35560a,a35561a,a35565a,a35566a,a35567a,a35571a,a35572a,a35575a,a35578a,a35579a,a35580a,a35584a,a35585a,a35589a,a35590a,a35591a,a35595a,a35596a,a35599a,a35602a,a35603a,a35604a,a35608a,a35609a,a35613a,a35614a,a35615a,a35619a,a35620a,a35623a,a35626a,a35627a,a35628a,a35632a,a35633a,a35637a,a35638a,a35639a,a35643a,a35644a,a35647a,a35650a,a35651a,a35652a,a35656a,a35657a,a35661a,a35662a,a35663a,a35667a,a35668a,a35671a,a35674a,a35675a,a35676a,a35680a,a35681a,a35685a,a35686a,a35687a,a35691a,a35692a,a35695a,a35698a,a35699a,a35700a,a35704a,a35705a,a35709a,a35710a,a35711a,a35715a,a35716a,a35719a,a35722a,a35723a,a35724a,a35728a,a35729a,a35733a,a35734a,a35735a,a35739a,a35740a,a35743a,a35746a,a35747a,a35748a,a35752a,a35753a,a35757a,a35758a,a35759a,a35763a,a35764a,a35767a,a35770a,a35771a,a35772a,a35776a,a35777a,a35781a,a35782a,a35783a,a35787a,a35788a,a35791a,a35794a,a35795a,a35796a,a35800a,a35801a,a35805a,a35806a,a35807a,a35811a,a35812a,a35815a,a35818a,a35819a,a35820a,a35824a,a35825a,a35829a,a35830a,a35831a,a35835a,a35836a,a35839a,a35842a,a35843a,a35844a,a35848a,a35849a,a35853a,a35854a,a35855a,a35859a,a35860a,a35863a,a35866a,a35867a,a35868a,a35872a,a35873a,a35877a,a35878a,a35879a,a35883a,a35884a,a35887a,a35890a,a35891a,a35892a,a35896a,a35897a,a35901a,a35902a,a35903a,a35907a,a35908a,a35911a,a35914a,a35915a,a35916a,a35920a,a35921a,a35925a,a35926a,a35927a,a35931a,a35932a,a35935a,a35938a,a35939a,a35940a,a35944a,a35945a,a35949a,a35950a,a35951a,a35955a,a35956a,a35959a,a35962a,a35963a,a35964a,a35968a,a35969a,a35973a,a35974a,a35975a,a35979a,a35980a,a35983a,a35986a,a35987a,a35988a,a35992a,a35993a,a35997a,a35998a,a35999a,a36003a,a36004a,a36007a,a36010a,a36011a,a36012a,a36016a,a36017a,a36021a,a36022a,a36023a,a36027a,a36028a,a36031a,a36034a,a36035a,a36036a,a36040a,a36041a,a36045a,a36046a,a36047a,a36051a,a36052a,a36055a,a36058a,a36059a,a36060a,a36064a,a36065a,a36069a,a36070a,a36071a,a36075a,a36076a,a36079a,a36082a,a36083a,a36084a,a36088a,a36089a,a36093a,a36094a,a36095a,a36099a,a36100a,a36103a,a36106a,a36107a,a36108a,a36112a,a36113a,a36117a,a36118a,a36119a,a36123a,a36124a,a36127a,a36130a,a36131a,a36132a,a36136a,a36137a,a36141a,a36142a,a36143a,a36147a,a36148a,a36151a,a36154a,a36155a,a36156a,a36160a,a36161a,a36165a,a36166a,a36167a,a36171a,a36172a,a36175a,a36178a,a36179a,a36180a,a36184a,a36185a,a36189a,a36190a,a36191a,a36195a,a36196a,a36199a,a36202a,a36203a,a36204a,a36208a,a36209a,a36213a,a36214a,a36215a,a36219a,a36220a,a36223a,a36226a,a36227a,a36228a,a36232a,a36233a,a36237a,a36238a,a36239a,a36243a,a36244a,a36247a,a36250a,a36251a,a36252a,a36256a,a36257a,a36261a,a36262a,a36263a,a36267a,a36268a,a36271a,a36274a,a36275a,a36276a,a36280a,a36281a,a36285a,a36286a,a36287a,a36291a,a36292a,a36295a,a36298a,a36299a,a36300a,a36304a,a36305a,a36309a,a36310a,a36311a,a36315a,a36316a,a36319a,a36322a,a36323a,a36324a,a36328a,a36329a,a36333a,a36334a,a36335a,a36339a,a36340a,a36343a,a36346a,a36347a,a36348a,a36352a,a36353a,a36357a,a36358a,a36359a,a36363a,a36364a,a36367a,a36370a,a36371a,a36372a,a36376a,a36377a,a36381a,a36382a,a36383a,a36387a,a36388a,a36391a,a36394a,a36395a,a36396a,a36400a,a36401a,a36405a,a36406a,a36407a,a36411a,a36412a,a36415a,a36418a,a36419a,a36420a,a36424a,a36425a,a36429a,a36430a,a36431a,a36435a,a36436a,a36439a,a36442a,a36443a,a36444a,a36448a,a36449a,a36453a,a36454a,a36455a,a36459a,a36460a,a36463a,a36466a,a36467a,a36468a,a36472a,a36473a,a36477a,a36478a,a36479a,a36483a,a36484a,a36487a,a36490a,a36491a,a36492a,a36496a,a36497a,a36501a,a36502a,a36503a,a36507a,a36508a,a36511a,a36514a,a36515a,a36516a,a36520a,a36521a,a36525a,a36526a,a36527a,a36531a,a36532a,a36535a,a36538a,a36539a,a36540a,a36544a,a36545a,a36549a,a36550a,a36551a,a36555a,a36556a,a36559a,a36562a,a36563a,a36564a,a36568a,a36569a,a36573a,a36574a,a36575a,a36579a,a36580a,a36583a,a36586a,a36587a,a36588a,a36592a,a36593a,a36597a,a36598a,a36599a,a36603a,a36604a,a36607a,a36610a,a36611a,a36612a,a36616a,a36617a,a36621a,a36622a,a36623a,a36627a,a36628a,a36631a,a36634a,a36635a,a36636a,a36640a,a36641a,a36645a,a36646a,a36647a,a36651a,a36652a,a36655a,a36658a,a36659a,a36660a,a36664a,a36665a,a36669a,a36670a,a36671a,a36675a,a36676a,a36679a,a36682a,a36683a,a36684a,a36688a,a36689a,a36693a,a36694a,a36695a,a36699a,a36700a,a36703a,a36706a,a36707a,a36708a,a36712a,a36713a,a36717a,a36718a,a36719a,a36723a,a36724a,a36727a,a36730a,a36731a,a36732a,a36736a,a36737a,a36741a,a36742a,a36743a,a36747a,a36748a,a36751a,a36754a,a36755a,a36756a,a36760a,a36761a,a36765a,a36766a,a36767a,a36771a,a36772a,a36775a,a36778a,a36779a,a36780a,a36784a,a36785a,a36789a,a36790a,a36791a,a36795a,a36796a,a36799a,a36802a,a36803a,a36804a,a36808a,a36809a,a36813a,a36814a,a36815a,a36819a,a36820a,a36823a,a36826a,a36827a,a36828a,a36832a,a36833a,a36837a,a36838a,a36839a,a36843a,a36844a,a36847a,a36850a,a36851a,a36852a,a36856a,a36857a,a36861a,a36862a,a36863a,a36867a,a36868a,a36871a,a36874a,a36875a,a36876a,a36880a,a36881a,a36885a,a36886a,a36887a,a36891a,a36892a,a36895a,a36898a,a36899a,a36900a,a36904a,a36905a,a36909a,a36910a,a36911a,a36915a,a36916a,a36919a,a36922a,a36923a,a36924a,a36928a,a36929a,a36933a,a36934a,a36935a,a36939a,a36940a,a36943a,a36946a,a36947a,a36948a,a36952a,a36953a,a36957a,a36958a,a36959a,a36963a,a36964a,a36967a,a36970a,a36971a,a36972a,a36976a,a36977a,a36981a,a36982a,a36983a,a36987a,a36988a,a36991a,a36994a,a36995a,a36996a,a37000a,a37001a,a37005a,a37006a,a37007a,a37011a,a37012a,a37015a,a37018a,a37019a,a37020a,a37024a,a37025a,a37029a,a37030a,a37031a,a37035a,a37036a,a37039a,a37042a,a37043a,a37044a,a37048a,a37049a,a37053a,a37054a,a37055a,a37059a,a37060a,a37063a,a37066a,a37067a,a37068a,a37072a,a37073a,a37077a,a37078a,a37079a,a37083a,a37084a,a37087a,a37090a,a37091a,a37092a,a37096a,a37097a,a37101a,a37102a,a37103a,a37107a,a37108a,a37111a,a37114a,a37115a,a37116a,a37120a,a37121a,a37125a,a37126a,a37127a,a37131a,a37132a,a37135a,a37138a,a37139a,a37140a,a37144a,a37145a,a37149a,a37150a,a37151a,a37155a,a37156a,a37159a,a37162a,a37163a,a37164a,a37168a,a37169a,a37173a,a37174a,a37175a,a37179a,a37180a,a37183a,a37186a,a37187a,a37188a,a37192a,a37193a,a37197a,a37198a,a37199a,a37203a,a37204a,a37207a,a37210a,a37211a,a37212a,a37216a,a37217a,a37221a,a37222a,a37223a,a37227a,a37228a,a37231a,a37234a,a37235a,a37236a,a37240a,a37241a,a37245a,a37246a,a37247a,a37251a,a37252a,a37255a,a37258a,a37259a,a37260a,a37264a,a37265a,a37269a,a37270a,a37271a,a37275a,a37276a,a37279a,a37282a,a37283a,a37284a,a37288a,a37289a,a37293a,a37294a,a37295a,a37299a,a37300a,a37303a,a37306a,a37307a,a37308a,a37312a,a37313a,a37317a,a37318a,a37319a,a37323a,a37324a,a37327a,a37330a,a37331a,a37332a,a37336a,a37337a,a37341a,a37342a,a37343a,a37347a,a37348a,a37351a,a37354a,a37355a,a37356a,a37360a,a37361a,a37365a,a37366a,a37367a,a37371a,a37372a,a37375a,a37378a,a37379a,a37380a,a37384a,a37385a,a37389a,a37390a,a37391a,a37395a,a37396a,a37399a,a37402a,a37403a,a37404a,a37408a,a37409a,a37413a,a37414a,a37415a,a37419a,a37420a,a37423a,a37426a,a37427a,a37428a,a37432a,a37433a,a37437a,a37438a,a37439a,a37443a,a37444a,a37447a,a37450a,a37451a,a37452a,a37456a,a37457a,a37461a,a37462a,a37463a,a37467a,a37468a,a37471a,a37474a,a37475a,a37476a,a37480a,a37481a,a37485a,a37486a,a37487a,a37491a,a37492a,a37495a,a37498a,a37499a,a37500a,a37504a,a37505a,a37509a,a37510a,a37511a,a37515a,a37516a,a37519a,a37522a,a37523a,a37524a,a37528a,a37529a,a37533a,a37534a,a37535a,a37539a,a37540a,a37543a,a37546a,a37547a,a37548a,a37552a,a37553a,a37557a,a37558a,a37559a,a37563a,a37564a,a37567a,a37570a,a37571a,a37572a,a37576a,a37577a,a37581a,a37582a,a37583a,a37587a,a37588a,a37591a,a37594a,a37595a,a37596a,a37600a,a37601a,a37605a,a37606a,a37607a,a37611a,a37612a,a37615a,a37618a,a37619a,a37620a,a37624a,a37625a,a37629a,a37630a,a37631a,a37635a,a37636a,a37639a,a37642a,a37643a,a37644a,a37648a,a37649a,a37653a,a37654a,a37655a,a37659a,a37660a,a37663a,a37666a,a37667a,a37668a,a37672a,a37673a,a37677a,a37678a,a37679a,a37683a,a37684a,a37687a,a37690a,a37691a,a37692a,a37696a,a37697a,a37701a,a37702a,a37703a,a37707a,a37708a,a37711a,a37714a,a37715a,a37716a,a37720a,a37721a,a37725a,a37726a,a37727a,a37731a,a37732a,a37735a,a37738a,a37739a,a37740a,a37744a,a37745a,a37749a,a37750a,a37751a,a37755a,a37756a,a37759a,a37762a,a37763a,a37764a,a37768a,a37769a,a37773a,a37774a,a37775a,a37779a,a37780a,a37783a,a37786a,a37787a,a37788a,a37792a,a37793a,a37797a,a37798a,a37799a,a37803a,a37804a,a37807a,a37810a,a37811a,a37812a,a37816a,a37817a,a37821a,a37822a,a37823a,a37827a,a37828a,a37831a,a37834a,a37835a,a37836a,a37840a,a37841a,a37845a,a37846a,a37847a,a37851a,a37852a,a37855a,a37858a,a37859a,a37860a,a37864a,a37865a,a37869a,a37870a,a37871a,a37875a,a37876a,a37879a,a37882a,a37883a,a37884a,a37888a,a37889a,a37893a,a37894a,a37895a,a37899a,a37900a,a37903a,a37906a,a37907a,a37908a,a37912a,a37913a,a37917a,a37918a,a37919a,a37923a,a37924a,a37927a,a37930a,a37931a,a37932a,a37936a,a37937a,a37941a,a37942a,a37943a,a37947a,a37948a,a37951a,a37954a,a37955a,a37956a,a37960a,a37961a,a37965a,a37966a,a37967a,a37971a,a37972a,a37975a,a37978a,a37979a,a37980a,a37984a,a37985a,a37989a,a37990a,a37991a,a37995a,a37996a,a37999a,a38002a,a38003a,a38004a,a38008a,a38009a,a38013a,a38014a,a38015a,a38019a,a38020a,a38023a,a38026a,a38027a,a38028a,a38032a,a38033a,a38037a,a38038a,a38039a,a38043a,a38044a,a38047a,a38050a,a38051a,a38052a,a38056a,a38057a,a38061a,a38062a,a38063a,a38067a,a38068a,a38071a,a38074a,a38075a,a38076a,a38080a,a38081a,a38085a,a38086a,a38087a,a38091a,a38092a,a38095a,a38098a,a38099a,a38100a,a38104a,a38105a,a38109a,a38110a,a38111a,a38115a,a38116a,a38119a,a38122a,a38123a,a38124a,a38128a,a38129a,a38133a,a38134a,a38135a,a38139a,a38140a,a38143a,a38146a,a38147a,a38148a,a38152a,a38153a,a38157a,a38158a,a38159a,a38163a,a38164a,a38167a,a38170a,a38171a,a38172a,a38176a,a38177a,a38181a,a38182a,a38183a,a38187a,a38188a,a38191a,a38194a,a38195a,a38196a,a38200a,a38201a,a38205a,a38206a,a38207a,a38211a,a38212a,a38215a,a38218a,a38219a,a38220a,a38224a,a38225a,a38229a,a38230a,a38231a,a38235a,a38236a,a38239a,a38242a,a38243a,a38244a,a38248a,a38249a,a38253a,a38254a,a38255a,a38259a,a38260a,a38263a,a38266a,a38267a,a38268a,a38272a,a38273a,a38277a,a38278a,a38279a,a38283a,a38284a,a38287a,a38290a,a38291a,a38292a,a38296a,a38297a,a38301a,a38302a,a38303a,a38307a,a38308a,a38311a,a38314a,a38315a,a38316a,a38320a,a38321a,a38325a,a38326a,a38327a,a38331a,a38332a,a38335a,a38338a,a38339a,a38340a,a38344a,a38345a,a38349a,a38350a,a38351a,a38355a,a38356a,a38359a,a38362a,a38363a,a38364a,a38368a,a38369a,a38373a,a38374a,a38375a,a38379a,a38380a,a38383a,a38386a,a38387a,a38388a,a38392a,a38393a,a38397a,a38398a,a38399a,a38403a,a38404a,a38407a,a38410a,a38411a,a38412a,a38416a,a38417a,a38421a,a38422a,a38423a,a38427a,a38428a,a38431a,a38434a,a38435a,a38436a,a38440a,a38441a,a38445a,a38446a,a38447a,a38451a,a38452a,a38455a,a38458a,a38459a,a38460a,a38464a,a38465a,a38469a,a38470a,a38471a,a38475a,a38476a,a38479a,a38482a,a38483a,a38484a,a38488a,a38489a,a38493a,a38494a,a38495a,a38499a,a38500a,a38503a,a38506a,a38507a,a38508a,a38512a,a38513a,a38517a,a38518a,a38519a,a38523a,a38524a,a38527a,a38530a,a38531a,a38532a,a38536a,a38537a,a38541a,a38542a,a38543a,a38547a,a38548a,a38551a,a38554a,a38555a,a38556a,a38560a,a38561a,a38565a,a38566a,a38567a,a38571a,a38572a,a38575a,a38578a,a38579a,a38580a,a38584a,a38585a,a38589a,a38590a,a38591a,a38595a,a38596a,a38599a,a38602a,a38603a,a38604a,a38608a,a38609a,a38613a,a38614a,a38615a,a38619a,a38620a,a38623a,a38626a,a38627a,a38628a,a38632a,a38633a,a38637a,a38638a,a38639a,a38643a,a38644a,a38647a,a38650a,a38651a,a38652a,a38656a,a38657a,a38661a,a38662a,a38663a,a38667a,a38668a,a38671a,a38674a,a38675a,a38676a,a38680a,a38681a,a38685a,a38686a,a38687a,a38691a,a38692a,a38695a,a38698a,a38699a,a38700a,a38704a,a38705a,a38709a,a38710a,a38711a,a38715a,a38716a,a38719a,a38722a,a38723a,a38724a,a38728a,a38729a,a38733a,a38734a,a38735a,a38739a,a38740a,a38743a,a38746a,a38747a,a38748a,a38752a,a38753a,a38757a,a38758a,a38759a,a38763a,a38764a,a38767a,a38770a,a38771a,a38772a,a38776a,a38777a,a38781a,a38782a,a38783a,a38787a,a38788a,a38791a,a38794a,a38795a,a38796a,a38800a,a38801a,a38805a,a38806a,a38807a,a38811a,a38812a,a38815a,a38818a,a38819a,a38820a,a38824a,a38825a,a38829a,a38830a,a38831a,a38835a,a38836a,a38839a,a38842a,a38843a,a38844a,a38848a,a38849a,a38853a,a38854a,a38855a,a38859a,a38860a,a38863a,a38866a,a38867a,a38868a,a38872a,a38873a,a38877a,a38878a,a38879a,a38883a,a38884a,a38887a,a38890a,a38891a,a38892a,a38896a,a38897a,a38901a,a38902a,a38903a,a38907a,a38908a,a38911a,a38914a,a38915a,a38916a,a38920a,a38921a,a38925a,a38926a,a38927a,a38931a,a38932a,a38935a,a38938a,a38939a,a38940a,a38944a,a38945a,a38949a,a38950a,a38951a,a38955a,a38956a,a38959a,a38962a,a38963a,a38964a,a38968a,a38969a,a38973a,a38974a,a38975a,a38979a,a38980a,a38983a,a38986a,a38987a,a38988a,a38992a,a38993a,a38997a,a38998a,a38999a,a39003a,a39004a,a39007a,a39010a,a39011a,a39012a,a39016a,a39017a,a39021a,a39022a,a39023a,a39027a,a39028a,a39031a,a39034a,a39035a,a39036a,a39040a,a39041a,a39045a,a39046a,a39047a,a39051a,a39052a,a39055a,a39058a,a39059a,a39060a,a39064a,a39065a,a39069a,a39070a,a39071a,a39075a,a39076a,a39079a,a39082a,a39083a,a39084a,a39088a,a39089a,a39093a,a39094a,a39095a,a39099a,a39100a,a39103a,a39106a,a39107a,a39108a,a39112a,a39113a,a39117a,a39118a,a39119a,a39123a,a39124a,a39127a,a39130a,a39131a,a39132a,a39136a,a39137a,a39141a,a39142a,a39143a,a39147a,a39148a,a39151a,a39154a,a39155a,a39156a,a39160a,a39161a,a39165a,a39166a,a39167a,a39171a,a39172a,a39175a,a39178a,a39179a,a39180a,a39184a,a39185a,a39189a,a39190a,a39191a,a39195a,a39196a,a39199a,a39202a,a39203a,a39204a,a39208a,a39209a,a39213a,a39214a,a39215a,a39219a,a39220a,a39223a,a39226a,a39227a,a39228a,a39232a,a39233a,a39237a,a39238a,a39239a,a39243a,a39244a,a39247a,a39250a,a39251a,a39252a,a39256a,a39257a,a39261a,a39262a,a39263a,a39267a,a39268a,a39271a,a39274a,a39275a,a39276a,a39280a,a39281a,a39285a,a39286a,a39287a,a39291a,a39292a,a39295a,a39298a,a39299a,a39300a,a39304a,a39305a,a39309a,a39310a,a39311a,a39315a,a39316a,a39319a,a39322a,a39323a,a39324a,a39328a,a39329a,a39333a,a39334a,a39335a,a39339a,a39340a,a39343a,a39346a,a39347a,a39348a,a39352a,a39353a,a39357a,a39358a,a39359a,a39363a,a39364a,a39367a,a39370a,a39371a,a39372a,a39376a,a39377a,a39381a,a39382a,a39383a,a39387a,a39388a,a39391a,a39394a,a39395a,a39396a,a39400a,a39401a,a39405a,a39406a,a39407a,a39411a,a39412a,a39415a,a39418a,a39419a,a39420a,a39424a,a39425a,a39429a,a39430a,a39431a,a39435a,a39436a,a39439a,a39442a,a39443a,a39444a,a39448a,a39449a,a39453a,a39454a,a39455a,a39459a,a39460a,a39463a,a39466a,a39467a,a39468a,a39472a,a39473a,a39477a,a39478a,a39479a,a39483a,a39484a,a39487a,a39490a,a39491a,a39492a,a39496a,a39497a,a39501a,a39502a,a39503a,a39507a,a39508a,a39511a,a39514a,a39515a,a39516a,a39520a,a39521a,a39525a,a39526a,a39527a,a39531a,a39532a,a39535a,a39538a,a39539a,a39540a,a39544a,a39545a,a39549a,a39550a,a39551a,a39555a,a39556a,a39559a,a39562a,a39563a,a39564a,a39568a,a39569a,a39573a,a39574a,a39575a,a39579a,a39580a,a39583a,a39586a,a39587a,a39588a,a39592a,a39593a,a39597a,a39598a,a39599a,a39603a,a39604a,a39607a,a39610a,a39611a,a39612a,a39616a,a39617a,a39621a,a39622a,a39623a,a39627a,a39628a,a39631a,a39634a,a39635a,a39636a,a39640a,a39641a,a39645a,a39646a,a39647a,a39651a,a39652a,a39655a,a39658a,a39659a,a39660a,a39664a,a39665a,a39669a,a39670a,a39671a,a39675a,a39676a,a39679a,a39682a,a39683a,a39684a,a39688a,a39689a,a39693a,a39694a,a39695a,a39699a,a39700a,a39703a,a39706a,a39707a,a39708a,a39712a,a39713a,a39717a,a39718a,a39719a,a39723a,a39724a,a39727a,a39730a,a39731a,a39732a,a39736a,a39737a,a39741a,a39742a,a39743a,a39747a,a39748a,a39751a,a39754a,a39755a,a39756a,a39760a,a39761a,a39765a,a39766a,a39767a,a39771a,a39772a,a39775a,a39778a,a39779a,a39780a,a39784a,a39785a,a39789a,a39790a,a39791a,a39795a,a39796a,a39799a,a39802a,a39803a,a39804a,a39808a,a39809a,a39813a,a39814a,a39815a,a39819a,a39820a,a39823a,a39826a,a39827a,a39828a,a39832a,a39833a,a39837a,a39838a,a39839a,a39843a,a39844a,a39847a,a39850a,a39851a,a39852a,a39856a,a39857a,a39861a,a39862a,a39863a,a39867a,a39868a,a39871a,a39874a,a39875a,a39876a,a39880a,a39881a,a39885a,a39886a,a39887a,a39891a,a39892a,a39895a,a39898a,a39899a,a39900a,a39904a,a39905a,a39909a,a39910a,a39911a,a39915a,a39916a,a39919a,a39922a,a39923a,a39924a,a39928a,a39929a,a39933a,a39934a,a39935a,a39939a,a39940a,a39943a,a39946a,a39947a,a39948a,a39952a,a39953a,a39957a,a39958a,a39959a,a39963a,a39964a,a39967a,a39970a,a39971a,a39972a,a39976a,a39977a,a39981a,a39982a,a39983a,a39987a,a39988a,a39991a,a39994a,a39995a,a39996a,a40000a,a40001a,a40005a,a40006a,a40007a,a40011a,a40012a,a40015a,a40018a,a40019a,a40020a,a40024a,a40025a,a40029a,a40030a,a40031a,a40035a,a40036a,a40039a,a40042a,a40043a,a40044a,a40048a,a40049a,a40053a,a40054a,a40055a,a40059a,a40060a,a40063a,a40066a,a40067a,a40068a,a40072a,a40073a,a40077a,a40078a,a40079a,a40083a,a40084a,a40087a,a40090a,a40091a,a40092a,a40096a,a40097a,a40101a,a40102a,a40103a,a40107a,a40108a,a40111a,a40114a,a40115a,a40116a,a40120a,a40121a,a40125a,a40126a,a40127a,a40131a,a40132a,a40135a,a40138a,a40139a,a40140a,a40144a,a40145a,a40149a,a40150a,a40151a,a40155a,a40156a,a40159a,a40162a,a40163a,a40164a,a40168a,a40169a,a40173a,a40174a,a40175a,a40179a,a40180a,a40183a,a40186a,a40187a,a40188a,a40192a,a40193a,a40197a,a40198a,a40199a,a40203a,a40204a,a40207a,a40210a,a40211a,a40212a,a40216a,a40217a,a40221a,a40222a,a40223a,a40227a,a40228a,a40231a,a40234a,a40235a,a40236a,a40240a,a40241a,a40245a,a40246a,a40247a,a40251a,a40252a,a40255a,a40258a,a40259a,a40260a,a40264a,a40265a,a40269a,a40270a,a40271a,a40275a,a40276a,a40279a,a40282a,a40283a,a40284a,a40288a,a40289a,a40293a,a40294a,a40295a,a40299a,a40300a,a40303a,a40306a,a40307a,a40308a,a40312a,a40313a,a40317a,a40318a,a40319a,a40323a,a40324a,a40327a,a40330a,a40331a,a40332a,a40336a,a40337a,a40341a,a40342a,a40343a,a40347a,a40348a,a40351a,a40354a,a40355a,a40356a,a40360a,a40361a,a40365a,a40366a,a40367a,a40371a,a40372a,a40375a,a40378a,a40379a,a40380a,a40384a,a40385a,a40389a,a40390a,a40391a,a40395a,a40396a,a40399a,a40402a,a40403a,a40404a,a40408a,a40409a,a40413a,a40414a,a40415a,a40419a,a40420a,a40423a,a40426a,a40427a,a40428a,a40432a,a40433a,a40437a,a40438a,a40439a,a40443a,a40444a,a40447a,a40450a,a40451a,a40452a,a40456a,a40457a,a40461a,a40462a,a40463a,a40467a,a40468a,a40471a,a40474a,a40475a,a40476a,a40480a,a40481a,a40485a,a40486a,a40487a,a40491a,a40492a,a40495a,a40498a,a40499a,a40500a,a40504a,a40505a,a40509a,a40510a,a40511a,a40515a,a40516a,a40519a,a40522a,a40523a,a40524a,a40528a,a40529a,a40533a,a40534a,a40535a,a40539a,a40540a,a40543a,a40546a,a40547a,a40548a,a40552a,a40553a,a40557a,a40558a,a40559a,a40563a,a40564a,a40567a,a40570a,a40571a,a40572a,a40576a,a40577a,a40581a,a40582a,a40583a,a40587a,a40588a,a40591a,a40594a,a40595a,a40596a,a40600a,a40601a,a40605a,a40606a,a40607a,a40611a,a40612a,a40615a,a40618a,a40619a,a40620a,a40624a,a40625a,a40629a,a40630a,a40631a,a40635a,a40636a,a40639a,a40642a,a40643a,a40644a,a40648a,a40649a,a40653a,a40654a,a40655a,a40659a,a40660a,a40663a,a40666a,a40667a,a40668a,a40672a,a40673a,a40677a,a40678a,a40679a,a40683a,a40684a,a40687a,a40690a,a40691a,a40692a,a40696a,a40697a,a40701a,a40702a,a40703a,a40707a,a40708a,a40711a,a40714a,a40715a,a40716a,a40720a,a40721a,a40725a,a40726a,a40727a,a40731a,a40732a,a40735a,a40738a,a40739a,a40740a,a40744a,a40745a,a40749a,a40750a,a40751a,a40755a,a40756a,a40759a,a40762a,a40763a,a40764a,a40768a,a40769a,a40773a,a40774a,a40775a,a40779a,a40780a,a40783a,a40786a,a40787a,a40788a,a40792a,a40793a,a40797a,a40798a,a40799a,a40803a,a40804a,a40807a,a40810a,a40811a,a40812a,a40816a,a40817a,a40821a,a40822a,a40823a,a40827a,a40828a,a40831a,a40834a,a40835a,a40836a,a40840a,a40841a,a40845a,a40846a,a40847a,a40851a,a40852a,a40855a,a40858a,a40859a,a40860a,a40864a,a40865a,a40869a,a40870a,a40871a,a40875a,a40876a,a40879a,a40882a,a40883a,a40884a,a40888a,a40889a,a40893a,a40894a,a40895a,a40899a,a40900a,a40903a,a40906a,a40907a,a40908a,a40912a,a40913a,a40917a,a40918a,a40919a,a40923a,a40924a,a40927a,a40930a,a40931a,a40932a,a40936a,a40937a,a40941a,a40942a,a40943a,a40947a,a40948a,a40951a,a40954a,a40955a,a40956a,a40960a,a40961a,a40965a,a40966a,a40967a,a40971a,a40972a,a40975a,a40978a,a40979a,a40980a,a40984a,a40985a,a40989a,a40990a,a40991a,a40995a,a40996a,a40999a,a41002a,a41003a,a41004a,a41008a,a41009a,a41013a,a41014a,a41015a,a41019a,a41020a,a41023a,a41026a,a41027a,a41028a,a41032a,a41033a,a41037a,a41038a,a41039a,a41043a,a41044a,a41047a,a41050a,a41051a,a41052a,a41056a,a41057a,a41061a,a41062a,a41063a,a41067a,a41068a,a41071a,a41074a,a41075a,a41076a,a41080a,a41081a,a41085a,a41086a,a41087a,a41091a,a41092a,a41095a,a41098a,a41099a,a41100a,a41104a,a41105a,a41109a,a41110a,a41111a,a41115a,a41116a,a41119a,a41122a,a41123a,a41124a,a41128a,a41129a,a41133a,a41134a,a41135a,a41139a,a41140a,a41143a,a41146a,a41147a,a41148a,a41152a,a41153a,a41157a,a41158a,a41159a,a41163a,a41164a,a41167a,a41170a,a41171a,a41172a,a41176a,a41177a,a41181a,a41182a,a41183a,a41187a,a41188a,a41191a,a41194a,a41195a,a41196a,a41200a,a41201a,a41205a,a41206a,a41207a,a41211a,a41212a,a41215a,a41218a,a41219a,a41220a,a41224a,a41225a,a41229a,a41230a,a41231a,a41235a,a41236a,a41239a,a41242a,a41243a,a41244a,a41248a,a41249a,a41253a,a41254a,a41255a,a41259a,a41260a,a41263a,a41266a,a41267a,a41268a,a41272a,a41273a,a41277a,a41278a,a41279a,a41283a,a41284a,a41287a,a41290a,a41291a,a41292a,a41296a,a41297a,a41301a,a41302a,a41303a,a41307a,a41308a,a41311a,a41314a,a41315a,a41316a,a41320a,a41321a,a41325a,a41326a,a41327a,a41331a,a41332a,a41335a,a41338a,a41339a,a41340a,a41344a,a41345a,a41349a,a41350a,a41351a,a41355a,a41356a,a41359a,a41362a,a41363a,a41364a,a41368a,a41369a,a41373a,a41374a,a41375a,a41379a,a41380a,a41383a,a41386a,a41387a,a41388a,a41392a,a41393a,a41397a,a41398a,a41399a,a41403a,a41404a,a41407a,a41410a,a41411a,a41412a,a41416a,a41417a,a41421a,a41422a,a41423a,a41427a,a41428a,a41431a,a41434a,a41435a,a41436a,a41440a,a41441a,a41445a,a41446a,a41447a,a41451a,a41452a,a41455a,a41458a,a41459a,a41460a,a41464a,a41465a,a41469a,a41470a,a41471a,a41475a,a41476a,a41479a,a41482a,a41483a,a41484a,a41488a,a41489a,a41493a,a41494a,a41495a,a41499a,a41500a,a41503a,a41506a,a41507a,a41508a,a41512a,a41513a,a41517a,a41518a,a41519a,a41523a,a41524a,a41527a,a41530a,a41531a,a41532a,a41536a,a41537a,a41541a,a41542a,a41543a,a41547a,a41548a,a41551a,a41554a,a41555a,a41556a,a41560a,a41561a,a41565a,a41566a,a41567a,a41571a,a41572a,a41575a,a41578a,a41579a,a41580a,a41584a,a41585a,a41589a,a41590a,a41591a,a41595a,a41596a,a41599a,a41602a,a41603a,a41604a,a41608a,a41609a,a41613a,a41614a,a41615a,a41619a,a41620a,a41623a,a41626a,a41627a,a41628a,a41632a,a41633a,a41637a,a41638a,a41639a,a41643a,a41644a,a41647a,a41650a,a41651a,a41652a,a41656a,a41657a,a41661a,a41662a,a41663a,a41667a,a41668a,a41671a,a41674a,a41675a,a41676a,a41680a,a41681a,a41685a,a41686a,a41687a,a41691a,a41692a,a41695a,a41698a,a41699a,a41700a,a41704a,a41705a,a41709a,a41710a,a41711a,a41715a,a41716a,a41719a,a41722a,a41723a,a41724a,a41728a,a41729a,a41733a,a41734a,a41735a,a41739a,a41740a,a41743a,a41746a,a41747a,a41748a,a41752a,a41753a,a41757a,a41758a,a41759a,a41763a,a41764a,a41767a,a41770a,a41771a,a41772a,a41776a,a41777a,a41781a,a41782a,a41783a,a41787a,a41788a,a41791a,a41794a,a41795a,a41796a,a41800a,a41801a,a41805a,a41806a,a41807a,a41811a,a41812a,a41815a,a41818a,a41819a,a41820a,a41824a,a41825a,a41829a,a41830a,a41831a,a41835a,a41836a,a41839a,a41842a,a41843a,a41844a,a41848a,a41849a,a41853a,a41854a,a41855a,a41859a,a41860a,a41863a,a41866a,a41867a,a41868a,a41872a,a41873a,a41877a,a41878a,a41879a,a41883a,a41884a,a41887a,a41890a,a41891a,a41892a,a41896a,a41897a,a41901a,a41902a,a41903a,a41907a,a41908a,a41911a,a41914a,a41915a,a41916a,a41920a,a41921a,a41925a,a41926a,a41927a,a41931a,a41932a,a41935a,a41938a,a41939a,a41940a,a41944a,a41945a,a41949a,a41950a,a41951a,a41955a,a41956a,a41959a,a41962a,a41963a,a41964a,a41968a,a41969a,a41973a,a41974a,a41975a,a41979a,a41980a,a41983a,a41986a,a41987a,a41988a,a41992a,a41993a,a41997a,a41998a,a41999a,a42003a,a42004a,a42007a,a42010a,a42011a,a42012a,a42016a,a42017a,a42021a,a42022a,a42023a,a42027a,a42028a,a42031a,a42034a,a42035a,a42036a,a42040a,a42041a,a42045a,a42046a,a42047a,a42051a,a42052a,a42055a,a42058a,a42059a,a42060a,a42064a,a42065a,a42069a,a42070a,a42071a,a42075a,a42076a,a42079a,a42082a,a42083a,a42084a,a42088a,a42089a,a42093a,a42094a,a42095a,a42099a,a42100a,a42103a,a42106a,a42107a,a42108a,a42112a,a42113a,a42117a,a42118a,a42119a,a42123a,a42124a,a42127a,a42130a,a42131a,a42132a,a42136a,a42137a,a42141a,a42142a,a42143a,a42147a,a42148a,a42151a,a42154a,a42155a,a42156a,a42160a,a42161a,a42165a,a42166a,a42167a,a42171a,a42172a,a42175a,a42178a,a42179a,a42180a,a42184a,a42185a,a42189a,a42190a,a42191a,a42195a,a42196a,a42199a,a42202a,a42203a,a42204a,a42208a,a42209a,a42213a,a42214a,a42215a,a42219a,a42220a,a42223a,a42226a,a42227a,a42228a,a42232a,a42233a,a42237a,a42238a,a42239a,a42243a,a42244a,a42247a,a42250a,a42251a,a42252a,a42256a,a42257a,a42261a,a42262a,a42263a,a42267a,a42268a,a42271a,a42274a,a42275a,a42276a,a42280a,a42281a,a42285a,a42286a,a42287a,a42291a,a42292a,a42295a,a42298a,a42299a,a42300a,a42304a,a42305a,a42309a,a42310a,a42311a,a42315a,a42316a,a42319a,a42322a,a42323a,a42324a,a42328a,a42329a,a42333a,a42334a,a42335a,a42339a,a42340a,a42343a,a42346a,a42347a,a42348a,a42352a,a42353a,a42357a,a42358a,a42359a,a42363a,a42364a,a42367a,a42370a,a42371a,a42372a,a42376a,a42377a,a42381a,a42382a,a42383a,a42387a,a42388a,a42391a,a42394a,a42395a,a42396a,a42400a,a42401a,a42405a,a42406a,a42407a,a42411a,a42412a,a42415a,a42418a,a42419a,a42420a,a42424a,a42425a,a42429a,a42430a,a42431a,a42435a,a42436a,a42439a,a42442a,a42443a,a42444a,a42448a,a42449a,a42453a,a42454a,a42455a,a42459a,a42460a,a42463a,a42466a,a42467a,a42468a,a42472a,a42473a,a42477a,a42478a,a42479a,a42483a,a42484a,a42487a,a42490a,a42491a,a42492a,a42496a,a42497a,a42500a,a42503a,a42504a,a42505a,a42509a,a42510a,a42513a,a42516a,a42517a,a42518a,a42522a,a42523a,a42526a,a42529a,a42530a,a42531a,a42535a,a42536a,a42539a,a42542a,a42543a,a42544a,a42548a,a42549a,a42552a,a42555a,a42556a,a42557a,a42561a,a42562a,a42565a,a42568a,a42569a,a42570a,a42574a,a42575a,a42578a,a42581a,a42582a,a42583a,a42587a,a42588a,a42591a,a42594a,a42595a,a42596a,a42600a,a42601a,a42604a,a42607a,a42608a,a42609a,a42613a,a42614a,a42617a,a42620a,a42621a,a42622a,a42626a,a42627a,a42630a,a42633a,a42634a,a42635a,a42639a,a42640a,a42643a,a42646a,a42647a,a42648a,a42652a,a42653a,a42656a,a42659a,a42660a,a42661a,a42665a,a42666a,a42669a,a42672a,a42673a,a42674a,a42678a,a42679a,a42682a,a42685a,a42686a,a42687a,a42691a,a42692a,a42695a,a42698a,a42699a,a42700a,a42704a,a42705a,a42708a,a42711a,a42712a,a42713a,a42717a,a42718a,a42721a,a42724a,a42725a,a42726a,a42730a,a42731a,a42734a,a42737a,a42738a,a42739a,a42743a,a42744a,a42747a,a42750a,a42751a,a42752a,a42756a,a42757a,a42760a,a42763a,a42764a,a42765a,a42769a,a42770a,a42773a,a42776a,a42777a,a42778a,a42782a,a42783a,a42786a,a42789a,a42790a,a42791a,a42795a,a42796a,a42799a,a42802a,a42803a,a42804a,a42808a,a42809a,a42812a,a42815a,a42816a,a42817a,a42821a,a42822a,a42825a,a42828a,a42829a,a42830a,a42834a,a42835a,a42838a,a42841a,a42842a,a42843a,a42847a,a42848a,a42851a,a42854a,a42855a,a42856a,a42860a,a42861a,a42864a,a42867a,a42868a,a42869a,a42873a,a42874a,a42877a,a42880a,a42881a,a42882a,a42886a,a42887a,a42890a,a42893a,a42894a,a42895a,a42899a,a42900a,a42903a,a42906a,a42907a,a42908a,a42912a,a42913a,a42916a,a42919a,a42920a,a42921a,a42925a,a42926a,a42929a,a42932a,a42933a,a42934a,a42938a,a42939a,a42942a,a42945a,a42946a,a42947a,a42951a,a42952a,a42955a,a42958a,a42959a,a42960a,a42964a,a42965a,a42968a,a42971a,a42972a,a42973a,a42977a,a42978a,a42981a,a42984a,a42985a,a42986a,a42990a,a42991a,a42994a,a42997a,a42998a,a42999a,a43003a,a43004a,a43007a,a43010a,a43011a,a43012a,a43016a,a43017a,a43020a,a43023a,a43024a,a43025a,a43029a,a43030a,a43033a,a43036a,a43037a,a43038a,a43042a,a43043a,a43046a,a43049a,a43050a,a43051a,a43055a,a43056a,a43059a,a43062a,a43063a,a43064a,a43068a,a43069a,a43072a,a43075a,a43076a,a43077a,a43081a,a43082a,a43085a,a43088a,a43089a,a43090a,a43094a,a43095a,a43098a,a43101a,a43102a,a43103a,a43107a,a43108a,a43111a,a43114a,a43115a,a43116a,a43120a,a43121a,a43124a,a43127a,a43128a,a43129a,a43133a,a43134a,a43137a,a43140a,a43141a,a43142a,a43146a,a43147a,a43150a,a43153a,a43154a,a43155a,a43159a,a43160a,a43163a,a43166a,a43167a,a43168a,a43172a,a43173a,a43176a,a43179a,a43180a,a43181a,a43185a,a43186a,a43189a,a43192a,a43193a,a43194a,a43198a,a43199a,a43202a,a43205a,a43206a,a43207a,a43211a,a43212a,a43215a,a43218a,a43219a,a43220a,a43224a,a43225a,a43228a,a43231a,a43232a,a43233a,a43237a,a43238a,a43241a,a43244a,a43245a,a43246a,a43250a,a43251a,a43254a,a43257a,a43258a,a43259a,a43263a,a43264a,a43267a,a43270a,a43271a,a43272a,a43276a,a43277a,a43280a,a43283a,a43284a,a43285a,a43289a,a43290a,a43293a,a43296a,a43297a,a43298a,a43302a,a43303a,a43306a,a43309a,a43310a,a43311a,a43315a,a43316a,a43319a,a43322a,a43323a,a43324a,a43328a,a43329a,a43332a,a43335a,a43336a,a43337a,a43341a,a43342a,a43345a,a43348a,a43349a,a43350a,a43354a,a43355a,a43358a,a43361a,a43362a,a43363a,a43367a,a43368a,a43371a,a43374a,a43375a,a43376a,a43380a,a43381a,a43384a,a43387a,a43388a,a43389a,a43393a,a43394a,a43397a,a43400a,a43401a,a43402a,a43406a,a43407a,a43410a,a43413a,a43414a,a43415a,a43419a,a43420a,a43423a,a43426a,a43427a,a43428a,a43432a,a43433a,a43436a,a43439a,a43440a,a43441a,a43445a,a43446a,a43449a,a43452a,a43453a,a43454a,a43458a,a43459a,a43462a,a43465a,a43466a,a43467a,a43471a,a43472a,a43475a,a43478a,a43479a,a43480a,a43484a,a43485a,a43488a,a43491a,a43492a,a43493a,a43497a,a43498a,a43501a,a43504a,a43505a,a43506a,a43510a,a43511a,a43514a,a43517a,a43518a,a43519a,a43523a,a43524a,a43527a,a43530a,a43531a,a43532a,a43536a,a43537a,a43540a,a43543a,a43544a,a43545a,a43549a,a43550a,a43553a,a43556a,a43557a,a43558a,a43562a,a43563a,a43566a,a43569a,a43570a,a43571a,a43575a,a43576a,a43579a,a43582a,a43583a,a43584a,a43588a,a43589a,a43592a,a43595a,a43596a,a43597a,a43601a,a43602a,a43605a,a43608a,a43609a,a43610a,a43614a,a43615a,a43618a,a43621a,a43622a,a43623a,a43627a,a43628a,a43631a,a43634a,a43635a,a43636a,a43640a,a43641a,a43644a,a43647a,a43648a,a43649a,a43653a,a43654a,a43657a,a43660a,a43661a,a43662a,a43666a,a43667a,a43670a,a43673a,a43674a,a43675a,a43679a,a43680a,a43683a,a43686a,a43687a,a43688a,a43692a,a43693a,a43696a,a43699a,a43700a,a43701a,a43705a,a43706a,a43709a,a43712a,a43713a,a43714a,a43718a,a43719a,a43722a,a43725a,a43726a,a43727a,a43731a,a43732a,a43735a,a43738a,a43739a,a43740a,a43744a,a43745a,a43748a,a43751a,a43752a,a43753a,a43757a,a43758a,a43761a,a43764a,a43765a,a43766a,a43770a,a43771a,a43774a,a43777a,a43778a,a43779a,a43783a,a43784a,a43787a,a43790a,a43791a,a43792a,a43796a,a43797a,a43800a,a43803a,a43804a,a43805a,a43809a,a43810a,a43813a,a43816a,a43817a,a43818a,a43822a,a43823a,a43826a,a43829a,a43830a,a43831a,a43835a,a43836a,a43839a,a43842a,a43843a,a43844a,a43848a,a43849a,a43852a,a43855a,a43856a,a43857a,a43861a,a43862a,a43865a,a43868a,a43869a,a43870a,a43874a,a43875a,a43878a,a43881a,a43882a,a43883a,a43887a,a43888a,a43891a,a43894a,a43895a,a43896a,a43900a,a43901a,a43904a,a43907a,a43908a,a43909a,a43913a,a43914a,a43917a,a43920a,a43921a,a43922a,a43926a,a43927a,a43930a,a43933a,a43934a,a43935a,a43939a,a43940a,a43943a,a43946a,a43947a,a43948a,a43952a,a43953a,a43956a,a43959a,a43960a,a43961a,a43965a,a43966a,a43969a,a43972a,a43973a,a43974a,a43978a,a43979a,a43982a,a43985a,a43986a,a43987a,a43991a,a43992a,a43995a,a43998a,a43999a,a44000a,a44004a,a44005a,a44008a,a44011a,a44012a,a44013a,a44017a,a44018a,a44021a,a44024a,a44025a,a44026a,a44030a,a44031a,a44034a,a44037a,a44038a,a44039a,a44043a,a44044a,a44047a,a44050a,a44051a,a44052a,a44056a,a44057a,a44060a,a44063a,a44064a,a44065a,a44069a,a44070a,a44073a,a44076a,a44077a,a44078a,a44082a,a44083a,a44086a,a44089a,a44090a,a44091a,a44095a,a44096a,a44099a,a44102a,a44103a,a44104a,a44108a,a44109a,a44112a,a44115a,a44116a,a44117a,a44121a,a44122a,a44125a,a44128a,a44129a,a44130a,a44134a,a44135a,a44138a,a44141a,a44142a,a44143a,a44147a,a44148a,a44151a,a44154a,a44155a,a44156a,a44160a,a44161a,a44164a,a44167a,a44168a,a44169a,a44173a,a44174a,a44177a,a44180a,a44181a,a44182a,a44186a,a44187a,a44190a,a44193a,a44194a,a44195a,a44199a,a44200a,a44203a,a44206a,a44207a,a44208a,a44212a,a44213a,a44216a,a44219a,a44220a,a44221a,a44225a,a44226a,a44229a,a44232a,a44233a,a44234a,a44238a,a44239a,a44242a,a44245a,a44246a,a44247a,a44251a,a44252a,a44255a,a44258a,a44259a,a44260a,a44264a,a44265a,a44268a,a44271a,a44272a,a44273a,a44277a,a44278a,a44281a,a44284a,a44285a,a44286a,a44290a,a44291a,a44294a,a44297a,a44298a,a44299a,a44303a,a44304a,a44307a,a44310a,a44311a,a44312a,a44316a,a44317a,a44320a,a44323a,a44324a,a44325a,a44329a,a44330a,a44333a,a44336a,a44337a,a44338a,a44342a,a44343a,a44346a,a44349a,a44350a,a44351a,a44355a,a44356a,a44359a,a44362a,a44363a,a44364a,a44368a,a44369a,a44372a,a44375a,a44376a,a44377a,a44381a,a44382a,a44385a,a44388a,a44389a,a44390a,a44394a,a44395a,a44398a,a44401a,a44402a,a44403a,a44407a,a44408a,a44411a,a44414a,a44415a,a44416a,a44420a,a44421a,a44424a,a44427a,a44428a,a44429a,a44433a,a44434a,a44437a,a44440a,a44441a,a44442a,a44446a,a44447a,a44450a,a44453a,a44454a,a44455a,a44459a,a44460a,a44463a,a44466a,a44467a,a44468a,a44472a,a44473a,a44476a,a44479a,a44480a,a44481a,a44485a,a44486a,a44489a,a44492a,a44493a,a44494a,a44498a,a44499a,a44502a,a44505a,a44506a,a44507a,a44511a,a44512a,a44515a,a44518a,a44519a,a44520a,a44524a,a44525a,a44528a,a44531a,a44532a,a44533a,a44537a,a44538a,a44541a,a44544a,a44545a,a44546a,a44550a,a44551a,a44554a,a44557a,a44558a,a44559a,a44563a,a44564a,a44567a,a44570a,a44571a,a44572a,a44576a,a44577a,a44580a,a44583a,a44584a,a44585a,a44589a,a44590a,a44593a,a44596a,a44597a,a44598a,a44602a,a44603a,a44606a,a44609a,a44610a,a44611a,a44615a,a44616a,a44619a,a44622a,a44623a,a44624a,a44628a,a44629a,a44632a,a44635a,a44636a,a44637a,a44641a,a44642a,a44645a,a44648a,a44649a,a44650a,a44654a,a44655a,a44658a,a44661a,a44662a,a44663a,a44667a,a44668a,a44671a,a44674a,a44675a,a44676a,a44680a,a44681a,a44684a,a44687a,a44688a,a44689a,a44693a,a44694a,a44697a,a44700a,a44701a,a44702a,a44706a,a44707a,a44710a,a44713a,a44714a,a44715a,a44719a,a44720a,a44723a,a44726a,a44727a,a44728a,a44732a,a44733a,a44736a,a44739a,a44740a,a44741a,a44745a,a44746a,a44749a,a44752a,a44753a,a44754a,a44758a,a44759a,a44762a,a44765a,a44766a,a44767a,a44771a,a44772a,a44775a,a44778a,a44779a,a44780a,a44784a,a44785a,a44788a,a44791a,a44792a,a44793a,a44797a,a44798a,a44801a,a44804a,a44805a,a44806a,a44810a,a44811a,a44814a,a44817a,a44818a,a44819a,a44823a,a44824a,a44827a,a44830a,a44831a,a44832a,a44836a,a44837a,a44840a,a44843a,a44844a,a44845a,a44849a,a44850a,a44853a,a44856a,a44857a,a44858a,a44862a,a44863a,a44866a,a44869a,a44870a,a44871a,a44875a,a44876a,a44879a,a44882a,a44883a,a44884a,a44888a,a44889a,a44892a,a44895a,a44896a,a44897a,a44901a,a44902a,a44905a,a44908a,a44909a,a44910a,a44914a,a44915a,a44918a,a44921a,a44922a,a44923a,a44927a,a44928a,a44931a,a44934a,a44935a,a44936a,a44940a,a44941a,a44944a,a44947a,a44948a,a44949a,a44953a,a44954a,a44957a,a44960a,a44961a,a44962a,a44966a,a44967a,a44970a,a44973a,a44974a,a44975a,a44979a,a44980a,a44983a,a44986a,a44987a,a44988a,a44992a,a44993a,a44996a,a44999a,a45000a,a45001a,a45005a,a45006a,a45009a,a45012a,a45013a,a45014a,a45018a,a45019a,a45022a,a45025a,a45026a,a45027a,a45031a,a45032a,a45035a,a45038a,a45039a,a45040a,a45044a,a45045a,a45048a,a45051a,a45052a,a45053a,a45057a,a45058a,a45061a,a45064a,a45065a,a45066a,a45070a,a45071a,a45074a,a45077a,a45078a,a45079a,a45083a,a45084a,a45087a,a45090a,a45091a,a45092a,a45096a,a45097a,a45100a,a45103a,a45104a,a45105a,a45109a,a45110a,a45113a,a45116a,a45117a,a45118a,a45122a,a45123a,a45126a,a45129a,a45130a,a45131a,a45135a,a45136a,a45139a,a45142a,a45143a,a45144a,a45148a,a45149a,a45152a,a45155a,a45156a,a45157a,a45161a,a45162a,a45165a,a45168a,a45169a,a45170a,a45174a,a45175a,a45178a,a45181a,a45182a,a45183a,a45187a,a45188a,a45191a,a45194a,a45195a,a45196a,a45200a,a45201a,a45204a,a45207a,a45208a,a45209a,a45213a,a45214a,a45217a,a45220a,a45221a,a45222a,a45226a,a45227a,a45230a,a45233a,a45234a,a45235a,a45239a,a45240a,a45243a,a45246a,a45247a,a45248a,a45252a,a45253a,a45256a,a45259a,a45260a,a45261a,a45265a,a45266a,a45269a,a45272a,a45273a,a45274a,a45278a,a45279a,a45282a,a45285a,a45286a,a45287a,a45291a,a45292a,a45295a,a45298a,a45299a,a45300a,a45304a,a45305a,a45308a,a45311a,a45312a,a45313a,a45317a,a45318a,a45321a,a45324a,a45325a,a45326a,a45330a,a45331a,a45334a,a45337a,a45338a,a45339a,a45343a,a45344a,a45347a,a45350a,a45351a,a45352a,a45356a,a45357a,a45360a,a45363a,a45364a,a45365a,a45369a,a45370a,a45373a,a45376a,a45377a,a45378a,a45382a,a45383a,a45386a,a45389a,a45390a,a45391a,a45395a,a45396a,a45399a,a45402a,a45403a,a45404a,a45408a,a45409a,a45412a,a45415a,a45416a,a45417a,a45421a,a45422a,a45425a,a45428a,a45429a,a45430a,a45434a,a45435a,a45438a,a45441a,a45442a,a45443a,a45447a,a45448a,a45451a,a45454a,a45455a,a45456a,a45460a,a45461a,a45464a,a45467a,a45468a,a45469a,a45473a,a45474a,a45477a,a45480a,a45481a,a45482a,a45486a,a45487a,a45490a,a45493a,a45494a,a45495a,a45499a,a45500a,a45503a,a45506a,a45507a,a45508a,a45512a,a45513a,a45516a,a45519a,a45520a,a45521a,a45525a,a45526a,a45529a,a45532a,a45533a,a45534a,a45538a,a45539a,a45542a,a45545a,a45546a,a45547a,a45551a,a45552a,a45555a,a45558a,a45559a,a45560a,a45564a,a45565a,a45568a,a45571a,a45572a,a45573a,a45577a,a45578a,a45581a,a45584a,a45585a,a45586a,a45590a,a45591a,a45594a,a45597a,a45598a,a45599a,a45603a,a45604a,a45607a,a45610a,a45611a,a45612a,a45616a,a45617a,a45620a,a45623a,a45624a,a45625a,a45629a,a45630a,a45633a,a45636a,a45637a,a45638a,a45642a,a45643a,a45646a,a45649a,a45650a,a45651a,a45655a,a45656a,a45659a,a45662a,a45663a,a45664a,a45668a,a45669a,a45672a,a45675a,a45676a,a45677a,a45681a,a45682a,a45685a,a45688a,a45689a,a45690a,a45694a,a45695a,a45698a,a45701a,a45702a,a45703a,a45707a,a45708a,a45711a,a45714a,a45715a,a45716a,a45720a,a45721a,a45724a,a45727a,a45728a,a45729a,a45733a,a45734a,a45737a,a45740a,a45741a,a45742a,a45746a,a45747a,a45750a,a45753a,a45754a,a45755a,a45759a,a45760a,a45763a,a45766a,a45767a,a45768a,a45772a,a45773a,a45776a,a45779a,a45780a,a45781a,a45785a,a45786a,a45789a,a45792a,a45793a,a45794a,a45798a,a45799a,a45802a,a45805a,a45806a,a45807a,a45811a,a45812a,a45815a,a45818a,a45819a,a45820a,a45824a,a45825a,a45828a,a45831a,a45832a,a45833a,a45837a,a45838a,a45841a,a45844a,a45845a,a45846a,a45850a,a45851a,a45854a,a45857a,a45858a,a45859a,a45863a,a45864a,a45867a,a45870a,a45871a,a45872a,a45876a,a45877a,a45880a,a45883a,a45884a,a45885a,a45889a,a45890a,a45893a,a45896a,a45897a,a45898a,a45902a,a45903a,a45906a,a45909a,a45910a,a45911a,a45915a,a45916a,a45919a,a45922a,a45923a,a45924a,a45928a,a45929a,a45932a,a45935a,a45936a,a45937a,a45941a,a45942a,a45945a,a45948a,a45949a,a45950a,a45954a,a45955a,a45958a,a45961a,a45962a,a45963a,a45967a,a45968a,a45971a,a45974a,a45975a,a45976a,a45980a,a45981a,a45984a,a45987a,a45988a,a45989a,a45993a,a45994a,a45997a,a46000a,a46001a,a46002a,a46006a,a46007a,a46010a,a46013a,a46014a,a46015a,a46019a,a46020a,a46023a,a46026a,a46027a,a46028a,a46032a,a46033a,a46036a,a46039a,a46040a,a46041a,a46045a,a46046a,a46049a,a46052a,a46053a,a46054a,a46058a,a46059a,a46062a,a46065a,a46066a,a46067a,a46071a,a46072a,a46075a,a46078a,a46079a,a46080a,a46084a,a46085a,a46088a,a46091a,a46092a,a46093a,a46097a,a46098a,a46101a,a46104a,a46105a,a46106a,a46110a,a46111a,a46114a,a46117a,a46118a,a46119a,a46123a,a46124a,a46127a,a46130a,a46131a,a46132a,a46136a,a46137a,a46140a,a46143a,a46144a,a46145a,a46149a,a46150a,a46153a,a46156a,a46157a,a46158a,a46162a,a46163a,a46166a,a46169a,a46170a,a46171a,a46175a,a46176a,a46179a,a46182a,a46183a,a46184a,a46188a,a46189a,a46192a,a46195a,a46196a,a46197a,a46201a,a46202a,a46205a,a46208a,a46209a,a46210a,a46214a,a46215a,a46218a,a46221a,a46222a,a46223a,a46227a,a46228a,a46231a,a46234a,a46235a,a46236a,a46240a,a46241a,a46244a,a46247a,a46248a,a46249a,a46253a,a46254a,a46257a,a46260a,a46261a,a46262a,a46266a,a46267a,a46270a,a46273a,a46274a,a46275a,a46279a,a46280a,a46283a,a46286a,a46287a,a46288a,a46292a,a46293a,a46296a,a46299a,a46300a,a46301a,a46305a,a46306a,a46309a,a46312a,a46313a,a46314a,a46318a,a46319a,a46322a,a46325a,a46326a,a46327a,a46331a,a46332a,a46335a,a46338a,a46339a,a46340a,a46344a,a46345a,a46348a,a46351a,a46352a,a46353a,a46357a,a46358a,a46361a,a46364a,a46365a,a46366a,a46370a,a46371a,a46374a,a46377a,a46378a,a46379a,a46383a,a46384a,a46387a,a46390a,a46391a,a46392a,a46396a,a46397a,a46400a,a46403a,a46404a,a46405a,a46409a,a46410a,a46413a,a46416a,a46417a,a46418a,a46422a,a46423a,a46426a,a46429a,a46430a,a46431a,a46435a,a46436a,a46439a,a46442a,a46443a,a46444a,a46448a,a46449a,a46452a,a46455a,a46456a,a46457a,a46461a,a46462a,a46465a,a46468a,a46469a,a46470a,a46474a,a46475a,a46478a,a46481a,a46482a,a46483a,a46487a,a46488a,a46491a,a46494a,a46495a,a46496a,a46500a,a46501a,a46504a,a46507a,a46508a,a46509a,a46513a,a46514a,a46517a,a46520a,a46521a,a46522a,a46526a,a46527a,a46530a,a46533a,a46534a,a46535a,a46539a,a46540a,a46543a,a46546a,a46547a,a46548a,a46552a,a46553a,a46556a,a46559a,a46560a,a46561a,a46565a,a46566a,a46569a,a46572a,a46573a,a46574a,a46578a,a46579a,a46582a,a46585a,a46586a,a46587a,a46591a,a46592a,a46595a,a46598a,a46599a,a46600a,a46604a,a46605a,a46608a,a46611a,a46612a,a46613a,a46617a,a46618a,a46621a,a46624a,a46625a,a46626a,a46630a,a46631a,a46634a,a46637a,a46638a,a46639a,a46643a,a46644a,a46647a,a46650a,a46651a,a46652a,a46656a,a46657a,a46660a,a46663a,a46664a,a46665a,a46669a,a46670a,a46673a,a46676a,a46677a,a46678a,a46682a,a46683a,a46686a,a46689a,a46690a,a46691a,a46695a,a46696a,a46699a,a46702a,a46703a,a46704a,a46708a,a46709a,a46712a,a46715a,a46716a,a46717a,a46721a,a46722a,a46725a,a46728a,a46729a,a46730a,a46734a,a46735a,a46738a,a46741a,a46742a,a46743a,a46747a,a46748a,a46751a,a46754a,a46755a,a46756a,a46760a,a46761a,a46764a,a46767a,a46768a,a46769a,a46773a,a46774a,a46777a,a46780a,a46781a,a46782a,a46786a,a46787a,a46790a,a46793a,a46794a,a46795a,a46799a,a46800a,a46803a,a46806a,a46807a,a46808a,a46812a,a46813a,a46816a,a46819a,a46820a,a46821a,a46825a,a46826a,a46829a,a46832a,a46833a,a46834a,a46838a,a46839a,a46842a,a46845a,a46846a,a46847a,a46851a,a46852a,a46855a,a46858a,a46859a,a46860a,a46864a,a46865a,a46868a,a46871a,a46872a,a46873a,a46877a,a46878a,a46881a,a46884a,a46885a,a46886a,a46890a,a46891a,a46894a,a46897a,a46898a,a46899a,a46903a,a46904a,a46907a,a46910a,a46911a,a46912a,a46916a,a46917a,a46920a,a46923a,a46924a,a46925a,a46929a,a46930a,a46933a,a46936a,a46937a,a46938a,a46942a,a46943a,a46946a,a46949a,a46950a,a46951a,a46955a,a46956a,a46959a,a46962a,a46963a,a46964a,a46968a,a46969a,a46972a,a46975a,a46976a,a46977a,a46981a,a46982a,a46985a,a46988a,a46989a,a46990a,a46994a,a46995a,a46998a,a47001a,a47002a,a47003a,a47007a,a47008a,a47011a,a47014a,a47015a,a47016a,a47020a,a47021a,a47024a,a47027a,a47028a,a47029a,a47033a,a47034a,a47037a,a47040a,a47041a,a47042a,a47046a,a47047a,a47050a,a47053a,a47054a,a47055a,a47059a,a47060a,a47063a,a47066a,a47067a,a47068a,a47072a,a47073a,a47076a,a47079a,a47080a,a47081a,a47085a,a47086a,a47089a,a47092a,a47093a,a47094a,a47098a,a47099a,a47102a,a47105a,a47106a,a47107a,a47111a,a47112a,a47115a,a47118a,a47119a,a47120a,a47124a,a47125a,a47128a,a47131a,a47132a,a47133a,a47137a,a47138a,a47141a,a47144a,a47145a,a47146a,a47150a,a47151a,a47154a,a47157a,a47158a,a47159a,a47163a,a47164a,a47167a,a47170a,a47171a,a47172a,a47176a,a47177a,a47180a,a47183a,a47184a,a47185a,a47189a,a47190a,a47193a,a47196a,a47197a,a47198a,a47202a,a47203a,a47206a,a47209a,a47210a,a47211a,a47215a,a47216a,a47219a,a47222a,a47223a,a47224a,a47228a,a47229a,a47232a,a47235a,a47236a,a47237a,a47241a,a47242a,a47245a,a47248a,a47249a,a47250a,a47254a,a47255a,a47258a,a47261a,a47262a,a47263a,a47267a,a47268a,a47271a,a47274a,a47275a,a47276a,a47280a,a47281a,a47284a,a47287a,a47288a,a47289a,a47293a,a47294a,a47297a,a47300a,a47301a,a47302a,a47306a,a47307a,a47310a,a47313a,a47314a,a47315a,a47319a,a47320a,a47323a,a47326a,a47327a,a47328a,a47332a,a47333a,a47336a,a47339a,a47340a,a47341a,a47345a,a47346a,a47349a,a47352a,a47353a,a47354a,a47358a,a47359a,a47362a,a47365a,a47366a,a47367a,a47371a,a47372a,a47375a,a47378a,a47379a,a47380a,a47384a,a47385a,a47388a,a47391a,a47392a,a47393a,a47397a,a47398a,a47401a,a47404a,a47405a,a47406a,a47410a,a47411a,a47414a,a47417a,a47418a,a47419a,a47423a,a47424a,a47427a,a47430a,a47431a,a47432a,a47436a,a47437a,a47440a,a47443a,a47444a,a47445a,a47449a,a47450a,a47453a,a47456a,a47457a,a47458a,a47462a,a47463a,a47466a,a47469a,a47470a,a47471a,a47475a,a47476a,a47479a,a47482a,a47483a,a47484a,a47488a,a47489a,a47492a,a47495a,a47496a,a47497a,a47501a,a47502a,a47505a,a47508a,a47509a,a47510a,a47514a,a47515a,a47518a,a47521a,a47522a,a47523a,a47527a,a47528a,a47531a,a47534a,a47535a,a47536a,a47540a,a47541a,a47544a,a47547a,a47548a,a47549a,a47553a,a47554a,a47557a,a47560a,a47561a,a47562a,a47566a,a47567a,a47570a,a47573a,a47574a,a47575a,a47579a,a47580a,a47583a,a47586a,a47587a,a47588a,a47592a,a47593a,a47596a,a47599a,a47600a,a47601a,a47605a,a47606a,a47609a,a47612a,a47613a,a47614a,a47618a,a47619a,a47622a,a47625a,a47626a,a47627a,a47631a,a47632a,a47635a,a47638a,a47639a,a47640a,a47644a,a47645a,a47648a,a47651a,a47652a,a47653a,a47657a,a47658a,a47661a,a47664a,a47665a,a47666a,a47670a,a47671a,a47674a,a47677a,a47678a,a47679a,a47683a,a47684a,a47687a,a47690a,a47691a,a47692a,a47696a,a47697a,a47700a,a47703a,a47704a,a47705a,a47709a,a47710a,a47713a,a47716a,a47717a,a47718a,a47722a,a47723a,a47726a,a47729a,a47730a,a47731a,a47735a,a47736a,a47739a,a47742a,a47743a,a47744a,a47748a,a47749a,a47752a,a47755a,a47756a,a47757a,a47761a,a47762a,a47765a,a47768a,a47769a,a47770a,a47774a,a47775a,a47778a,a47781a,a47782a,a47783a,a47787a,a47788a,a47791a,a47794a,a47795a,a47796a,a47800a,a47801a,a47804a,a47807a,a47808a,a47809a,a47813a,a47814a,a47817a,a47820a,a47821a,a47822a,a47826a,a47827a,a47830a,a47833a,a47834a,a47835a,a47839a,a47840a,a47843a,a47846a,a47847a,a47848a,a47852a,a47853a,a47856a,a47859a,a47860a,a47861a,a47865a,a47866a,a47869a,a47872a,a47873a,a47874a,a47878a,a47879a,a47882a,a47885a,a47886a,a47887a,a47891a,a47892a,a47895a,a47898a,a47899a,a47900a,a47904a,a47905a,a47908a,a47911a,a47912a,a47913a,a47917a,a47918a,a47921a,a47924a,a47925a,a47926a,a47930a,a47931a,a47934a,a47937a,a47938a,a47939a,a47943a,a47944a,a47947a,a47950a,a47951a,a47952a,a47956a,a47957a,a47960a,a47963a,a47964a,a47965a,a47969a,a47970a,a47973a,a47976a,a47977a,a47978a,a47982a,a47983a,a47986a,a47989a,a47990a,a47991a,a47995a,a47996a,a47999a,a48002a,a48003a,a48004a,a48008a,a48009a,a48012a,a48015a,a48016a,a48017a,a48021a,a48022a,a48025a,a48028a,a48029a,a48030a,a48034a,a48035a,a48038a,a48041a,a48042a,a48043a,a48047a,a48048a,a48051a,a48054a,a48055a,a48056a,a48060a,a48061a,a48064a,a48067a,a48068a,a48069a,a48073a,a48074a,a48077a,a48080a,a48081a,a48082a,a48086a,a48087a,a48090a,a48093a,a48094a,a48095a,a48099a,a48100a,a48103a,a48106a,a48107a,a48108a,a48112a,a48113a,a48116a,a48119a,a48120a,a48121a,a48125a,a48126a,a48129a,a48132a,a48133a,a48134a,a48138a,a48139a,a48142a,a48145a,a48146a,a48147a,a48151a,a48152a,a48155a,a48158a,a48159a,a48160a,a48164a,a48165a,a48168a,a48171a,a48172a,a48173a,a48177a,a48178a,a48181a,a48184a,a48185a,a48186a,a48190a,a48191a,a48194a,a48197a,a48198a,a48199a,a48203a,a48204a,a48207a,a48210a,a48211a,a48212a,a48216a,a48217a,a48220a,a48223a,a48224a,a48225a,a48229a,a48230a,a48233a,a48236a,a48237a,a48238a,a48242a,a48243a,a48246a,a48249a,a48250a,a48251a,a48255a,a48256a,a48259a,a48262a,a48263a,a48264a,a48268a,a48269a,a48272a,a48275a,a48276a,a48277a,a48281a,a48282a,a48285a,a48288a,a48289a,a48290a,a48294a,a48295a,a48298a,a48301a,a48302a,a48303a,a48307a,a48308a,a48311a,a48314a,a48315a,a48316a,a48320a,a48321a,a48324a,a48327a,a48328a,a48329a,a48333a,a48334a,a48337a,a48340a,a48341a,a48342a,a48346a,a48347a,a48350a,a48353a,a48354a,a48355a,a48359a,a48360a,a48363a,a48366a,a48367a,a48368a,a48372a,a48373a,a48376a,a48379a,a48380a,a48381a,a48385a,a48386a,a48389a,a48392a,a48393a,a48394a,a48398a,a48399a,a48402a,a48405a,a48406a,a48407a,a48411a,a48412a,a48415a,a48418a,a48419a,a48420a,a48424a,a48425a,a48428a,a48431a,a48432a,a48433a,a48437a,a48438a,a48441a,a48444a,a48445a,a48446a,a48450a,a48451a,a48454a,a48457a,a48458a,a48459a,a48463a,a48464a,a48467a,a48470a,a48471a,a48472a,a48476a,a48477a,a48480a,a48483a,a48484a,a48485a,a48489a,a48490a,a48493a,a48496a,a48497a,a48498a,a48502a,a48503a,a48506a,a48509a,a48510a,a48511a,a48515a,a48516a,a48519a,a48522a,a48523a,a48524a,a48528a,a48529a,a48532a,a48535a,a48536a,a48537a,a48541a,a48542a,a48545a,a48548a,a48549a,a48550a,a48554a,a48555a,a48558a,a48561a,a48562a,a48563a,a48567a,a48568a,a48571a,a48574a,a48575a,a48576a,a48580a,a48581a,a48584a,a48587a,a48588a,a48589a,a48593a,a48594a,a48597a,a48600a,a48601a,a48602a,a48606a,a48607a,a48610a,a48613a,a48614a,a48615a,a48619a,a48620a,a48623a,a48626a,a48627a,a48628a,a48632a,a48633a,a48636a,a48639a,a48640a,a48641a,a48645a,a48646a,a48649a,a48652a,a48653a,a48654a,a48658a,a48659a,a48662a,a48665a,a48666a,a48667a,a48671a,a48672a,a48675a,a48678a,a48679a,a48680a,a48684a,a48685a,a48688a,a48691a,a48692a,a48693a,a48697a,a48698a,a48701a,a48704a,a48705a,a48706a,a48710a,a48711a,a48714a,a48717a,a48718a,a48719a,a48723a,a48724a,a48727a,a48730a,a48731a,a48732a,a48736a,a48737a,a48740a,a48743a,a48744a,a48745a,a48749a,a48750a,a48753a,a48756a,a48757a,a48758a,a48762a,a48763a,a48766a,a48769a,a48770a,a48771a,a48775a,a48776a,a48779a,a48782a,a48783a,a48784a,a48788a,a48789a,a48792a,a48795a,a48796a,a48797a,a48801a,a48802a,a48805a,a48808a,a48809a,a48810a,a48814a,a48815a,a48818a,a48821a,a48822a,a48823a,a48827a,a48828a,a48831a,a48834a,a48835a,a48836a,a48840a,a48841a,a48844a,a48847a,a48848a,a48849a,a48853a,a48854a,a48857a,a48860a,a48861a,a48862a,a48866a,a48867a,a48870a,a48873a,a48874a,a48875a,a48879a,a48880a,a48883a,a48886a,a48887a,a48888a,a48892a,a48893a,a48896a,a48899a,a48900a,a48901a,a48905a,a48906a,a48909a,a48912a,a48913a,a48914a,a48918a,a48919a,a48922a,a48925a,a48926a,a48927a,a48931a,a48932a,a48935a,a48938a,a48939a,a48940a,a48944a,a48945a,a48948a,a48951a,a48952a,a48953a,a48957a,a48958a,a48961a,a48964a,a48965a,a48966a,a48970a,a48971a,a48974a,a48977a,a48978a,a48979a,a48983a,a48984a,a48987a,a48990a,a48991a,a48992a,a48996a,a48997a,a49000a,a49003a,a49004a,a49005a,a49009a,a49010a,a49013a,a49016a,a49017a,a49018a,a49022a,a49023a,a49026a,a49029a,a49030a,a49031a,a49035a,a49036a,a49039a,a49042a,a49043a,a49044a,a49048a,a49049a,a49052a,a49055a,a49056a,a49057a,a49061a,a49062a,a49065a,a49068a,a49069a,a49070a,a49074a,a49075a,a49078a,a49081a,a49082a,a49083a,a49087a,a49088a,a49091a,a49094a,a49095a,a49096a,a49100a,a49101a,a49104a,a49107a,a49108a,a49109a,a49113a,a49114a,a49117a,a49120a,a49121a,a49122a,a49126a,a49127a,a49130a,a49133a,a49134a,a49135a,a49139a,a49140a,a49143a,a49146a,a49147a,a49148a,a49152a,a49153a,a49156a,a49159a,a49160a,a49161a,a49165a,a49166a,a49169a,a49172a,a49173a,a49174a,a49178a,a49179a,a49182a,a49185a,a49186a,a49187a,a49191a,a49192a,a49195a,a49198a,a49199a,a49200a,a49204a,a49205a,a49208a,a49211a,a49212a,a49213a,a49217a,a49218a,a49221a,a49224a,a49225a,a49226a,a49230a,a49231a,a49234a,a49237a,a49238a,a49239a,a49243a,a49244a,a49247a,a49250a,a49251a,a49252a,a49256a,a49257a,a49260a,a49263a,a49264a,a49265a,a49269a,a49270a,a49273a,a49276a,a49277a,a49278a,a49282a,a49283a,a49286a,a49289a,a49290a,a49291a,a49295a,a49296a,a49299a,a49302a,a49303a,a49304a,a49308a,a49309a,a49312a,a49315a,a49316a,a49317a,a49321a,a49322a,a49325a,a49328a,a49329a,a49330a,a49334a,a49335a,a49338a,a49341a,a49342a,a49343a,a49347a,a49348a,a49351a,a49354a,a49355a,a49356a,a49360a,a49361a,a49364a,a49367a,a49368a,a49369a,a49373a,a49374a,a49377a,a49380a,a49381a,a49382a,a49386a,a49387a,a49390a,a49393a,a49394a,a49395a,a49399a,a49400a,a49403a,a49406a,a49407a,a49408a,a49412a,a49413a,a49416a,a49419a,a49420a,a49421a,a49425a,a49426a,a49429a,a49432a,a49433a,a49434a,a49438a,a49439a,a49442a,a49445a,a49446a,a49447a,a49451a,a49452a,a49455a,a49458a,a49459a,a49460a,a49464a,a49465a,a49468a,a49471a,a49472a,a49473a,a49477a,a49478a,a49481a,a49484a,a49485a,a49486a,a49490a,a49491a,a49494a,a49497a,a49498a,a49499a,a49503a,a49504a,a49507a,a49510a,a49511a,a49512a,a49516a,a49517a,a49520a,a49523a,a49524a,a49525a,a49529a,a49530a,a49533a,a49536a,a49537a,a49538a,a49542a,a49543a,a49546a,a49549a,a49550a,a49551a,a49555a,a49556a,a49559a,a49562a,a49563a,a49564a,a49568a,a49569a,a49572a,a49575a,a49576a,a49577a,a49581a,a49582a,a49585a,a49588a,a49589a,a49590a,a49594a,a49595a,a49598a,a49601a,a49602a,a49603a,a49607a,a49608a,a49611a,a49614a,a49615a,a49616a,a49620a,a49621a,a49624a,a49627a,a49628a,a49629a,a49633a,a49634a,a49637a,a49640a,a49641a,a49642a,a49646a,a49647a,a49650a,a49653a,a49654a,a49655a,a49659a,a49660a,a49663a,a49666a,a49667a,a49668a,a49672a,a49673a,a49676a,a49679a,a49680a,a49681a,a49685a,a49686a,a49689a,a49692a,a49693a,a49694a,a49698a,a49699a,a49702a,a49705a,a49706a,a49707a,a49711a,a49712a,a49715a,a49718a,a49719a,a49720a,a49724a,a49725a,a49728a,a49731a,a49732a,a49733a,a49737a,a49738a,a49741a,a49744a,a49745a,a49746a,a49750a,a49751a,a49754a,a49757a,a49758a,a49759a,a49763a,a49764a,a49767a,a49770a,a49771a,a49772a,a49776a,a49777a,a49780a,a49783a,a49784a,a49785a,a49789a,a49790a,a49793a,a49796a,a49797a,a49798a,a49802a,a49803a,a49806a,a49809a,a49810a,a49811a,a49815a,a49816a,a49819a,a49822a,a49823a,a49824a,a49828a,a49829a,a49832a,a49835a,a49836a,a49837a,a49841a,a49842a,a49845a,a49848a,a49849a,a49850a,a49854a,a49855a,a49858a,a49861a,a49862a,a49863a,a49867a,a49868a,a49871a,a49874a,a49875a,a49876a,a49880a,a49881a,a49884a,a49887a,a49888a,a49889a,a49893a,a49894a,a49897a,a49900a,a49901a,a49902a,a49906a,a49907a,a49910a,a49913a,a49914a,a49915a,a49919a,a49920a,a49923a,a49926a,a49927a,a49928a,a49932a,a49933a,a49936a,a49939a,a49940a,a49941a,a49945a,a49946a,a49949a,a49952a,a49953a,a49954a,a49958a,a49959a,a49962a,a49965a,a49966a,a49967a,a49971a,a49972a,a49975a,a49978a,a49979a,a49980a,a49984a,a49985a,a49988a,a49991a,a49992a,a49993a,a49997a,a49998a,a50001a,a50004a,a50005a,a50006a,a50010a,a50011a,a50014a,a50017a,a50018a,a50019a,a50023a,a50024a,a50027a,a50030a,a50031a,a50032a,a50036a,a50037a,a50040a,a50043a,a50044a,a50045a,a50049a,a50050a,a50053a,a50056a,a50057a,a50058a,a50062a,a50063a,a50066a,a50069a,a50070a,a50071a,a50075a,a50076a,a50079a,a50082a,a50083a,a50084a,a50088a,a50089a,a50092a,a50095a,a50096a,a50097a,a50101a,a50102a,a50105a,a50108a,a50109a,a50110a,a50114a,a50115a,a50118a,a50121a,a50122a,a50123a,a50127a,a50128a,a50131a,a50134a,a50135a,a50136a,a50140a,a50141a,a50144a,a50147a,a50148a,a50149a,a50153a,a50154a,a50157a,a50160a,a50161a,a50162a,a50166a,a50167a,a50170a,a50173a,a50174a,a50175a,a50179a,a50180a,a50183a,a50186a,a50187a,a50188a,a50192a,a50193a,a50196a,a50199a,a50200a,a50201a,a50205a,a50206a,a50209a,a50212a,a50213a,a50214a,a50218a,a50219a,a50222a,a50225a,a50226a,a50227a,a50231a,a50232a,a50235a,a50238a,a50239a,a50240a,a50244a,a50245a,a50248a,a50251a,a50252a,a50253a,a50257a,a50258a,a50261a,a50264a,a50265a,a50266a,a50270a,a50271a,a50274a,a50277a,a50278a,a50279a,a50283a,a50284a,a50287a,a50290a,a50291a,a50292a,a50296a,a50297a,a50300a,a50303a,a50304a,a50305a,a50309a,a50310a,a50313a,a50316a,a50317a,a50318a,a50322a,a50323a,a50326a,a50329a,a50330a,a50331a,a50335a,a50336a,a50339a,a50342a,a50343a,a50344a,a50348a,a50349a,a50352a,a50355a,a50356a,a50357a,a50361a,a50362a,a50365a,a50368a,a50369a,a50370a,a50374a,a50375a,a50378a,a50381a,a50382a,a50383a,a50387a,a50388a,a50391a,a50394a,a50395a,a50396a,a50400a,a50401a,a50404a,a50407a,a50408a,a50409a,a50413a,a50414a,a50417a,a50420a,a50421a,a50422a,a50426a,a50427a,a50430a,a50433a,a50434a,a50435a,a50439a,a50440a,a50443a,a50446a,a50447a,a50448a,a50452a,a50453a,a50456a,a50459a,a50460a,a50461a,a50465a,a50466a,a50469a,a50472a,a50473a,a50474a,a50478a,a50479a,a50482a,a50485a,a50486a,a50487a,a50491a,a50492a,a50495a,a50498a,a50499a,a50500a,a50504a,a50505a,a50508a,a50511a,a50512a,a50513a,a50517a,a50518a,a50521a,a50524a,a50525a,a50526a,a50530a,a50531a,a50534a,a50537a,a50538a,a50539a,a50543a,a50544a,a50547a,a50550a,a50551a,a50552a,a50556a,a50557a,a50560a,a50563a,a50564a,a50565a,a50569a,a50570a,a50573a,a50576a,a50577a,a50578a,a50582a,a50583a,a50586a,a50589a,a50590a,a50591a,a50595a,a50596a,a50599a,a50602a,a50603a,a50604a,a50608a,a50609a,a50612a,a50615a,a50616a,a50617a,a50621a,a50622a,a50625a,a50628a,a50629a,a50630a,a50634a,a50635a,a50638a,a50641a,a50642a,a50643a,a50647a,a50648a,a50651a,a50654a,a50655a,a50656a,a50660a,a50661a,a50664a,a50667a,a50668a,a50669a,a50673a,a50674a,a50677a,a50680a,a50681a,a50682a,a50686a,a50687a,a50690a,a50693a,a50694a,a50695a,a50699a,a50700a,a50703a,a50706a,a50707a,a50708a,a50712a,a50713a,a50716a,a50719a,a50720a,a50721a,a50725a,a50726a,a50729a,a50732a,a50733a,a50734a,a50738a,a50739a,a50742a,a50745a,a50746a,a50747a,a50751a,a50752a,a50755a,a50758a,a50759a,a50760a,a50764a,a50765a,a50768a,a50771a,a50772a,a50773a,a50777a,a50778a,a50781a,a50784a,a50785a,a50786a,a50790a,a50791a,a50794a,a50797a,a50798a,a50799a,a50803a,a50804a,a50807a,a50810a,a50811a,a50812a,a50816a,a50817a,a50820a,a50823a,a50824a,a50825a,a50829a,a50830a,a50833a,a50836a,a50837a,a50838a,a50842a,a50843a,a50846a,a50849a,a50850a,a50851a,a50855a,a50856a,a50859a,a50862a,a50863a,a50864a,a50868a,a50869a,a50872a,a50875a,a50876a,a50877a,a50881a,a50882a,a50885a,a50888a,a50889a,a50890a,a50894a,a50895a,a50898a,a50901a,a50902a,a50903a,a50907a,a50908a,a50911a,a50914a,a50915a,a50916a,a50920a,a50921a,a50924a,a50927a,a50928a,a50929a,a50933a,a50934a,a50937a,a50940a,a50941a,a50942a,a50946a,a50947a,a50950a,a50953a,a50954a,a50955a,a50959a,a50960a,a50963a,a50966a,a50967a,a50968a,a50972a,a50973a,a50976a,a50979a,a50980a,a50981a,a50985a,a50986a,a50989a,a50992a,a50993a,a50994a,a50998a,a50999a,a51002a,a51005a,a51006a,a51007a,a51011a,a51012a,a51015a,a51018a,a51019a,a51020a,a51024a,a51025a,a51028a,a51031a,a51032a,a51033a,a51037a,a51038a,a51041a,a51044a,a51045a,a51046a,a51050a,a51051a,a51054a,a51057a,a51058a,a51059a,a51063a,a51064a,a51067a,a51070a,a51071a,a51072a,a51076a,a51077a,a51080a,a51083a,a51084a,a51085a,a51089a,a51090a,a51093a,a51096a,a51097a,a51098a,a51102a,a51103a,a51106a,a51109a,a51110a,a51111a,a51115a,a51116a,a51119a,a51122a,a51123a,a51124a,a51128a,a51129a,a51132a,a51135a,a51136a,a51137a,a51141a,a51142a,a51145a,a51148a,a51149a,a51150a,a51154a,a51155a,a51158a,a51161a,a51162a,a51163a,a51167a,a51168a,a51171a,a51174a,a51175a,a51176a,a51180a,a51181a,a51184a,a51187a,a51188a,a51189a,a51193a,a51194a,a51197a,a51200a,a51201a,a51202a,a51206a,a51207a,a51210a,a51213a,a51214a,a51215a,a51219a,a51220a,a51223a,a51226a,a51227a,a51228a,a51232a,a51233a,a51236a,a51239a,a51240a,a51241a,a51245a,a51246a,a51249a,a51252a,a51253a,a51254a,a51258a,a51259a,a51262a,a51265a,a51266a,a51267a,a51271a,a51272a,a51275a,a51278a,a51279a,a51280a,a51284a,a51285a,a51288a,a51291a,a51292a,a51293a,a51297a,a51298a,a51301a,a51304a,a51305a,a51306a,a51310a,a51311a,a51314a,a51317a,a51318a,a51319a,a51323a,a51324a,a51327a,a51330a,a51331a,a51332a,a51336a,a51337a,a51340a,a51343a,a51344a,a51345a,a51349a,a51350a,a51353a,a51356a,a51357a,a51358a,a51362a,a51363a,a51366a,a51369a,a51370a,a51371a,a51375a,a51376a,a51379a,a51382a,a51383a,a51384a,a51388a,a51389a,a51392a,a51395a,a51396a,a51397a,a51401a,a51402a,a51405a,a51408a,a51409a,a51410a,a51414a,a51415a,a51418a,a51421a,a51422a,a51423a,a51427a,a51428a,a51431a,a51434a,a51435a,a51436a,a51440a,a51441a,a51444a,a51447a,a51448a,a51449a,a51453a,a51454a,a51457a,a51460a,a51461a,a51462a,a51466a,a51467a,a51470a,a51473a,a51474a,a51475a,a51479a,a51480a,a51483a,a51486a,a51487a,a51488a,a51492a,a51493a,a51496a,a51499a,a51500a,a51501a,a51505a,a51506a,a51509a,a51512a,a51513a,a51514a,a51518a,a51519a,a51522a,a51525a,a51526a,a51527a,a51531a,a51532a,a51535a,a51538a,a51539a,a51540a,a51544a,a51545a,a51548a,a51551a,a51552a,a51553a,a51557a,a51558a,a51561a,a51564a,a51565a,a51566a,a51570a,a51571a,a51574a,a51577a,a51578a,a51579a,a51583a,a51584a,a51587a,a51590a,a51591a,a51592a,a51596a,a51597a,a51600a,a51603a,a51604a,a51605a,a51609a,a51610a,a51613a,a51616a,a51617a,a51618a,a51622a,a51623a,a51626a,a51629a,a51630a,a51631a,a51635a,a51636a,a51639a,a51642a,a51643a,a51644a,a51648a,a51649a,a51652a,a51655a,a51656a,a51657a,a51661a,a51662a,a51665a,a51668a,a51669a,a51670a,a51674a,a51675a,a51678a,a51681a,a51682a,a51683a,a51687a,a51688a,a51691a,a51694a,a51695a,a51696a,a51700a,a51701a,a51704a,a51707a,a51708a,a51709a,a51713a,a51714a,a51717a,a51720a,a51721a,a51722a,a51726a,a51727a,a51730a,a51733a,a51734a,a51735a,a51739a,a51740a,a51743a,a51746a,a51747a,a51748a,a51752a,a51753a,a51756a,a51759a,a51760a,a51761a,a51765a,a51766a,a51769a,a51772a,a51773a,a51774a,a51778a,a51779a,a51782a,a51785a,a51786a,a51787a,a51791a,a51792a,a51795a,a51798a,a51799a,a51800a,a51804a,a51805a,a51808a,a51811a,a51812a,a51813a,a51817a,a51818a,a51821a,a51824a,a51825a,a51826a,a51830a,a51831a,a51834a,a51837a,a51838a,a51839a,a51843a,a51844a,a51847a,a51850a,a51851a,a51852a,a51856a,a51857a,a51860a,a51863a,a51864a,a51865a,a51869a,a51870a,a51873a,a51876a,a51877a,a51878a,a51882a,a51883a,a51886a,a51889a,a51890a,a51891a,a51895a,a51896a,a51899a,a51902a,a51903a,a51904a,a51908a,a51909a,a51912a,a51915a,a51916a,a51917a,a51921a,a51922a,a51925a,a51928a,a51929a,a51930a,a51934a,a51935a,a51938a,a51941a,a51942a,a51943a,a51947a,a51948a,a51951a,a51954a,a51955a,a51956a,a51960a,a51961a,a51964a,a51967a,a51968a,a51969a,a51973a,a51974a,a51977a,a51980a,a51981a,a51982a,a51986a,a51987a,a51990a,a51993a,a51994a,a51995a,a51999a,a52000a,a52003a,a52006a,a52007a,a52008a,a52012a,a52013a,a52016a,a52019a,a52020a,a52021a,a52025a,a52026a,a52029a,a52032a,a52033a,a52034a,a52038a,a52039a,a52042a,a52045a,a52046a,a52047a,a52051a,a52052a,a52055a,a52058a,a52059a,a52060a,a52064a,a52065a,a52068a,a52071a,a52072a,a52073a,a52077a,a52078a,a52081a,a52084a,a52085a,a52086a,a52090a,a52091a,a52094a,a52097a,a52098a,a52099a,a52103a,a52104a,a52107a,a52110a,a52111a,a52112a,a52116a,a52117a,a52120a,a52123a,a52124a,a52125a,a52129a,a52130a,a52133a,a52136a,a52137a,a52138a,a52142a,a52143a,a52146a,a52149a,a52150a,a52151a,a52155a,a52156a,a52159a,a52162a,a52163a,a52164a,a52168a,a52169a,a52172a,a52175a,a52176a,a52177a,a52181a,a52182a,a52185a,a52188a,a52189a,a52190a,a52194a,a52195a,a52198a,a52201a,a52202a,a52203a,a52207a,a52208a,a52211a,a52214a,a52215a,a52216a,a52220a,a52221a,a52224a,a52227a,a52228a,a52229a,a52233a,a52234a,a52237a,a52240a,a52241a,a52242a,a52246a,a52247a,a52250a,a52253a,a52254a,a52255a,a52259a,a52260a,a52263a,a52266a,a52267a,a52268a,a52272a,a52273a,a52276a,a52279a,a52280a,a52281a,a52285a,a52286a,a52289a,a52292a,a52293a,a52294a,a52298a,a52299a,a52302a,a52305a,a52306a,a52307a,a52311a,a52312a,a52315a,a52318a,a52319a,a52320a,a52324a,a52325a,a52328a,a52331a,a52332a,a52333a,a52337a,a52338a,a52341a,a52344a,a52345a,a52346a,a52350a,a52351a,a52354a,a52357a,a52358a,a52359a,a52363a,a52364a,a52367a,a52370a,a52371a,a52372a,a52376a,a52377a,a52380a,a52383a,a52384a,a52385a,a52389a,a52390a,a52393a,a52396a,a52397a,a52398a,a52402a,a52403a,a52406a,a52409a,a52410a,a52411a,a52415a,a52416a,a52419a,a52422a,a52423a,a52424a,a52428a,a52429a,a52432a,a52435a,a52436a,a52437a,a52441a,a52442a,a52445a,a52448a,a52449a,a52450a,a52454a,a52455a,a52458a,a52461a,a52462a,a52463a,a52467a,a52468a,a52471a,a52474a,a52475a,a52476a,a52480a,a52481a,a52484a,a52487a,a52488a,a52489a,a52493a,a52494a,a52497a,a52500a,a52501a,a52502a,a52506a,a52507a,a52510a,a52513a,a52514a,a52515a,a52519a,a52520a,a52523a,a52526a,a52527a,a52528a,a52532a,a52533a,a52536a,a52539a,a52540a,a52541a,a52545a,a52546a,a52549a,a52552a,a52553a,a52554a,a52558a,a52559a,a52562a,a52565a,a52566a,a52567a,a52571a,a52572a,a52575a,a52578a,a52579a,a52580a,a52584a,a52585a,a52588a,a52591a,a52592a,a52593a,a52597a,a52598a,a52601a,a52604a,a52605a,a52606a,a52610a,a52611a,a52614a,a52617a,a52618a,a52619a,a52623a,a52624a,a52627a,a52630a,a52631a,a52632a,a52636a,a52637a,a52640a,a52643a,a52644a,a52645a,a52649a,a52650a,a52653a,a52656a,a52657a,a52658a,a52662a,a52663a,a52666a,a52669a,a52670a,a52671a,a52675a,a52676a,a52679a,a52682a,a52683a,a52684a,a52688a,a52689a,a52692a,a52695a,a52696a,a52697a,a52701a,a52702a,a52705a,a52708a,a52709a,a52710a,a52714a,a52715a,a52718a,a52721a,a52722a,a52723a,a52727a,a52728a,a52731a,a52734a,a52735a,a52736a,a52740a,a52741a,a52744a,a52747a,a52748a,a52749a,a52753a,a52754a,a52757a,a52760a,a52761a,a52762a,a52766a,a52767a,a52770a,a52773a,a52774a,a52775a,a52779a,a52780a,a52783a,a52786a,a52787a,a52788a,a52792a,a52793a,a52796a,a52799a,a52800a,a52801a,a52805a,a52806a,a52809a,a52812a,a52813a,a52814a,a52818a,a52819a,a52822a,a52825a,a52826a,a52827a,a52831a,a52832a,a52835a,a52838a,a52839a,a52840a,a52844a,a52845a,a52848a,a52851a,a52852a,a52853a,a52857a,a52858a,a52861a,a52864a,a52865a,a52866a,a52870a,a52871a,a52874a,a52877a,a52878a,a52879a,a52883a,a52884a,a52887a,a52890a,a52891a,a52892a,a52896a,a52897a,a52900a,a52903a,a52904a,a52905a,a52909a,a52910a,a52913a,a52916a,a52917a,a52918a,a52922a,a52923a,a52926a,a52929a,a52930a,a52931a,a52935a,a52936a,a52939a,a52942a,a52943a,a52944a,a52948a,a52949a,a52952a,a52955a,a52956a,a52957a,a52961a,a52962a,a52965a,a52968a,a52969a,a52970a,a52974a,a52975a,a52978a,a52981a,a52982a,a52983a,a52987a,a52988a,a52991a,a52994a,a52995a,a52996a,a53000a,a53001a,a53004a,a53007a,a53008a,a53009a,a53013a,a53014a,a53017a,a53020a,a53021a,a53022a,a53026a,a53027a,a53030a,a53033a,a53034a,a53035a,a53039a,a53040a,a53043a,a53046a,a53047a,a53048a,a53052a,a53053a,a53056a,a53059a,a53060a,a53061a,a53065a,a53066a,a53069a,a53072a,a53073a,a53074a,a53078a,a53079a,a53082a,a53085a,a53086a,a53087a,a53091a,a53092a,a53095a,a53098a,a53099a,a53100a,a53104a,a53105a,a53108a,a53111a,a53112a,a53113a,a53117a,a53118a,a53121a,a53124a,a53125a,a53126a,a53130a,a53131a,a53134a,a53137a,a53138a,a53139a,a53143a,a53144a,a53147a,a53150a,a53151a,a53152a,a53156a,a53157a,a53160a,a53163a,a53164a,a53165a,a53169a,a53170a,a53173a,a53176a,a53177a,a53178a,a53182a,a53183a,a53186a,a53189a,a53190a,a53191a,a53195a,a53196a,a53199a,a53202a,a53203a,a53204a,a53208a,a53209a,a53212a,a53215a,a53216a,a53217a,a53221a,a53222a,a53225a,a53228a,a53229a,a53230a,a53234a,a53235a,a53238a,a53241a,a53242a,a53243a,a53247a,a53248a,a53251a,a53254a,a53255a,a53256a,a53260a,a53261a,a53264a,a53267a,a53268a,a53269a,a53273a,a53274a,a53277a,a53280a,a53281a,a53282a,a53286a,a53287a,a53290a,a53293a,a53294a,a53295a,a53299a,a53300a,a53303a,a53306a,a53307a,a53308a,a53312a,a53313a,a53316a,a53319a,a53320a,a53321a,a53325a,a53326a,a53329a,a53332a,a53333a,a53334a,a53338a,a53339a,a53342a,a53345a,a53346a,a53347a,a53351a,a53352a,a53355a,a53358a,a53359a,a53360a,a53364a,a53365a,a53368a,a53371a,a53372a,a53373a,a53377a,a53378a,a53381a,a53384a,a53385a,a53386a,a53390a,a53391a,a53394a,a53397a,a53398a,a53399a,a53403a,a53404a,a53407a,a53410a,a53411a,a53412a,a53416a,a53417a,a53420a,a53423a,a53424a,a53425a,a53429a,a53430a,a53433a,a53436a,a53437a,a53438a,a53442a,a53443a,a53446a,a53449a,a53450a,a53451a,a53455a,a53456a,a53459a,a53462a,a53463a,a53464a,a53468a,a53469a,a53472a,a53475a,a53476a,a53477a,a53481a,a53482a,a53485a,a53488a,a53489a,a53490a,a53494a,a53495a,a53498a,a53501a,a53502a,a53503a,a53507a,a53508a,a53511a,a53514a,a53515a,a53516a,a53520a,a53521a,a53524a,a53527a,a53528a,a53529a,a53533a,a53534a,a53537a,a53540a,a53541a,a53542a,a53546a,a53547a,a53550a,a53553a,a53554a,a53555a,a53559a,a53560a,a53563a,a53566a,a53567a,a53568a,a53572a,a53573a,a53576a,a53579a,a53580a,a53581a,a53585a,a53586a,a53589a,a53592a,a53593a,a53594a,a53598a,a53599a,a53602a,a53605a,a53606a,a53607a,a53611a,a53612a,a53615a,a53618a,a53619a,a53620a,a53624a,a53625a,a53628a,a53631a,a53632a,a53633a,a53637a,a53638a,a53641a,a53644a,a53645a,a53646a,a53650a,a53651a,a53654a,a53657a,a53658a,a53659a,a53663a,a53664a,a53667a,a53670a,a53671a,a53672a,a53676a,a53677a,a53680a,a53683a,a53684a,a53685a,a53689a,a53690a,a53693a,a53696a,a53697a,a53698a,a53702a,a53703a,a53706a,a53709a,a53710a,a53711a,a53715a,a53716a,a53719a,a53722a,a53723a,a53724a,a53728a,a53729a,a53732a,a53735a,a53736a,a53737a,a53741a,a53742a,a53745a,a53748a,a53749a,a53750a,a53754a,a53755a,a53758a,a53761a,a53762a,a53763a,a53767a,a53768a,a53771a,a53774a,a53775a,a53776a,a53780a,a53781a,a53784a,a53787a,a53788a,a53789a,a53793a,a53794a,a53797a,a53800a,a53801a,a53802a,a53806a,a53807a,a53810a,a53813a,a53814a,a53815a,a53819a,a53820a,a53823a,a53826a,a53827a,a53828a,a53832a,a53833a,a53836a,a53839a,a53840a,a53841a,a53845a,a53846a,a53849a,a53852a,a53853a,a53854a,a53858a,a53859a,a53862a,a53865a,a53866a,a53867a,a53871a,a53872a,a53875a,a53878a,a53879a,a53880a,a53884a,a53885a,a53888a,a53891a,a53892a,a53893a,a53897a,a53898a,a53901a,a53904a,a53905a,a53906a,a53910a,a53911a,a53914a,a53917a,a53918a,a53919a,a53923a,a53924a,a53927a,a53930a,a53931a,a53932a,a53936a,a53937a,a53940a,a53943a,a53944a,a53945a,a53949a,a53950a,a53953a,a53956a,a53957a,a53958a,a53962a,a53963a,a53966a,a53969a,a53970a,a53971a,a53975a,a53976a,a53979a,a53982a,a53983a,a53984a,a53988a,a53989a,a53992a,a53995a,a53996a,a53997a,a54001a,a54002a,a54005a,a54008a,a54009a,a54010a,a54014a,a54015a,a54018a,a54021a,a54022a,a54023a,a54027a,a54028a,a54031a,a54034a,a54035a,a54036a,a54040a,a54041a,a54044a,a54047a,a54048a,a54049a,a54053a,a54054a,a54057a,a54060a,a54061a,a54062a,a54066a,a54067a,a54070a,a54073a,a54074a,a54075a,a54079a,a54080a,a54083a,a54086a,a54087a,a54088a,a54092a,a54093a,a54096a,a54099a,a54100a,a54101a,a54105a,a54106a,a54109a,a54112a,a54113a,a54114a,a54118a,a54119a,a54122a,a54125a,a54126a,a54127a,a54131a,a54132a,a54135a,a54138a,a54139a,a54140a,a54144a,a54145a,a54148a,a54151a,a54152a,a54153a,a54157a,a54158a,a54161a,a54164a,a54165a,a54166a,a54170a,a54171a,a54174a,a54177a,a54178a,a54179a,a54183a,a54184a,a54187a,a54190a,a54191a,a54192a,a54196a,a54197a,a54200a,a54203a,a54204a,a54205a,a54209a,a54210a,a54213a,a54216a,a54217a,a54218a,a54222a,a54223a,a54226a,a54229a,a54230a,a54231a,a54235a,a54236a,a54239a,a54242a,a54243a,a54244a,a54248a,a54249a,a54252a,a54255a,a54256a,a54257a,a54261a,a54262a,a54265a,a54268a,a54269a,a54270a,a54274a,a54275a,a54278a,a54281a,a54282a,a54283a,a54287a,a54288a,a54291a,a54294a,a54295a,a54296a,a54300a,a54301a,a54304a,a54307a,a54308a,a54309a,a54313a,a54314a,a54317a,a54320a,a54321a,a54322a,a54326a,a54327a,a54330a,a54333a,a54334a,a54335a,a54339a,a54340a,a54343a,a54346a,a54347a,a54348a,a54352a,a54353a,a54356a,a54359a,a54360a,a54361a,a54365a,a54366a,a54369a,a54372a,a54373a,a54374a,a54378a,a54379a,a54382a,a54385a,a54386a,a54387a,a54391a,a54392a,a54395a,a54398a,a54399a,a54400a,a54404a,a54405a,a54408a,a54411a,a54412a,a54413a,a54417a,a54418a,a54421a,a54424a,a54425a,a54426a,a54430a,a54431a,a54434a,a54437a,a54438a,a54439a,a54443a,a54444a,a54447a,a54450a,a54451a,a54452a,a54456a,a54457a,a54460a,a54463a,a54464a,a54465a,a54469a,a54470a,a54473a,a54476a,a54477a,a54478a,a54482a,a54483a,a54486a,a54489a,a54490a,a54491a,a54495a,a54496a,a54499a,a54502a,a54503a,a54504a,a54508a,a54509a,a54512a,a54515a,a54516a,a54517a,a54521a,a54522a,a54525a,a54528a,a54529a,a54530a,a54534a,a54535a,a54538a,a54541a,a54542a,a54543a,a54547a,a54548a,a54551a,a54554a,a54555a,a54556a,a54560a,a54561a,a54564a,a54567a,a54568a,a54569a,a54573a,a54574a,a54577a,a54580a,a54581a,a54582a,a54586a,a54587a,a54590a,a54593a,a54594a,a54595a,a54599a,a54600a,a54603a,a54606a,a54607a,a54608a,a54612a,a54613a,a54616a,a54619a,a54620a,a54621a,a54625a,a54626a,a54629a,a54632a,a54633a,a54634a,a54638a,a54639a,a54642a,a54645a,a54646a,a54647a,a54651a,a54652a,a54655a,a54658a,a54659a,a54660a,a54664a,a54665a,a54668a,a54671a,a54672a,a54673a,a54677a,a54678a,a54681a,a54684a,a54685a,a54686a,a54690a,a54691a,a54694a,a54697a,a54698a,a54699a,a54703a,a54704a,a54707a,a54710a,a54711a,a54712a,a54716a,a54717a,a54720a,a54723a,a54724a,a54725a,a54729a,a54730a,a54733a,a54736a,a54737a,a54738a,a54742a,a54743a,a54746a,a54749a,a54750a,a54751a,a54755a,a54756a,a54759a,a54762a,a54763a,a54764a,a54768a,a54769a,a54772a,a54775a,a54776a,a54777a,a54781a,a54782a,a54785a,a54788a,a54789a,a54790a,a54794a,a54795a,a54798a,a54801a,a54802a,a54803a,a54807a,a54808a,a54811a,a54814a,a54815a,a54816a,a54820a,a54821a,a54824a,a54827a,a54828a,a54829a,a54833a,a54834a,a54837a,a54840a,a54841a,a54842a,a54846a,a54847a,a54850a,a54853a,a54854a,a54855a,a54859a,a54860a,a54863a,a54866a,a54867a,a54868a,a54872a,a54873a,a54876a,a54879a,a54880a,a54881a,a54885a,a54886a,a54889a,a54892a,a54893a,a54894a,a54898a,a54899a,a54902a,a54905a,a54906a,a54907a,a54911a,a54912a,a54915a,a54918a,a54919a,a54920a,a54924a,a54925a,a54928a,a54931a,a54932a,a54933a,a54937a,a54938a,a54941a,a54944a,a54945a,a54946a,a54950a,a54951a,a54954a,a54957a,a54958a,a54959a,a54963a,a54964a,a54967a,a54970a,a54971a,a54972a,a54976a,a54977a,a54980a,a54983a,a54984a,a54985a,a54989a,a54990a,a54993a,a54996a,a54997a,a54998a,a55002a,a55003a,a55006a,a55009a,a55010a,a55011a,a55015a,a55016a,a55019a,a55022a,a55023a,a55024a,a55028a,a55029a,a55032a,a55035a,a55036a,a55037a,a55041a,a55042a,a55045a,a55048a,a55049a,a55050a,a55054a,a55055a,a55058a,a55061a,a55062a,a55063a,a55067a,a55068a,a55071a,a55074a,a55075a,a55076a,a55080a,a55081a,a55084a,a55087a,a55088a,a55089a,a55093a,a55094a,a55097a,a55100a,a55101a,a55102a,a55106a,a55107a,a55110a,a55113a,a55114a,a55115a,a55119a,a55120a,a55123a,a55126a,a55127a,a55128a,a55132a,a55133a,a55136a,a55139a,a55140a,a55141a,a55145a,a55146a,a55149a,a55152a,a55153a,a55154a,a55158a,a55159a,a55162a,a55165a,a55166a,a55167a,a55171a,a55172a,a55175a,a55178a,a55179a,a55180a,a55184a,a55185a,a55188a,a55191a,a55192a,a55193a,a55197a,a55198a,a55201a,a55204a,a55205a,a55206a,a55210a,a55211a,a55214a,a55217a,a55218a,a55219a,a55223a,a55224a,a55227a,a55230a,a55231a,a55232a,a55236a,a55237a,a55240a,a55243a,a55244a,a55245a,a55249a,a55250a,a55253a,a55256a,a55257a,a55258a,a55262a,a55263a,a55266a,a55269a,a55270a,a55271a,a55275a,a55276a,a55279a,a55282a,a55283a,a55284a,a55288a,a55289a,a55292a,a55295a,a55296a,a55297a,a55301a,a55302a,a55305a,a55308a,a55309a,a55310a,a55314a,a55315a,a55318a,a55321a,a55322a,a55323a,a55327a,a55328a,a55331a,a55334a,a55335a,a55336a,a55340a,a55341a,a55344a,a55347a,a55348a,a55349a,a55353a,a55354a,a55357a,a55360a,a55361a,a55362a,a55366a,a55367a,a55370a,a55373a,a55374a,a55375a,a55379a,a55380a,a55383a,a55386a,a55387a,a55388a,a55392a,a55393a,a55396a,a55399a,a55400a,a55401a,a55405a,a55406a,a55409a,a55412a,a55413a,a55414a,a55418a,a55419a,a55422a,a55425a,a55426a,a55427a,a55431a,a55432a,a55435a,a55438a,a55439a,a55440a,a55444a,a55445a,a55448a,a55451a,a55452a,a55453a,a55457a,a55458a,a55461a,a55464a,a55465a,a55466a,a55470a,a55471a,a55474a,a55477a,a55478a,a55479a,a55483a,a55484a,a55487a,a55490a,a55491a,a55492a,a55496a,a55497a,a55500a,a55503a,a55504a,a55505a,a55509a,a55510a,a55513a,a55516a,a55517a,a55518a,a55522a,a55523a,a55526a,a55529a,a55530a,a55531a,a55535a,a55536a,a55539a,a55542a,a55543a,a55544a,a55548a,a55549a,a55552a,a55555a,a55556a,a55557a,a55561a,a55562a,a55565a,a55568a,a55569a,a55570a,a55574a,a55575a,a55578a,a55581a,a55582a,a55583a,a55587a,a55588a,a55591a,a55594a,a55595a,a55596a,a55600a,a55601a,a55604a,a55607a,a55608a,a55609a,a55613a,a55614a,a55617a,a55620a,a55621a,a55622a,a55626a,a55627a,a55630a,a55633a,a55634a,a55635a,a55639a,a55640a,a55643a,a55646a,a55647a,a55648a,a55652a,a55653a,a55656a,a55659a,a55660a,a55661a,a55665a,a55666a,a55669a,a55672a,a55673a,a55674a,a55678a,a55679a,a55682a,a55685a,a55686a,a55687a,a55691a,a55692a,a55695a,a55698a,a55699a,a55700a,a55704a,a55705a,a55708a,a55711a,a55712a,a55713a,a55717a,a55718a,a55721a,a55724a,a55725a,a55726a,a55730a,a55731a,a55734a,a55737a,a55738a,a55739a,a55743a,a55744a,a55747a,a55750a,a55751a,a55752a,a55756a,a55757a,a55760a,a55763a,a55764a,a55765a,a55769a,a55770a,a55773a,a55776a,a55777a,a55778a,a55782a,a55783a,a55786a,a55789a,a55790a,a55791a,a55795a,a55796a,a55799a,a55802a,a55803a,a55804a,a55808a,a55809a,a55812a,a55815a,a55816a,a55817a,a55821a,a55822a,a55825a,a55828a,a55829a,a55830a,a55834a,a55835a,a55838a,a55841a,a55842a,a55843a,a55847a,a55848a,a55851a,a55854a,a55855a,a55856a,a55860a,a55861a,a55864a,a55867a,a55868a,a55869a,a55873a,a55874a,a55877a,a55880a,a55881a,a55882a,a55886a,a55887a,a55890a,a55893a,a55894a,a55895a,a55899a,a55900a,a55903a,a55906a,a55907a,a55908a,a55912a,a55913a,a55916a,a55919a,a55920a,a55921a,a55925a,a55926a,a55929a,a55932a,a55933a,a55934a,a55938a,a55939a,a55942a,a55945a,a55946a,a55947a,a55951a,a55952a,a55955a,a55958a,a55959a,a55960a,a55964a,a55965a,a55968a,a55971a,a55972a,a55973a,a55977a,a55978a,a55981a,a55984a,a55985a,a55986a,a55990a,a55991a,a55994a,a55997a,a55998a,a55999a,a56003a,a56004a,a56007a,a56010a,a56011a,a56012a,a56016a,a56017a,a56020a,a56023a,a56024a,a56025a,a56029a,a56030a,a56033a,a56036a,a56037a,a56038a,a56042a,a56043a,a56046a,a56049a,a56050a,a56051a,a56055a,a56056a,a56059a,a56062a,a56063a,a56064a,a56068a,a56069a,a56072a,a56075a,a56076a,a56077a,a56081a,a56082a,a56085a,a56088a,a56089a,a56090a,a56094a,a56095a,a56098a,a56101a,a56102a,a56103a,a56107a,a56108a,a56111a,a56114a,a56115a,a56116a,a56120a,a56121a,a56124a,a56127a,a56128a,a56129a,a56133a,a56134a,a56137a,a56140a,a56141a,a56142a,a56146a,a56147a,a56150a,a56153a,a56154a,a56155a,a56159a,a56160a,a56163a,a56166a,a56167a,a56168a,a56172a,a56173a,a56176a,a56179a,a56180a,a56181a,a56185a,a56186a,a56189a,a56192a,a56193a,a56194a,a56198a,a56199a,a56202a,a56205a,a56206a,a56207a,a56211a,a56212a,a56215a,a56218a,a56219a,a56220a,a56224a,a56225a,a56228a,a56231a,a56232a,a56233a,a56237a,a56238a,a56241a,a56244a,a56245a,a56246a,a56250a,a56251a,a56254a,a56257a,a56258a,a56259a,a56263a,a56264a,a56267a,a56270a,a56271a,a56272a,a56276a,a56277a,a56280a,a56283a,a56284a,a56285a,a56289a,a56290a,a56293a,a56296a,a56297a,a56298a,a56302a,a56303a,a56306a,a56309a,a56310a,a56311a,a56315a,a56316a,a56319a,a56322a,a56323a,a56324a,a56328a,a56329a,a56332a,a56335a,a56336a,a56337a,a56341a,a56342a,a56345a,a56348a,a56349a,a56350a,a56354a,a56355a,a56358a,a56361a,a56362a,a56363a,a56367a,a56368a,a56371a,a56374a,a56375a,a56376a,a56380a,a56381a,a56384a,a56387a,a56388a,a56389a,a56393a,a56394a,a56397a,a56400a,a56401a,a56402a,a56406a,a56407a,a56410a,a56413a,a56414a,a56415a,a56419a,a56420a,a56423a,a56426a,a56427a,a56428a,a56432a,a56433a,a56436a,a56439a,a56440a,a56441a,a56445a,a56446a,a56449a,a56452a,a56453a,a56454a,a56458a,a56459a,a56462a,a56465a,a56466a,a56467a,a56471a,a56472a,a56475a,a56478a,a56479a,a56480a,a56484a,a56485a,a56488a,a56491a,a56492a,a56493a,a56497a,a56498a,a56501a,a56504a,a56505a,a56506a,a56510a,a56511a,a56514a,a56517a,a56518a,a56519a,a56523a,a56524a,a56527a,a56530a,a56531a,a56532a,a56536a,a56537a,a56540a,a56543a,a56544a,a56545a,a56549a,a56550a,a56553a,a56556a,a56557a,a56558a,a56562a,a56563a,a56566a,a56569a,a56570a,a56571a,a56575a,a56576a,a56579a,a56582a,a56583a,a56584a,a56588a,a56589a,a56592a,a56595a,a56596a,a56597a,a56601a,a56602a,a56605a,a56608a,a56609a,a56610a,a56614a,a56615a,a56618a,a56621a,a56622a,a56623a,a56627a,a56628a,a56631a,a56634a,a56635a,a56636a,a56640a,a56641a,a56644a,a56647a,a56648a,a56649a,a56653a,a56654a,a56657a,a56660a,a56661a,a56662a,a56666a,a56667a,a56670a,a56673a,a56674a,a56675a,a56679a,a56680a,a56683a,a56686a,a56687a,a56688a,a56692a,a56693a,a56696a,a56699a,a56700a,a56701a,a56705a,a56706a,a56709a,a56712a,a56713a,a56714a,a56718a,a56719a,a56722a,a56725a,a56726a,a56727a,a56731a,a56732a,a56735a,a56738a,a56739a,a56740a,a56744a,a56745a,a56748a,a56751a,a56752a,a56753a,a56757a,a56758a,a56761a,a56764a,a56765a,a56766a,a56770a,a56771a,a56774a,a56777a,a56778a,a56779a,a56783a,a56784a,a56787a,a56790a,a56791a,a56792a,a56796a,a56797a,a56800a,a56803a,a56804a,a56805a,a56809a,a56810a,a56813a,a56816a,a56817a,a56818a,a56822a,a56823a,a56826a,a56829a,a56830a,a56831a,a56835a,a56836a,a56839a,a56842a,a56843a,a56844a,a56848a,a56849a,a56852a,a56855a,a56856a,a56857a,a56861a,a56862a,a56865a,a56868a,a56869a,a56870a,a56874a,a56875a,a56878a,a56881a,a56882a,a56883a,a56887a,a56888a,a56891a,a56894a,a56895a,a56896a,a56900a,a56901a,a56904a,a56907a,a56908a,a56909a,a56913a,a56914a,a56917a,a56920a,a56921a,a56922a,a56926a,a56927a,a56930a,a56933a,a56934a,a56935a,a56939a,a56940a,a56943a,a56946a,a56947a,a56948a,a56952a,a56953a,a56956a,a56959a,a56960a,a56961a,a56965a,a56966a,a56969a,a56972a,a56973a,a56974a,a56978a,a56979a,a56982a,a56985a,a56986a,a56987a,a56991a,a56992a,a56995a,a56998a,a56999a,a57000a,a57004a,a57005a,a57008a,a57011a,a57012a,a57013a,a57017a,a57018a,a57021a,a57024a,a57025a,a57026a,a57030a,a57031a,a57034a,a57037a,a57038a,a57039a,a57043a,a57044a,a57047a,a57050a,a57051a,a57052a,a57056a,a57057a,a57060a,a57063a,a57064a,a57065a,a57069a,a57070a,a57073a,a57076a,a57077a,a57078a,a57082a,a57083a,a57086a,a57089a,a57090a,a57091a,a57095a,a57096a,a57099a,a57102a,a57103a,a57104a,a57108a,a57109a,a57112a,a57115a,a57116a,a57117a,a57121a,a57122a,a57125a,a57128a,a57129a,a57130a,a57134a,a57135a,a57138a,a57141a,a57142a,a57143a,a57147a,a57148a,a57151a,a57154a,a57155a,a57156a,a57160a,a57161a,a57164a,a57167a,a57168a,a57169a,a57173a,a57174a,a57177a,a57180a,a57181a,a57182a,a57186a,a57187a,a57190a,a57193a,a57194a,a57195a,a57199a,a57200a,a57203a,a57206a,a57207a,a57208a,a57212a,a57213a,a57216a,a57219a,a57220a,a57221a,a57225a,a57226a,a57229a,a57232a,a57233a,a57234a,a57238a,a57239a,a57242a,a57245a,a57246a,a57247a,a57251a,a57252a,a57255a,a57258a,a57259a,a57260a,a57264a,a57265a,a57268a,a57271a,a57272a,a57273a,a57277a,a57278a,a57281a,a57284a,a57285a,a57286a,a57290a,a57291a,a57294a,a57297a,a57298a,a57299a,a57303a,a57304a,a57307a,a57310a,a57311a,a57312a,a57316a,a57317a,a57320a,a57323a,a57324a,a57325a,a57329a,a57330a,a57333a,a57336a,a57337a,a57338a,a57342a,a57343a,a57346a,a57349a,a57350a,a57351a,a57355a,a57356a,a57359a,a57362a,a57363a,a57364a,a57368a,a57369a,a57372a,a57375a,a57376a,a57377a,a57381a,a57382a,a57385a,a57388a,a57389a,a57390a,a57394a,a57395a,a57398a,a57401a,a57402a,a57403a,a57407a,a57408a,a57411a,a57414a,a57415a,a57416a,a57420a,a57421a,a57424a,a57427a,a57428a,a57429a,a57433a,a57434a,a57437a,a57440a,a57441a,a57442a,a57446a,a57447a,a57450a,a57453a,a57454a,a57455a,a57459a,a57460a,a57463a,a57466a,a57467a,a57468a,a57472a,a57473a,a57476a,a57479a,a57480a,a57481a,a57485a,a57486a,a57489a,a57492a,a57493a,a57494a,a57498a,a57499a,a57502a,a57505a,a57506a,a57507a,a57511a,a57512a,a57515a,a57518a,a57519a,a57520a,a57524a,a57525a,a57528a,a57531a,a57532a,a57533a,a57537a,a57538a,a57541a,a57544a,a57545a,a57546a,a57550a,a57551a,a57554a,a57557a,a57558a,a57559a,a57563a,a57564a,a57567a,a57570a,a57571a,a57572a,a57576a,a57577a,a57580a,a57583a,a57584a,a57585a,a57589a,a57590a,a57593a,a57596a,a57597a,a57598a,a57602a,a57603a,a57606a,a57609a,a57610a,a57611a,a57615a,a57616a,a57619a,a57622a,a57623a,a57624a,a57628a,a57629a,a57632a,a57635a,a57636a,a57637a,a57641a,a57642a,a57645a,a57648a,a57649a,a57650a,a57654a,a57655a,a57658a,a57661a,a57662a,a57663a,a57667a,a57668a,a57671a,a57674a,a57675a,a57676a,a57680a,a57681a,a57684a,a57687a,a57688a,a57689a,a57693a,a57694a,a57697a,a57700a,a57701a,a57702a,a57706a,a57707a,a57710a,a57713a,a57714a,a57715a,a57719a,a57720a,a57723a,a57726a,a57727a,a57728a,a57732a,a57733a,a57736a,a57739a,a57740a,a57741a,a57745a,a57746a,a57749a,a57752a,a57753a,a57754a,a57758a,a57759a,a57762a,a57765a,a57766a,a57767a,a57771a,a57772a,a57775a,a57778a,a57779a,a57780a,a57784a,a57785a,a57788a,a57791a,a57792a,a57793a,a57797a,a57798a,a57801a,a57804a,a57805a,a57806a,a57810a,a57811a,a57814a,a57817a,a57818a,a57819a,a57823a,a57824a,a57827a,a57830a,a57831a,a57832a,a57836a,a57837a,a57840a,a57843a,a57844a,a57845a,a57849a,a57850a,a57853a,a57856a,a57857a,a57858a,a57862a,a57863a,a57866a,a57869a,a57870a,a57871a,a57875a,a57876a,a57879a,a57882a,a57883a,a57884a,a57888a,a57889a,a57892a,a57895a,a57896a,a57897a,a57901a,a57902a,a57905a,a57908a,a57909a,a57910a,a57914a,a57915a,a57918a,a57921a,a57922a,a57923a,a57927a,a57928a,a57931a,a57934a,a57935a,a57936a,a57940a,a57941a,a57944a,a57947a,a57948a,a57949a,a57953a,a57954a,a57957a,a57960a,a57961a,a57962a,a57966a,a57967a,a57970a,a57973a,a57974a,a57975a,a57979a,a57980a,a57983a,a57986a,a57987a,a57988a,a57992a,a57993a,a57996a,a57999a,a58000a,a58001a,a58005a,a58006a,a58009a,a58012a,a58013a,a58014a,a58018a,a58019a,a58022a,a58025a,a58026a,a58027a,a58031a,a58032a,a58035a,a58038a,a58039a,a58040a,a58044a,a58045a,a58048a,a58051a,a58052a,a58053a,a58057a,a58058a,a58061a,a58064a,a58065a,a58066a,a58070a,a58071a,a58074a,a58077a,a58078a,a58079a,a58083a,a58084a,a58087a,a58090a,a58091a,a58092a,a58096a,a58097a,a58100a,a58103a,a58104a,a58105a,a58109a,a58110a,a58113a,a58116a,a58117a,a58118a,a58122a,a58123a,a58126a,a58129a,a58130a,a58131a,a58135a,a58136a,a58139a,a58142a,a58143a,a58144a,a58148a,a58149a,a58152a,a58155a,a58156a,a58157a,a58161a,a58162a,a58165a,a58168a,a58169a,a58170a,a58174a,a58175a,a58178a,a58181a,a58182a,a58183a,a58187a,a58188a,a58191a,a58194a,a58195a,a58196a,a58200a,a58201a,a58204a,a58207a,a58208a,a58209a,a58213a,a58214a,a58217a,a58220a,a58221a,a58222a,a58226a,a58227a,a58230a,a58233a,a58234a,a58235a,a58239a,a58240a,a58243a,a58246a,a58247a,a58248a,a58252a,a58253a,a58256a,a58259a,a58260a,a58261a,a58265a,a58266a,a58269a,a58272a,a58273a,a58274a,a58278a,a58279a,a58282a,a58285a,a58286a,a58287a,a58291a,a58292a,a58295a,a58298a,a58299a,a58300a,a58304a,a58305a,a58308a,a58311a,a58312a,a58313a,a58317a,a58318a,a58321a,a58324a,a58325a,a58326a,a58330a,a58331a,a58334a,a58337a,a58338a,a58339a,a58343a,a58344a,a58347a,a58350a,a58351a,a58352a,a58356a,a58357a,a58360a,a58363a,a58364a,a58365a,a58369a,a58370a,a58373a,a58376a,a58377a,a58378a,a58382a,a58383a,a58386a,a58389a,a58390a,a58391a,a58395a,a58396a,a58399a,a58402a,a58403a,a58404a,a58408a,a58409a,a58412a,a58415a,a58416a,a58417a,a58421a,a58422a,a58425a,a58428a,a58429a,a58430a,a58434a,a58435a,a58438a,a58441a,a58442a,a58443a,a58447a,a58448a,a58451a,a58454a,a58455a,a58456a,a58460a,a58461a,a58464a,a58467a,a58468a,a58469a,a58473a,a58474a,a58477a,a58480a,a58481a,a58482a,a58486a,a58487a,a58490a,a58493a,a58494a,a58495a,a58499a,a58500a,a58503a,a58506a,a58507a,a58508a,a58512a,a58513a,a58516a,a58519a,a58520a,a58521a,a58525a,a58526a,a58529a,a58532a,a58533a,a58534a,a58538a,a58539a,a58542a,a58545a,a58546a,a58547a,a58551a,a58552a,a58555a,a58558a,a58559a,a58560a,a58564a,a58565a,a58568a,a58571a,a58572a,a58573a,a58577a,a58578a,a58581a,a58584a,a58585a,a58586a,a58590a,a58591a,a58594a,a58597a,a58598a,a58599a,a58603a,a58604a,a58607a,a58610a,a58611a,a58612a,a58616a,a58617a,a58620a,a58623a,a58624a,a58625a,a58629a,a58630a,a58633a,a58636a,a58637a,a58638a,a58642a,a58643a,a58646a,a58649a,a58650a,a58651a,a58655a,a58656a,a58659a,a58662a,a58663a,a58664a,a58668a,a58669a,a58672a,a58675a,a58676a,a58677a,a58681a,a58682a,a58685a,a58688a,a58689a,a58690a,a58694a,a58695a,a58698a,a58701a,a58702a,a58703a,a58707a,a58708a,a58711a,a58714a,a58715a,a58716a,a58720a,a58721a,a58724a,a58727a,a58728a,a58729a,a58733a,a58734a,a58737a,a58740a,a58741a,a58742a,a58746a,a58747a,a58750a,a58753a,a58754a,a58755a,a58759a,a58760a,a58763a,a58766a,a58767a,a58768a,a58772a,a58773a,a58776a,a58779a,a58780a,a58781a,a58785a,a58786a,a58789a,a58792a,a58793a,a58794a,a58798a,a58799a,a58802a,a58805a,a58806a,a58807a,a58811a,a58812a,a58815a,a58818a,a58819a,a58820a,a58824a,a58825a,a58828a,a58831a,a58832a,a58833a,a58837a,a58838a,a58841a,a58844a,a58845a,a58846a,a58850a,a58851a,a58854a,a58857a,a58858a,a58859a,a58863a,a58864a,a58867a,a58870a,a58871a,a58872a,a58876a,a58877a,a58880a,a58883a,a58884a,a58885a,a58889a,a58890a,a58893a,a58896a,a58897a,a58898a,a58902a,a58903a,a58906a,a58909a,a58910a,a58911a,a58915a,a58916a,a58919a,a58922a,a58923a,a58924a,a58928a,a58929a,a58932a,a58935a,a58936a,a58937a,a58941a,a58942a,a58945a,a58948a,a58949a,a58950a,a58954a,a58955a,a58958a,a58961a,a58962a,a58963a,a58967a,a58968a,a58971a,a58974a,a58975a,a58976a,a58980a,a58981a,a58984a,a58987a,a58988a,a58989a,a58993a,a58994a,a58997a,a59000a,a59001a,a59002a,a59006a,a59007a,a59010a,a59013a,a59014a,a59015a,a59019a,a59020a,a59023a,a59026a,a59027a,a59028a,a59032a,a59033a,a59036a,a59039a,a59040a,a59041a,a59045a,a59046a,a59049a,a59052a,a59053a,a59054a,a59058a,a59059a,a59062a,a59065a,a59066a,a59067a,a59071a,a59072a,a59075a,a59078a,a59079a,a59080a,a59084a,a59085a,a59088a,a59091a,a59092a,a59093a,a59097a,a59098a,a59101a,a59104a,a59105a,a59106a,a59110a,a59111a,a59114a,a59117a,a59118a,a59119a,a59123a,a59124a,a59127a,a59130a,a59131a,a59132a,a59136a,a59137a,a59140a,a59143a,a59144a,a59145a,a59149a,a59150a,a59153a,a59156a,a59157a,a59158a,a59162a,a59163a,a59166a,a59169a,a59170a,a59171a,a59175a,a59176a,a59179a,a59182a,a59183a,a59184a,a59188a,a59189a,a59192a,a59195a,a59196a,a59197a,a59201a,a59202a,a59205a,a59208a,a59209a,a59210a,a59214a,a59215a,a59218a,a59221a,a59222a,a59223a,a59227a,a59228a,a59231a,a59234a,a59235a,a59236a,a59240a,a59241a,a59244a,a59247a,a59248a,a59249a,a59253a,a59254a,a59257a,a59260a,a59261a,a59262a,a59266a,a59267a,a59270a,a59273a,a59274a,a59275a,a59279a,a59280a,a59283a,a59286a,a59287a,a59288a,a59292a,a59293a,a59296a,a59299a,a59300a,a59301a,a59305a,a59306a,a59309a,a59312a,a59313a,a59314a,a59318a,a59319a,a59322a,a59325a,a59326a,a59327a,a59331a,a59332a,a59335a,a59338a,a59339a,a59340a,a59344a,a59345a,a59348a,a59351a,a59352a,a59353a,a59357a,a59358a,a59361a,a59364a,a59365a,a59366a,a59370a,a59371a,a59374a,a59377a,a59378a,a59379a,a59383a,a59384a,a59387a,a59390a,a59391a,a59392a,a59396a,a59397a,a59400a,a59403a,a59404a,a59405a,a59409a,a59410a,a59413a,a59416a,a59417a,a59418a,a59422a,a59423a,a59426a,a59429a,a59430a,a59431a,a59435a,a59436a,a59439a,a59442a,a59443a,a59444a,a59448a,a59449a,a59452a,a59455a,a59456a,a59457a,a59461a,a59462a,a59465a,a59468a,a59469a,a59470a,a59474a,a59475a,a59478a,a59481a,a59482a,a59483a,a59487a,a59488a,a59491a,a59494a,a59495a,a59496a,a59500a,a59501a,a59504a,a59507a,a59508a,a59509a,a59513a,a59514a,a59517a,a59520a,a59521a,a59522a,a59526a,a59527a,a59530a,a59533a,a59534a,a59535a,a59539a,a59540a,a59543a,a59546a,a59547a,a59548a,a59552a,a59553a,a59556a,a59559a,a59560a,a59561a,a59565a,a59566a,a59569a,a59572a,a59573a,a59574a,a59578a,a59579a,a59582a,a59585a,a59586a,a59587a,a59591a,a59592a,a59595a,a59598a,a59599a,a59600a,a59604a,a59605a,a59608a,a59611a,a59612a,a59613a,a59617a,a59618a,a59621a,a59624a,a59625a,a59626a,a59630a,a59631a,a59634a,a59637a,a59638a,a59639a,a59643a,a59644a,a59647a,a59650a,a59651a,a59652a,a59656a,a59657a,a59660a,a59663a,a59664a,a59665a,a59669a,a59670a,a59673a,a59676a,a59677a,a59678a,a59682a,a59683a,a59686a,a59689a,a59690a,a59691a,a59695a,a59696a,a59699a,a59702a,a59703a,a59704a,a59708a,a59709a,a59712a,a59715a,a59716a,a59717a,a59721a,a59722a,a59725a,a59728a,a59729a,a59730a,a59734a,a59735a,a59738a,a59741a,a59742a,a59743a,a59747a,a59748a,a59751a,a59754a,a59755a,a59756a,a59760a,a59761a,a59764a,a59767a,a59768a,a59769a,a59773a,a59774a,a59777a,a59780a,a59781a,a59782a,a59786a,a59787a,a59790a,a59793a,a59794a,a59795a,a59799a,a59800a,a59803a,a59806a,a59807a,a59808a,a59812a,a59813a,a59816a,a59819a,a59820a,a59821a,a59825a,a59826a,a59829a,a59832a,a59833a,a59834a,a59838a,a59839a,a59842a,a59845a,a59846a,a59847a,a59851a,a59852a,a59855a,a59858a,a59859a,a59860a,a59864a,a59865a,a59868a,a59871a,a59872a,a59873a,a59877a,a59878a,a59881a,a59884a,a59885a,a59886a,a59890a,a59891a,a59894a,a59897a,a59898a,a59899a,a59903a,a59904a,a59907a,a59910a,a59911a,a59912a,a59916a,a59917a,a59920a,a59923a,a59924a,a59925a,a59929a,a59930a,a59933a,a59936a,a59937a,a59938a,a59942a,a59943a,a59946a,a59949a,a59950a,a59951a,a59955a,a59956a,a59959a,a59962a,a59963a,a59964a,a59968a,a59969a,a59972a,a59975a,a59976a,a59977a,a59981a,a59982a,a59985a,a59988a,a59989a,a59990a,a59994a,a59995a,a59998a,a60001a,a60002a,a60003a,a60007a,a60008a,a60011a,a60014a,a60015a,a60016a,a60020a,a60021a,a60024a,a60027a,a60028a,a60029a,a60033a,a60034a,a60037a,a60040a,a60041a,a60042a,a60046a,a60047a,a60050a,a60053a,a60054a,a60055a,a60059a,a60060a,a60063a,a60066a,a60067a,a60068a,a60072a,a60073a,a60076a,a60079a,a60080a,a60081a,a60085a,a60086a,a60089a,a60092a,a60093a,a60094a,a60098a,a60099a,a60102a,a60105a,a60106a,a60107a,a60111a,a60112a,a60115a,a60118a,a60119a,a60120a,a60124a,a60125a,a60128a,a60131a,a60132a,a60133a,a60137a,a60138a,a60141a,a60144a,a60145a,a60146a,a60150a,a60151a,a60154a,a60157a,a60158a,a60159a,a60163a,a60164a,a60167a,a60170a,a60171a,a60172a,a60176a,a60177a,a60180a,a60183a,a60184a,a60185a,a60189a,a60190a,a60193a,a60196a,a60197a,a60198a,a60202a,a60203a,a60206a,a60209a,a60210a,a60211a,a60215a,a60216a,a60219a,a60222a,a60223a,a60224a,a60228a,a60229a,a60232a,a60235a,a60236a,a60237a,a60241a,a60242a,a60245a,a60248a,a60249a,a60250a,a60254a,a60255a,a60258a,a60261a,a60262a,a60263a,a60267a,a60268a,a60271a,a60274a,a60275a,a60276a,a60280a,a60281a,a60284a,a60287a,a60288a,a60289a,a60292a,a60295a,a60296a,a60299a,a60302a,a60303a,a60304a,a60308a,a60309a,a60312a,a60315a,a60316a,a60317a,a60320a,a60323a,a60324a,a60327a,a60330a,a60331a,a60332a,a60336a,a60337a,a60340a,a60343a,a60344a,a60345a,a60348a,a60351a,a60352a,a60355a,a60358a,a60359a,a60360a,a60364a,a60365a,a60368a,a60371a,a60372a,a60373a,a60376a,a60379a,a60380a,a60383a,a60386a,a60387a,a60388a,a60392a,a60393a,a60396a,a60399a,a60400a,a60401a,a60404a,a60407a,a60408a,a60411a,a60414a,a60415a,a60416a,a60420a,a60421a,a60424a,a60427a,a60428a,a60429a,a60432a,a60435a,a60436a,a60439a,a60442a,a60443a,a60444a,a60448a,a60449a,a60452a,a60455a,a60456a,a60457a,a60460a,a60463a,a60464a,a60467a,a60470a,a60471a,a60472a,a60476a,a60477a,a60480a,a60483a,a60484a,a60485a,a60488a,a60491a,a60492a,a60495a,a60498a,a60499a,a60500a,a60504a,a60505a,a60508a,a60511a,a60512a,a60513a,a60516a,a60519a,a60520a,a60523a,a60526a,a60527a,a60528a,a60532a,a60533a,a60536a,a60539a,a60540a,a60541a,a60544a,a60547a,a60548a,a60551a,a60554a,a60555a,a60556a,a60560a,a60561a,a60564a,a60567a,a60568a,a60569a,a60572a,a60575a,a60576a,a60579a,a60582a,a60583a,a60584a,a60588a,a60589a,a60592a,a60595a,a60596a,a60597a,a60600a,a60603a,a60604a,a60607a,a60610a,a60611a,a60612a,a60616a,a60617a,a60620a,a60623a,a60624a,a60625a,a60628a,a60631a,a60632a,a60635a,a60638a,a60639a,a60640a,a60644a,a60645a,a60648a,a60651a,a60652a,a60653a,a60656a,a60659a,a60660a,a60663a,a60666a,a60667a,a60668a,a60672a,a60673a,a60676a,a60679a,a60680a,a60681a,a60684a,a60687a,a60688a,a60691a,a60694a,a60695a,a60696a,a60700a,a60701a,a60704a,a60707a,a60708a,a60709a,a60712a,a60715a,a60716a,a60719a,a60722a,a60723a,a60724a,a60728a,a60729a,a60732a,a60735a,a60736a,a60737a,a60740a,a60743a,a60744a,a60747a,a60750a,a60751a,a60752a,a60756a,a60757a,a60760a,a60763a,a60764a,a60765a,a60768a,a60771a,a60772a,a60775a,a60778a,a60779a,a60780a,a60784a,a60785a,a60788a,a60791a,a60792a,a60793a,a60796a,a60799a,a60800a,a60803a,a60806a,a60807a,a60808a,a60812a,a60813a,a60816a,a60819a,a60820a,a60821a,a60824a,a60827a,a60828a,a60831a,a60834a,a60835a,a60836a,a60840a,a60841a,a60844a,a60847a,a60848a,a60849a,a60852a,a60855a,a60856a,a60859a,a60862a,a60863a,a60864a,a60868a,a60869a,a60872a,a60875a,a60876a,a60877a,a60880a,a60883a,a60884a,a60887a,a60890a,a60891a,a60892a,a60896a,a60897a,a60900a,a60903a,a60904a,a60905a,a60908a,a60911a,a60912a,a60915a,a60918a,a60919a,a60920a,a60924a,a60925a,a60928a,a60931a,a60932a,a60933a,a60936a,a60939a,a60940a,a60943a,a60946a,a60947a,a60948a,a60952a,a60953a,a60956a,a60959a,a60960a,a60961a,a60964a,a60967a,a60968a,a60971a,a60974a,a60975a,a60976a,a60980a,a60981a,a60984a,a60987a,a60988a,a60989a,a60992a,a60995a,a60996a,a60999a,a61002a,a61003a,a61004a,a61008a,a61009a,a61012a,a61015a,a61016a,a61017a,a61020a,a61023a,a61024a,a61027a,a61030a,a61031a,a61032a,a61036a,a61037a,a61040a,a61043a,a61044a,a61045a,a61048a,a61051a,a61052a,a61055a,a61058a,a61059a,a61060a,a61064a,a61065a,a61068a,a61071a,a61072a,a61073a,a61076a,a61079a,a61080a,a61083a,a61086a,a61087a,a61088a,a61092a,a61093a,a61096a,a61099a,a61100a,a61101a,a61104a,a61107a,a61108a,a61111a,a61114a,a61115a,a61116a,a61120a,a61121a,a61124a,a61127a,a61128a,a61129a,a61132a,a61135a,a61136a,a61139a,a61142a,a61143a,a61144a,a61148a,a61149a,a61152a,a61155a,a61156a,a61157a,a61160a,a61163a,a61164a,a61167a,a61170a,a61171a,a61172a,a61176a,a61177a,a61180a,a61183a,a61184a,a61185a,a61188a,a61191a,a61192a,a61195a,a61198a,a61199a,a61200a,a61204a,a61205a,a61208a,a61211a,a61212a,a61213a,a61216a,a61219a,a61220a,a61223a,a61226a,a61227a,a61228a,a61232a,a61233a,a61236a,a61239a,a61240a,a61241a,a61244a,a61247a,a61248a,a61251a,a61254a,a61255a,a61256a,a61260a,a61261a,a61264a,a61267a,a61268a,a61269a,a61272a,a61275a,a61276a,a61279a,a61282a,a61283a,a61284a,a61288a,a61289a,a61292a,a61295a,a61296a,a61297a,a61300a,a61303a,a61304a,a61307a,a61310a,a61311a,a61312a,a61316a,a61317a,a61320a,a61323a,a61324a,a61325a,a61328a,a61331a,a61332a,a61335a,a61338a,a61339a,a61340a,a61344a,a61345a,a61348a,a61351a,a61352a,a61353a,a61356a,a61359a,a61360a,a61363a,a61366a,a61367a,a61368a,a61372a,a61373a,a61376a,a61379a,a61380a,a61381a,a61384a,a61387a,a61388a,a61391a,a61394a,a61395a,a61396a,a61400a,a61401a,a61404a,a61407a,a61408a,a61409a,a61412a,a61415a,a61416a,a61419a,a61422a,a61423a,a61424a,a61428a,a61429a,a61432a,a61435a,a61436a,a61437a,a61440a,a61443a,a61444a,a61447a,a61450a,a61451a,a61452a,a61456a,a61457a,a61460a,a61463a,a61464a,a61465a,a61468a,a61471a,a61472a,a61475a,a61478a,a61479a,a61480a,a61484a,a61485a,a61488a,a61491a,a61492a,a61493a,a61496a,a61499a,a61500a,a61503a,a61506a,a61507a,a61508a,a61512a,a61513a,a61516a,a61519a,a61520a,a61521a,a61524a,a61527a,a61528a,a61531a,a61534a,a61535a,a61536a,a61540a,a61541a,a61544a,a61547a,a61548a,a61549a,a61552a,a61555a,a61556a,a61559a,a61562a,a61563a,a61564a,a61568a,a61569a,a61572a,a61575a,a61576a,a61577a,a61580a,a61583a,a61584a,a61587a,a61590a,a61591a,a61592a,a61596a,a61597a,a61600a,a61603a,a61604a,a61605a,a61608a,a61611a,a61612a,a61615a,a61618a,a61619a,a61620a,a61624a,a61625a,a61628a,a61631a,a61632a,a61633a,a61636a,a61639a,a61640a,a61643a,a61646a,a61647a,a61648a,a61652a,a61653a,a61656a,a61659a,a61660a,a61661a,a61664a,a61667a,a61668a,a61671a,a61674a,a61675a,a61676a,a61680a,a61681a,a61684a,a61687a,a61688a,a61689a,a61692a,a61695a,a61696a,a61699a,a61702a,a61703a,a61704a,a61708a,a61709a,a61712a,a61715a,a61716a,a61717a,a61720a,a61723a,a61724a,a61727a,a61730a,a61731a,a61732a,a61736a,a61737a,a61740a,a61743a,a61744a,a61745a,a61748a,a61751a,a61752a,a61755a,a61758a,a61759a,a61760a,a61764a,a61765a,a61768a,a61771a,a61772a,a61773a,a61776a,a61779a,a61780a,a61783a,a61786a,a61787a,a61788a,a61792a,a61793a,a61796a,a61799a,a61800a,a61801a,a61804a,a61807a,a61808a,a61811a,a61814a,a61815a,a61816a,a61820a,a61821a,a61824a,a61827a,a61828a,a61829a,a61832a,a61835a,a61836a,a61839a,a61842a,a61843a,a61844a,a61848a,a61849a,a61852a,a61855a,a61856a,a61857a,a61860a,a61863a,a61864a,a61867a,a61870a,a61871a,a61872a,a61876a,a61877a,a61880a,a61883a,a61884a,a61885a,a61888a,a61891a,a61892a,a61895a,a61898a,a61899a,a61900a,a61904a,a61905a,a61908a,a61911a,a61912a,a61913a,a61916a,a61919a,a61920a,a61923a,a61926a,a61927a,a61928a,a61932a,a61933a,a61936a,a61939a,a61940a,a61941a,a61944a,a61947a,a61948a,a61951a,a61954a,a61955a,a61956a,a61960a,a61961a,a61964a,a61967a,a61968a,a61969a,a61972a,a61975a,a61976a,a61979a,a61982a,a61983a,a61984a,a61988a,a61989a,a61992a,a61995a,a61996a,a61997a,a62000a,a62003a,a62004a,a62007a,a62010a,a62011a,a62012a,a62016a,a62017a,a62020a,a62023a,a62024a,a62025a,a62028a,a62031a,a62032a,a62035a,a62038a,a62039a,a62040a,a62044a,a62045a,a62048a,a62051a,a62052a,a62053a,a62056a,a62059a,a62060a,a62063a,a62066a,a62067a,a62068a,a62072a,a62073a,a62076a,a62079a,a62080a,a62081a,a62084a,a62087a,a62088a,a62091a,a62094a,a62095a,a62096a,a62100a,a62101a,a62104a,a62107a,a62108a,a62109a,a62112a,a62115a,a62116a,a62119a,a62122a,a62123a,a62124a,a62128a,a62129a,a62132a,a62135a,a62136a,a62137a,a62140a,a62143a,a62144a,a62147a,a62150a,a62151a,a62152a,a62156a,a62157a,a62160a,a62163a,a62164a,a62165a,a62168a,a62171a,a62172a,a62175a,a62178a,a62179a,a62180a,a62184a,a62185a,a62188a,a62191a,a62192a,a62193a,a62196a,a62199a,a62200a,a62203a,a62206a,a62207a,a62208a,a62212a,a62213a,a62216a,a62219a,a62220a,a62221a,a62224a,a62227a,a62228a,a62231a,a62234a,a62235a,a62236a,a62240a,a62241a,a62244a,a62247a,a62248a,a62249a,a62252a,a62255a,a62256a,a62259a,a62262a,a62263a,a62264a,a62268a,a62269a,a62272a,a62275a,a62276a,a62277a,a62280a,a62283a,a62284a,a62287a,a62290a,a62291a,a62292a,a62296a,a62297a,a62300a,a62303a,a62304a,a62305a,a62308a,a62311a,a62312a,a62315a,a62318a,a62319a,a62320a,a62324a,a62325a,a62328a,a62331a,a62332a,a62333a,a62336a,a62339a,a62340a,a62343a,a62346a,a62347a,a62348a,a62352a,a62353a,a62356a,a62359a,a62360a,a62361a,a62364a,a62367a,a62368a,a62371a,a62374a,a62375a,a62376a,a62380a,a62381a,a62384a,a62387a,a62388a,a62389a,a62392a,a62395a,a62396a,a62399a,a62402a,a62403a,a62404a,a62408a,a62409a,a62412a,a62415a,a62416a,a62417a,a62420a,a62423a,a62424a,a62427a,a62430a,a62431a,a62432a,a62436a,a62437a,a62440a,a62443a,a62444a,a62445a,a62448a,a62451a,a62452a,a62455a,a62458a,a62459a,a62460a,a62464a,a62465a,a62468a,a62471a,a62472a,a62473a,a62476a,a62479a,a62480a,a62483a,a62486a,a62487a,a62488a,a62492a,a62493a,a62496a,a62499a,a62500a,a62501a,a62504a,a62507a,a62508a,a62511a,a62514a,a62515a,a62516a,a62520a,a62521a,a62524a,a62527a,a62528a,a62529a,a62532a,a62535a,a62536a,a62539a,a62542a,a62543a,a62544a,a62548a,a62549a,a62552a,a62555a,a62556a,a62557a,a62560a,a62563a,a62564a,a62567a,a62570a,a62571a,a62572a,a62576a,a62577a,a62580a,a62583a,a62584a,a62585a,a62588a,a62591a,a62592a,a62595a,a62598a,a62599a,a62600a,a62604a,a62605a,a62608a,a62611a,a62612a,a62613a,a62616a,a62619a,a62620a,a62623a,a62626a,a62627a,a62628a,a62632a,a62633a,a62636a,a62639a,a62640a,a62641a,a62644a,a62647a,a62648a,a62651a,a62654a,a62655a,a62656a,a62660a,a62661a,a62664a,a62667a,a62668a,a62669a,a62672a,a62675a,a62676a,a62679a,a62682a,a62683a,a62684a,a62688a,a62689a,a62692a,a62695a,a62696a,a62697a,a62700a,a62703a,a62704a,a62707a,a62710a,a62711a,a62712a,a62716a,a62717a,a62720a,a62723a,a62724a,a62725a,a62728a,a62731a,a62732a,a62735a,a62738a,a62739a,a62740a,a62744a,a62745a,a62748a,a62751a,a62752a,a62753a,a62756a,a62759a,a62760a,a62763a,a62766a,a62767a,a62768a,a62772a,a62773a,a62776a,a62779a,a62780a,a62781a,a62784a,a62787a,a62788a,a62791a,a62794a,a62795a,a62796a,a62800a,a62801a,a62804a,a62807a,a62808a,a62809a,a62812a,a62815a,a62816a,a62819a,a62822a,a62823a,a62824a,a62828a,a62829a,a62832a,a62835a,a62836a,a62837a,a62840a,a62843a,a62844a,a62847a,a62850a,a62851a,a62852a,a62856a,a62857a,a62860a,a62863a,a62864a,a62865a,a62868a,a62871a,a62872a,a62875a,a62878a,a62879a,a62880a,a62884a,a62885a,a62888a,a62891a,a62892a,a62893a,a62896a,a62899a,a62900a,a62903a,a62906a,a62907a,a62908a,a62912a,a62913a,a62916a,a62919a,a62920a,a62921a,a62924a,a62927a,a62928a,a62931a,a62934a,a62935a,a62936a,a62940a,a62941a,a62944a,a62947a,a62948a,a62949a,a62952a,a62955a,a62956a,a62959a,a62962a,a62963a,a62964a,a62968a,a62969a,a62972a,a62975a,a62976a,a62977a,a62980a,a62983a,a62984a,a62987a,a62990a,a62991a,a62992a,a62996a,a62997a,a63000a,a63003a,a63004a,a63005a,a63008a,a63011a,a63012a,a63015a,a63018a,a63019a,a63020a,a63024a,a63025a,a63028a,a63031a,a63032a,a63033a,a63036a,a63039a,a63040a,a63043a,a63046a,a63047a,a63048a,a63052a,a63053a,a63056a,a63059a,a63060a,a63061a,a63064a,a63067a,a63068a,a63071a,a63074a,a63075a,a63076a,a63080a,a63081a,a63084a,a63087a,a63088a,a63089a,a63092a,a63095a,a63096a,a63099a,a63102a,a63103a,a63104a,a63108a,a63109a,a63112a,a63115a,a63116a,a63117a,a63120a,a63123a,a63124a,a63127a,a63130a,a63131a,a63132a,a63136a,a63137a,a63140a,a63143a,a63144a,a63145a,a63148a,a63151a,a63152a,a63155a,a63158a,a63159a,a63160a,a63164a,a63165a,a63168a,a63171a,a63172a,a63173a,a63176a,a63179a,a63180a,a63183a,a63186a,a63187a,a63188a,a63192a,a63193a,a63196a,a63199a,a63200a,a63201a,a63204a,a63207a,a63208a,a63211a,a63214a,a63215a,a63216a,a63220a,a63221a,a63224a,a63227a,a63228a,a63229a,a63232a,a63235a,a63236a,a63239a,a63242a,a63243a,a63244a,a63248a,a63249a,a63252a,a63255a,a63256a,a63257a,a63260a,a63263a,a63264a,a63267a,a63270a,a63271a,a63272a,a63276a,a63277a,a63280a,a63283a,a63284a,a63285a,a63288a,a63291a,a63292a,a63295a,a63298a,a63299a,a63300a,a63304a,a63305a,a63308a,a63311a,a63312a,a63313a,a63316a,a63319a,a63320a,a63323a,a63326a,a63327a,a63328a,a63332a,a63333a,a63336a,a63339a,a63340a,a63341a,a63344a,a63347a,a63348a,a63351a,a63354a,a63355a,a63356a,a63360a,a63361a,a63364a,a63367a,a63368a,a63369a,a63372a,a63375a,a63376a,a63379a,a63382a,a63383a,a63384a,a63388a,a63389a,a63392a,a63395a,a63396a,a63397a,a63400a,a63403a,a63404a,a63407a,a63410a,a63411a,a63412a,a63416a,a63417a,a63420a,a63423a,a63424a,a63425a,a63428a,a63431a,a63432a,a63435a,a63438a,a63439a,a63440a,a63444a,a63445a,a63448a,a63451a,a63452a,a63453a,a63456a,a63459a,a63460a,a63463a,a63466a,a63467a,a63468a,a63472a,a63473a,a63476a,a63479a,a63480a,a63481a,a63484a,a63487a,a63488a,a63491a,a63494a,a63495a,a63496a,a63500a,a63501a,a63504a,a63507a,a63508a,a63509a,a63512a,a63515a,a63516a,a63519a,a63522a,a63523a,a63524a,a63528a,a63529a,a63532a,a63535a,a63536a,a63537a,a63540a,a63543a,a63544a,a63547a,a63550a,a63551a,a63552a,a63556a,a63557a,a63560a,a63563a,a63564a,a63565a,a63568a,a63571a,a63572a,a63575a,a63578a,a63579a,a63580a,a63584a,a63585a,a63588a,a63591a,a63592a,a63593a,a63596a,a63599a,a63600a,a63603a,a63606a,a63607a,a63608a,a63612a,a63613a,a63616a,a63619a,a63620a,a63621a,a63624a,a63627a,a63628a,a63631a,a63634a,a63635a,a63636a,a63640a,a63641a,a63644a,a63647a,a63648a,a63649a,a63652a,a63655a,a63656a,a63659a,a63662a,a63663a,a63664a,a63668a,a63669a,a63672a,a63675a,a63676a,a63677a,a63680a,a63683a,a63684a,a63687a,a63690a,a63691a,a63692a,a63696a,a63697a,a63700a,a63703a,a63704a,a63705a,a63708a,a63711a,a63712a,a63715a,a63718a,a63719a,a63720a,a63724a,a63725a,a63728a,a63731a,a63732a,a63733a,a63736a,a63739a,a63740a,a63743a,a63746a,a63747a,a63748a,a63752a,a63753a,a63756a,a63759a,a63760a,a63761a,a63764a,a63767a,a63768a,a63771a,a63774a,a63775a,a63776a,a63780a,a63781a,a63784a,a63787a,a63788a,a63789a,a63792a,a63795a,a63796a,a63799a,a63802a,a63803a,a63804a,a63808a,a63809a,a63812a,a63815a,a63816a,a63817a,a63820a,a63823a,a63824a,a63827a,a63830a,a63831a,a63832a,a63836a,a63837a,a63840a,a63843a,a63844a,a63845a,a63848a,a63851a,a63852a,a63855a,a63858a,a63859a,a63860a,a63864a,a63865a,a63868a,a63871a,a63872a,a63873a,a63876a,a63879a,a63880a,a63883a,a63886a,a63887a,a63888a,a63892a,a63893a,a63896a,a63899a,a63900a,a63901a,a63904a,a63907a,a63908a,a63911a,a63914a,a63915a,a63916a,a63920a,a63921a,a63924a,a63927a,a63928a,a63929a,a63932a,a63935a,a63936a,a63939a,a63942a,a63943a,a63944a,a63948a,a63949a,a63952a,a63955a,a63956a,a63957a,a63960a,a63963a,a63964a,a63967a,a63970a,a63971a,a63972a,a63976a,a63977a,a63980a,a63983a,a63984a,a63985a,a63988a,a63991a,a63992a,a63995a,a63998a,a63999a,a64000a,a64004a,a64005a,a64008a,a64011a,a64012a,a64013a,a64016a,a64019a,a64020a,a64023a,a64026a,a64027a,a64028a,a64032a,a64033a,a64036a,a64039a,a64040a,a64041a,a64044a,a64047a,a64048a,a64051a,a64054a,a64055a,a64056a,a64060a,a64061a,a64064a,a64067a,a64068a,a64069a,a64072a,a64075a,a64076a,a64079a,a64082a,a64083a,a64084a,a64088a,a64089a,a64092a,a64095a,a64096a,a64097a,a64100a,a64103a,a64104a,a64107a,a64110a,a64111a,a64112a,a64116a,a64117a,a64120a,a64123a,a64124a,a64125a,a64128a,a64131a,a64132a,a64135a,a64138a,a64139a,a64140a,a64144a,a64145a,a64148a,a64151a,a64152a,a64153a,a64156a,a64159a,a64160a,a64163a,a64166a,a64167a,a64168a,a64172a,a64173a,a64176a,a64179a,a64180a,a64181a,a64184a,a64187a,a64188a,a64191a,a64194a,a64195a,a64196a,a64200a,a64201a,a64204a,a64207a,a64208a,a64209a,a64212a,a64215a,a64216a,a64219a,a64222a,a64223a,a64224a,a64228a,a64229a,a64232a,a64235a,a64236a,a64237a,a64240a,a64243a,a64244a,a64247a,a64250a,a64251a,a64252a,a64256a,a64257a,a64260a,a64263a,a64264a,a64265a,a64268a,a64271a,a64272a,a64275a,a64278a,a64279a,a64280a,a64284a,a64285a,a64288a,a64291a,a64292a,a64293a,a64296a,a64299a,a64300a,a64303a,a64306a,a64307a,a64308a,a64312a,a64313a,a64316a,a64319a,a64320a,a64321a,a64324a,a64327a,a64328a,a64331a,a64334a,a64335a,a64336a,a64340a,a64341a,a64344a,a64347a,a64348a,a64349a,a64352a,a64355a,a64356a,a64359a,a64362a,a64363a,a64364a,a64368a,a64369a,a64372a,a64375a,a64376a,a64377a,a64380a,a64383a,a64384a,a64387a,a64390a,a64391a,a64392a,a64396a,a64397a,a64400a,a64403a,a64404a,a64405a,a64408a,a64411a,a64412a,a64415a,a64418a,a64419a,a64420a,a64424a,a64425a,a64428a,a64431a,a64432a,a64433a,a64436a,a64439a,a64440a,a64443a,a64446a,a64447a,a64448a,a64452a,a64453a,a64456a,a64459a,a64460a,a64461a,a64464a,a64467a,a64468a,a64471a,a64474a,a64475a,a64476a,a64480a,a64481a,a64484a,a64487a,a64488a,a64489a,a64492a,a64495a,a64496a,a64499a,a64502a,a64503a,a64504a,a64508a,a64509a,a64512a,a64515a,a64516a,a64517a,a64520a,a64523a,a64524a,a64527a,a64530a,a64531a,a64532a,a64536a,a64537a,a64540a,a64543a,a64544a,a64545a,a64548a,a64551a,a64552a,a64555a,a64558a,a64559a,a64560a,a64564a,a64565a,a64568a,a64571a,a64572a,a64573a,a64576a,a64579a,a64580a,a64583a,a64586a,a64587a,a64588a,a64592a,a64593a,a64596a,a64599a,a64600a,a64601a,a64604a,a64607a,a64608a,a64611a,a64614a,a64615a,a64616a,a64620a,a64621a,a64624a,a64627a,a64628a,a64629a,a64632a,a64635a,a64636a,a64639a,a64642a,a64643a,a64644a,a64648a,a64649a,a64652a,a64655a,a64656a,a64657a,a64660a,a64663a,a64664a,a64667a,a64670a,a64671a,a64672a,a64676a,a64677a,a64680a,a64683a,a64684a,a64685a,a64688a,a64691a,a64692a,a64695a,a64698a,a64699a,a64700a,a64704a,a64705a,a64708a,a64711a,a64712a,a64713a,a64716a,a64719a,a64720a,a64723a,a64726a,a64727a,a64728a,a64732a,a64733a,a64736a,a64739a,a64740a,a64741a,a64744a,a64747a,a64748a,a64751a,a64754a,a64755a,a64756a,a64760a,a64761a,a64764a,a64767a,a64768a,a64769a,a64772a,a64775a,a64776a,a64779a,a64782a,a64783a,a64784a,a64788a,a64789a,a64792a,a64795a,a64796a,a64797a,a64800a,a64803a,a64804a,a64807a,a64810a,a64811a,a64812a,a64816a,a64817a,a64820a,a64823a,a64824a,a64825a,a64828a,a64831a,a64832a,a64835a,a64838a,a64839a,a64840a,a64844a,a64845a,a64848a,a64851a,a64852a,a64853a,a64856a,a64859a,a64860a,a64863a,a64866a,a64867a,a64868a,a64872a,a64873a,a64876a,a64879a,a64880a,a64881a,a64884a,a64887a,a64888a,a64891a,a64894a,a64895a,a64896a,a64900a,a64901a,a64904a,a64907a,a64908a,a64909a,a64912a,a64915a,a64916a,a64919a,a64922a,a64923a,a64924a,a64928a,a64929a,a64932a,a64935a,a64936a,a64937a,a64940a,a64943a,a64944a,a64947a,a64950a,a64951a,a64952a,a64956a,a64957a,a64960a,a64963a,a64964a,a64965a,a64968a,a64971a,a64972a,a64975a,a64978a,a64979a,a64980a,a64984a,a64985a,a64988a,a64991a,a64992a,a64993a,a64996a,a64999a,a65000a,a65003a,a65006a,a65007a,a65008a,a65012a,a65013a,a65016a,a65019a,a65020a,a65021a,a65024a,a65027a,a65028a,a65031a,a65034a,a65035a,a65036a,a65040a,a65041a,a65044a,a65047a,a65048a,a65049a,a65052a,a65055a,a65056a,a65059a,a65062a,a65063a,a65064a,a65068a,a65069a,a65072a,a65075a,a65076a,a65077a,a65080a,a65083a,a65084a,a65087a,a65090a,a65091a,a65092a,a65096a,a65097a,a65100a,a65103a,a65104a,a65105a,a65108a,a65111a,a65112a,a65115a,a65118a,a65119a,a65120a,a65124a,a65125a,a65128a,a65131a,a65132a,a65133a,a65136a,a65139a,a65140a,a65143a,a65146a,a65147a,a65148a,a65152a,a65153a,a65156a,a65159a,a65160a,a65161a,a65164a,a65167a,a65168a,a65171a,a65174a,a65175a,a65176a,a65180a,a65181a,a65184a,a65187a,a65188a,a65189a,a65192a,a65195a,a65196a,a65199a,a65202a,a65203a,a65204a,a65208a,a65209a,a65212a,a65215a,a65216a,a65217a,a65220a,a65223a,a65224a,a65227a,a65230a,a65231a,a65232a,a65236a,a65237a,a65240a,a65243a,a65244a,a65245a,a65248a,a65251a,a65252a,a65255a,a65258a,a65259a,a65260a,a65264a,a65265a,a65268a,a65271a,a65272a,a65273a,a65276a,a65279a,a65280a,a65283a,a65286a,a65287a,a65288a,a65292a,a65293a,a65296a,a65299a,a65300a,a65301a,a65304a,a65307a,a65308a,a65311a,a65314a,a65315a,a65316a,a65320a,a65321a,a65324a,a65327a,a65328a,a65329a,a65332a,a65335a,a65336a,a65339a,a65342a,a65343a,a65344a,a65348a,a65349a,a65352a,a65355a,a65356a,a65357a,a65360a,a65363a,a65364a,a65367a,a65370a,a65371a,a65372a,a65376a,a65377a,a65380a,a65383a,a65384a,a65385a,a65388a,a65391a,a65392a,a65395a,a65398a,a65399a,a65400a,a65404a,a65405a,a65408a,a65411a,a65412a,a65413a,a65416a,a65419a,a65420a,a65423a,a65426a,a65427a,a65428a,a65432a,a65433a,a65436a,a65439a,a65440a,a65441a,a65444a,a65447a,a65448a,a65451a,a65454a,a65455a,a65456a,a65460a,a65461a,a65464a,a65467a,a65468a,a65469a,a65472a,a65475a,a65476a,a65479a,a65482a,a65483a,a65484a,a65488a,a65489a,a65492a,a65495a,a65496a,a65497a,a65500a,a65503a,a65504a,a65507a,a65510a,a65511a,a65512a,a65516a,a65517a,a65520a,a65523a,a65524a,a65525a,a65528a,a65531a,a65532a,a65535a,a65538a,a65539a,a65540a,a65544a,a65545a,a65548a,a65551a,a65552a,a65553a,a65556a,a65559a,a65560a,a65563a,a65566a,a65567a,a65568a,a65572a,a65573a,a65576a,a65579a,a65580a,a65581a,a65584a,a65587a,a65588a,a65591a,a65594a,a65595a,a65596a,a65600a,a65601a,a65604a,a65607a,a65608a,a65609a,a65612a,a65615a,a65616a,a65619a,a65622a,a65623a,a65624a,a65628a,a65629a,a65632a,a65635a,a65636a,a65637a,a65640a,a65643a,a65644a,a65647a,a65650a,a65651a,a65652a,a65656a,a65657a,a65660a,a65663a,a65664a,a65665a,a65668a,a65671a,a65672a,a65675a,a65678a,a65679a,a65680a,a65684a,a65685a,a65688a,a65691a,a65692a,a65693a,a65696a,a65699a,a65700a,a65703a,a65706a,a65707a,a65708a,a65712a,a65713a,a65716a,a65719a,a65720a,a65721a,a65724a,a65727a,a65728a,a65731a,a65734a,a65735a,a65736a,a65740a,a65741a,a65744a,a65747a,a65748a,a65749a,a65752a,a65755a,a65756a,a65759a,a65762a,a65763a,a65764a,a65768a,a65769a,a65772a,a65775a,a65776a,a65777a,a65780a,a65783a,a65784a,a65787a,a65790a,a65791a,a65792a,a65796a,a65797a,a65800a,a65803a,a65804a,a65805a,a65808a,a65811a,a65812a,a65815a,a65818a,a65819a,a65820a,a65824a,a65825a,a65828a,a65831a,a65832a,a65833a,a65836a,a65839a,a65840a,a65843a,a65846a,a65847a,a65848a,a65852a,a65853a,a65856a,a65859a,a65860a,a65861a,a65864a,a65867a,a65868a,a65871a,a65874a,a65875a,a65876a,a65880a,a65881a,a65884a,a65887a,a65888a,a65889a,a65892a,a65895a,a65896a,a65899a,a65902a,a65903a,a65904a,a65908a,a65909a,a65912a,a65915a,a65916a,a65917a,a65920a,a65923a,a65924a,a65927a,a65930a,a65931a,a65932a,a65936a,a65937a,a65940a,a65943a,a65944a,a65945a,a65948a,a65951a,a65952a,a65955a,a65958a,a65959a,a65960a,a65964a,a65965a,a65968a,a65971a,a65972a,a65973a,a65976a,a65979a,a65980a,a65983a,a65986a,a65987a,a65988a,a65992a,a65993a,a65996a,a65999a,a66000a,a66001a,a66004a,a66007a,a66008a,a66011a,a66014a,a66015a,a66016a,a66020a,a66021a,a66024a,a66027a,a66028a,a66029a,a66032a,a66035a,a66036a,a66039a,a66042a,a66043a,a66044a,a66048a,a66049a,a66052a,a66055a,a66056a,a66057a,a66060a,a66063a,a66064a,a66067a,a66070a,a66071a,a66072a,a66076a,a66077a,a66080a,a66083a,a66084a,a66085a,a66088a,a66091a,a66092a,a66095a,a66098a,a66099a,a66100a,a66104a,a66105a,a66108a,a66111a,a66112a,a66113a,a66116a,a66119a,a66120a,a66123a,a66126a,a66127a,a66128a,a66132a,a66133a,a66136a,a66139a,a66140a,a66141a,a66144a,a66147a,a66148a,a66151a,a66154a,a66155a,a66156a,a66160a,a66161a,a66164a,a66167a,a66168a,a66169a,a66172a,a66175a,a66176a,a66179a,a66182a,a66183a,a66184a,a66188a,a66189a,a66192a,a66195a,a66196a,a66197a,a66200a,a66203a,a66204a,a66207a,a66210a,a66211a,a66212a,a66216a,a66217a,a66220a,a66223a,a66224a,a66225a,a66228a,a66231a,a66232a,a66235a,a66238a,a66239a,a66240a,a66244a,a66245a,a66248a,a66251a,a66252a,a66253a,a66256a,a66259a,a66260a,a66263a,a66266a,a66267a,a66268a,a66272a,a66273a,a66276a,a66279a,a66280a,a66281a,a66284a,a66287a,a66288a,a66291a,a66294a,a66295a,a66296a,a66300a,a66301a,a66304a,a66307a,a66308a,a66309a,a66312a,a66315a,a66316a,a66319a,a66322a,a66323a,a66324a,a66328a,a66329a,a66332a,a66335a,a66336a,a66337a,a66340a,a66343a,a66344a,a66347a,a66350a,a66351a,a66352a,a66356a,a66357a,a66360a,a66363a,a66364a,a66365a,a66368a,a66371a,a66372a,a66375a,a66378a,a66379a,a66380a,a66384a,a66385a,a66388a,a66391a,a66392a,a66393a,a66396a,a66399a,a66400a,a66403a,a66406a,a66407a,a66408a,a66412a,a66413a,a66416a,a66419a,a66420a,a66421a,a66424a,a66427a,a66428a,a66431a,a66434a,a66435a,a66436a,a66440a,a66441a,a66444a,a66447a,a66448a,a66449a,a66452a,a66455a,a66456a,a66459a,a66462a,a66463a,a66464a,a66468a,a66469a,a66472a,a66475a,a66476a,a66477a,a66480a,a66483a,a66484a,a66487a,a66490a,a66491a,a66492a,a66496a,a66497a,a66500a,a66503a,a66504a,a66505a,a66508a,a66511a,a66512a,a66515a,a66518a,a66519a,a66520a,a66524a,a66525a,a66528a,a66531a,a66532a,a66533a,a66536a,a66539a,a66540a,a66543a,a66546a,a66547a,a66548a,a66552a,a66553a,a66556a,a66559a,a66560a,a66561a,a66564a,a66567a,a66568a,a66571a,a66574a,a66575a,a66576a,a66580a,a66581a,a66584a,a66587a,a66588a,a66589a,a66592a,a66595a,a66596a,a66599a,a66602a,a66603a,a66604a,a66608a,a66609a,a66612a,a66615a,a66616a,a66617a,a66620a,a66623a,a66624a,a66627a,a66630a,a66631a,a66632a,a66636a,a66637a,a66640a,a66643a,a66644a,a66645a,a66648a,a66651a,a66652a,a66655a,a66658a,a66659a,a66660a,a66664a,a66665a,a66668a,a66671a,a66672a,a66673a,a66676a,a66679a,a66680a,a66683a,a66686a,a66687a,a66688a,a66692a,a66693a,a66696a,a66699a,a66700a,a66701a,a66704a,a66707a,a66708a,a66711a,a66714a,a66715a,a66716a,a66720a,a66721a,a66724a,a66727a,a66728a,a66729a,a66732a,a66735a,a66736a,a66739a,a66742a,a66743a,a66744a,a66748a,a66749a,a66752a,a66755a,a66756a,a66757a,a66760a,a66763a,a66764a,a66767a,a66770a,a66771a,a66772a,a66776a,a66777a,a66780a,a66783a,a66784a,a66785a,a66788a,a66791a,a66792a,a66795a,a66798a,a66799a,a66800a,a66804a,a66805a,a66808a,a66811a,a66812a,a66813a,a66816a,a66819a,a66820a,a66823a,a66826a,a66827a,a66828a,a66832a,a66833a,a66836a,a66839a,a66840a,a66841a,a66844a,a66847a,a66848a,a66851a,a66854a,a66855a,a66856a,a66860a,a66861a,a66864a,a66867a,a66868a,a66869a,a66872a,a66875a,a66876a,a66879a,a66882a,a66883a,a66884a,a66888a,a66889a,a66892a,a66895a,a66896a,a66897a,a66900a,a66903a,a66904a,a66907a,a66910a,a66911a,a66912a,a66916a,a66917a,a66920a,a66923a,a66924a,a66925a,a66928a,a66931a,a66932a,a66935a,a66938a,a66939a,a66940a,a66944a,a66945a,a66948a,a66951a,a66952a,a66953a,a66956a,a66959a,a66960a,a66963a,a66966a,a66967a,a66968a,a66972a,a66973a,a66976a,a66979a,a66980a,a66981a,a66984a,a66987a,a66988a,a66991a,a66994a,a66995a,a66996a,a67000a,a67001a,a67004a,a67007a,a67008a,a67009a,a67012a,a67015a,a67016a,a67019a,a67022a,a67023a,a67024a,a67028a,a67029a,a67032a,a67035a,a67036a,a67037a,a67040a,a67043a,a67044a,a67047a,a67050a,a67051a,a67052a,a67056a,a67057a,a67060a,a67063a,a67064a,a67065a,a67068a,a67071a,a67072a,a67075a,a67078a,a67079a,a67080a,a67084a,a67085a,a67088a,a67091a,a67092a,a67093a,a67096a,a67099a,a67100a,a67103a,a67106a,a67107a,a67108a,a67112a,a67113a,a67116a,a67119a,a67120a,a67121a,a67124a,a67127a,a67128a,a67131a,a67134a,a67135a,a67136a,a67140a,a67141a,a67144a,a67147a,a67148a,a67149a,a67152a,a67155a,a67156a,a67159a,a67162a,a67163a,a67164a,a67168a,a67169a,a67172a,a67175a,a67176a,a67177a,a67180a,a67183a,a67184a,a67187a,a67190a,a67191a,a67192a,a67196a,a67197a,a67200a,a67203a,a67204a,a67205a,a67208a,a67211a,a67212a,a67215a,a67218a,a67219a,a67220a,a67224a,a67225a,a67228a,a67231a,a67232a,a67233a,a67236a,a67239a,a67240a,a67243a,a67246a,a67247a,a67248a,a67252a,a67253a,a67256a,a67259a,a67260a,a67261a,a67264a,a67267a,a67268a,a67271a,a67274a,a67275a,a67276a,a67280a,a67281a,a67284a,a67287a,a67288a,a67289a,a67292a,a67295a,a67296a,a67299a,a67302a,a67303a,a67304a,a67308a,a67309a,a67312a,a67315a,a67316a,a67317a,a67320a,a67323a,a67324a,a67327a,a67330a,a67331a,a67332a,a67336a,a67337a,a67340a,a67343a,a67344a,a67345a,a67348a,a67351a,a67352a,a67355a,a67358a,a67359a,a67360a,a67364a,a67365a,a67368a,a67371a,a67372a,a67373a,a67376a,a67379a,a67380a,a67383a,a67386a,a67387a,a67388a,a67392a,a67393a,a67396a,a67399a,a67400a,a67401a,a67404a,a67407a,a67408a,a67411a,a67414a,a67415a,a67416a,a67420a,a67421a,a67424a,a67427a,a67428a,a67429a,a67432a,a67435a,a67436a,a67439a,a67442a,a67443a,a67444a,a67448a,a67449a,a67452a,a67455a,a67456a,a67457a,a67460a,a67463a,a67464a,a67467a,a67470a,a67471a,a67472a,a67476a,a67477a,a67480a,a67483a,a67484a,a67485a,a67488a,a67491a,a67492a,a67495a,a67498a,a67499a,a67500a,a67504a,a67505a,a67508a,a67511a,a67512a,a67513a,a67516a,a67519a,a67520a,a67523a,a67526a,a67527a,a67528a,a67532a,a67533a,a67536a,a67539a,a67540a,a67541a,a67544a,a67547a,a67548a,a67551a,a67554a,a67555a,a67556a,a67560a,a67561a,a67564a,a67567a,a67568a,a67569a,a67572a,a67575a,a67576a,a67579a,a67582a,a67583a,a67584a,a67588a,a67589a,a67592a,a67595a,a67596a,a67597a,a67600a,a67603a,a67604a,a67607a,a67610a,a67611a,a67612a,a67616a,a67617a,a67620a,a67623a,a67624a,a67625a,a67628a,a67631a,a67632a,a67635a,a67638a,a67639a,a67640a,a67644a,a67645a,a67648a,a67651a,a67652a,a67653a,a67656a,a67659a,a67660a,a67663a,a67666a,a67667a,a67668a,a67672a,a67673a,a67676a,a67679a,a67680a,a67681a,a67684a,a67687a,a67688a,a67691a,a67694a,a67695a,a67696a,a67700a,a67701a,a67704a,a67707a,a67708a,a67709a,a67712a,a67715a,a67716a,a67719a,a67722a,a67723a,a67724a,a67728a,a67729a,a67732a,a67735a,a67736a,a67737a,a67740a,a67743a,a67744a,a67747a,a67750a,a67751a,a67752a,a67756a,a67757a,a67760a,a67763a,a67764a,a67765a,a67768a,a67771a,a67772a,a67775a,a67778a,a67779a,a67780a,a67784a,a67785a,a67788a,a67791a,a67792a,a67793a,a67796a,a67799a,a67800a,a67803a,a67806a,a67807a,a67808a,a67812a,a67813a,a67816a,a67819a,a67820a,a67821a,a67824a,a67827a,a67828a,a67831a,a67834a,a67835a,a67836a,a67840a,a67841a,a67844a,a67847a,a67848a,a67849a,a67852a,a67855a,a67856a,a67859a,a67862a,a67863a,a67864a,a67868a,a67869a,a67872a,a67875a,a67876a,a67877a,a67880a,a67883a,a67884a,a67887a,a67890a,a67891a,a67892a,a67896a,a67897a,a67900a,a67903a,a67904a,a67905a,a67908a,a67911a,a67912a,a67915a,a67918a,a67919a,a67920a,a67924a,a67925a,a67928a,a67931a,a67932a,a67933a,a67936a,a67939a,a67940a,a67943a,a67946a,a67947a,a67948a,a67952a,a67953a,a67956a,a67959a,a67960a,a67961a,a67964a,a67967a,a67968a,a67971a,a67974a,a67975a,a67976a,a67980a,a67981a,a67984a,a67987a,a67988a,a67989a,a67992a,a67995a,a67996a,a67999a,a68002a,a68003a,a68004a,a68008a,a68009a,a68012a,a68015a,a68016a,a68017a,a68020a,a68023a,a68024a,a68027a,a68030a,a68031a,a68032a,a68036a,a68037a,a68040a,a68043a,a68044a,a68045a,a68048a,a68051a,a68052a,a68055a,a68058a,a68059a,a68060a,a68064a,a68065a,a68068a,a68071a,a68072a,a68073a,a68076a,a68079a,a68080a,a68083a,a68086a,a68087a,a68088a,a68092a,a68093a,a68096a,a68099a,a68100a,a68101a,a68104a,a68107a,a68108a,a68111a,a68114a,a68115a,a68116a,a68120a,a68121a,a68124a,a68127a,a68128a,a68129a,a68132a,a68135a,a68136a,a68139a,a68142a,a68143a,a68144a,a68148a,a68149a,a68152a,a68155a,a68156a,a68157a,a68160a,a68163a,a68164a,a68167a,a68170a,a68171a,a68172a,a68176a,a68177a,a68180a,a68183a,a68184a,a68185a,a68188a,a68191a,a68192a,a68195a,a68198a,a68199a,a68200a,a68204a,a68205a,a68208a,a68211a,a68212a,a68213a,a68216a,a68219a,a68220a,a68223a,a68226a,a68227a,a68228a,a68232a,a68233a,a68236a,a68239a,a68240a,a68241a,a68244a,a68247a,a68248a,a68251a,a68254a,a68255a,a68256a,a68260a,a68261a,a68264a,a68267a,a68268a,a68269a,a68272a,a68275a,a68276a,a68279a,a68282a,a68283a,a68284a,a68288a,a68289a,a68292a,a68295a,a68296a,a68297a,a68300a,a68303a,a68304a,a68307a,a68310a,a68311a,a68312a,a68316a,a68317a,a68320a,a68323a,a68324a,a68325a,a68328a,a68331a,a68332a,a68335a,a68338a,a68339a,a68340a,a68344a,a68345a,a68348a,a68351a,a68352a,a68353a,a68356a,a68359a,a68360a,a68363a,a68366a,a68367a,a68368a,a68372a,a68373a,a68376a,a68379a,a68380a,a68381a,a68384a,a68387a,a68388a,a68391a,a68394a,a68395a,a68396a,a68400a,a68401a,a68404a,a68407a,a68408a,a68409a,a68412a,a68415a,a68416a,a68419a,a68422a,a68423a,a68424a,a68428a,a68429a,a68432a,a68435a,a68436a,a68437a,a68440a,a68443a,a68444a,a68447a,a68450a,a68451a,a68452a,a68456a,a68457a,a68460a,a68463a,a68464a,a68465a,a68468a,a68471a,a68472a,a68475a,a68478a,a68479a,a68480a,a68484a,a68485a,a68488a,a68491a,a68492a,a68493a,a68496a,a68499a,a68500a,a68503a,a68506a,a68507a,a68508a,a68512a,a68513a,a68516a,a68519a,a68520a,a68521a,a68524a,a68527a,a68528a,a68531a,a68534a,a68535a,a68536a,a68540a,a68541a,a68544a,a68547a,a68548a,a68549a,a68552a,a68555a,a68556a,a68559a,a68562a,a68563a,a68564a,a68568a,a68569a,a68572a,a68575a,a68576a,a68577a,a68580a,a68583a,a68584a,a68587a,a68590a,a68591a,a68592a,a68596a,a68597a,a68600a,a68603a,a68604a,a68605a,a68608a,a68611a,a68612a,a68615a,a68618a,a68619a,a68620a,a68624a,a68625a,a68628a,a68631a,a68632a,a68633a,a68636a,a68639a,a68640a,a68643a,a68646a,a68647a,a68648a,a68652a,a68653a,a68656a,a68659a,a68660a,a68661a,a68664a,a68667a,a68668a,a68671a,a68674a,a68675a,a68676a,a68680a,a68681a,a68684a,a68687a,a68688a,a68689a,a68692a,a68695a,a68696a,a68699a,a68702a,a68703a,a68704a,a68708a,a68709a,a68712a,a68715a,a68716a,a68717a,a68720a,a68723a,a68724a,a68727a,a68730a,a68731a,a68732a,a68736a,a68737a,a68740a,a68743a,a68744a,a68745a,a68748a,a68751a,a68752a,a68755a,a68758a,a68759a,a68760a,a68764a,a68765a,a68768a,a68771a,a68772a,a68773a,a68776a,a68779a,a68780a,a68783a,a68786a,a68787a,a68788a,a68792a,a68793a,a68796a,a68799a,a68800a,a68801a,a68804a,a68807a,a68808a,a68811a,a68814a,a68815a,a68816a,a68820a,a68821a,a68824a,a68827a,a68828a,a68829a,a68832a,a68835a,a68836a,a68839a,a68842a,a68843a,a68844a,a68848a,a68849a,a68852a,a68855a,a68856a,a68857a,a68860a,a68863a,a68864a,a68867a,a68870a,a68871a,a68872a,a68876a,a68877a,a68880a,a68883a,a68884a,a68885a,a68888a,a68891a,a68892a,a68895a,a68898a,a68899a,a68900a,a68904a,a68905a,a68908a,a68911a,a68912a,a68913a,a68916a,a68919a,a68920a,a68923a,a68926a,a68927a,a68928a,a68932a,a68933a,a68936a,a68939a,a68940a,a68941a,a68944a,a68947a,a68948a,a68951a,a68954a,a68955a,a68956a,a68960a,a68961a,a68964a,a68967a,a68968a,a68969a,a68972a,a68975a,a68976a,a68979a,a68982a,a68983a,a68984a,a68988a,a68989a,a68992a,a68995a,a68996a,a68997a,a69000a,a69003a,a69004a,a69007a,a69010a,a69011a,a69012a,a69016a,a69017a,a69020a,a69023a,a69024a,a69025a,a69028a,a69031a,a69032a,a69035a,a69038a,a69039a,a69040a,a69044a,a69045a,a69048a,a69051a,a69052a,a69053a,a69056a,a69059a,a69060a,a69063a,a69066a,a69067a,a69068a,a69072a,a69073a,a69076a,a69079a,a69080a,a69081a,a69084a,a69087a,a69088a,a69091a,a69094a,a69095a,a69096a,a69100a,a69101a,a69104a,a69107a,a69108a,a69109a,a69112a,a69115a,a69116a,a69119a,a69122a,a69123a,a69124a,a69128a,a69129a,a69132a,a69135a,a69136a,a69137a,a69140a,a69143a,a69144a,a69147a,a69150a,a69151a,a69152a,a69156a,a69157a,a69160a,a69163a,a69164a,a69165a,a69168a,a69171a,a69172a,a69175a,a69178a,a69179a,a69180a,a69184a,a69185a,a69188a,a69191a,a69192a,a69193a,a69196a,a69199a,a69200a,a69203a,a69206a,a69207a,a69208a,a69212a,a69213a,a69216a,a69219a,a69220a,a69221a,a69224a,a69227a,a69228a,a69231a,a69234a,a69235a,a69236a,a69240a,a69241a,a69244a,a69247a,a69248a,a69249a,a69252a,a69255a,a69256a,a69259a,a69262a,a69263a,a69264a,a69268a,a69269a,a69272a,a69275a,a69276a,a69277a,a69280a,a69283a,a69284a,a69287a,a69290a,a69291a,a69292a,a69296a,a69297a,a69300a,a69303a,a69304a,a69305a,a69308a,a69311a,a69312a,a69315a,a69318a,a69319a,a69320a,a69324a,a69325a,a69328a,a69331a,a69332a,a69333a,a69336a,a69339a,a69340a,a69343a,a69346a,a69347a,a69348a,a69352a,a69353a,a69356a,a69359a,a69360a,a69361a,a69364a,a69367a,a69368a,a69371a,a69374a,a69375a,a69376a,a69380a,a69381a,a69384a,a69387a,a69388a,a69389a,a69392a,a69395a,a69396a,a69399a,a69402a,a69403a,a69404a,a69408a,a69409a,a69412a,a69415a,a69416a,a69417a,a69420a,a69423a,a69424a,a69427a,a69430a,a69431a,a69432a,a69436a,a69437a,a69440a,a69443a,a69444a,a69445a,a69448a,a69451a,a69452a,a69455a,a69458a,a69459a,a69460a,a69464a,a69465a,a69468a,a69471a,a69472a,a69473a,a69476a,a69479a,a69480a,a69483a,a69486a,a69487a,a69488a,a69492a,a69493a,a69496a,a69499a,a69500a,a69501a,a69504a,a69507a,a69508a,a69511a,a69514a,a69515a,a69516a,a69520a,a69521a,a69524a,a69527a,a69528a,a69529a,a69532a,a69535a,a69536a,a69539a,a69542a,a69543a,a69544a,a69548a,a69549a,a69552a,a69555a,a69556a,a69557a,a69560a,a69563a,a69564a,a69567a,a69570a,a69571a,a69572a,a69576a,a69577a,a69580a,a69583a,a69584a,a69585a,a69588a,a69591a,a69592a,a69595a,a69598a,a69599a,a69600a,a69604a,a69605a,a69608a,a69611a,a69612a,a69613a,a69616a,a69619a,a69620a,a69623a,a69626a,a69627a,a69628a,a69632a,a69633a,a69636a,a69639a,a69640a,a69641a,a69644a,a69647a,a69648a,a69651a,a69654a,a69655a,a69656a,a69660a,a69661a,a69664a,a69667a,a69668a,a69669a,a69672a,a69675a,a69676a,a69679a,a69682a,a69683a,a69684a,a69688a,a69689a,a69692a,a69695a,a69696a,a69697a,a69700a,a69703a,a69704a,a69707a,a69710a,a69711a,a69712a,a69716a,a69717a,a69720a,a69723a,a69724a,a69725a,a69728a,a69731a,a69732a,a69735a,a69738a,a69739a,a69740a,a69744a,a69745a,a69748a,a69751a,a69752a,a69753a,a69756a,a69759a,a69760a,a69763a,a69766a,a69767a,a69768a,a69772a,a69773a,a69776a,a69779a,a69780a,a69781a,a69784a,a69787a,a69788a,a69791a,a69794a,a69795a,a69796a,a69800a,a69801a,a69804a,a69807a,a69808a,a69809a,a69812a,a69815a,a69816a,a69819a,a69822a,a69823a,a69824a,a69828a,a69829a,a69832a,a69835a,a69836a,a69837a,a69840a,a69843a,a69844a,a69847a,a69850a,a69851a,a69852a,a69856a,a69857a,a69860a,a69863a,a69864a,a69865a,a69868a,a69871a,a69872a,a69875a,a69878a,a69879a,a69880a,a69884a,a69885a,a69888a,a69891a,a69892a,a69893a,a69896a,a69899a,a69900a,a69903a,a69906a,a69907a,a69908a,a69912a,a69913a,a69916a,a69919a,a69920a,a69921a,a69924a,a69927a,a69928a,a69931a,a69934a,a69935a,a69936a,a69940a,a69941a,a69944a,a69947a,a69948a,a69949a,a69952a,a69955a,a69956a,a69959a,a69962a,a69963a,a69964a,a69968a,a69969a,a69972a,a69975a,a69976a,a69977a,a69980a,a69983a,a69984a,a69987a,a69990a,a69991a,a69992a,a69996a,a69997a,a70000a,a70003a,a70004a,a70005a,a70008a,a70011a,a70012a,a70015a,a70018a,a70019a,a70020a,a70024a,a70025a,a70028a,a70031a,a70032a,a70033a,a70036a,a70039a,a70040a,a70043a,a70046a,a70047a,a70048a,a70052a,a70053a,a70056a,a70059a,a70060a,a70061a,a70064a,a70067a,a70068a,a70071a,a70074a,a70075a,a70076a,a70080a,a70081a,a70084a,a70087a,a70088a,a70089a,a70092a,a70095a,a70096a,a70099a,a70102a,a70103a,a70104a,a70108a,a70109a,a70112a,a70115a,a70116a,a70117a,a70120a,a70123a,a70124a,a70127a,a70130a,a70131a,a70132a,a70136a,a70137a,a70140a,a70143a,a70144a,a70145a,a70148a,a70151a,a70152a,a70155a,a70158a,a70159a,a70160a,a70164a,a70165a,a70168a,a70171a,a70172a,a70173a,a70176a,a70179a,a70180a,a70183a,a70186a,a70187a,a70188a,a70192a,a70193a,a70196a,a70199a,a70200a,a70201a,a70204a,a70207a,a70208a,a70211a,a70214a,a70215a,a70216a,a70220a,a70221a,a70224a,a70227a,a70228a,a70229a,a70232a,a70235a,a70236a,a70239a,a70242a,a70243a,a70244a,a70248a,a70249a,a70252a,a70255a,a70256a,a70257a,a70260a,a70263a,a70264a,a70267a,a70270a,a70271a,a70272a,a70276a,a70277a,a70280a,a70283a,a70284a,a70285a,a70288a,a70291a,a70292a,a70295a,a70298a,a70299a,a70300a,a70304a,a70305a,a70308a,a70311a,a70312a,a70313a,a70316a,a70319a,a70320a,a70323a,a70326a,a70327a,a70328a,a70332a,a70333a,a70336a,a70339a,a70340a,a70341a,a70344a,a70347a,a70348a,a70351a,a70354a,a70355a,a70356a,a70360a,a70361a,a70364a,a70367a,a70368a,a70369a,a70372a,a70375a,a70376a,a70379a,a70382a,a70383a,a70384a,a70388a,a70389a,a70392a,a70395a,a70396a,a70397a,a70400a,a70403a,a70404a,a70407a,a70410a,a70411a,a70412a,a70416a,a70417a,a70420a,a70423a,a70424a,a70425a,a70428a,a70431a,a70432a,a70435a,a70438a,a70439a,a70440a,a70444a,a70445a,a70448a,a70451a,a70452a,a70453a,a70456a,a70459a,a70460a,a70463a,a70466a,a70467a,a70468a,a70472a,a70473a,a70476a,a70479a,a70480a,a70481a,a70484a,a70487a,a70488a,a70491a,a70494a,a70495a,a70496a,a70500a,a70501a,a70504a,a70507a,a70508a,a70509a,a70512a,a70515a,a70516a,a70519a,a70522a,a70523a,a70524a,a70528a,a70529a,a70532a,a70535a,a70536a,a70537a,a70540a,a70543a,a70544a,a70547a,a70550a,a70551a,a70552a,a70556a,a70557a,a70560a,a70563a,a70564a,a70565a,a70568a,a70571a,a70572a,a70575a,a70578a,a70579a,a70580a,a70584a,a70585a,a70588a,a70591a,a70592a,a70593a,a70596a,a70599a,a70600a,a70603a,a70606a,a70607a,a70608a,a70612a,a70613a,a70616a,a70619a,a70620a,a70621a,a70624a,a70627a,a70628a,a70631a,a70634a,a70635a,a70636a,a70640a,a70641a,a70644a,a70647a,a70648a,a70649a,a70652a,a70655a,a70656a,a70659a,a70662a,a70663a,a70664a,a70668a,a70669a,a70672a,a70675a,a70676a,a70677a,a70680a,a70683a,a70684a,a70687a,a70690a,a70691a,a70692a,a70696a,a70697a,a70700a,a70703a,a70704a,a70705a,a70708a,a70711a,a70712a,a70715a,a70718a,a70719a,a70720a,a70724a,a70725a,a70728a,a70731a,a70732a,a70733a,a70736a,a70739a,a70740a,a70743a,a70746a,a70747a,a70748a,a70752a,a70753a,a70756a,a70759a,a70760a,a70761a,a70764a,a70767a,a70768a,a70771a,a70774a,a70775a,a70776a,a70780a,a70781a,a70784a,a70787a,a70788a,a70789a,a70792a,a70795a,a70796a,a70799a,a70802a,a70803a,a70804a,a70808a,a70809a,a70812a,a70815a,a70816a,a70817a,a70820a,a70823a,a70824a,a70827a,a70830a,a70831a,a70832a,a70836a,a70837a,a70840a,a70843a,a70844a,a70845a,a70848a,a70851a,a70852a,a70855a,a70858a,a70859a,a70860a,a70864a,a70865a,a70868a,a70871a,a70872a,a70873a,a70876a,a70879a,a70880a,a70883a,a70886a,a70887a,a70888a,a70892a,a70893a,a70896a,a70899a,a70900a,a70901a,a70904a,a70907a,a70908a,a70911a,a70914a,a70915a,a70916a,a70920a,a70921a,a70924a,a70927a,a70928a,a70929a,a70932a,a70935a,a70936a,a70939a,a70942a,a70943a,a70944a,a70948a,a70949a,a70952a,a70955a,a70956a,a70957a,a70960a,a70963a,a70964a,a70967a,a70970a,a70971a,a70972a,a70976a,a70977a,a70980a,a70983a,a70984a,a70985a,a70988a,a70991a,a70992a,a70995a,a70998a,a70999a,a71000a,a71004a,a71005a,a71008a,a71011a,a71012a,a71013a,a71016a,a71019a,a71020a,a71023a,a71026a,a71027a,a71028a,a71032a,a71033a,a71036a,a71039a,a71040a,a71041a,a71044a,a71047a,a71048a,a71051a,a71054a,a71055a,a71056a,a71060a,a71061a,a71064a,a71067a,a71068a,a71069a,a71072a,a71075a,a71076a,a71079a,a71082a,a71083a,a71084a,a71088a,a71089a,a71092a,a71095a,a71096a,a71097a,a71100a,a71103a,a71104a,a71107a,a71110a,a71111a,a71112a,a71116a,a71117a,a71120a,a71123a,a71124a,a71125a,a71128a,a71131a,a71132a,a71135a,a71138a,a71139a,a71140a,a71144a,a71145a,a71148a,a71151a,a71152a,a71153a,a71156a,a71159a,a71160a,a71163a,a71166a,a71167a,a71168a,a71172a,a71173a,a71176a,a71179a,a71180a,a71181a,a71184a,a71187a,a71188a,a71191a,a71194a,a71195a,a71196a,a71200a,a71201a,a71204a,a71207a,a71208a,a71209a,a71212a,a71215a,a71216a,a71219a,a71222a,a71223a,a71224a,a71228a,a71229a,a71232a,a71235a,a71236a,a71237a,a71240a,a71243a,a71244a,a71247a,a71250a,a71251a,a71252a,a71256a,a71257a,a71260a,a71263a,a71264a,a71265a,a71268a,a71271a,a71272a,a71275a,a71278a,a71279a,a71280a,a71284a,a71285a,a71288a,a71291a,a71292a,a71293a,a71296a,a71299a,a71300a,a71303a,a71306a,a71307a,a71308a,a71312a,a71313a,a71316a,a71319a,a71320a,a71321a,a71324a,a71327a,a71328a,a71331a,a71334a,a71335a,a71336a,a71340a,a71341a,a71344a,a71347a,a71348a,a71349a,a71352a,a71355a,a71356a,a71359a,a71362a,a71363a,a71364a,a71368a,a71369a,a71372a,a71375a,a71376a,a71377a,a71380a,a71383a,a71384a,a71387a,a71390a,a71391a,a71392a,a71396a,a71397a,a71400a,a71403a,a71404a,a71405a,a71408a,a71411a,a71412a,a71415a,a71418a,a71419a,a71420a,a71424a,a71425a,a71428a,a71431a,a71432a,a71433a,a71436a,a71439a,a71440a,a71443a,a71446a,a71447a,a71448a,a71452a,a71453a,a71456a,a71459a,a71460a,a71461a,a71464a,a71467a,a71468a,a71471a,a71474a,a71475a,a71476a,a71480a,a71481a,a71484a,a71487a,a71488a,a71489a,a71492a,a71495a,a71496a,a71499a,a71502a,a71503a,a71504a,a71508a,a71509a,a71512a,a71515a,a71516a,a71517a,a71520a,a71523a,a71524a,a71527a,a71530a,a71531a,a71532a,a71536a,a71537a,a71540a,a71543a,a71544a,a71545a,a71548a,a71551a,a71552a,a71555a,a71558a,a71559a,a71560a,a71564a,a71565a,a71568a,a71571a,a71572a,a71573a,a71576a,a71579a,a71580a,a71583a,a71586a,a71587a,a71588a,a71592a,a71593a,a71596a,a71599a,a71600a,a71601a,a71604a,a71607a,a71608a,a71611a,a71614a,a71615a,a71616a,a71620a,a71621a,a71624a,a71627a,a71628a,a71629a,a71632a,a71635a,a71636a,a71639a,a71642a,a71643a,a71644a,a71648a,a71649a,a71652a,a71655a,a71656a,a71657a,a71660a,a71663a,a71664a,a71667a,a71670a,a71671a,a71672a,a71676a,a71677a,a71680a,a71683a,a71684a,a71685a,a71688a,a71691a,a71692a,a71695a,a71698a,a71699a,a71700a,a71704a,a71705a,a71708a,a71711a,a71712a,a71713a,a71716a,a71719a,a71720a,a71723a,a71726a,a71727a,a71728a,a71732a,a71733a,a71736a,a71739a,a71740a,a71741a,a71744a,a71747a,a71748a,a71751a,a71754a,a71755a,a71756a,a71760a,a71761a,a71764a,a71767a,a71768a,a71769a,a71772a,a71775a,a71776a,a71779a,a71782a,a71783a,a71784a,a71788a,a71789a,a71792a,a71795a,a71796a,a71797a,a71800a,a71803a,a71804a,a71807a,a71810a,a71811a,a71812a,a71816a,a71817a,a71820a,a71823a,a71824a,a71825a,a71828a,a71831a,a71832a,a71835a,a71838a,a71839a,a71840a,a71844a,a71845a,a71848a,a71851a,a71852a,a71853a,a71856a,a71859a,a71860a,a71863a,a71866a,a71867a,a71868a,a71872a,a71873a,a71876a,a71879a,a71880a,a71881a,a71884a,a71887a,a71888a,a71891a,a71894a,a71895a,a71896a,a71900a,a71901a,a71904a,a71907a,a71908a,a71909a,a71912a,a71915a,a71916a,a71919a,a71922a,a71923a,a71924a,a71928a,a71929a,a71932a,a71935a,a71936a,a71937a,a71940a,a71943a,a71944a,a71947a,a71950a,a71951a,a71952a,a71956a,a71957a,a71960a,a71963a,a71964a,a71965a,a71968a,a71971a,a71972a,a71975a,a71978a,a71979a,a71980a,a71984a,a71985a,a71988a,a71991a,a71992a,a71993a,a71996a,a71999a,a72000a,a72003a,a72006a,a72007a,a72008a,a72012a,a72013a,a72016a,a72019a,a72020a,a72021a,a72024a,a72027a,a72028a,a72031a,a72034a,a72035a,a72036a,a72040a,a72041a,a72044a,a72047a,a72048a,a72049a,a72052a,a72055a,a72056a,a72059a,a72062a,a72063a,a72064a,a72068a,a72069a,a72072a,a72075a,a72076a,a72077a,a72080a,a72083a,a72084a,a72087a,a72090a,a72091a,a72092a,a72096a,a72097a,a72100a,a72103a,a72104a,a72105a,a72108a,a72111a,a72112a,a72115a,a72118a,a72119a,a72120a,a72124a,a72125a,a72128a,a72131a,a72132a,a72133a,a72136a,a72139a,a72140a,a72143a,a72146a,a72147a,a72148a,a72152a,a72153a,a72156a,a72159a,a72160a,a72161a,a72164a,a72167a,a72168a,a72171a,a72174a,a72175a,a72176a,a72180a,a72181a,a72184a,a72187a,a72188a,a72189a,a72192a,a72195a,a72196a,a72199a,a72202a,a72203a,a72204a,a72208a,a72209a,a72212a,a72215a,a72216a,a72217a,a72220a,a72223a,a72224a,a72227a,a72230a,a72231a,a72232a,a72236a,a72237a,a72240a,a72243a,a72244a,a72245a,a72248a,a72251a,a72252a,a72255a,a72258a,a72259a,a72260a,a72264a,a72265a,a72268a,a72271a,a72272a,a72273a,a72276a,a72279a,a72280a,a72283a,a72286a,a72287a,a72288a,a72292a,a72293a,a72296a,a72299a,a72300a,a72301a,a72304a,a72307a,a72308a,a72311a,a72314a,a72315a,a72316a,a72320a,a72321a,a72324a,a72327a,a72328a,a72329a,a72332a,a72335a,a72336a,a72339a,a72342a,a72343a,a72344a,a72348a,a72349a,a72352a,a72355a,a72356a,a72357a,a72360a,a72363a,a72364a,a72367a,a72370a,a72371a,a72372a,a72376a,a72377a,a72380a,a72383a,a72384a,a72385a,a72388a,a72391a,a72392a,a72395a,a72398a,a72399a,a72400a,a72404a,a72405a,a72408a,a72411a,a72412a,a72413a,a72416a,a72419a,a72420a,a72423a,a72426a,a72427a,a72428a,a72432a,a72433a,a72436a,a72439a,a72440a,a72441a,a72444a,a72447a,a72448a,a72451a,a72454a,a72455a,a72456a,a72460a,a72461a,a72464a,a72467a,a72468a,a72469a,a72472a,a72475a,a72476a,a72479a,a72482a,a72483a,a72484a,a72488a,a72489a,a72492a,a72495a,a72496a,a72497a,a72500a,a72503a,a72504a,a72507a,a72510a,a72511a,a72512a,a72516a,a72517a,a72520a,a72523a,a72524a,a72525a,a72528a,a72531a,a72532a,a72535a,a72538a,a72539a,a72540a,a72544a,a72545a,a72548a,a72551a,a72552a,a72553a,a72556a,a72559a,a72560a,a72563a,a72566a,a72567a,a72568a,a72572a,a72573a,a72576a,a72579a,a72580a,a72581a,a72584a,a72587a,a72588a,a72591a,a72594a,a72595a,a72596a,a72600a,a72601a,a72604a,a72607a,a72608a,a72609a,a72612a,a72615a,a72616a,a72619a,a72622a,a72623a,a72624a,a72628a,a72629a,a72632a,a72635a,a72636a,a72637a,a72640a,a72643a,a72644a,a72647a,a72650a,a72651a,a72652a,a72656a,a72657a,a72660a,a72663a,a72664a,a72665a,a72668a,a72671a,a72672a,a72675a,a72678a,a72679a,a72680a,a72684a,a72685a,a72688a,a72691a,a72692a,a72693a,a72696a,a72699a,a72700a,a72703a,a72706a,a72707a,a72708a,a72712a,a72713a,a72716a,a72719a,a72720a,a72721a,a72724a,a72727a,a72728a,a72731a,a72734a,a72735a,a72736a,a72740a,a72741a,a72744a,a72747a,a72748a,a72749a,a72752a,a72755a,a72756a,a72759a,a72762a,a72763a,a72764a,a72768a,a72769a,a72772a,a72775a,a72776a,a72777a,a72780a,a72783a,a72784a,a72787a,a72790a,a72791a,a72792a,a72796a,a72797a,a72800a,a72803a,a72804a,a72805a,a72808a,a72811a,a72812a,a72815a,a72818a,a72819a,a72820a,a72824a,a72825a,a72828a,a72831a,a72832a,a72833a,a72836a,a72839a,a72840a,a72843a,a72846a,a72847a,a72848a,a72852a,a72853a,a72856a,a72859a,a72860a,a72861a,a72864a,a72867a,a72868a,a72871a,a72874a,a72875a,a72876a,a72880a,a72881a,a72884a,a72887a,a72888a,a72889a,a72892a,a72895a,a72896a,a72899a,a72902a,a72903a,a72904a,a72908a,a72909a,a72912a,a72915a,a72916a,a72917a,a72920a,a72923a,a72924a,a72927a,a72930a,a72931a,a72932a,a72936a,a72937a,a72940a,a72943a,a72944a,a72945a,a72948a,a72951a,a72952a,a72955a,a72958a,a72959a,a72960a,a72964a,a72965a,a72968a,a72971a,a72972a,a72973a,a72976a,a72979a,a72980a,a72983a,a72986a,a72987a,a72988a,a72992a,a72993a,a72996a,a72999a,a73000a,a73001a,a73004a,a73007a,a73008a,a73011a,a73014a,a73015a,a73016a,a73020a,a73021a,a73024a,a73027a,a73028a,a73029a,a73032a,a73035a,a73036a,a73039a,a73042a,a73043a,a73044a,a73048a,a73049a,a73052a,a73055a,a73056a,a73057a,a73060a,a73063a,a73064a,a73067a,a73070a,a73071a,a73072a,a73076a,a73077a,a73080a,a73083a,a73084a,a73085a,a73088a,a73091a,a73092a,a73095a,a73098a,a73099a,a73100a,a73104a,a73105a,a73108a,a73111a,a73112a,a73113a,a73116a,a73119a,a73120a,a73123a,a73126a,a73127a,a73128a,a73132a,a73133a,a73136a,a73139a,a73140a,a73141a,a73144a,a73147a,a73148a,a73151a,a73154a,a73155a,a73156a,a73160a,a73161a,a73164a,a73167a,a73168a,a73169a,a73172a,a73175a,a73176a,a73179a,a73182a,a73183a,a73184a,a73188a,a73189a,a73192a,a73195a,a73196a,a73197a,a73200a,a73203a,a73204a,a73207a,a73210a,a73211a,a73212a,a73216a,a73217a,a73220a,a73223a,a73224a,a73225a,a73228a,a73231a,a73232a,a73235a,a73238a,a73239a,a73240a,a73244a,a73245a,a73248a,a73251a,a73252a,a73253a,a73256a,a73259a,a73260a,a73263a,a73266a,a73267a,a73268a,a73272a,a73273a,a73276a,a73279a,a73280a,a73281a,a73284a,a73287a,a73288a,a73291a,a73294a,a73295a,a73296a,a73300a,a73301a,a73304a,a73307a,a73308a,a73309a,a73312a,a73315a,a73316a,a73319a,a73322a,a73323a,a73324a,a73328a,a73329a,a73332a,a73335a,a73336a,a73337a,a73340a,a73343a,a73344a,a73347a,a73350a,a73351a,a73352a,a73356a,a73357a,a73360a,a73363a,a73364a,a73365a,a73368a,a73371a,a73372a,a73375a,a73378a,a73379a,a73380a,a73384a,a73385a,a73388a,a73391a,a73392a,a73393a,a73396a,a73399a,a73400a,a73403a,a73406a,a73407a,a73408a,a73412a,a73413a,a73416a,a73419a,a73420a,a73421a,a73424a,a73427a,a73428a,a73431a,a73434a,a73435a,a73436a,a73440a,a73441a,a73444a,a73447a,a73448a,a73449a,a73452a,a73455a,a73456a,a73459a,a73462a,a73463a,a73464a,a73468a,a73469a,a73472a,a73475a,a73476a,a73477a,a73480a,a73483a,a73484a,a73487a,a73490a,a73491a,a73492a,a73496a,a73497a,a73500a,a73503a,a73504a,a73505a,a73508a,a73511a,a73512a,a73515a,a73518a,a73519a,a73520a,a73524a,a73525a,a73528a,a73531a,a73532a,a73533a,a73536a,a73539a,a73540a,a73543a,a73546a,a73547a,a73548a,a73552a,a73553a,a73556a,a73559a,a73560a,a73561a,a73564a,a73567a,a73568a,a73571a,a73574a,a73575a,a73576a,a73580a,a73581a,a73584a,a73587a,a73588a,a73589a,a73592a,a73595a,a73596a,a73599a,a73602a,a73603a,a73604a,a73608a,a73609a,a73612a,a73615a,a73616a,a73617a,a73620a,a73623a,a73624a,a73627a,a73630a,a73631a,a73632a,a73636a,a73637a,a73640a,a73643a,a73644a,a73645a,a73648a,a73651a,a73652a,a73655a,a73658a,a73659a,a73660a,a73664a,a73665a,a73668a,a73671a,a73672a,a73673a,a73676a,a73679a,a73680a,a73683a,a73686a,a73687a,a73688a,a73692a,a73693a,a73696a,a73699a,a73700a,a73701a,a73704a,a73707a,a73708a,a73711a,a73714a,a73715a,a73716a,a73720a,a73721a,a73724a,a73727a,a73728a,a73729a,a73732a,a73735a,a73736a,a73739a,a73742a,a73743a,a73744a,a73748a,a73749a,a73752a,a73755a,a73756a,a73757a,a73760a,a73763a,a73764a,a73767a,a73770a,a73771a,a73772a,a73776a,a73777a,a73780a,a73783a,a73784a,a73785a,a73788a,a73791a,a73792a,a73795a,a73798a,a73799a,a73800a,a73804a,a73805a,a73808a,a73811a,a73812a,a73813a,a73816a,a73819a,a73820a,a73823a,a73826a,a73827a,a73828a,a73832a,a73833a,a73836a,a73839a,a73840a,a73841a,a73844a,a73847a,a73848a,a73851a,a73854a,a73855a,a73856a,a73860a,a73861a,a73864a,a73867a,a73868a,a73869a,a73872a,a73875a,a73876a,a73879a,a73882a,a73883a,a73884a,a73888a,a73889a,a73892a,a73895a,a73896a,a73897a,a73900a,a73903a,a73904a,a73907a,a73910a,a73911a,a73912a,a73916a,a73917a,a73920a,a73923a,a73924a,a73925a,a73928a,a73931a,a73932a,a73935a,a73938a,a73939a,a73940a,a73944a,a73945a,a73948a,a73951a,a73952a,a73953a,a73956a,a73959a,a73960a,a73963a,a73966a,a73967a,a73968a,a73972a,a73973a,a73976a,a73979a,a73980a,a73981a,a73984a,a73987a,a73988a,a73991a,a73994a,a73995a,a73996a,a74000a,a74001a,a74004a,a74007a,a74008a,a74009a,a74012a,a74015a,a74016a,a74019a,a74022a,a74023a,a74024a,a74028a,a74029a,a74032a,a74035a,a74036a,a74037a,a74040a,a74043a,a74044a,a74047a,a74050a,a74051a,a74052a,a74056a,a74057a,a74060a,a74063a,a74064a,a74065a,a74068a,a74071a,a74072a,a74075a,a74078a,a74079a,a74080a,a74084a,a74085a,a74088a,a74091a,a74092a,a74093a,a74096a,a74099a,a74100a,a74103a,a74106a,a74107a,a74108a,a74112a,a74113a,a74116a,a74119a,a74120a,a74121a,a74124a,a74127a,a74128a,a74131a,a74134a,a74135a,a74136a,a74140a,a74141a,a74144a,a74147a,a74148a,a74149a,a74152a,a74155a,a74156a,a74159a,a74162a,a74163a,a74164a,a74168a,a74169a,a74172a,a74175a,a74176a,a74177a,a74180a,a74183a,a74184a,a74187a,a74190a,a74191a,a74192a,a74196a,a74197a,a74200a,a74203a,a74204a,a74205a,a74208a,a74211a,a74212a,a74215a,a74218a,a74219a,a74220a,a74224a,a74225a,a74228a,a74231a,a74232a,a74233a,a74236a,a74239a,a74240a,a74243a,a74246a,a74247a,a74248a,a74252a,a74253a,a74256a,a74259a,a74260a,a74261a,a74264a,a74267a,a74268a,a74271a,a74274a,a74275a,a74276a,a74280a,a74281a,a74284a,a74287a,a74288a,a74289a,a74292a,a74295a,a74296a,a74299a,a74302a,a74303a,a74304a,a74308a,a74309a,a74312a,a74315a,a74316a,a74317a,a74320a,a74323a,a74324a,a74327a,a74330a,a74331a,a74332a,a74336a,a74337a,a74340a,a74343a,a74344a,a74345a,a74348a,a74351a,a74352a,a74355a,a74358a,a74359a,a74360a,a74364a,a74365a,a74368a,a74371a,a74372a,a74373a,a74376a,a74379a,a74380a,a74383a,a74386a,a74387a,a74388a,a74392a,a74393a,a74396a,a74399a,a74400a,a74401a,a74404a,a74407a,a74408a,a74411a,a74414a,a74415a,a74416a,a74420a,a74421a,a74424a,a74427a,a74428a,a74429a,a74432a,a74435a,a74436a,a74439a,a74442a,a74443a,a74444a,a74448a,a74449a,a74452a,a74455a,a74456a,a74457a,a74460a,a74463a,a74464a,a74467a,a74470a,a74471a,a74472a,a74476a,a74477a,a74480a,a74483a,a74484a,a74485a,a74488a,a74491a,a74492a,a74495a,a74498a,a74499a,a74500a,a74504a,a74505a,a74508a,a74511a,a74512a,a74513a,a74516a,a74519a,a74520a,a74523a,a74526a,a74527a,a74528a,a74532a,a74533a,a74536a,a74539a,a74540a,a74541a,a74544a,a74547a,a74548a,a74551a,a74554a,a74555a,a74556a,a74560a,a74561a,a74564a,a74567a,a74568a,a74569a,a74572a,a74575a,a74576a,a74579a,a74582a,a74583a,a74584a,a74588a,a74589a,a74592a,a74595a,a74596a,a74597a,a74600a,a74603a,a74604a,a74607a,a74610a,a74611a,a74612a,a74616a,a74617a,a74620a,a74623a,a74624a,a74625a,a74628a,a74631a,a74632a,a74635a,a74638a,a74639a,a74640a,a74644a,a74645a,a74648a,a74651a,a74652a,a74653a,a74656a,a74659a,a74660a,a74663a,a74666a,a74667a,a74668a,a74672a,a74673a,a74676a,a74679a,a74680a,a74681a,a74684a,a74687a,a74688a,a74691a,a74694a,a74695a,a74696a,a74700a,a74701a,a74704a,a74707a,a74708a,a74709a,a74712a,a74715a,a74716a,a74719a,a74722a,a74723a,a74724a,a74728a,a74729a,a74732a,a74735a,a74736a,a74737a,a74740a,a74743a,a74744a,a74747a,a74750a,a74751a,a74752a,a74756a,a74757a,a74760a,a74763a,a74764a,a74765a,a74768a,a74771a,a74772a,a74775a,a74778a,a74779a,a74780a,a74784a,a74785a,a74788a,a74791a,a74792a,a74793a,a74796a,a74799a,a74800a,a74803a,a74806a,a74807a,a74808a,a74812a,a74813a,a74816a,a74819a,a74820a,a74821a,a74824a,a74827a,a74828a,a74831a,a74834a,a74835a,a74836a,a74840a,a74841a,a74844a,a74847a,a74848a,a74849a,a74852a,a74855a,a74856a,a74859a,a74862a,a74863a,a74864a,a74868a,a74869a,a74872a,a74875a,a74876a,a74877a,a74880a,a74883a,a74884a,a74887a,a74890a,a74891a,a74892a,a74896a,a74897a,a74900a,a74903a,a74904a,a74905a,a74908a,a74911a,a74912a,a74915a,a74918a,a74919a,a74920a,a74924a,a74925a,a74928a,a74931a,a74932a,a74933a,a74936a,a74939a,a74940a,a74943a,a74946a,a74947a,a74948a,a74952a,a74953a,a74956a,a74959a,a74960a,a74961a,a74964a,a74967a,a74968a,a74971a,a74974a,a74975a,a74976a,a74980a,a74981a,a74984a,a74987a,a74988a,a74989a,a74992a,a74995a,a74996a,a74999a,a75002a,a75003a,a75004a,a75008a,a75009a,a75012a,a75015a,a75016a,a75017a,a75020a,a75023a,a75024a,a75027a,a75030a,a75031a,a75032a,a75036a,a75037a,a75040a,a75043a,a75044a,a75045a,a75048a,a75051a,a75052a,a75055a,a75058a,a75059a,a75060a,a75064a,a75065a,a75068a,a75071a,a75072a,a75073a,a75076a,a75079a,a75080a,a75083a,a75086a,a75087a,a75088a,a75092a,a75093a,a75096a,a75099a,a75100a,a75101a,a75104a,a75107a,a75108a,a75111a,a75114a,a75115a,a75116a,a75120a,a75121a,a75124a,a75127a,a75128a,a75129a,a75132a,a75135a,a75136a,a75139a,a75142a,a75143a,a75144a,a75148a,a75149a,a75152a,a75155a,a75156a,a75157a,a75160a,a75163a,a75164a,a75167a,a75170a,a75171a,a75172a,a75175a,a75178a,a75179a,a75182a,a75185a,a75186a,a75187a,a75190a,a75193a,a75194a,a75197a,a75200a,a75201a,a75202a,a75205a,a75208a,a75209a,a75212a,a75215a,a75216a,a75217a,a75220a,a75223a,a75224a,a75227a,a75230a,a75231a,a75232a,a75235a,a75238a,a75239a,a75242a,a75245a,a75246a,a75247a,a75250a,a75253a,a75254a,a75257a,a75260a,a75261a,a75262a,a75265a,a75268a,a75269a,a75272a,a75275a,a75276a,a75277a,a75280a,a75283a,a75284a,a75287a,a75290a,a75291a,a75292a,a75295a,a75298a,a75299a,a75302a,a75305a,a75306a,a75307a,a75310a,a75313a,a75314a,a75317a,a75320a,a75321a,a75322a,a75325a,a75328a,a75329a,a75332a,a75335a,a75336a,a75337a,a75340a,a75343a,a75344a,a75347a,a75350a,a75351a,a75352a,a75355a,a75358a,a75359a,a75362a,a75365a,a75366a,a75367a,a75370a,a75373a,a75374a,a75377a,a75380a,a75381a,a75382a,a75385a,a75388a,a75389a,a75392a,a75395a,a75396a,a75397a,a75400a,a75403a,a75404a,a75407a,a75410a,a75411a,a75412a,a75415a,a75418a,a75419a,a75422a,a75425a,a75426a,a75427a,a75430a,a75433a,a75434a,a75437a,a75440a,a75441a,a75442a,a75445a,a75448a,a75449a,a75452a,a75455a,a75456a,a75457a,a75460a,a75463a,a75464a,a75467a,a75470a,a75471a,a75472a,a75475a,a75478a,a75479a,a75482a,a75485a,a75486a,a75487a,a75490a,a75493a,a75494a,a75497a,a75500a,a75501a,a75502a,a75505a,a75508a,a75509a,a75512a,a75515a,a75516a,a75517a,a75520a,a75523a,a75524a,a75527a,a75530a,a75531a,a75532a,a75535a,a75538a,a75539a,a75542a,a75545a,a75546a,a75547a,a75550a,a75553a,a75554a,a75557a,a75560a,a75561a,a75562a,a75565a,a75568a,a75569a,a75572a,a75575a,a75576a,a75577a,a75580a,a75583a,a75584a,a75587a,a75590a,a75591a,a75592a,a75595a,a75598a,a75599a,a75602a,a75605a,a75606a,a75607a,a75610a,a75613a,a75614a,a75617a,a75620a,a75621a,a75622a,a75625a,a75628a,a75629a,a75632a,a75635a,a75636a,a75637a,a75640a,a75643a,a75644a,a75647a,a75650a,a75651a,a75652a,a75655a,a75658a,a75659a,a75662a,a75665a,a75666a,a75667a,a75670a,a75673a,a75674a,a75677a,a75680a,a75681a,a75682a,a75685a,a75688a,a75689a,a75692a,a75695a,a75696a,a75697a,a75700a,a75703a,a75704a,a75707a,a75710a,a75711a,a75712a,a75715a,a75718a,a75719a,a75722a,a75725a,a75726a,a75727a,a75730a,a75733a,a75734a,a75737a,a75740a,a75741a,a75742a,a75745a,a75748a,a75749a,a75752a,a75755a,a75756a,a75757a,a75760a,a75763a,a75764a,a75767a,a75770a,a75771a,a75772a,a75775a,a75778a,a75779a,a75782a,a75785a,a75786a,a75787a,a75790a,a75793a,a75794a,a75797a,a75800a,a75801a,a75802a,a75805a,a75808a,a75809a,a75812a,a75815a,a75816a,a75817a,a75820a,a75823a,a75824a,a75827a,a75830a,a75831a,a75832a,a75835a,a75838a,a75839a,a75842a,a75845a,a75846a,a75847a,a75850a,a75853a,a75854a,a75857a,a75860a,a75861a,a75862a,a75865a,a75868a,a75869a,a75872a,a75875a,a75876a,a75877a,a75880a,a75883a,a75884a,a75887a,a75890a,a75891a,a75892a,a75895a,a75898a,a75899a,a75902a,a75905a,a75906a,a75907a,a75910a,a75913a,a75914a,a75917a,a75920a,a75921a,a75922a,a75925a,a75928a,a75929a,a75932a,a75935a,a75936a,a75937a,a75940a,a75943a,a75944a,a75947a,a75950a,a75951a,a75952a,a75955a,a75958a,a75959a,a75962a,a75965a,a75966a,a75967a,a75970a,a75973a,a75974a,a75977a,a75980a,a75981a,a75982a,a75985a,a75988a,a75989a,a75992a,a75995a,a75996a,a75997a,a76000a,a76003a,a76004a,a76007a,a76010a,a76011a,a76012a,a76015a,a76018a,a76019a,a76022a,a76025a,a76026a,a76027a,a76030a,a76033a,a76034a,a76037a,a76040a,a76041a,a76042a,a76045a,a76048a,a76049a,a76052a,a76055a,a76056a,a76057a,a76060a,a76063a,a76064a,a76067a,a76070a,a76071a,a76072a,a76075a,a76078a,a76079a,a76082a,a76085a,a76086a,a76087a,a76090a,a76093a,a76094a,a76097a,a76100a,a76101a,a76102a,a76105a,a76108a,a76109a,a76112a,a76115a,a76116a,a76117a,a76120a,a76123a,a76124a,a76127a,a76130a,a76131a,a76132a,a76135a,a76138a,a76139a,a76142a,a76145a,a76146a,a76147a,a76150a,a76153a,a76154a,a76157a,a76160a,a76161a,a76162a,a76165a,a76168a,a76169a,a76172a,a76175a,a76176a,a76177a,a76180a,a76183a,a76184a,a76187a,a76190a,a76191a,a76192a,a76195a,a76198a,a76199a,a76202a,a76205a,a76206a,a76207a,a76210a,a76213a,a76214a,a76217a,a76220a,a76221a,a76222a,a76225a,a76228a,a76229a,a76232a,a76235a,a76236a,a76237a,a76240a,a76243a,a76244a,a76247a,a76250a,a76251a,a76252a,a76255a,a76258a,a76259a,a76262a,a76265a,a76266a,a76267a,a76270a,a76273a,a76274a,a76277a,a76280a,a76281a,a76282a,a76285a,a76288a,a76289a,a76292a,a76295a,a76296a,a76297a,a76300a,a76303a,a76304a,a76307a,a76310a,a76311a,a76312a,a76315a,a76318a,a76319a,a76322a,a76325a,a76326a,a76327a,a76330a,a76333a,a76334a,a76337a,a76340a,a76341a,a76342a,a76345a,a76348a,a76349a,a76352a,a76355a,a76356a,a76357a,a76360a,a76363a,a76364a,a76367a,a76370a,a76371a,a76372a,a76375a,a76378a,a76379a,a76382a,a76385a,a76386a,a76387a,a76390a,a76393a,a76394a,a76397a,a76400a,a76401a,a76402a,a76405a,a76408a,a76409a,a76412a,a76415a,a76416a,a76417a,a76420a,a76423a,a76424a,a76427a,a76430a,a76431a,a76432a,a76435a,a76438a,a76439a,a76442a,a76445a,a76446a,a76447a,a76450a,a76453a,a76454a,a76457a,a76460a,a76461a,a76462a,a76465a,a76468a,a76469a,a76472a,a76475a,a76476a,a76477a,a76480a,a76483a,a76484a,a76487a,a76490a,a76491a,a76492a,a76495a,a76498a,a76499a,a76502a,a76505a,a76506a,a76507a,a76510a,a76513a,a76514a,a76517a,a76520a,a76521a,a76522a,a76525a,a76528a,a76529a,a76532a,a76535a,a76536a,a76537a,a76540a,a76543a,a76544a,a76547a,a76550a,a76551a,a76552a,a76555a,a76558a,a76559a,a76562a,a76565a,a76566a,a76567a,a76570a,a76573a,a76574a,a76577a,a76580a,a76581a,a76582a,a76585a,a76588a,a76589a,a76592a,a76595a,a76596a,a76597a,a76600a,a76603a,a76604a,a76607a,a76610a,a76611a,a76612a,a76615a,a76618a,a76619a,a76622a,a76625a,a76626a,a76627a,a76630a,a76633a,a76634a,a76637a,a76640a,a76641a,a76642a,a76645a,a76648a,a76649a,a76652a,a76655a,a76656a,a76657a,a76660a,a76663a,a76664a,a76667a,a76670a,a76671a,a76672a,a76675a,a76678a,a76679a,a76682a,a76685a,a76686a,a76687a,a76690a,a76693a,a76694a,a76697a,a76700a,a76701a,a76702a,a76705a,a76708a,a76709a,a76712a,a76715a,a76716a,a76717a,a76720a,a76723a,a76724a,a76727a,a76730a,a76731a,a76732a,a76735a,a76738a,a76739a,a76742a,a76745a,a76746a,a76747a,a76750a,a76753a,a76754a,a76757a,a76760a,a76761a,a76762a,a76765a,a76768a,a76769a,a76772a,a76775a,a76776a,a76777a,a76780a,a76783a,a76784a,a76787a,a76790a,a76791a,a76792a,a76795a,a76798a,a76799a,a76802a,a76805a,a76806a,a76807a,a76810a,a76813a,a76814a,a76817a,a76820a,a76821a,a76822a,a76825a,a76828a,a76829a,a76832a,a76835a,a76836a,a76837a,a76840a,a76843a,a76844a,a76847a,a76850a,a76851a,a76852a,a76855a,a76858a,a76859a,a76862a,a76865a,a76866a,a76867a,a76870a,a76873a,a76874a,a76877a,a76880a,a76881a,a76882a,a76885a,a76888a,a76889a,a76892a,a76895a,a76896a,a76897a,a76900a,a76903a,a76904a,a76907a,a76910a,a76911a,a76912a,a76915a,a76918a,a76919a,a76922a,a76925a,a76926a,a76927a,a76930a,a76933a,a76934a,a76937a,a76940a,a76941a,a76942a,a76945a,a76948a,a76949a,a76952a,a76955a,a76956a,a76957a,a76960a,a76963a,a76964a,a76967a,a76970a,a76971a,a76972a,a76975a,a76978a,a76979a,a76982a,a76985a,a76986a,a76987a,a76990a,a76993a,a76994a,a76997a,a77000a,a77001a,a77002a,a77005a,a77008a,a77009a,a77012a,a77015a,a77016a,a77017a,a77020a,a77023a,a77024a,a77027a,a77030a,a77031a,a77032a,a77035a,a77038a,a77039a,a77042a,a77045a,a77046a,a77047a,a77050a,a77053a,a77054a,a77057a,a77060a,a77061a,a77062a,a77065a,a77068a,a77069a,a77072a,a77075a,a77076a,a77077a,a77080a,a77083a,a77084a,a77087a,a77090a,a77091a,a77092a,a77095a,a77098a,a77099a,a77102a,a77105a,a77106a,a77107a,a77110a,a77113a,a77114a,a77117a,a77120a,a77121a,a77122a,a77125a,a77128a,a77129a,a77132a,a77135a,a77136a,a77137a,a77140a,a77143a,a77144a,a77147a,a77150a,a77151a,a77152a,a77155a,a77158a,a77159a,a77162a,a77165a,a77166a,a77167a,a77170a,a77173a,a77174a,a77177a,a77180a,a77181a,a77182a,a77185a,a77188a,a77189a,a77192a,a77195a,a77196a,a77197a,a77200a,a77203a,a77204a,a77207a,a77210a,a77211a,a77212a,a77215a,a77218a,a77219a,a77222a,a77225a,a77226a,a77227a,a77230a,a77233a,a77234a,a77237a,a77240a,a77241a,a77242a,a77245a,a77248a,a77249a,a77252a,a77255a,a77256a,a77257a,a77260a,a77263a,a77264a,a77267a,a77270a,a77271a,a77272a,a77275a,a77278a,a77279a,a77282a,a77285a,a77286a,a77287a,a77290a,a77293a,a77294a,a77297a,a77300a,a77301a,a77302a,a77305a,a77308a,a77309a,a77312a,a77315a,a77316a,a77317a,a77320a,a77323a,a77324a,a77327a,a77330a,a77331a,a77332a,a77335a,a77338a,a77339a,a77342a,a77345a,a77346a,a77347a,a77350a,a77353a,a77354a,a77357a,a77360a,a77361a,a77362a,a77365a,a77368a,a77369a,a77372a,a77375a,a77376a,a77377a,a77380a,a77383a,a77384a,a77387a,a77390a,a77391a,a77392a,a77395a,a77398a,a77399a,a77402a,a77405a,a77406a,a77407a,a77410a,a77413a,a77414a,a77417a,a77420a,a77421a,a77422a,a77425a,a77428a,a77429a,a77432a,a77435a,a77436a,a77437a,a77440a,a77443a,a77444a,a77447a,a77450a,a77451a,a77452a,a77455a,a77458a,a77459a,a77462a,a77465a,a77466a,a77467a,a77470a,a77473a,a77474a,a77477a,a77480a,a77481a,a77482a,a77485a,a77488a,a77489a,a77492a,a77495a,a77496a,a77497a,a77500a,a77503a,a77504a,a77507a,a77510a,a77511a,a77512a,a77515a,a77518a,a77519a,a77522a,a77525a,a77526a,a77527a,a77530a,a77533a,a77534a,a77537a,a77540a,a77541a,a77542a,a77545a,a77548a,a77549a,a77552a,a77555a,a77556a,a77557a,a77560a,a77563a,a77564a,a77567a,a77570a,a77571a,a77572a,a77575a,a77578a,a77579a,a77582a,a77585a,a77586a,a77587a,a77590a,a77593a,a77594a,a77597a,a77600a,a77601a,a77602a,a77605a,a77608a,a77609a,a77612a,a77615a,a77616a,a77617a,a77620a,a77623a,a77624a,a77627a,a77630a,a77631a,a77632a,a77635a,a77638a,a77639a,a77642a,a77645a,a77646a,a77647a,a77650a,a77653a,a77654a,a77657a,a77660a,a77661a,a77662a,a77665a,a77668a,a77669a,a77672a,a77675a,a77676a,a77677a,a77680a,a77683a,a77684a,a77687a,a77690a,a77691a,a77692a,a77695a,a77698a,a77699a,a77702a,a77705a,a77706a,a77707a,a77710a,a77713a,a77714a,a77717a,a77720a,a77721a,a77722a,a77725a,a77728a,a77729a,a77732a,a77735a,a77736a,a77737a,a77740a,a77743a,a77744a,a77747a,a77750a,a77751a,a77752a,a77755a,a77758a,a77759a,a77762a,a77765a,a77766a,a77767a,a77770a,a77773a,a77774a,a77777a,a77780a,a77781a,a77782a,a77785a,a77788a,a77789a,a77792a,a77795a,a77796a,a77797a,a77800a,a77803a,a77804a,a77807a,a77810a,a77811a,a77812a,a77815a,a77818a,a77819a,a77822a,a77825a,a77826a,a77827a,a77830a,a77833a,a77834a,a77837a,a77840a,a77841a,a77842a,a77845a,a77848a,a77849a,a77852a,a77855a,a77856a,a77857a,a77860a,a77863a,a77864a,a77867a,a77870a,a77871a,a77872a,a77875a,a77878a,a77879a,a77882a,a77885a,a77886a,a77887a,a77890a,a77893a,a77894a,a77897a,a77900a,a77901a,a77902a,a77905a,a77908a,a77909a,a77912a,a77915a,a77916a,a77917a,a77920a,a77923a,a77924a,a77927a,a77930a,a77931a,a77932a,a77935a,a77938a,a77939a,a77942a,a77945a,a77946a,a77947a,a77950a,a77953a,a77954a,a77957a,a77960a,a77961a,a77962a,a77965a,a77968a,a77969a,a77972a,a77975a,a77976a,a77977a,a77980a,a77983a,a77984a,a77987a,a77990a,a77991a,a77992a,a77995a,a77998a,a77999a,a78002a,a78005a,a78006a,a78007a,a78010a,a78013a,a78014a,a78017a,a78020a,a78021a,a78022a,a78025a,a78028a,a78029a,a78032a,a78035a,a78036a,a78037a,a78040a,a78043a,a78044a,a78047a,a78050a,a78051a,a78052a,a78055a,a78058a,a78059a,a78062a,a78065a,a78066a,a78067a,a78070a,a78073a,a78074a,a78077a,a78080a,a78081a,a78082a,a78085a,a78088a,a78089a,a78092a,a78095a,a78096a,a78097a,a78100a,a78103a,a78104a,a78107a,a78110a,a78111a,a78112a,a78115a,a78118a,a78119a,a78122a,a78125a,a78126a,a78127a,a78130a,a78133a,a78134a,a78137a,a78140a,a78141a,a78142a,a78145a,a78148a,a78149a,a78152a,a78155a,a78156a,a78157a,a78160a,a78163a,a78164a,a78167a,a78170a,a78171a,a78172a,a78175a,a78178a,a78179a,a78182a,a78185a,a78186a,a78187a,a78190a,a78193a,a78194a,a78197a,a78200a,a78201a,a78202a,a78205a,a78208a,a78209a,a78212a,a78215a,a78216a,a78217a,a78220a,a78223a,a78224a,a78227a,a78230a,a78231a,a78232a,a78235a,a78238a,a78239a,a78242a,a78245a,a78246a,a78247a,a78250a,a78253a,a78254a,a78257a,a78260a,a78261a,a78262a,a78265a,a78268a,a78269a,a78272a,a78275a,a78276a,a78277a,a78280a,a78283a,a78284a,a78287a,a78290a,a78291a,a78292a,a78295a,a78298a,a78299a,a78302a,a78305a,a78306a,a78307a,a78310a,a78313a,a78314a,a78317a,a78320a,a78321a,a78322a,a78325a,a78328a,a78329a,a78332a,a78335a,a78336a,a78337a,a78340a,a78343a,a78344a,a78347a,a78350a,a78351a,a78352a,a78355a,a78358a,a78359a,a78362a,a78365a,a78366a,a78367a,a78370a,a78373a,a78374a,a78377a,a78380a,a78381a,a78382a,a78385a,a78388a,a78389a,a78392a,a78395a,a78396a,a78397a,a78400a,a78403a,a78404a,a78407a,a78410a,a78411a,a78412a,a78415a,a78418a,a78419a,a78422a,a78425a,a78426a,a78427a,a78430a,a78433a,a78434a,a78437a,a78440a,a78441a,a78442a,a78445a,a78448a,a78449a,a78452a,a78455a,a78456a,a78457a,a78460a,a78463a,a78464a,a78467a,a78470a,a78471a,a78472a,a78475a,a78478a,a78479a,a78482a,a78485a,a78486a,a78487a,a78490a,a78493a,a78494a,a78497a,a78500a,a78501a,a78502a,a78505a,a78508a,a78509a,a78512a,a78515a,a78516a,a78517a,a78520a,a78523a,a78524a,a78527a,a78530a,a78531a,a78532a,a78535a,a78538a,a78539a,a78542a,a78545a,a78546a,a78547a,a78550a,a78553a,a78554a,a78557a,a78560a,a78561a,a78562a,a78565a,a78568a,a78569a,a78572a,a78575a,a78576a,a78577a,a78580a,a78583a,a78584a,a78587a,a78590a,a78591a,a78592a,a78595a,a78598a,a78599a,a78602a,a78605a,a78606a,a78607a,a78610a,a78613a,a78614a,a78617a,a78620a,a78621a,a78622a,a78625a,a78628a,a78629a,a78632a,a78635a,a78636a,a78637a,a78640a,a78643a,a78644a,a78647a,a78650a,a78651a,a78652a,a78655a,a78658a,a78659a,a78662a,a78665a,a78666a,a78667a,a78670a,a78673a,a78674a,a78677a,a78680a,a78681a,a78682a,a78685a,a78688a,a78689a,a78692a,a78695a,a78696a,a78697a,a78700a,a78703a,a78704a,a78707a,a78710a,a78711a,a78712a,a78715a,a78718a,a78719a,a78722a,a78725a,a78726a,a78727a,a78730a,a78733a,a78734a,a78737a,a78740a,a78741a,a78742a,a78745a,a78748a,a78749a,a78752a,a78755a,a78756a,a78757a,a78760a,a78763a,a78764a,a78767a,a78770a,a78771a,a78772a,a78775a,a78778a,a78779a,a78782a,a78785a,a78786a,a78787a,a78790a,a78793a,a78794a,a78797a,a78800a,a78801a,a78802a,a78805a,a78808a,a78809a,a78812a,a78815a,a78816a,a78817a,a78820a,a78823a,a78824a,a78827a,a78830a,a78831a,a78832a,a78835a,a78838a,a78839a,a78842a,a78845a,a78846a,a78847a,a78850a,a78853a,a78854a,a78857a,a78860a,a78861a,a78862a,a78865a,a78868a,a78869a,a78872a,a78875a,a78876a,a78877a,a78880a,a78883a,a78884a,a78887a,a78890a,a78891a,a78892a,a78895a,a78898a,a78899a,a78902a,a78905a,a78906a,a78907a,a78910a,a78913a,a78914a,a78917a,a78920a,a78921a,a78922a,a78925a,a78928a,a78929a,a78932a,a78935a,a78936a,a78937a,a78940a,a78943a,a78944a,a78947a,a78950a,a78951a,a78952a,a78955a,a78958a,a78959a,a78962a,a78965a,a78966a,a78967a,a78970a,a78973a,a78974a,a78977a,a78980a,a78981a,a78982a,a78985a,a78988a,a78989a,a78992a,a78995a,a78996a,a78997a,a79000a,a79003a,a79004a,a79007a,a79010a,a79011a,a79012a,a79015a,a79018a,a79019a,a79022a,a79025a,a79026a,a79027a,a79030a,a79033a,a79034a,a79037a,a79040a,a79041a,a79042a,a79045a,a79048a,a79049a,a79052a,a79055a,a79056a,a79057a,a79060a,a79063a,a79064a,a79067a,a79070a,a79071a,a79072a,a79075a,a79078a,a79079a,a79082a,a79085a,a79086a,a79087a,a79090a,a79093a,a79094a,a79097a,a79100a,a79101a,a79102a,a79105a,a79108a,a79109a,a79112a,a79115a,a79116a,a79117a,a79120a,a79123a,a79124a,a79127a,a79130a,a79131a,a79132a,a79135a,a79138a,a79139a,a79142a,a79145a,a79146a,a79147a,a79150a,a79153a,a79154a,a79157a,a79160a,a79161a,a79162a,a79165a,a79168a,a79169a,a79172a,a79175a,a79176a,a79177a,a79180a,a79183a,a79184a,a79187a,a79190a,a79191a,a79192a,a79195a,a79198a,a79199a,a79202a,a79205a,a79206a,a79207a,a79210a,a79213a,a79214a,a79217a,a79220a,a79221a,a79222a,a79225a,a79228a,a79229a,a79232a,a79235a,a79236a,a79237a,a79240a,a79243a,a79244a,a79247a,a79250a,a79251a,a79252a,a79255a,a79258a,a79259a,a79262a,a79265a,a79266a,a79267a,a79270a,a79273a,a79274a,a79277a,a79280a,a79281a,a79282a,a79285a,a79288a,a79289a,a79292a,a79295a,a79296a,a79297a,a79300a,a79303a,a79304a,a79307a,a79310a,a79311a,a79312a,a79315a,a79318a,a79319a,a79322a,a79325a,a79326a,a79327a,a79330a,a79333a,a79334a,a79337a,a79340a,a79341a,a79342a,a79345a,a79348a,a79349a,a79352a,a79355a,a79356a,a79357a,a79360a,a79363a,a79364a,a79367a,a79370a,a79371a,a79372a,a79375a,a79378a,a79379a,a79382a,a79385a,a79386a,a79387a,a79390a,a79393a,a79394a,a79397a,a79400a,a79401a,a79402a,a79405a,a79408a,a79409a,a79412a,a79415a,a79416a,a79417a,a79420a,a79423a,a79424a,a79427a,a79430a,a79431a,a79432a,a79435a,a79438a,a79439a,a79442a,a79445a,a79446a,a79447a,a79450a,a79453a,a79454a,a79457a,a79460a,a79461a,a79462a,a79465a,a79468a,a79469a,a79472a,a79475a,a79476a,a79477a,a79480a,a79483a,a79484a,a79487a,a79490a,a79491a,a79492a,a79495a,a79498a,a79499a,a79502a,a79505a,a79506a,a79507a,a79510a,a79513a,a79514a,a79517a,a79520a,a79521a,a79522a,a79525a,a79528a,a79529a,a79532a,a79535a,a79536a,a79537a,a79540a,a79543a,a79544a,a79547a,a79550a,a79551a,a79552a,a79555a,a79558a,a79559a,a79562a,a79565a,a79566a,a79567a,a79570a,a79573a,a79574a,a79577a,a79580a,a79581a,a79582a,a79585a,a79588a,a79589a,a79592a,a79595a,a79596a,a79597a,a79600a,a79603a,a79604a,a79607a,a79610a,a79611a,a79612a,a79615a,a79618a,a79619a,a79622a,a79625a,a79626a,a79627a,a79630a,a79633a,a79634a,a79637a,a79640a,a79641a,a79642a,a79645a,a79648a,a79649a,a79652a,a79655a,a79656a,a79657a,a79660a,a79663a,a79664a,a79667a,a79670a,a79671a,a79672a,a79675a,a79678a,a79679a,a79682a,a79685a,a79686a,a79687a,a79690a,a79693a,a79694a,a79697a,a79700a,a79701a,a79702a,a79705a,a79708a,a79709a,a79712a,a79715a,a79716a,a79717a,a79720a,a79723a,a79724a,a79727a,a79730a,a79731a,a79732a,a79735a,a79738a,a79739a,a79742a,a79745a,a79746a,a79747a,a79750a,a79753a,a79754a,a79757a,a79760a,a79761a,a79762a,a79765a,a79768a,a79769a,a79772a,a79775a,a79776a,a79777a,a79780a,a79783a,a79784a,a79787a,a79790a,a79791a,a79792a,a79795a,a79798a,a79799a,a79802a,a79805a,a79806a,a79807a,a79810a,a79813a,a79814a,a79817a,a79820a,a79821a,a79822a,a79825a,a79828a,a79829a,a79832a,a79835a,a79836a,a79837a,a79840a,a79843a,a79844a,a79847a,a79850a,a79851a,a79852a,a79855a,a79858a,a79859a,a79862a,a79865a,a79866a,a79867a,a79870a,a79873a,a79874a,a79877a,a79880a,a79881a,a79882a,a79885a,a79888a,a79889a,a79892a,a79895a,a79896a,a79897a,a79900a,a79903a,a79904a,a79907a,a79910a,a79911a,a79912a,a79915a,a79918a,a79919a,a79922a,a79925a,a79926a,a79927a,a79930a,a79933a,a79934a,a79937a,a79940a,a79941a,a79942a,a79945a,a79948a,a79949a,a79952a,a79955a,a79956a,a79957a,a79960a,a79963a,a79964a,a79967a,a79970a,a79971a,a79972a,a79975a,a79978a,a79979a,a79982a,a79985a,a79986a,a79987a,a79990a,a79993a,a79994a,a79997a,a80000a,a80001a,a80002a,a80005a,a80008a,a80009a,a80012a,a80015a,a80016a,a80017a,a80020a,a80023a,a80024a,a80027a,a80030a,a80031a,a80032a,a80035a,a80038a,a80039a,a80042a,a80045a,a80046a,a80047a,a80050a,a80053a,a80054a,a80057a,a80060a,a80061a,a80062a,a80065a,a80068a,a80069a,a80072a,a80075a,a80076a,a80077a,a80080a,a80083a,a80084a,a80087a,a80090a,a80091a,a80092a,a80095a,a80098a,a80099a,a80102a,a80105a,a80106a,a80107a,a80110a,a80113a,a80114a,a80117a,a80120a,a80121a,a80122a,a80125a,a80128a,a80129a,a80132a,a80135a,a80136a,a80137a,a80140a,a80143a,a80144a,a80147a,a80150a,a80151a,a80152a,a80155a,a80158a,a80159a,a80162a,a80165a,a80166a,a80167a,a80170a,a80173a,a80174a,a80177a,a80180a,a80181a,a80182a,a80185a,a80188a,a80189a,a80192a,a80195a,a80196a,a80197a,a80200a,a80203a,a80204a,a80207a,a80210a,a80211a,a80212a,a80215a,a80218a,a80219a,a80222a,a80225a,a80226a,a80227a,a80230a,a80233a,a80234a,a80237a,a80240a,a80241a,a80242a,a80245a,a80248a,a80249a,a80252a,a80255a,a80256a,a80257a,a80260a,a80263a,a80264a,a80267a,a80270a,a80271a,a80272a,a80275a,a80278a,a80279a,a80282a,a80285a,a80286a,a80287a,a80290a,a80293a,a80294a,a80297a,a80300a,a80301a,a80302a,a80305a,a80308a,a80309a,a80312a,a80315a,a80316a,a80317a,a80320a,a80323a,a80324a,a80327a,a80330a,a80331a,a80332a,a80335a,a80338a,a80339a,a80342a,a80345a,a80346a,a80347a,a80350a,a80353a,a80354a,a80357a,a80360a,a80361a,a80362a,a80365a,a80368a,a80369a,a80372a,a80375a,a80376a,a80377a,a80380a,a80383a,a80384a,a80387a,a80390a,a80391a,a80392a,a80395a,a80398a,a80399a,a80402a,a80405a,a80406a,a80407a,a80410a,a80413a,a80414a,a80417a,a80420a,a80421a,a80422a,a80425a,a80428a,a80429a,a80432a,a80435a,a80436a,a80437a,a80440a,a80443a,a80444a,a80447a,a80450a,a80451a,a80452a,a80455a,a80458a,a80459a,a80462a,a80465a,a80466a,a80467a,a80470a,a80473a,a80474a,a80477a,a80480a,a80481a,a80482a,a80485a,a80488a,a80489a,a80492a,a80495a,a80496a,a80497a,a80500a,a80503a,a80504a,a80507a,a80510a,a80511a,a80512a,a80515a,a80518a,a80519a,a80522a,a80525a,a80526a,a80527a,a80530a,a80533a,a80534a,a80537a,a80540a,a80541a,a80542a,a80545a,a80548a,a80549a,a80552a,a80555a,a80556a,a80557a,a80560a,a80563a,a80564a,a80567a,a80570a,a80571a,a80572a,a80575a,a80578a,a80579a,a80582a,a80585a,a80586a,a80587a,a80590a,a80593a,a80594a,a80597a,a80600a,a80601a,a80602a,a80605a,a80608a,a80609a,a80612a,a80615a,a80616a,a80617a,a80620a,a80623a,a80624a,a80627a,a80630a,a80631a,a80632a,a80635a,a80638a,a80639a,a80642a,a80645a,a80646a,a80647a,a80650a,a80653a,a80654a,a80657a,a80660a,a80661a,a80662a,a80665a,a80668a,a80669a,a80672a,a80675a,a80676a,a80677a,a80680a,a80683a,a80684a,a80687a,a80690a,a80691a,a80692a,a80695a,a80698a,a80699a,a80702a,a80705a,a80706a,a80707a,a80710a,a80713a,a80714a,a80717a,a80720a,a80721a,a80722a,a80725a,a80728a,a80729a,a80732a,a80735a,a80736a,a80737a,a80740a,a80743a,a80744a,a80747a,a80750a,a80751a,a80752a,a80755a,a80758a,a80759a,a80762a,a80765a,a80766a,a80767a,a80770a,a80773a,a80774a,a80777a,a80780a,a80781a,a80782a,a80785a,a80788a,a80789a,a80792a,a80795a,a80796a,a80797a,a80800a,a80803a,a80804a,a80807a,a80810a,a80811a,a80812a,a80815a,a80818a,a80819a,a80822a,a80825a,a80826a,a80827a,a80830a,a80833a,a80834a,a80837a,a80840a,a80841a,a80842a,a80845a,a80848a,a80849a,a80852a,a80855a,a80856a,a80857a,a80860a,a80863a,a80864a,a80867a,a80870a,a80871a,a80872a,a80875a,a80878a,a80879a,a80882a,a80885a,a80886a,a80887a,a80890a,a80893a,a80894a,a80897a,a80900a,a80901a,a80902a,a80905a,a80908a,a80909a,a80912a,a80915a,a80916a,a80917a,a80920a,a80923a,a80924a,a80927a,a80930a,a80931a,a80932a,a80935a,a80938a,a80939a,a80942a,a80945a,a80946a,a80947a,a80950a,a80953a,a80954a,a80957a,a80960a,a80961a,a80962a,a80965a,a80968a,a80969a,a80972a,a80975a,a80976a,a80977a,a80980a,a80983a,a80984a,a80987a,a80990a,a80991a,a80992a,a80995a,a80998a,a80999a,a81002a,a81005a,a81006a,a81007a,a81010a,a81013a,a81014a,a81017a,a81020a,a81021a,a81022a,a81025a,a81028a,a81029a,a81032a,a81035a,a81036a,a81037a,a81040a,a81043a,a81044a,a81047a,a81050a,a81051a,a81052a,a81055a,a81058a,a81059a,a81062a,a81065a,a81066a,a81067a,a81070a,a81073a,a81074a,a81077a,a81080a,a81081a,a81082a,a81085a,a81088a,a81089a,a81092a,a81095a,a81096a,a81097a,a81100a,a81103a,a81104a,a81107a,a81110a,a81111a,a81112a,a81115a,a81118a,a81119a,a81122a,a81125a,a81126a,a81127a,a81130a,a81133a,a81134a,a81137a,a81140a,a81141a,a81142a,a81145a,a81148a,a81149a,a81152a,a81155a,a81156a,a81157a,a81160a,a81163a,a81164a,a81167a,a81170a,a81171a,a81172a,a81175a,a81178a,a81179a,a81182a,a81185a,a81186a,a81187a,a81190a,a81193a,a81194a,a81197a,a81200a,a81201a,a81202a,a81205a,a81208a,a81209a,a81212a,a81215a,a81216a,a81217a,a81220a,a81223a,a81224a,a81227a,a81230a,a81231a,a81232a,a81235a,a81238a,a81239a,a81242a,a81245a,a81246a,a81247a,a81250a,a81253a,a81254a,a81257a,a81260a,a81261a,a81262a,a81265a,a81268a,a81269a,a81272a,a81275a,a81276a,a81277a,a81280a,a81283a,a81284a,a81287a,a81290a,a81291a,a81292a,a81295a,a81298a,a81299a,a81302a,a81305a,a81306a,a81307a,a81310a,a81313a,a81314a,a81317a,a81320a,a81321a,a81322a,a81325a,a81328a,a81329a,a81332a,a81335a,a81336a,a81337a,a81340a,a81343a,a81344a,a81347a,a81350a,a81351a,a81352a,a81355a,a81358a,a81359a,a81362a,a81365a,a81366a,a81367a,a81370a,a81373a,a81374a,a81377a,a81380a,a81381a,a81382a,a81385a,a81388a,a81389a,a81392a,a81395a,a81396a,a81397a,a81400a,a81403a,a81404a,a81407a,a81410a,a81411a,a81412a,a81415a,a81418a,a81419a,a81422a,a81425a,a81426a,a81427a,a81430a,a81433a,a81434a,a81437a,a81440a,a81441a,a81442a,a81445a,a81448a,a81449a,a81452a,a81455a,a81456a,a81457a,a81460a,a81463a,a81464a,a81467a,a81470a,a81471a,a81472a,a81475a,a81478a,a81479a,a81482a,a81485a,a81486a,a81487a,a81490a,a81493a,a81494a,a81497a,a81500a,a81501a,a81502a,a81505a,a81508a,a81509a,a81512a,a81515a,a81516a,a81517a,a81520a,a81523a,a81524a,a81527a,a81530a,a81531a,a81532a,a81535a,a81538a,a81539a,a81542a,a81545a,a81546a,a81547a,a81550a,a81553a,a81554a,a81557a,a81560a,a81561a,a81562a,a81565a,a81568a,a81569a,a81572a,a81575a,a81576a,a81577a,a81580a,a81583a,a81584a,a81587a,a81590a,a81591a,a81592a,a81595a,a81598a,a81599a,a81602a,a81605a,a81606a,a81607a,a81610a,a81613a,a81614a,a81617a,a81620a,a81621a,a81622a,a81625a,a81628a,a81629a,a81632a,a81635a,a81636a,a81637a,a81640a,a81643a,a81644a,a81647a,a81650a,a81651a,a81652a,a81655a,a81658a,a81659a,a81662a,a81665a,a81666a,a81667a,a81670a,a81673a,a81674a,a81677a,a81680a,a81681a,a81682a,a81685a,a81688a,a81689a,a81692a,a81695a,a81696a,a81697a,a81700a,a81703a,a81704a,a81707a,a81710a,a81711a,a81712a,a81715a,a81718a,a81719a,a81722a,a81725a,a81726a,a81727a,a81730a,a81733a,a81734a,a81737a,a81740a,a81741a,a81742a,a81745a,a81748a,a81749a,a81752a,a81755a,a81756a,a81757a,a81760a,a81763a,a81764a,a81767a,a81770a,a81771a,a81772a,a81775a,a81778a,a81779a,a81782a,a81785a,a81786a,a81787a,a81790a,a81793a,a81794a,a81797a,a81800a,a81801a,a81802a,a81805a,a81808a,a81809a,a81812a,a81815a,a81816a,a81817a,a81820a,a81823a,a81824a,a81827a,a81830a,a81831a,a81832a,a81835a,a81838a,a81839a,a81842a,a81845a,a81846a,a81847a,a81850a,a81853a,a81854a,a81857a,a81860a,a81861a,a81862a,a81865a,a81868a,a81869a,a81872a,a81875a,a81876a,a81877a,a81880a,a81883a,a81884a,a81887a,a81890a,a81891a,a81892a,a81895a,a81898a,a81899a,a81902a,a81905a,a81906a,a81907a,a81910a,a81913a,a81914a,a81917a,a81920a,a81921a,a81922a,a81925a,a81928a,a81929a,a81932a,a81935a,a81936a,a81937a,a81940a,a81943a,a81944a,a81947a,a81950a,a81951a,a81952a,a81955a,a81958a,a81959a,a81962a,a81965a,a81966a,a81967a,a81970a,a81973a,a81974a,a81977a,a81980a,a81981a,a81982a,a81985a,a81988a,a81989a,a81992a,a81995a,a81996a,a81997a,a82000a,a82003a,a82004a,a82007a,a82010a,a82011a,a82012a,a82015a,a82018a,a82019a,a82022a,a82025a,a82026a,a82027a,a82030a,a82033a,a82034a,a82037a,a82040a,a82041a,a82042a,a82045a,a82048a,a82049a,a82052a,a82055a,a82056a,a82057a,a82060a,a82063a,a82064a,a82067a,a82070a,a82071a,a82072a,a82075a,a82078a,a82079a,a82082a,a82085a,a82086a,a82087a,a82090a,a82093a,a82094a,a82097a,a82100a,a82101a,a82102a,a82105a,a82108a,a82109a,a82112a,a82115a,a82116a,a82117a,a82120a,a82123a,a82124a,a82127a,a82130a,a82131a,a82132a,a82135a,a82138a,a82139a,a82142a,a82145a,a82146a,a82147a,a82150a,a82153a,a82154a,a82157a,a82160a,a82161a,a82162a,a82165a,a82168a,a82169a,a82172a,a82175a,a82176a,a82177a,a82180a,a82183a,a82184a,a82187a,a82190a,a82191a,a82192a,a82195a,a82198a,a82199a,a82202a,a82205a,a82206a,a82207a,a82210a,a82213a,a82214a,a82217a,a82220a,a82221a,a82222a,a82225a,a82228a,a82229a,a82232a,a82235a,a82236a,a82237a,a82240a,a82243a,a82244a,a82247a,a82250a,a82251a,a82252a,a82255a,a82258a,a82259a,a82262a,a82265a,a82266a,a82267a,a82270a,a82273a,a82274a,a82277a,a82280a,a82281a,a82282a,a82285a,a82288a,a82289a,a82292a,a82295a,a82296a,a82297a,a82300a,a82303a,a82304a,a82307a,a82310a,a82311a,a82312a,a82315a,a82318a,a82319a,a82322a,a82325a,a82326a,a82327a,a82330a,a82333a,a82334a,a82337a,a82340a,a82341a,a82342a,a82345a,a82348a,a82349a,a82352a,a82355a,a82356a,a82357a,a82360a,a82363a,a82364a,a82367a,a82370a,a82371a,a82372a,a82375a,a82378a,a82379a,a82382a,a82385a,a82386a,a82387a,a82390a,a82393a,a82394a,a82397a,a82400a,a82401a,a82402a,a82405a,a82408a,a82409a,a82412a,a82415a,a82416a,a82417a,a82420a,a82423a,a82424a,a82427a,a82430a,a82431a,a82432a,a82435a,a82438a,a82439a,a82442a,a82445a,a82446a,a82447a,a82450a,a82453a,a82454a,a82457a,a82460a,a82461a,a82462a,a82465a,a82468a,a82469a,a82472a,a82475a,a82476a,a82477a,a82480a,a82483a,a82484a,a82487a,a82490a,a82491a,a82492a,a82495a,a82498a,a82499a,a82502a,a82505a,a82506a,a82507a,a82510a,a82513a,a82514a,a82517a,a82520a,a82521a,a82522a,a82525a,a82528a,a82529a,a82532a,a82535a,a82536a,a82537a,a82540a,a82543a,a82544a,a82547a,a82550a,a82551a,a82552a,a82555a,a82558a,a82559a,a82562a,a82565a,a82566a,a82567a,a82570a,a82573a,a82574a,a82577a,a82580a,a82581a,a82582a,a82585a,a82588a,a82589a,a82592a,a82595a,a82596a,a82597a,a82600a,a82603a,a82604a,a82607a,a82610a,a82611a,a82612a,a82615a,a82618a,a82619a,a82622a,a82625a,a82626a,a82627a,a82630a,a82633a,a82634a,a82637a,a82640a,a82641a,a82642a,a82645a,a82648a,a82649a,a82652a,a82655a,a82656a,a82657a,a82660a,a82663a,a82664a,a82667a,a82670a,a82671a,a82672a,a82675a,a82678a,a82679a,a82682a,a82685a,a82686a,a82687a,a82690a,a82693a,a82694a,a82697a,a82700a,a82701a,a82702a,a82705a,a82708a,a82709a,a82712a,a82715a,a82716a,a82717a,a82720a,a82723a,a82724a,a82727a,a82730a,a82731a,a82732a,a82735a,a82738a,a82739a,a82742a,a82745a,a82746a,a82747a,a82750a,a82753a,a82754a,a82757a,a82760a,a82761a,a82762a,a82765a,a82768a,a82769a,a82772a,a82775a,a82776a,a82777a,a82780a,a82783a,a82784a,a82787a,a82790a,a82791a,a82792a,a82795a,a82798a,a82799a,a82802a,a82805a,a82806a,a82807a,a82810a,a82813a,a82814a,a82817a,a82820a,a82821a,a82822a,a82825a,a82828a,a82829a,a82832a,a82835a,a82836a,a82837a,a82840a,a82843a,a82844a,a82847a,a82850a,a82851a,a82852a,a82855a,a82858a,a82859a,a82862a,a82865a,a82866a,a82867a,a82870a,a82873a,a82874a,a82877a,a82880a,a82881a,a82882a,a82885a,a82888a,a82889a,a82892a,a82895a,a82896a,a82897a,a82900a,a82903a,a82904a,a82907a,a82910a,a82911a,a82912a,a82915a,a82918a,a82919a,a82922a,a82925a,a82926a,a82927a,a82930a,a82933a,a82934a,a82937a,a82940a,a82941a,a82942a,a82945a,a82948a,a82949a,a82952a,a82955a,a82956a,a82957a,a82960a,a82963a,a82964a,a82967a,a82970a,a82971a,a82972a,a82975a,a82978a,a82979a,a82982a,a82985a,a82986a,a82987a,a82990a,a82993a,a82994a,a82997a,a83000a,a83001a,a83002a,a83005a,a83008a,a83009a,a83012a,a83015a,a83016a,a83017a,a83020a,a83023a,a83024a,a83027a,a83030a,a83031a,a83032a,a83035a,a83038a,a83039a,a83042a,a83045a,a83046a,a83047a,a83050a,a83053a,a83054a,a83057a,a83060a,a83061a,a83062a,a83065a,a83068a,a83069a,a83072a,a83075a,a83076a,a83077a,a83080a,a83083a,a83084a,a83087a,a83090a,a83091a,a83092a,a83095a,a83098a,a83099a,a83102a,a83105a,a83106a,a83107a,a83110a,a83113a,a83114a,a83117a,a83120a,a83121a,a83122a,a83125a,a83128a,a83129a,a83132a,a83135a,a83136a,a83137a,a83140a,a83143a,a83144a,a83147a,a83150a,a83151a,a83152a,a83155a,a83158a,a83159a,a83162a,a83165a,a83166a,a83167a,a83170a,a83173a,a83174a,a83177a,a83180a,a83181a,a83182a,a83185a,a83188a,a83189a,a83192a,a83195a,a83196a,a83197a,a83200a,a83203a,a83204a,a83207a,a83210a,a83211a,a83212a,a83215a,a83218a,a83219a,a83222a,a83225a,a83226a,a83227a,a83230a,a83233a,a83234a,a83237a,a83240a,a83241a,a83242a,a83245a,a83248a,a83249a,a83252a,a83255a,a83256a,a83257a,a83260a,a83263a,a83264a,a83267a,a83270a,a83271a,a83272a,a83275a,a83278a,a83279a,a83282a,a83285a,a83286a,a83287a,a83290a,a83293a,a83294a,a83297a,a83300a,a83301a,a83302a,a83305a,a83308a,a83309a,a83312a,a83315a,a83316a,a83317a,a83320a,a83323a,a83324a,a83327a,a83330a,a83331a,a83332a,a83335a,a83338a,a83339a,a83342a,a83345a,a83346a,a83347a,a83350a,a83353a,a83354a,a83357a,a83360a,a83361a,a83362a,a83365a,a83368a,a83369a,a83372a,a83375a,a83376a,a83377a,a83380a,a83383a,a83384a,a83387a,a83390a,a83391a,a83392a,a83395a,a83398a,a83399a,a83402a,a83405a,a83406a,a83407a,a83410a,a83413a,a83414a,a83417a,a83420a,a83421a,a83422a,a83425a,a83428a,a83429a,a83432a,a83435a,a83436a,a83437a,a83440a,a83443a,a83444a,a83447a,a83450a,a83451a,a83452a,a83455a,a83458a,a83459a,a83462a,a83465a,a83466a,a83467a,a83470a,a83473a,a83474a,a83477a,a83480a,a83481a,a83482a,a83485a,a83488a,a83489a,a83492a,a83495a,a83496a,a83497a,a83500a,a83503a,a83504a,a83507a,a83510a,a83511a,a83512a,a83515a,a83518a,a83519a,a83522a,a83525a,a83526a,a83527a,a83530a,a83533a,a83534a,a83537a,a83540a,a83541a,a83542a,a83545a,a83548a,a83549a,a83552a,a83555a,a83556a,a83557a,a83560a,a83563a,a83564a,a83567a,a83570a,a83571a,a83572a,a83575a,a83578a,a83579a,a83582a,a83585a,a83586a,a83587a,a83590a,a83593a,a83594a,a83597a,a83600a,a83601a,a83602a,a83605a,a83608a,a83609a,a83612a,a83615a,a83616a,a83617a,a83620a,a83623a,a83624a,a83627a,a83630a,a83631a,a83632a,a83635a,a83638a,a83639a,a83642a,a83645a,a83646a,a83647a,a83650a,a83653a,a83654a,a83657a,a83660a,a83661a,a83662a,a83665a,a83668a,a83669a,a83672a,a83675a,a83676a,a83677a,a83680a,a83683a,a83684a,a83687a,a83690a,a83691a,a83692a,a83695a,a83698a,a83699a,a83702a,a83705a,a83706a,a83707a,a83710a,a83713a,a83714a,a83717a,a83720a,a83721a,a83722a,a83725a,a83728a,a83729a,a83732a,a83735a,a83736a,a83737a,a83740a,a83743a,a83744a,a83747a,a83750a,a83751a,a83752a,a83755a,a83758a,a83759a,a83762a,a83765a,a83766a,a83767a,a83770a,a83773a,a83774a,a83777a,a83780a,a83781a,a83782a,a83785a,a83788a,a83789a,a83792a,a83795a,a83796a,a83797a,a83800a,a83803a,a83804a,a83807a,a83810a,a83811a,a83812a,a83815a,a83818a,a83819a,a83822a,a83825a,a83826a,a83827a,a83830a,a83833a,a83834a,a83837a,a83840a,a83841a,a83842a,a83845a,a83848a,a83849a,a83852a,a83855a,a83856a,a83857a,a83860a,a83863a,a83864a,a83867a,a83870a,a83871a,a83872a,a83875a,a83878a,a83879a,a83882a,a83885a,a83886a,a83887a,a83890a,a83893a,a83894a,a83897a,a83900a,a83901a,a83902a,a83905a,a83908a,a83909a,a83912a,a83915a,a83916a,a83917a,a83920a,a83923a,a83924a,a83927a,a83930a,a83931a,a83932a,a83935a,a83938a,a83939a,a83942a,a83945a,a83946a,a83947a,a83950a,a83953a,a83954a,a83957a,a83960a,a83961a,a83962a,a83965a,a83968a,a83969a,a83972a,a83975a,a83976a,a83977a,a83980a,a83983a,a83984a,a83987a,a83990a,a83991a,a83992a,a83995a,a83998a,a83999a,a84002a,a84005a,a84006a,a84007a,a84010a,a84013a,a84014a,a84017a,a84020a,a84021a,a84022a,a84025a,a84028a,a84029a,a84032a,a84035a,a84036a,a84037a,a84040a,a84043a,a84044a,a84047a,a84050a,a84051a,a84052a,a84055a,a84058a,a84059a,a84062a,a84065a,a84066a,a84067a,a84070a,a84073a,a84074a,a84077a,a84080a,a84081a,a84082a,a84085a,a84088a,a84089a,a84092a,a84095a,a84096a,a84097a,a84100a,a84103a,a84104a,a84107a,a84110a,a84111a,a84112a,a84115a,a84118a,a84119a,a84122a,a84125a,a84126a,a84127a,a84130a,a84133a,a84134a,a84137a,a84140a,a84141a,a84142a,a84145a,a84148a,a84149a,a84152a,a84155a,a84156a,a84157a,a84160a,a84163a,a84164a,a84167a,a84170a,a84171a,a84172a,a84175a,a84178a,a84179a,a84182a,a84185a,a84186a,a84187a,a84190a,a84193a,a84194a,a84197a,a84200a,a84201a,a84202a,a84205a,a84208a,a84209a,a84212a,a84215a,a84216a,a84217a,a84220a,a84223a,a84224a,a84227a,a84230a,a84231a,a84232a,a84235a,a84238a,a84239a,a84242a,a84245a,a84246a,a84247a,a84250a,a84253a,a84254a,a84257a,a84260a,a84261a,a84262a,a84265a,a84268a,a84269a,a84272a,a84275a,a84276a,a84277a,a84280a,a84283a,a84284a,a84287a,a84290a,a84291a,a84292a,a84295a,a84298a,a84299a,a84302a,a84305a,a84306a,a84307a,a84310a,a84313a,a84314a,a84317a,a84320a,a84321a,a84322a,a84325a,a84328a,a84329a,a84332a,a84335a,a84336a,a84337a,a84340a,a84343a,a84344a,a84347a,a84350a,a84351a,a84352a,a84355a,a84358a,a84359a,a84362a,a84365a,a84366a,a84367a,a84370a,a84373a,a84374a,a84377a,a84380a,a84381a,a84382a,a84385a,a84388a,a84389a,a84392a,a84395a,a84396a,a84397a,a84400a,a84403a,a84404a,a84407a,a84410a,a84411a,a84412a,a84415a,a84418a,a84419a,a84422a,a84425a,a84426a,a84427a,a84430a,a84433a,a84434a,a84437a,a84440a,a84441a,a84442a,a84445a,a84448a,a84449a,a84452a,a84455a,a84456a,a84457a,a84460a,a84463a,a84464a,a84467a,a84470a,a84471a,a84472a,a84475a,a84478a,a84479a,a84482a,a84485a,a84486a,a84487a,a84490a,a84493a,a84494a,a84497a,a84500a,a84501a,a84502a,a84505a,a84508a,a84509a,a84512a,a84515a,a84516a,a84517a,a84520a,a84523a,a84524a,a84527a,a84530a,a84531a,a84532a,a84535a,a84538a,a84539a,a84542a,a84545a,a84546a,a84547a,a84550a,a84553a,a84554a,a84557a,a84560a,a84561a,a84562a,a84565a,a84568a,a84569a,a84572a,a84575a,a84576a,a84577a,a84580a,a84583a,a84584a,a84587a,a84590a,a84591a,a84592a,a84595a,a84598a,a84599a,a84602a,a84605a,a84606a,a84607a,a84610a,a84613a,a84614a,a84617a,a84620a,a84621a,a84622a,a84625a,a84628a,a84629a,a84632a,a84635a,a84636a,a84637a,a84640a,a84643a,a84644a,a84647a,a84650a,a84651a,a84652a,a84655a,a84658a,a84659a,a84662a,a84665a,a84666a,a84667a,a84670a,a84673a,a84674a,a84677a,a84680a,a84681a,a84682a,a84685a,a84688a,a84689a,a84692a,a84695a,a84696a,a84697a,a84700a,a84703a,a84704a,a84707a,a84710a,a84711a,a84712a,a84715a,a84718a,a84719a,a84722a,a84725a,a84726a,a84727a,a84730a,a84733a,a84734a,a84737a,a84740a,a84741a,a84742a,a84745a,a84748a,a84749a,a84752a,a84755a,a84756a,a84757a,a84760a,a84763a,a84764a,a84767a,a84770a,a84771a,a84772a,a84775a,a84778a,a84779a,a84782a,a84785a,a84786a,a84787a,a84790a,a84793a,a84794a,a84797a,a84800a,a84801a,a84802a,a84805a,a84808a,a84809a,a84812a,a84815a,a84816a,a84817a,a84820a,a84823a,a84824a,a84827a,a84830a,a84831a,a84832a,a84835a,a84838a,a84839a,a84842a,a84845a,a84846a,a84847a,a84850a,a84853a,a84854a,a84857a,a84860a,a84861a,a84862a,a84865a,a84868a,a84869a,a84872a,a84875a,a84876a,a84877a,a84880a,a84883a,a84884a,a84887a,a84890a,a84891a,a84892a,a84895a,a84898a,a84899a,a84902a,a84905a,a84906a,a84907a,a84910a,a84913a,a84914a,a84917a,a84920a,a84921a,a84922a,a84925a,a84928a,a84929a,a84932a,a84935a,a84936a,a84937a,a84940a,a84943a,a84944a,a84947a,a84950a,a84951a,a84952a,a84955a,a84958a,a84959a,a84962a,a84965a,a84966a,a84967a,a84970a,a84973a,a84974a,a84977a,a84981a,a84982a,a84983a,a84984a,a84987a,a84990a,a84991a,a84994a,a84997a,a84998a,a84999a,a85002a,a85005a,a85006a,a85009a,a85013a,a85014a,a85015a,a85016a,a85019a,a85022a,a85023a,a85026a,a85029a,a85030a,a85031a,a85034a,a85037a,a85038a,a85041a,a85045a,a85046a,a85047a,a85048a,a85051a,a85054a,a85055a,a85058a,a85061a,a85062a,a85063a,a85066a,a85069a,a85070a,a85073a,a85077a,a85078a,a85079a,a85080a,a85083a,a85086a,a85087a,a85090a,a85093a,a85094a,a85095a,a85098a,a85101a,a85102a,a85105a,a85109a,a85110a,a85111a,a85112a,a85115a,a85118a,a85119a,a85122a,a85125a,a85126a,a85127a,a85130a,a85133a,a85134a,a85137a,a85141a,a85142a,a85143a,a85144a,a85147a,a85150a,a85151a,a85154a,a85157a,a85158a,a85159a,a85162a,a85165a,a85166a,a85169a,a85173a,a85174a,a85175a,a85176a,a85179a,a85182a,a85183a,a85186a,a85189a,a85190a,a85191a,a85194a,a85197a,a85198a,a85201a,a85205a,a85206a,a85207a,a85208a,a85211a,a85214a,a85215a,a85218a,a85221a,a85222a,a85223a,a85226a,a85229a,a85230a,a85233a,a85237a,a85238a,a85239a,a85240a,a85243a,a85246a,a85247a,a85250a,a85253a,a85254a,a85255a,a85258a,a85261a,a85262a,a85265a,a85269a,a85270a,a85271a,a85272a,a85275a,a85278a,a85279a,a85282a,a85285a,a85286a,a85287a,a85290a,a85293a,a85294a,a85297a,a85301a,a85302a,a85303a,a85304a,a85307a,a85310a,a85311a,a85314a,a85317a,a85318a,a85319a,a85322a,a85325a,a85326a,a85329a,a85333a,a85334a,a85335a,a85336a,a85339a,a85342a,a85343a,a85346a,a85349a,a85350a,a85351a,a85354a,a85357a,a85358a,a85361a,a85365a,a85366a,a85367a,a85368a,a85371a,a85374a,a85375a,a85378a,a85381a,a85382a,a85383a,a85386a,a85389a,a85390a,a85393a,a85397a,a85398a,a85399a,a85400a,a85403a,a85406a,a85407a,a85410a,a85413a,a85414a,a85415a,a85418a,a85421a,a85422a,a85425a,a85429a,a85430a,a85431a,a85432a,a85435a,a85438a,a85439a,a85442a,a85445a,a85446a,a85447a,a85450a,a85453a,a85454a,a85457a,a85461a,a85462a,a85463a,a85464a,a85467a,a85470a,a85471a,a85474a,a85477a,a85478a,a85479a,a85482a,a85485a,a85486a,a85489a,a85493a,a85494a,a85495a,a85496a,a85499a,a85502a,a85503a,a85506a,a85509a,a85510a,a85511a,a85514a,a85517a,a85518a,a85521a,a85525a,a85526a,a85527a,a85528a,a85531a,a85534a,a85535a,a85538a,a85541a,a85542a,a85543a,a85546a,a85549a,a85550a,a85553a,a85557a,a85558a,a85559a,a85560a,a85563a,a85566a,a85567a,a85570a,a85573a,a85574a,a85575a,a85578a,a85581a,a85582a,a85585a,a85589a,a85590a,a85591a,a85592a,a85595a,a85598a,a85599a,a85602a,a85605a,a85606a,a85607a,a85610a,a85613a,a85614a,a85617a,a85621a,a85622a,a85623a,a85624a,a85627a,a85630a,a85631a,a85634a,a85637a,a85638a,a85639a,a85642a,a85645a,a85646a,a85649a,a85653a,a85654a,a85655a,a85656a,a85659a,a85662a,a85663a,a85666a,a85669a,a85670a,a85671a,a85674a,a85677a,a85678a,a85681a,a85685a,a85686a,a85687a,a85688a,a85691a,a85694a,a85695a,a85698a,a85701a,a85702a,a85703a,a85706a,a85709a,a85710a,a85713a,a85717a,a85718a,a85719a,a85720a,a85723a,a85726a,a85727a,a85730a,a85733a,a85734a,a85735a,a85738a,a85741a,a85742a,a85745a,a85749a,a85750a,a85751a,a85752a,a85755a,a85758a,a85759a,a85762a,a85765a,a85766a,a85767a,a85770a,a85773a,a85774a,a85777a,a85781a,a85782a,a85783a,a85784a,a85787a,a85790a,a85791a,a85794a,a85797a,a85798a,a85799a,a85802a,a85805a,a85806a,a85809a,a85813a,a85814a,a85815a,a85816a,a85819a,a85822a,a85823a,a85826a,a85829a,a85830a,a85831a,a85834a,a85837a,a85838a,a85841a,a85845a,a85846a,a85847a,a85848a,a85851a,a85854a,a85855a,a85858a,a85861a,a85862a,a85863a,a85866a,a85869a,a85870a,a85873a,a85877a,a85878a,a85879a,a85880a,a85883a,a85886a,a85887a,a85890a,a85893a,a85894a,a85895a,a85898a,a85901a,a85902a,a85905a,a85909a,a85910a,a85911a,a85912a,a85915a,a85918a,a85919a,a85922a,a85925a,a85926a,a85927a,a85930a,a85933a,a85934a,a85937a,a85941a,a85942a,a85943a,a85944a,a85947a,a85950a,a85951a,a85954a,a85957a,a85958a,a85959a,a85962a,a85965a,a85966a,a85969a,a85973a,a85974a,a85975a,a85976a,a85979a,a85982a,a85983a,a85986a,a85989a,a85990a,a85991a,a85994a,a85997a,a85998a,a86001a,a86005a,a86006a,a86007a,a86008a,a86011a,a86014a,a86015a,a86018a,a86021a,a86022a,a86023a,a86026a,a86029a,a86030a,a86033a,a86037a,a86038a,a86039a,a86040a,a86043a,a86046a,a86047a,a86050a,a86053a,a86054a,a86055a,a86058a,a86061a,a86062a,a86065a,a86069a,a86070a,a86071a,a86072a,a86075a,a86078a,a86079a,a86082a,a86085a,a86086a,a86087a,a86090a,a86093a,a86094a,a86097a,a86101a,a86102a,a86103a,a86104a,a86107a,a86110a,a86111a,a86114a,a86117a,a86118a,a86119a,a86122a,a86125a,a86126a,a86129a,a86133a,a86134a,a86135a,a86136a,a86139a,a86142a,a86143a,a86146a,a86149a,a86150a,a86151a,a86154a,a86157a,a86158a,a86161a,a86165a,a86166a,a86167a,a86168a,a86171a,a86174a,a86175a,a86178a,a86181a,a86182a,a86183a,a86186a,a86189a,a86190a,a86193a,a86197a,a86198a,a86199a,a86200a,a86203a,a86206a,a86207a,a86210a,a86213a,a86214a,a86215a,a86218a,a86221a,a86222a,a86225a,a86229a,a86230a,a86231a,a86232a,a86235a,a86238a,a86239a,a86242a,a86245a,a86246a,a86247a,a86250a,a86253a,a86254a,a86257a,a86261a,a86262a,a86263a,a86264a,a86267a,a86270a,a86271a,a86274a,a86277a,a86278a,a86279a,a86282a,a86285a,a86286a,a86289a,a86293a,a86294a,a86295a,a86296a,a86299a,a86302a,a86303a,a86306a,a86309a,a86310a,a86311a,a86314a,a86317a,a86318a,a86321a,a86325a,a86326a,a86327a,a86328a,a86331a,a86334a,a86335a,a86338a,a86341a,a86342a,a86343a,a86346a,a86349a,a86350a,a86353a,a86357a,a86358a,a86359a,a86360a,a86363a,a86366a,a86367a,a86370a,a86373a,a86374a,a86375a,a86378a,a86381a,a86382a,a86385a,a86389a,a86390a,a86391a,a86392a,a86395a,a86398a,a86399a,a86402a,a86405a,a86406a,a86407a,a86410a,a86413a,a86414a,a86417a,a86421a,a86422a,a86423a,a86424a,a86427a,a86430a,a86431a,a86434a,a86437a,a86438a,a86439a,a86442a,a86445a,a86446a,a86449a,a86453a,a86454a,a86455a,a86456a,a86459a,a86462a,a86463a,a86466a,a86469a,a86470a,a86471a,a86474a,a86477a,a86478a,a86481a,a86485a,a86486a,a86487a,a86488a,a86491a,a86494a,a86495a,a86498a,a86501a,a86502a,a86503a,a86506a,a86509a,a86510a,a86513a,a86517a,a86518a,a86519a,a86520a,a86523a,a86526a,a86527a,a86530a,a86533a,a86534a,a86535a,a86538a,a86541a,a86542a,a86545a,a86549a,a86550a,a86551a,a86552a,a86555a,a86558a,a86559a,a86562a,a86565a,a86566a,a86567a,a86570a,a86573a,a86574a,a86577a,a86581a,a86582a,a86583a,a86584a,a86587a,a86590a,a86591a,a86594a,a86597a,a86598a,a86599a,a86602a,a86605a,a86606a,a86609a,a86613a,a86614a,a86615a,a86616a,a86619a,a86622a,a86623a,a86626a,a86629a,a86630a,a86631a,a86634a,a86637a,a86638a,a86641a,a86645a,a86646a,a86647a,a86648a,a86651a,a86654a,a86655a,a86658a,a86661a,a86662a,a86663a,a86666a,a86669a,a86670a,a86673a,a86677a,a86678a,a86679a,a86680a,a86683a,a86686a,a86687a,a86690a,a86693a,a86694a,a86695a,a86698a,a86701a,a86702a,a86705a,a86709a,a86710a,a86711a,a86712a,a86715a,a86718a,a86719a,a86722a,a86725a,a86726a,a86727a,a86730a,a86733a,a86734a,a86737a,a86741a,a86742a,a86743a,a86744a,a86747a,a86750a,a86751a,a86754a,a86757a,a86758a,a86759a,a86762a,a86765a,a86766a,a86769a,a86773a,a86774a,a86775a,a86776a,a86779a,a86782a,a86783a,a86786a,a86789a,a86790a,a86791a,a86794a,a86797a,a86798a,a86801a,a86805a,a86806a,a86807a,a86808a,a86811a,a86814a,a86815a,a86818a,a86821a,a86822a,a86823a,a86826a,a86829a,a86830a,a86833a,a86837a,a86838a,a86839a,a86840a,a86843a,a86846a,a86847a,a86850a,a86853a,a86854a,a86855a,a86858a,a86861a,a86862a,a86865a,a86869a,a86870a,a86871a,a86872a,a86875a,a86878a,a86879a,a86882a,a86885a,a86886a,a86887a,a86890a,a86893a,a86894a,a86897a,a86901a,a86902a,a86903a,a86904a,a86907a,a86910a,a86911a,a86914a,a86917a,a86918a,a86919a,a86922a,a86925a,a86926a,a86929a,a86933a,a86934a,a86935a,a86936a,a86939a,a86942a,a86943a,a86946a,a86949a,a86950a,a86951a,a86954a,a86957a,a86958a,a86961a,a86965a,a86966a,a86967a,a86968a,a86971a,a86974a,a86975a,a86978a,a86981a,a86982a,a86983a,a86986a,a86989a,a86990a,a86993a,a86997a,a86998a,a86999a,a87000a,a87003a,a87006a,a87007a,a87010a,a87013a,a87014a,a87015a,a87018a,a87021a,a87022a,a87025a,a87029a,a87030a,a87031a,a87032a,a87035a,a87038a,a87039a,a87042a,a87045a,a87046a,a87047a,a87050a,a87053a,a87054a,a87057a,a87061a,a87062a,a87063a,a87064a,a87067a,a87070a,a87071a,a87074a,a87077a,a87078a,a87079a,a87082a,a87085a,a87086a,a87089a,a87093a,a87094a,a87095a,a87096a,a87099a,a87102a,a87103a,a87106a,a87109a,a87110a,a87111a,a87114a,a87117a,a87118a,a87121a,a87125a,a87126a,a87127a,a87128a,a87131a,a87134a,a87135a,a87138a,a87141a,a87142a,a87143a,a87146a,a87149a,a87150a,a87153a,a87157a,a87158a,a87159a,a87160a,a87163a,a87166a,a87167a,a87170a,a87173a,a87174a,a87175a,a87178a,a87181a,a87182a,a87185a,a87189a,a87190a,a87191a,a87192a,a87195a,a87198a,a87199a,a87202a,a87205a,a87206a,a87207a,a87210a,a87213a,a87214a,a87217a,a87221a,a87222a,a87223a,a87224a,a87227a,a87230a,a87231a,a87234a,a87237a,a87238a,a87239a,a87242a,a87245a,a87246a,a87249a,a87253a,a87254a,a87255a,a87256a,a87259a,a87262a,a87263a,a87266a,a87269a,a87270a,a87271a,a87274a,a87277a,a87278a,a87281a,a87285a,a87286a,a87287a,a87288a,a87291a,a87294a,a87295a,a87298a,a87301a,a87302a,a87303a,a87306a,a87309a,a87310a,a87313a,a87317a,a87318a,a87319a,a87320a,a87323a,a87326a,a87327a,a87330a,a87333a,a87334a,a87335a,a87338a,a87341a,a87342a,a87345a,a87349a,a87350a,a87351a,a87352a,a87355a,a87358a,a87359a,a87362a,a87365a,a87366a,a87367a,a87370a,a87373a,a87374a,a87377a,a87381a,a87382a,a87383a,a87384a,a87387a,a87390a,a87391a,a87394a,a87397a,a87398a,a87399a,a87402a,a87405a,a87406a,a87409a,a87413a,a87414a,a87415a,a87416a,a87419a,a87422a,a87423a,a87426a,a87429a,a87430a,a87431a,a87434a,a87437a,a87438a,a87441a,a87445a,a87446a,a87447a,a87448a,a87451a,a87454a,a87455a,a87458a,a87461a,a87462a,a87463a,a87466a,a87469a,a87470a,a87473a,a87477a,a87478a,a87479a,a87480a,a87483a,a87486a,a87487a,a87490a,a87493a,a87494a,a87495a,a87498a,a87501a,a87502a,a87505a,a87509a,a87510a,a87511a,a87512a,a87515a,a87518a,a87519a,a87522a,a87525a,a87526a,a87527a,a87530a,a87533a,a87534a,a87537a,a87541a,a87542a,a87543a,a87544a,a87547a,a87550a,a87551a,a87554a,a87557a,a87558a,a87559a,a87562a,a87565a,a87566a,a87569a,a87573a,a87574a,a87575a,a87576a,a87579a,a87582a,a87583a,a87586a,a87589a,a87590a,a87591a,a87594a,a87597a,a87598a,a87601a,a87605a,a87606a,a87607a,a87608a,a87611a,a87614a,a87615a,a87618a,a87621a,a87622a,a87623a,a87626a,a87629a,a87630a,a87633a,a87637a,a87638a,a87639a,a87640a,a87643a,a87646a,a87647a,a87650a,a87653a,a87654a,a87655a,a87658a,a87661a,a87662a,a87665a,a87669a,a87670a,a87671a,a87672a,a87675a,a87678a,a87679a,a87682a,a87685a,a87686a,a87687a,a87690a,a87693a,a87694a,a87697a,a87701a,a87702a,a87703a,a87704a,a87707a,a87710a,a87711a,a87714a,a87717a,a87718a,a87719a,a87722a,a87725a,a87726a,a87729a,a87733a,a87734a,a87735a,a87736a,a87739a,a87742a,a87743a,a87746a,a87749a,a87750a,a87751a,a87754a,a87757a,a87758a,a87761a,a87765a,a87766a,a87767a,a87768a,a87771a,a87774a,a87775a,a87778a,a87781a,a87782a,a87783a,a87786a,a87789a,a87790a,a87793a,a87797a,a87798a,a87799a,a87800a,a87803a,a87806a,a87807a,a87810a,a87813a,a87814a,a87815a,a87818a,a87821a,a87822a,a87825a,a87829a,a87830a,a87831a,a87832a,a87835a,a87838a,a87839a,a87842a,a87845a,a87846a,a87847a,a87850a,a87853a,a87854a,a87857a,a87861a,a87862a,a87863a,a87864a,a87867a,a87870a,a87871a,a87874a,a87877a,a87878a,a87879a,a87882a,a87885a,a87886a,a87889a,a87893a,a87894a,a87895a,a87896a,a87899a,a87902a,a87903a,a87906a,a87909a,a87910a,a87911a,a87914a,a87917a,a87918a,a87921a,a87925a,a87926a,a87927a,a87928a,a87931a,a87934a,a87935a,a87938a,a87941a,a87942a,a87943a,a87946a,a87949a,a87950a,a87953a,a87957a,a87958a,a87959a,a87960a,a87963a,a87966a,a87967a,a87970a,a87973a,a87974a,a87975a,a87978a,a87981a,a87982a,a87985a,a87989a,a87990a,a87991a,a87992a,a87995a,a87998a,a87999a,a88002a,a88005a,a88006a,a88007a,a88010a,a88013a,a88014a,a88017a,a88021a,a88022a,a88023a,a88024a,a88027a,a88030a,a88031a,a88034a,a88037a,a88038a,a88039a,a88042a,a88045a,a88046a,a88049a,a88053a,a88054a,a88055a,a88056a,a88059a,a88062a,a88063a,a88066a,a88069a,a88070a,a88071a,a88074a,a88077a,a88078a,a88081a,a88085a,a88086a,a88087a,a88088a,a88091a,a88094a,a88095a,a88098a,a88101a,a88102a,a88103a,a88106a,a88109a,a88110a,a88113a,a88117a,a88118a,a88119a,a88120a,a88123a,a88126a,a88127a,a88130a,a88133a,a88134a,a88135a,a88138a,a88141a,a88142a,a88145a,a88149a,a88150a,a88151a,a88152a,a88155a,a88158a,a88159a,a88162a,a88165a,a88166a,a88167a,a88170a,a88173a,a88174a,a88177a,a88181a,a88182a,a88183a,a88184a,a88187a,a88190a,a88191a,a88194a,a88197a,a88198a,a88199a,a88202a,a88205a,a88206a,a88209a,a88213a,a88214a,a88215a,a88216a,a88219a,a88222a,a88223a,a88226a,a88229a,a88230a,a88231a,a88234a,a88237a,a88238a,a88241a,a88245a,a88246a,a88247a,a88248a,a88251a,a88254a,a88255a,a88258a,a88261a,a88262a,a88263a,a88266a,a88269a,a88270a,a88273a,a88277a,a88278a,a88279a,a88280a,a88283a,a88286a,a88287a,a88290a,a88294a,a88295a,a88296a,a88297a,a88300a,a88303a,a88304a,a88307a,a88311a,a88312a,a88313a,a88314a,a88317a,a88320a,a88321a,a88324a,a88328a,a88329a,a88330a,a88331a,a88334a,a88337a,a88338a,a88341a,a88345a,a88346a,a88347a,a88348a,a88351a,a88354a,a88355a,a88358a,a88362a,a88363a,a88364a,a88365a,a88368a,a88371a,a88372a,a88375a,a88379a,a88380a,a88381a,a88382a,a88385a,a88388a,a88389a,a88392a,a88396a,a88397a,a88398a,a88399a,a88402a,a88405a,a88406a,a88409a,a88413a,a88414a,a88415a,a88416a,a88419a,a88422a,a88423a,a88426a,a88430a,a88431a,a88432a,a88433a,a88436a,a88439a,a88440a,a88443a,a88447a,a88448a,a88449a,a88450a,a88453a,a88456a,a88457a,a88460a,a88464a,a88465a,a88466a,a88467a,a88470a,a88473a,a88474a,a88477a,a88481a,a88482a,a88483a,a88484a,a88487a,a88490a,a88491a,a88494a,a88498a,a88499a,a88500a,a88501a,a88504a,a88507a,a88508a,a88511a,a88515a,a88516a,a88517a,a88518a,a88521a,a88524a,a88525a,a88528a,a88532a,a88533a,a88534a,a88535a,a88538a,a88541a,a88542a,a88545a,a88549a,a88550a,a88551a,a88552a,a88555a,a88558a,a88559a,a88562a,a88566a,a88567a,a88568a,a88569a,a88572a,a88575a,a88576a,a88579a,a88583a,a88584a,a88585a,a88586a,a88589a,a88592a,a88593a,a88596a,a88600a,a88601a,a88602a,a88603a,a88606a,a88609a,a88610a,a88613a,a88617a,a88618a,a88619a,a88620a,a88623a,a88626a,a88627a,a88630a,a88634a,a88635a,a88636a,a88637a,a88640a,a88643a,a88644a,a88647a,a88651a,a88652a,a88653a,a88654a,a88657a,a88660a,a88661a,a88664a,a88668a,a88669a,a88670a,a88671a,a88674a,a88677a,a88678a,a88681a,a88685a,a88686a,a88687a,a88688a: std_logic;
begin

A105 <=( a9520a ) or ( a6347a );
 a1a <=( a88688a  and  a88671a );
 a2a <=( a88654a  and  a88637a );
 a3a <=( a88620a  and  a88603a );
 a4a <=( a88586a  and  a88569a );
 a5a <=( a88552a  and  a88535a );
 a6a <=( a88518a  and  a88501a );
 a7a <=( a88484a  and  a88467a );
 a8a <=( a88450a  and  a88433a );
 a9a <=( a88416a  and  a88399a );
 a10a <=( a88382a  and  a88365a );
 a11a <=( a88348a  and  a88331a );
 a12a <=( a88314a  and  a88297a );
 a13a <=( a88280a  and  a88263a );
 a14a <=( a88248a  and  a88231a );
 a15a <=( a88216a  and  a88199a );
 a16a <=( a88184a  and  a88167a );
 a17a <=( a88152a  and  a88135a );
 a18a <=( a88120a  and  a88103a );
 a19a <=( a88088a  and  a88071a );
 a20a <=( a88056a  and  a88039a );
 a21a <=( a88024a  and  a88007a );
 a22a <=( a87992a  and  a87975a );
 a23a <=( a87960a  and  a87943a );
 a24a <=( a87928a  and  a87911a );
 a25a <=( a87896a  and  a87879a );
 a26a <=( a87864a  and  a87847a );
 a27a <=( a87832a  and  a87815a );
 a28a <=( a87800a  and  a87783a );
 a29a <=( a87768a  and  a87751a );
 a30a <=( a87736a  and  a87719a );
 a31a <=( a87704a  and  a87687a );
 a32a <=( a87672a  and  a87655a );
 a33a <=( a87640a  and  a87623a );
 a34a <=( a87608a  and  a87591a );
 a35a <=( a87576a  and  a87559a );
 a36a <=( a87544a  and  a87527a );
 a37a <=( a87512a  and  a87495a );
 a38a <=( a87480a  and  a87463a );
 a39a <=( a87448a  and  a87431a );
 a40a <=( a87416a  and  a87399a );
 a41a <=( a87384a  and  a87367a );
 a42a <=( a87352a  and  a87335a );
 a43a <=( a87320a  and  a87303a );
 a44a <=( a87288a  and  a87271a );
 a45a <=( a87256a  and  a87239a );
 a46a <=( a87224a  and  a87207a );
 a47a <=( a87192a  and  a87175a );
 a48a <=( a87160a  and  a87143a );
 a49a <=( a87128a  and  a87111a );
 a50a <=( a87096a  and  a87079a );
 a51a <=( a87064a  and  a87047a );
 a52a <=( a87032a  and  a87015a );
 a53a <=( a87000a  and  a86983a );
 a54a <=( a86968a  and  a86951a );
 a55a <=( a86936a  and  a86919a );
 a56a <=( a86904a  and  a86887a );
 a57a <=( a86872a  and  a86855a );
 a58a <=( a86840a  and  a86823a );
 a59a <=( a86808a  and  a86791a );
 a60a <=( a86776a  and  a86759a );
 a61a <=( a86744a  and  a86727a );
 a62a <=( a86712a  and  a86695a );
 a63a <=( a86680a  and  a86663a );
 a64a <=( a86648a  and  a86631a );
 a65a <=( a86616a  and  a86599a );
 a66a <=( a86584a  and  a86567a );
 a67a <=( a86552a  and  a86535a );
 a68a <=( a86520a  and  a86503a );
 a69a <=( a86488a  and  a86471a );
 a70a <=( a86456a  and  a86439a );
 a71a <=( a86424a  and  a86407a );
 a72a <=( a86392a  and  a86375a );
 a73a <=( a86360a  and  a86343a );
 a74a <=( a86328a  and  a86311a );
 a75a <=( a86296a  and  a86279a );
 a76a <=( a86264a  and  a86247a );
 a77a <=( a86232a  and  a86215a );
 a78a <=( a86200a  and  a86183a );
 a79a <=( a86168a  and  a86151a );
 a80a <=( a86136a  and  a86119a );
 a81a <=( a86104a  and  a86087a );
 a82a <=( a86072a  and  a86055a );
 a83a <=( a86040a  and  a86023a );
 a84a <=( a86008a  and  a85991a );
 a85a <=( a85976a  and  a85959a );
 a86a <=( a85944a  and  a85927a );
 a87a <=( a85912a  and  a85895a );
 a88a <=( a85880a  and  a85863a );
 a89a <=( a85848a  and  a85831a );
 a90a <=( a85816a  and  a85799a );
 a91a <=( a85784a  and  a85767a );
 a92a <=( a85752a  and  a85735a );
 a93a <=( a85720a  and  a85703a );
 a94a <=( a85688a  and  a85671a );
 a95a <=( a85656a  and  a85639a );
 a96a <=( a85624a  and  a85607a );
 a97a <=( a85592a  and  a85575a );
 a98a <=( a85560a  and  a85543a );
 a99a <=( a85528a  and  a85511a );
 a100a <=( a85496a  and  a85479a );
 a101a <=( a85464a  and  a85447a );
 a102a <=( a85432a  and  a85415a );
 a103a <=( a85400a  and  a85383a );
 a104a <=( a85368a  and  a85351a );
 a105a <=( a85336a  and  a85319a );
 a106a <=( a85304a  and  a85287a );
 a107a <=( a85272a  and  a85255a );
 a108a <=( a85240a  and  a85223a );
 a109a <=( a85208a  and  a85191a );
 a110a <=( a85176a  and  a85159a );
 a111a <=( a85144a  and  a85127a );
 a112a <=( a85112a  and  a85095a );
 a113a <=( a85080a  and  a85063a );
 a114a <=( a85048a  and  a85031a );
 a115a <=( a85016a  and  a84999a );
 a116a <=( a84984a  and  a84967a );
 a117a <=( a84952a  and  a84937a );
 a118a <=( a84922a  and  a84907a );
 a119a <=( a84892a  and  a84877a );
 a120a <=( a84862a  and  a84847a );
 a121a <=( a84832a  and  a84817a );
 a122a <=( a84802a  and  a84787a );
 a123a <=( a84772a  and  a84757a );
 a124a <=( a84742a  and  a84727a );
 a125a <=( a84712a  and  a84697a );
 a126a <=( a84682a  and  a84667a );
 a127a <=( a84652a  and  a84637a );
 a128a <=( a84622a  and  a84607a );
 a129a <=( a84592a  and  a84577a );
 a130a <=( a84562a  and  a84547a );
 a131a <=( a84532a  and  a84517a );
 a132a <=( a84502a  and  a84487a );
 a133a <=( a84472a  and  a84457a );
 a134a <=( a84442a  and  a84427a );
 a135a <=( a84412a  and  a84397a );
 a136a <=( a84382a  and  a84367a );
 a137a <=( a84352a  and  a84337a );
 a138a <=( a84322a  and  a84307a );
 a139a <=( a84292a  and  a84277a );
 a140a <=( a84262a  and  a84247a );
 a141a <=( a84232a  and  a84217a );
 a142a <=( a84202a  and  a84187a );
 a143a <=( a84172a  and  a84157a );
 a144a <=( a84142a  and  a84127a );
 a145a <=( a84112a  and  a84097a );
 a146a <=( a84082a  and  a84067a );
 a147a <=( a84052a  and  a84037a );
 a148a <=( a84022a  and  a84007a );
 a149a <=( a83992a  and  a83977a );
 a150a <=( a83962a  and  a83947a );
 a151a <=( a83932a  and  a83917a );
 a152a <=( a83902a  and  a83887a );
 a153a <=( a83872a  and  a83857a );
 a154a <=( a83842a  and  a83827a );
 a155a <=( a83812a  and  a83797a );
 a156a <=( a83782a  and  a83767a );
 a157a <=( a83752a  and  a83737a );
 a158a <=( a83722a  and  a83707a );
 a159a <=( a83692a  and  a83677a );
 a160a <=( a83662a  and  a83647a );
 a161a <=( a83632a  and  a83617a );
 a162a <=( a83602a  and  a83587a );
 a163a <=( a83572a  and  a83557a );
 a164a <=( a83542a  and  a83527a );
 a165a <=( a83512a  and  a83497a );
 a166a <=( a83482a  and  a83467a );
 a167a <=( a83452a  and  a83437a );
 a168a <=( a83422a  and  a83407a );
 a169a <=( a83392a  and  a83377a );
 a170a <=( a83362a  and  a83347a );
 a171a <=( a83332a  and  a83317a );
 a172a <=( a83302a  and  a83287a );
 a173a <=( a83272a  and  a83257a );
 a174a <=( a83242a  and  a83227a );
 a175a <=( a83212a  and  a83197a );
 a176a <=( a83182a  and  a83167a );
 a177a <=( a83152a  and  a83137a );
 a178a <=( a83122a  and  a83107a );
 a179a <=( a83092a  and  a83077a );
 a180a <=( a83062a  and  a83047a );
 a181a <=( a83032a  and  a83017a );
 a182a <=( a83002a  and  a82987a );
 a183a <=( a82972a  and  a82957a );
 a184a <=( a82942a  and  a82927a );
 a185a <=( a82912a  and  a82897a );
 a186a <=( a82882a  and  a82867a );
 a187a <=( a82852a  and  a82837a );
 a188a <=( a82822a  and  a82807a );
 a189a <=( a82792a  and  a82777a );
 a190a <=( a82762a  and  a82747a );
 a191a <=( a82732a  and  a82717a );
 a192a <=( a82702a  and  a82687a );
 a193a <=( a82672a  and  a82657a );
 a194a <=( a82642a  and  a82627a );
 a195a <=( a82612a  and  a82597a );
 a196a <=( a82582a  and  a82567a );
 a197a <=( a82552a  and  a82537a );
 a198a <=( a82522a  and  a82507a );
 a199a <=( a82492a  and  a82477a );
 a200a <=( a82462a  and  a82447a );
 a201a <=( a82432a  and  a82417a );
 a202a <=( a82402a  and  a82387a );
 a203a <=( a82372a  and  a82357a );
 a204a <=( a82342a  and  a82327a );
 a205a <=( a82312a  and  a82297a );
 a206a <=( a82282a  and  a82267a );
 a207a <=( a82252a  and  a82237a );
 a208a <=( a82222a  and  a82207a );
 a209a <=( a82192a  and  a82177a );
 a210a <=( a82162a  and  a82147a );
 a211a <=( a82132a  and  a82117a );
 a212a <=( a82102a  and  a82087a );
 a213a <=( a82072a  and  a82057a );
 a214a <=( a82042a  and  a82027a );
 a215a <=( a82012a  and  a81997a );
 a216a <=( a81982a  and  a81967a );
 a217a <=( a81952a  and  a81937a );
 a218a <=( a81922a  and  a81907a );
 a219a <=( a81892a  and  a81877a );
 a220a <=( a81862a  and  a81847a );
 a221a <=( a81832a  and  a81817a );
 a222a <=( a81802a  and  a81787a );
 a223a <=( a81772a  and  a81757a );
 a224a <=( a81742a  and  a81727a );
 a225a <=( a81712a  and  a81697a );
 a226a <=( a81682a  and  a81667a );
 a227a <=( a81652a  and  a81637a );
 a228a <=( a81622a  and  a81607a );
 a229a <=( a81592a  and  a81577a );
 a230a <=( a81562a  and  a81547a );
 a231a <=( a81532a  and  a81517a );
 a232a <=( a81502a  and  a81487a );
 a233a <=( a81472a  and  a81457a );
 a234a <=( a81442a  and  a81427a );
 a235a <=( a81412a  and  a81397a );
 a236a <=( a81382a  and  a81367a );
 a237a <=( a81352a  and  a81337a );
 a238a <=( a81322a  and  a81307a );
 a239a <=( a81292a  and  a81277a );
 a240a <=( a81262a  and  a81247a );
 a241a <=( a81232a  and  a81217a );
 a242a <=( a81202a  and  a81187a );
 a243a <=( a81172a  and  a81157a );
 a244a <=( a81142a  and  a81127a );
 a245a <=( a81112a  and  a81097a );
 a246a <=( a81082a  and  a81067a );
 a247a <=( a81052a  and  a81037a );
 a248a <=( a81022a  and  a81007a );
 a249a <=( a80992a  and  a80977a );
 a250a <=( a80962a  and  a80947a );
 a251a <=( a80932a  and  a80917a );
 a252a <=( a80902a  and  a80887a );
 a253a <=( a80872a  and  a80857a );
 a254a <=( a80842a  and  a80827a );
 a255a <=( a80812a  and  a80797a );
 a256a <=( a80782a  and  a80767a );
 a257a <=( a80752a  and  a80737a );
 a258a <=( a80722a  and  a80707a );
 a259a <=( a80692a  and  a80677a );
 a260a <=( a80662a  and  a80647a );
 a261a <=( a80632a  and  a80617a );
 a262a <=( a80602a  and  a80587a );
 a263a <=( a80572a  and  a80557a );
 a264a <=( a80542a  and  a80527a );
 a265a <=( a80512a  and  a80497a );
 a266a <=( a80482a  and  a80467a );
 a267a <=( a80452a  and  a80437a );
 a268a <=( a80422a  and  a80407a );
 a269a <=( a80392a  and  a80377a );
 a270a <=( a80362a  and  a80347a );
 a271a <=( a80332a  and  a80317a );
 a272a <=( a80302a  and  a80287a );
 a273a <=( a80272a  and  a80257a );
 a274a <=( a80242a  and  a80227a );
 a275a <=( a80212a  and  a80197a );
 a276a <=( a80182a  and  a80167a );
 a277a <=( a80152a  and  a80137a );
 a278a <=( a80122a  and  a80107a );
 a279a <=( a80092a  and  a80077a );
 a280a <=( a80062a  and  a80047a );
 a281a <=( a80032a  and  a80017a );
 a282a <=( a80002a  and  a79987a );
 a283a <=( a79972a  and  a79957a );
 a284a <=( a79942a  and  a79927a );
 a285a <=( a79912a  and  a79897a );
 a286a <=( a79882a  and  a79867a );
 a287a <=( a79852a  and  a79837a );
 a288a <=( a79822a  and  a79807a );
 a289a <=( a79792a  and  a79777a );
 a290a <=( a79762a  and  a79747a );
 a291a <=( a79732a  and  a79717a );
 a292a <=( a79702a  and  a79687a );
 a293a <=( a79672a  and  a79657a );
 a294a <=( a79642a  and  a79627a );
 a295a <=( a79612a  and  a79597a );
 a296a <=( a79582a  and  a79567a );
 a297a <=( a79552a  and  a79537a );
 a298a <=( a79522a  and  a79507a );
 a299a <=( a79492a  and  a79477a );
 a300a <=( a79462a  and  a79447a );
 a301a <=( a79432a  and  a79417a );
 a302a <=( a79402a  and  a79387a );
 a303a <=( a79372a  and  a79357a );
 a304a <=( a79342a  and  a79327a );
 a305a <=( a79312a  and  a79297a );
 a306a <=( a79282a  and  a79267a );
 a307a <=( a79252a  and  a79237a );
 a308a <=( a79222a  and  a79207a );
 a309a <=( a79192a  and  a79177a );
 a310a <=( a79162a  and  a79147a );
 a311a <=( a79132a  and  a79117a );
 a312a <=( a79102a  and  a79087a );
 a313a <=( a79072a  and  a79057a );
 a314a <=( a79042a  and  a79027a );
 a315a <=( a79012a  and  a78997a );
 a316a <=( a78982a  and  a78967a );
 a317a <=( a78952a  and  a78937a );
 a318a <=( a78922a  and  a78907a );
 a319a <=( a78892a  and  a78877a );
 a320a <=( a78862a  and  a78847a );
 a321a <=( a78832a  and  a78817a );
 a322a <=( a78802a  and  a78787a );
 a323a <=( a78772a  and  a78757a );
 a324a <=( a78742a  and  a78727a );
 a325a <=( a78712a  and  a78697a );
 a326a <=( a78682a  and  a78667a );
 a327a <=( a78652a  and  a78637a );
 a328a <=( a78622a  and  a78607a );
 a329a <=( a78592a  and  a78577a );
 a330a <=( a78562a  and  a78547a );
 a331a <=( a78532a  and  a78517a );
 a332a <=( a78502a  and  a78487a );
 a333a <=( a78472a  and  a78457a );
 a334a <=( a78442a  and  a78427a );
 a335a <=( a78412a  and  a78397a );
 a336a <=( a78382a  and  a78367a );
 a337a <=( a78352a  and  a78337a );
 a338a <=( a78322a  and  a78307a );
 a339a <=( a78292a  and  a78277a );
 a340a <=( a78262a  and  a78247a );
 a341a <=( a78232a  and  a78217a );
 a342a <=( a78202a  and  a78187a );
 a343a <=( a78172a  and  a78157a );
 a344a <=( a78142a  and  a78127a );
 a345a <=( a78112a  and  a78097a );
 a346a <=( a78082a  and  a78067a );
 a347a <=( a78052a  and  a78037a );
 a348a <=( a78022a  and  a78007a );
 a349a <=( a77992a  and  a77977a );
 a350a <=( a77962a  and  a77947a );
 a351a <=( a77932a  and  a77917a );
 a352a <=( a77902a  and  a77887a );
 a353a <=( a77872a  and  a77857a );
 a354a <=( a77842a  and  a77827a );
 a355a <=( a77812a  and  a77797a );
 a356a <=( a77782a  and  a77767a );
 a357a <=( a77752a  and  a77737a );
 a358a <=( a77722a  and  a77707a );
 a359a <=( a77692a  and  a77677a );
 a360a <=( a77662a  and  a77647a );
 a361a <=( a77632a  and  a77617a );
 a362a <=( a77602a  and  a77587a );
 a363a <=( a77572a  and  a77557a );
 a364a <=( a77542a  and  a77527a );
 a365a <=( a77512a  and  a77497a );
 a366a <=( a77482a  and  a77467a );
 a367a <=( a77452a  and  a77437a );
 a368a <=( a77422a  and  a77407a );
 a369a <=( a77392a  and  a77377a );
 a370a <=( a77362a  and  a77347a );
 a371a <=( a77332a  and  a77317a );
 a372a <=( a77302a  and  a77287a );
 a373a <=( a77272a  and  a77257a );
 a374a <=( a77242a  and  a77227a );
 a375a <=( a77212a  and  a77197a );
 a376a <=( a77182a  and  a77167a );
 a377a <=( a77152a  and  a77137a );
 a378a <=( a77122a  and  a77107a );
 a379a <=( a77092a  and  a77077a );
 a380a <=( a77062a  and  a77047a );
 a381a <=( a77032a  and  a77017a );
 a382a <=( a77002a  and  a76987a );
 a383a <=( a76972a  and  a76957a );
 a384a <=( a76942a  and  a76927a );
 a385a <=( a76912a  and  a76897a );
 a386a <=( a76882a  and  a76867a );
 a387a <=( a76852a  and  a76837a );
 a388a <=( a76822a  and  a76807a );
 a389a <=( a76792a  and  a76777a );
 a390a <=( a76762a  and  a76747a );
 a391a <=( a76732a  and  a76717a );
 a392a <=( a76702a  and  a76687a );
 a393a <=( a76672a  and  a76657a );
 a394a <=( a76642a  and  a76627a );
 a395a <=( a76612a  and  a76597a );
 a396a <=( a76582a  and  a76567a );
 a397a <=( a76552a  and  a76537a );
 a398a <=( a76522a  and  a76507a );
 a399a <=( a76492a  and  a76477a );
 a400a <=( a76462a  and  a76447a );
 a401a <=( a76432a  and  a76417a );
 a402a <=( a76402a  and  a76387a );
 a403a <=( a76372a  and  a76357a );
 a404a <=( a76342a  and  a76327a );
 a405a <=( a76312a  and  a76297a );
 a406a <=( a76282a  and  a76267a );
 a407a <=( a76252a  and  a76237a );
 a408a <=( a76222a  and  a76207a );
 a409a <=( a76192a  and  a76177a );
 a410a <=( a76162a  and  a76147a );
 a411a <=( a76132a  and  a76117a );
 a412a <=( a76102a  and  a76087a );
 a413a <=( a76072a  and  a76057a );
 a414a <=( a76042a  and  a76027a );
 a415a <=( a76012a  and  a75997a );
 a416a <=( a75982a  and  a75967a );
 a417a <=( a75952a  and  a75937a );
 a418a <=( a75922a  and  a75907a );
 a419a <=( a75892a  and  a75877a );
 a420a <=( a75862a  and  a75847a );
 a421a <=( a75832a  and  a75817a );
 a422a <=( a75802a  and  a75787a );
 a423a <=( a75772a  and  a75757a );
 a424a <=( a75742a  and  a75727a );
 a425a <=( a75712a  and  a75697a );
 a426a <=( a75682a  and  a75667a );
 a427a <=( a75652a  and  a75637a );
 a428a <=( a75622a  and  a75607a );
 a429a <=( a75592a  and  a75577a );
 a430a <=( a75562a  and  a75547a );
 a431a <=( a75532a  and  a75517a );
 a432a <=( a75502a  and  a75487a );
 a433a <=( a75472a  and  a75457a );
 a434a <=( a75442a  and  a75427a );
 a435a <=( a75412a  and  a75397a );
 a436a <=( a75382a  and  a75367a );
 a437a <=( a75352a  and  a75337a );
 a438a <=( a75322a  and  a75307a );
 a439a <=( a75292a  and  a75277a );
 a440a <=( a75262a  and  a75247a );
 a441a <=( a75232a  and  a75217a );
 a442a <=( a75202a  and  a75187a );
 a443a <=( a75172a  and  a75157a );
 a444a <=( a75144a  and  a75129a );
 a445a <=( a75116a  and  a75101a );
 a446a <=( a75088a  and  a75073a );
 a447a <=( a75060a  and  a75045a );
 a448a <=( a75032a  and  a75017a );
 a449a <=( a75004a  and  a74989a );
 a450a <=( a74976a  and  a74961a );
 a451a <=( a74948a  and  a74933a );
 a452a <=( a74920a  and  a74905a );
 a453a <=( a74892a  and  a74877a );
 a454a <=( a74864a  and  a74849a );
 a455a <=( a74836a  and  a74821a );
 a456a <=( a74808a  and  a74793a );
 a457a <=( a74780a  and  a74765a );
 a458a <=( a74752a  and  a74737a );
 a459a <=( a74724a  and  a74709a );
 a460a <=( a74696a  and  a74681a );
 a461a <=( a74668a  and  a74653a );
 a462a <=( a74640a  and  a74625a );
 a463a <=( a74612a  and  a74597a );
 a464a <=( a74584a  and  a74569a );
 a465a <=( a74556a  and  a74541a );
 a466a <=( a74528a  and  a74513a );
 a467a <=( a74500a  and  a74485a );
 a468a <=( a74472a  and  a74457a );
 a469a <=( a74444a  and  a74429a );
 a470a <=( a74416a  and  a74401a );
 a471a <=( a74388a  and  a74373a );
 a472a <=( a74360a  and  a74345a );
 a473a <=( a74332a  and  a74317a );
 a474a <=( a74304a  and  a74289a );
 a475a <=( a74276a  and  a74261a );
 a476a <=( a74248a  and  a74233a );
 a477a <=( a74220a  and  a74205a );
 a478a <=( a74192a  and  a74177a );
 a479a <=( a74164a  and  a74149a );
 a480a <=( a74136a  and  a74121a );
 a481a <=( a74108a  and  a74093a );
 a482a <=( a74080a  and  a74065a );
 a483a <=( a74052a  and  a74037a );
 a484a <=( a74024a  and  a74009a );
 a485a <=( a73996a  and  a73981a );
 a486a <=( a73968a  and  a73953a );
 a487a <=( a73940a  and  a73925a );
 a488a <=( a73912a  and  a73897a );
 a489a <=( a73884a  and  a73869a );
 a490a <=( a73856a  and  a73841a );
 a491a <=( a73828a  and  a73813a );
 a492a <=( a73800a  and  a73785a );
 a493a <=( a73772a  and  a73757a );
 a494a <=( a73744a  and  a73729a );
 a495a <=( a73716a  and  a73701a );
 a496a <=( a73688a  and  a73673a );
 a497a <=( a73660a  and  a73645a );
 a498a <=( a73632a  and  a73617a );
 a499a <=( a73604a  and  a73589a );
 a500a <=( a73576a  and  a73561a );
 a501a <=( a73548a  and  a73533a );
 a502a <=( a73520a  and  a73505a );
 a503a <=( a73492a  and  a73477a );
 a504a <=( a73464a  and  a73449a );
 a505a <=( a73436a  and  a73421a );
 a506a <=( a73408a  and  a73393a );
 a507a <=( a73380a  and  a73365a );
 a508a <=( a73352a  and  a73337a );
 a509a <=( a73324a  and  a73309a );
 a510a <=( a73296a  and  a73281a );
 a511a <=( a73268a  and  a73253a );
 a512a <=( a73240a  and  a73225a );
 a513a <=( a73212a  and  a73197a );
 a514a <=( a73184a  and  a73169a );
 a515a <=( a73156a  and  a73141a );
 a516a <=( a73128a  and  a73113a );
 a517a <=( a73100a  and  a73085a );
 a518a <=( a73072a  and  a73057a );
 a519a <=( a73044a  and  a73029a );
 a520a <=( a73016a  and  a73001a );
 a521a <=( a72988a  and  a72973a );
 a522a <=( a72960a  and  a72945a );
 a523a <=( a72932a  and  a72917a );
 a524a <=( a72904a  and  a72889a );
 a525a <=( a72876a  and  a72861a );
 a526a <=( a72848a  and  a72833a );
 a527a <=( a72820a  and  a72805a );
 a528a <=( a72792a  and  a72777a );
 a529a <=( a72764a  and  a72749a );
 a530a <=( a72736a  and  a72721a );
 a531a <=( a72708a  and  a72693a );
 a532a <=( a72680a  and  a72665a );
 a533a <=( a72652a  and  a72637a );
 a534a <=( a72624a  and  a72609a );
 a535a <=( a72596a  and  a72581a );
 a536a <=( a72568a  and  a72553a );
 a537a <=( a72540a  and  a72525a );
 a538a <=( a72512a  and  a72497a );
 a539a <=( a72484a  and  a72469a );
 a540a <=( a72456a  and  a72441a );
 a541a <=( a72428a  and  a72413a );
 a542a <=( a72400a  and  a72385a );
 a543a <=( a72372a  and  a72357a );
 a544a <=( a72344a  and  a72329a );
 a545a <=( a72316a  and  a72301a );
 a546a <=( a72288a  and  a72273a );
 a547a <=( a72260a  and  a72245a );
 a548a <=( a72232a  and  a72217a );
 a549a <=( a72204a  and  a72189a );
 a550a <=( a72176a  and  a72161a );
 a551a <=( a72148a  and  a72133a );
 a552a <=( a72120a  and  a72105a );
 a553a <=( a72092a  and  a72077a );
 a554a <=( a72064a  and  a72049a );
 a555a <=( a72036a  and  a72021a );
 a556a <=( a72008a  and  a71993a );
 a557a <=( a71980a  and  a71965a );
 a558a <=( a71952a  and  a71937a );
 a559a <=( a71924a  and  a71909a );
 a560a <=( a71896a  and  a71881a );
 a561a <=( a71868a  and  a71853a );
 a562a <=( a71840a  and  a71825a );
 a563a <=( a71812a  and  a71797a );
 a564a <=( a71784a  and  a71769a );
 a565a <=( a71756a  and  a71741a );
 a566a <=( a71728a  and  a71713a );
 a567a <=( a71700a  and  a71685a );
 a568a <=( a71672a  and  a71657a );
 a569a <=( a71644a  and  a71629a );
 a570a <=( a71616a  and  a71601a );
 a571a <=( a71588a  and  a71573a );
 a572a <=( a71560a  and  a71545a );
 a573a <=( a71532a  and  a71517a );
 a574a <=( a71504a  and  a71489a );
 a575a <=( a71476a  and  a71461a );
 a576a <=( a71448a  and  a71433a );
 a577a <=( a71420a  and  a71405a );
 a578a <=( a71392a  and  a71377a );
 a579a <=( a71364a  and  a71349a );
 a580a <=( a71336a  and  a71321a );
 a581a <=( a71308a  and  a71293a );
 a582a <=( a71280a  and  a71265a );
 a583a <=( a71252a  and  a71237a );
 a584a <=( a71224a  and  a71209a );
 a585a <=( a71196a  and  a71181a );
 a586a <=( a71168a  and  a71153a );
 a587a <=( a71140a  and  a71125a );
 a588a <=( a71112a  and  a71097a );
 a589a <=( a71084a  and  a71069a );
 a590a <=( a71056a  and  a71041a );
 a591a <=( a71028a  and  a71013a );
 a592a <=( a71000a  and  a70985a );
 a593a <=( a70972a  and  a70957a );
 a594a <=( a70944a  and  a70929a );
 a595a <=( a70916a  and  a70901a );
 a596a <=( a70888a  and  a70873a );
 a597a <=( a70860a  and  a70845a );
 a598a <=( a70832a  and  a70817a );
 a599a <=( a70804a  and  a70789a );
 a600a <=( a70776a  and  a70761a );
 a601a <=( a70748a  and  a70733a );
 a602a <=( a70720a  and  a70705a );
 a603a <=( a70692a  and  a70677a );
 a604a <=( a70664a  and  a70649a );
 a605a <=( a70636a  and  a70621a );
 a606a <=( a70608a  and  a70593a );
 a607a <=( a70580a  and  a70565a );
 a608a <=( a70552a  and  a70537a );
 a609a <=( a70524a  and  a70509a );
 a610a <=( a70496a  and  a70481a );
 a611a <=( a70468a  and  a70453a );
 a612a <=( a70440a  and  a70425a );
 a613a <=( a70412a  and  a70397a );
 a614a <=( a70384a  and  a70369a );
 a615a <=( a70356a  and  a70341a );
 a616a <=( a70328a  and  a70313a );
 a617a <=( a70300a  and  a70285a );
 a618a <=( a70272a  and  a70257a );
 a619a <=( a70244a  and  a70229a );
 a620a <=( a70216a  and  a70201a );
 a621a <=( a70188a  and  a70173a );
 a622a <=( a70160a  and  a70145a );
 a623a <=( a70132a  and  a70117a );
 a624a <=( a70104a  and  a70089a );
 a625a <=( a70076a  and  a70061a );
 a626a <=( a70048a  and  a70033a );
 a627a <=( a70020a  and  a70005a );
 a628a <=( a69992a  and  a69977a );
 a629a <=( a69964a  and  a69949a );
 a630a <=( a69936a  and  a69921a );
 a631a <=( a69908a  and  a69893a );
 a632a <=( a69880a  and  a69865a );
 a633a <=( a69852a  and  a69837a );
 a634a <=( a69824a  and  a69809a );
 a635a <=( a69796a  and  a69781a );
 a636a <=( a69768a  and  a69753a );
 a637a <=( a69740a  and  a69725a );
 a638a <=( a69712a  and  a69697a );
 a639a <=( a69684a  and  a69669a );
 a640a <=( a69656a  and  a69641a );
 a641a <=( a69628a  and  a69613a );
 a642a <=( a69600a  and  a69585a );
 a643a <=( a69572a  and  a69557a );
 a644a <=( a69544a  and  a69529a );
 a645a <=( a69516a  and  a69501a );
 a646a <=( a69488a  and  a69473a );
 a647a <=( a69460a  and  a69445a );
 a648a <=( a69432a  and  a69417a );
 a649a <=( a69404a  and  a69389a );
 a650a <=( a69376a  and  a69361a );
 a651a <=( a69348a  and  a69333a );
 a652a <=( a69320a  and  a69305a );
 a653a <=( a69292a  and  a69277a );
 a654a <=( a69264a  and  a69249a );
 a655a <=( a69236a  and  a69221a );
 a656a <=( a69208a  and  a69193a );
 a657a <=( a69180a  and  a69165a );
 a658a <=( a69152a  and  a69137a );
 a659a <=( a69124a  and  a69109a );
 a660a <=( a69096a  and  a69081a );
 a661a <=( a69068a  and  a69053a );
 a662a <=( a69040a  and  a69025a );
 a663a <=( a69012a  and  a68997a );
 a664a <=( a68984a  and  a68969a );
 a665a <=( a68956a  and  a68941a );
 a666a <=( a68928a  and  a68913a );
 a667a <=( a68900a  and  a68885a );
 a668a <=( a68872a  and  a68857a );
 a669a <=( a68844a  and  a68829a );
 a670a <=( a68816a  and  a68801a );
 a671a <=( a68788a  and  a68773a );
 a672a <=( a68760a  and  a68745a );
 a673a <=( a68732a  and  a68717a );
 a674a <=( a68704a  and  a68689a );
 a675a <=( a68676a  and  a68661a );
 a676a <=( a68648a  and  a68633a );
 a677a <=( a68620a  and  a68605a );
 a678a <=( a68592a  and  a68577a );
 a679a <=( a68564a  and  a68549a );
 a680a <=( a68536a  and  a68521a );
 a681a <=( a68508a  and  a68493a );
 a682a <=( a68480a  and  a68465a );
 a683a <=( a68452a  and  a68437a );
 a684a <=( a68424a  and  a68409a );
 a685a <=( a68396a  and  a68381a );
 a686a <=( a68368a  and  a68353a );
 a687a <=( a68340a  and  a68325a );
 a688a <=( a68312a  and  a68297a );
 a689a <=( a68284a  and  a68269a );
 a690a <=( a68256a  and  a68241a );
 a691a <=( a68228a  and  a68213a );
 a692a <=( a68200a  and  a68185a );
 a693a <=( a68172a  and  a68157a );
 a694a <=( a68144a  and  a68129a );
 a695a <=( a68116a  and  a68101a );
 a696a <=( a68088a  and  a68073a );
 a697a <=( a68060a  and  a68045a );
 a698a <=( a68032a  and  a68017a );
 a699a <=( a68004a  and  a67989a );
 a700a <=( a67976a  and  a67961a );
 a701a <=( a67948a  and  a67933a );
 a702a <=( a67920a  and  a67905a );
 a703a <=( a67892a  and  a67877a );
 a704a <=( a67864a  and  a67849a );
 a705a <=( a67836a  and  a67821a );
 a706a <=( a67808a  and  a67793a );
 a707a <=( a67780a  and  a67765a );
 a708a <=( a67752a  and  a67737a );
 a709a <=( a67724a  and  a67709a );
 a710a <=( a67696a  and  a67681a );
 a711a <=( a67668a  and  a67653a );
 a712a <=( a67640a  and  a67625a );
 a713a <=( a67612a  and  a67597a );
 a714a <=( a67584a  and  a67569a );
 a715a <=( a67556a  and  a67541a );
 a716a <=( a67528a  and  a67513a );
 a717a <=( a67500a  and  a67485a );
 a718a <=( a67472a  and  a67457a );
 a719a <=( a67444a  and  a67429a );
 a720a <=( a67416a  and  a67401a );
 a721a <=( a67388a  and  a67373a );
 a722a <=( a67360a  and  a67345a );
 a723a <=( a67332a  and  a67317a );
 a724a <=( a67304a  and  a67289a );
 a725a <=( a67276a  and  a67261a );
 a726a <=( a67248a  and  a67233a );
 a727a <=( a67220a  and  a67205a );
 a728a <=( a67192a  and  a67177a );
 a729a <=( a67164a  and  a67149a );
 a730a <=( a67136a  and  a67121a );
 a731a <=( a67108a  and  a67093a );
 a732a <=( a67080a  and  a67065a );
 a733a <=( a67052a  and  a67037a );
 a734a <=( a67024a  and  a67009a );
 a735a <=( a66996a  and  a66981a );
 a736a <=( a66968a  and  a66953a );
 a737a <=( a66940a  and  a66925a );
 a738a <=( a66912a  and  a66897a );
 a739a <=( a66884a  and  a66869a );
 a740a <=( a66856a  and  a66841a );
 a741a <=( a66828a  and  a66813a );
 a742a <=( a66800a  and  a66785a );
 a743a <=( a66772a  and  a66757a );
 a744a <=( a66744a  and  a66729a );
 a745a <=( a66716a  and  a66701a );
 a746a <=( a66688a  and  a66673a );
 a747a <=( a66660a  and  a66645a );
 a748a <=( a66632a  and  a66617a );
 a749a <=( a66604a  and  a66589a );
 a750a <=( a66576a  and  a66561a );
 a751a <=( a66548a  and  a66533a );
 a752a <=( a66520a  and  a66505a );
 a753a <=( a66492a  and  a66477a );
 a754a <=( a66464a  and  a66449a );
 a755a <=( a66436a  and  a66421a );
 a756a <=( a66408a  and  a66393a );
 a757a <=( a66380a  and  a66365a );
 a758a <=( a66352a  and  a66337a );
 a759a <=( a66324a  and  a66309a );
 a760a <=( a66296a  and  a66281a );
 a761a <=( a66268a  and  a66253a );
 a762a <=( a66240a  and  a66225a );
 a763a <=( a66212a  and  a66197a );
 a764a <=( a66184a  and  a66169a );
 a765a <=( a66156a  and  a66141a );
 a766a <=( a66128a  and  a66113a );
 a767a <=( a66100a  and  a66085a );
 a768a <=( a66072a  and  a66057a );
 a769a <=( a66044a  and  a66029a );
 a770a <=( a66016a  and  a66001a );
 a771a <=( a65988a  and  a65973a );
 a772a <=( a65960a  and  a65945a );
 a773a <=( a65932a  and  a65917a );
 a774a <=( a65904a  and  a65889a );
 a775a <=( a65876a  and  a65861a );
 a776a <=( a65848a  and  a65833a );
 a777a <=( a65820a  and  a65805a );
 a778a <=( a65792a  and  a65777a );
 a779a <=( a65764a  and  a65749a );
 a780a <=( a65736a  and  a65721a );
 a781a <=( a65708a  and  a65693a );
 a782a <=( a65680a  and  a65665a );
 a783a <=( a65652a  and  a65637a );
 a784a <=( a65624a  and  a65609a );
 a785a <=( a65596a  and  a65581a );
 a786a <=( a65568a  and  a65553a );
 a787a <=( a65540a  and  a65525a );
 a788a <=( a65512a  and  a65497a );
 a789a <=( a65484a  and  a65469a );
 a790a <=( a65456a  and  a65441a );
 a791a <=( a65428a  and  a65413a );
 a792a <=( a65400a  and  a65385a );
 a793a <=( a65372a  and  a65357a );
 a794a <=( a65344a  and  a65329a );
 a795a <=( a65316a  and  a65301a );
 a796a <=( a65288a  and  a65273a );
 a797a <=( a65260a  and  a65245a );
 a798a <=( a65232a  and  a65217a );
 a799a <=( a65204a  and  a65189a );
 a800a <=( a65176a  and  a65161a );
 a801a <=( a65148a  and  a65133a );
 a802a <=( a65120a  and  a65105a );
 a803a <=( a65092a  and  a65077a );
 a804a <=( a65064a  and  a65049a );
 a805a <=( a65036a  and  a65021a );
 a806a <=( a65008a  and  a64993a );
 a807a <=( a64980a  and  a64965a );
 a808a <=( a64952a  and  a64937a );
 a809a <=( a64924a  and  a64909a );
 a810a <=( a64896a  and  a64881a );
 a811a <=( a64868a  and  a64853a );
 a812a <=( a64840a  and  a64825a );
 a813a <=( a64812a  and  a64797a );
 a814a <=( a64784a  and  a64769a );
 a815a <=( a64756a  and  a64741a );
 a816a <=( a64728a  and  a64713a );
 a817a <=( a64700a  and  a64685a );
 a818a <=( a64672a  and  a64657a );
 a819a <=( a64644a  and  a64629a );
 a820a <=( a64616a  and  a64601a );
 a821a <=( a64588a  and  a64573a );
 a822a <=( a64560a  and  a64545a );
 a823a <=( a64532a  and  a64517a );
 a824a <=( a64504a  and  a64489a );
 a825a <=( a64476a  and  a64461a );
 a826a <=( a64448a  and  a64433a );
 a827a <=( a64420a  and  a64405a );
 a828a <=( a64392a  and  a64377a );
 a829a <=( a64364a  and  a64349a );
 a830a <=( a64336a  and  a64321a );
 a831a <=( a64308a  and  a64293a );
 a832a <=( a64280a  and  a64265a );
 a833a <=( a64252a  and  a64237a );
 a834a <=( a64224a  and  a64209a );
 a835a <=( a64196a  and  a64181a );
 a836a <=( a64168a  and  a64153a );
 a837a <=( a64140a  and  a64125a );
 a838a <=( a64112a  and  a64097a );
 a839a <=( a64084a  and  a64069a );
 a840a <=( a64056a  and  a64041a );
 a841a <=( a64028a  and  a64013a );
 a842a <=( a64000a  and  a63985a );
 a843a <=( a63972a  and  a63957a );
 a844a <=( a63944a  and  a63929a );
 a845a <=( a63916a  and  a63901a );
 a846a <=( a63888a  and  a63873a );
 a847a <=( a63860a  and  a63845a );
 a848a <=( a63832a  and  a63817a );
 a849a <=( a63804a  and  a63789a );
 a850a <=( a63776a  and  a63761a );
 a851a <=( a63748a  and  a63733a );
 a852a <=( a63720a  and  a63705a );
 a853a <=( a63692a  and  a63677a );
 a854a <=( a63664a  and  a63649a );
 a855a <=( a63636a  and  a63621a );
 a856a <=( a63608a  and  a63593a );
 a857a <=( a63580a  and  a63565a );
 a858a <=( a63552a  and  a63537a );
 a859a <=( a63524a  and  a63509a );
 a860a <=( a63496a  and  a63481a );
 a861a <=( a63468a  and  a63453a );
 a862a <=( a63440a  and  a63425a );
 a863a <=( a63412a  and  a63397a );
 a864a <=( a63384a  and  a63369a );
 a865a <=( a63356a  and  a63341a );
 a866a <=( a63328a  and  a63313a );
 a867a <=( a63300a  and  a63285a );
 a868a <=( a63272a  and  a63257a );
 a869a <=( a63244a  and  a63229a );
 a870a <=( a63216a  and  a63201a );
 a871a <=( a63188a  and  a63173a );
 a872a <=( a63160a  and  a63145a );
 a873a <=( a63132a  and  a63117a );
 a874a <=( a63104a  and  a63089a );
 a875a <=( a63076a  and  a63061a );
 a876a <=( a63048a  and  a63033a );
 a877a <=( a63020a  and  a63005a );
 a878a <=( a62992a  and  a62977a );
 a879a <=( a62964a  and  a62949a );
 a880a <=( a62936a  and  a62921a );
 a881a <=( a62908a  and  a62893a );
 a882a <=( a62880a  and  a62865a );
 a883a <=( a62852a  and  a62837a );
 a884a <=( a62824a  and  a62809a );
 a885a <=( a62796a  and  a62781a );
 a886a <=( a62768a  and  a62753a );
 a887a <=( a62740a  and  a62725a );
 a888a <=( a62712a  and  a62697a );
 a889a <=( a62684a  and  a62669a );
 a890a <=( a62656a  and  a62641a );
 a891a <=( a62628a  and  a62613a );
 a892a <=( a62600a  and  a62585a );
 a893a <=( a62572a  and  a62557a );
 a894a <=( a62544a  and  a62529a );
 a895a <=( a62516a  and  a62501a );
 a896a <=( a62488a  and  a62473a );
 a897a <=( a62460a  and  a62445a );
 a898a <=( a62432a  and  a62417a );
 a899a <=( a62404a  and  a62389a );
 a900a <=( a62376a  and  a62361a );
 a901a <=( a62348a  and  a62333a );
 a902a <=( a62320a  and  a62305a );
 a903a <=( a62292a  and  a62277a );
 a904a <=( a62264a  and  a62249a );
 a905a <=( a62236a  and  a62221a );
 a906a <=( a62208a  and  a62193a );
 a907a <=( a62180a  and  a62165a );
 a908a <=( a62152a  and  a62137a );
 a909a <=( a62124a  and  a62109a );
 a910a <=( a62096a  and  a62081a );
 a911a <=( a62068a  and  a62053a );
 a912a <=( a62040a  and  a62025a );
 a913a <=( a62012a  and  a61997a );
 a914a <=( a61984a  and  a61969a );
 a915a <=( a61956a  and  a61941a );
 a916a <=( a61928a  and  a61913a );
 a917a <=( a61900a  and  a61885a );
 a918a <=( a61872a  and  a61857a );
 a919a <=( a61844a  and  a61829a );
 a920a <=( a61816a  and  a61801a );
 a921a <=( a61788a  and  a61773a );
 a922a <=( a61760a  and  a61745a );
 a923a <=( a61732a  and  a61717a );
 a924a <=( a61704a  and  a61689a );
 a925a <=( a61676a  and  a61661a );
 a926a <=( a61648a  and  a61633a );
 a927a <=( a61620a  and  a61605a );
 a928a <=( a61592a  and  a61577a );
 a929a <=( a61564a  and  a61549a );
 a930a <=( a61536a  and  a61521a );
 a931a <=( a61508a  and  a61493a );
 a932a <=( a61480a  and  a61465a );
 a933a <=( a61452a  and  a61437a );
 a934a <=( a61424a  and  a61409a );
 a935a <=( a61396a  and  a61381a );
 a936a <=( a61368a  and  a61353a );
 a937a <=( a61340a  and  a61325a );
 a938a <=( a61312a  and  a61297a );
 a939a <=( a61284a  and  a61269a );
 a940a <=( a61256a  and  a61241a );
 a941a <=( a61228a  and  a61213a );
 a942a <=( a61200a  and  a61185a );
 a943a <=( a61172a  and  a61157a );
 a944a <=( a61144a  and  a61129a );
 a945a <=( a61116a  and  a61101a );
 a946a <=( a61088a  and  a61073a );
 a947a <=( a61060a  and  a61045a );
 a948a <=( a61032a  and  a61017a );
 a949a <=( a61004a  and  a60989a );
 a950a <=( a60976a  and  a60961a );
 a951a <=( a60948a  and  a60933a );
 a952a <=( a60920a  and  a60905a );
 a953a <=( a60892a  and  a60877a );
 a954a <=( a60864a  and  a60849a );
 a955a <=( a60836a  and  a60821a );
 a956a <=( a60808a  and  a60793a );
 a957a <=( a60780a  and  a60765a );
 a958a <=( a60752a  and  a60737a );
 a959a <=( a60724a  and  a60709a );
 a960a <=( a60696a  and  a60681a );
 a961a <=( a60668a  and  a60653a );
 a962a <=( a60640a  and  a60625a );
 a963a <=( a60612a  and  a60597a );
 a964a <=( a60584a  and  a60569a );
 a965a <=( a60556a  and  a60541a );
 a966a <=( a60528a  and  a60513a );
 a967a <=( a60500a  and  a60485a );
 a968a <=( a60472a  and  a60457a );
 a969a <=( a60444a  and  a60429a );
 a970a <=( a60416a  and  a60401a );
 a971a <=( a60388a  and  a60373a );
 a972a <=( a60360a  and  a60345a );
 a973a <=( a60332a  and  a60317a );
 a974a <=( a60304a  and  a60289a );
 a975a <=( a60276a  and  a60263a );
 a976a <=( a60250a  and  a60237a );
 a977a <=( a60224a  and  a60211a );
 a978a <=( a60198a  and  a60185a );
 a979a <=( a60172a  and  a60159a );
 a980a <=( a60146a  and  a60133a );
 a981a <=( a60120a  and  a60107a );
 a982a <=( a60094a  and  a60081a );
 a983a <=( a60068a  and  a60055a );
 a984a <=( a60042a  and  a60029a );
 a985a <=( a60016a  and  a60003a );
 a986a <=( a59990a  and  a59977a );
 a987a <=( a59964a  and  a59951a );
 a988a <=( a59938a  and  a59925a );
 a989a <=( a59912a  and  a59899a );
 a990a <=( a59886a  and  a59873a );
 a991a <=( a59860a  and  a59847a );
 a992a <=( a59834a  and  a59821a );
 a993a <=( a59808a  and  a59795a );
 a994a <=( a59782a  and  a59769a );
 a995a <=( a59756a  and  a59743a );
 a996a <=( a59730a  and  a59717a );
 a997a <=( a59704a  and  a59691a );
 a998a <=( a59678a  and  a59665a );
 a999a <=( a59652a  and  a59639a );
 a1000a <=( a59626a  and  a59613a );
 a1001a <=( a59600a  and  a59587a );
 a1002a <=( a59574a  and  a59561a );
 a1003a <=( a59548a  and  a59535a );
 a1004a <=( a59522a  and  a59509a );
 a1005a <=( a59496a  and  a59483a );
 a1006a <=( a59470a  and  a59457a );
 a1007a <=( a59444a  and  a59431a );
 a1008a <=( a59418a  and  a59405a );
 a1009a <=( a59392a  and  a59379a );
 a1010a <=( a59366a  and  a59353a );
 a1011a <=( a59340a  and  a59327a );
 a1012a <=( a59314a  and  a59301a );
 a1013a <=( a59288a  and  a59275a );
 a1014a <=( a59262a  and  a59249a );
 a1015a <=( a59236a  and  a59223a );
 a1016a <=( a59210a  and  a59197a );
 a1017a <=( a59184a  and  a59171a );
 a1018a <=( a59158a  and  a59145a );
 a1019a <=( a59132a  and  a59119a );
 a1020a <=( a59106a  and  a59093a );
 a1021a <=( a59080a  and  a59067a );
 a1022a <=( a59054a  and  a59041a );
 a1023a <=( a59028a  and  a59015a );
 a1024a <=( a59002a  and  a58989a );
 a1025a <=( a58976a  and  a58963a );
 a1026a <=( a58950a  and  a58937a );
 a1027a <=( a58924a  and  a58911a );
 a1028a <=( a58898a  and  a58885a );
 a1029a <=( a58872a  and  a58859a );
 a1030a <=( a58846a  and  a58833a );
 a1031a <=( a58820a  and  a58807a );
 a1032a <=( a58794a  and  a58781a );
 a1033a <=( a58768a  and  a58755a );
 a1034a <=( a58742a  and  a58729a );
 a1035a <=( a58716a  and  a58703a );
 a1036a <=( a58690a  and  a58677a );
 a1037a <=( a58664a  and  a58651a );
 a1038a <=( a58638a  and  a58625a );
 a1039a <=( a58612a  and  a58599a );
 a1040a <=( a58586a  and  a58573a );
 a1041a <=( a58560a  and  a58547a );
 a1042a <=( a58534a  and  a58521a );
 a1043a <=( a58508a  and  a58495a );
 a1044a <=( a58482a  and  a58469a );
 a1045a <=( a58456a  and  a58443a );
 a1046a <=( a58430a  and  a58417a );
 a1047a <=( a58404a  and  a58391a );
 a1048a <=( a58378a  and  a58365a );
 a1049a <=( a58352a  and  a58339a );
 a1050a <=( a58326a  and  a58313a );
 a1051a <=( a58300a  and  a58287a );
 a1052a <=( a58274a  and  a58261a );
 a1053a <=( a58248a  and  a58235a );
 a1054a <=( a58222a  and  a58209a );
 a1055a <=( a58196a  and  a58183a );
 a1056a <=( a58170a  and  a58157a );
 a1057a <=( a58144a  and  a58131a );
 a1058a <=( a58118a  and  a58105a );
 a1059a <=( a58092a  and  a58079a );
 a1060a <=( a58066a  and  a58053a );
 a1061a <=( a58040a  and  a58027a );
 a1062a <=( a58014a  and  a58001a );
 a1063a <=( a57988a  and  a57975a );
 a1064a <=( a57962a  and  a57949a );
 a1065a <=( a57936a  and  a57923a );
 a1066a <=( a57910a  and  a57897a );
 a1067a <=( a57884a  and  a57871a );
 a1068a <=( a57858a  and  a57845a );
 a1069a <=( a57832a  and  a57819a );
 a1070a <=( a57806a  and  a57793a );
 a1071a <=( a57780a  and  a57767a );
 a1072a <=( a57754a  and  a57741a );
 a1073a <=( a57728a  and  a57715a );
 a1074a <=( a57702a  and  a57689a );
 a1075a <=( a57676a  and  a57663a );
 a1076a <=( a57650a  and  a57637a );
 a1077a <=( a57624a  and  a57611a );
 a1078a <=( a57598a  and  a57585a );
 a1079a <=( a57572a  and  a57559a );
 a1080a <=( a57546a  and  a57533a );
 a1081a <=( a57520a  and  a57507a );
 a1082a <=( a57494a  and  a57481a );
 a1083a <=( a57468a  and  a57455a );
 a1084a <=( a57442a  and  a57429a );
 a1085a <=( a57416a  and  a57403a );
 a1086a <=( a57390a  and  a57377a );
 a1087a <=( a57364a  and  a57351a );
 a1088a <=( a57338a  and  a57325a );
 a1089a <=( a57312a  and  a57299a );
 a1090a <=( a57286a  and  a57273a );
 a1091a <=( a57260a  and  a57247a );
 a1092a <=( a57234a  and  a57221a );
 a1093a <=( a57208a  and  a57195a );
 a1094a <=( a57182a  and  a57169a );
 a1095a <=( a57156a  and  a57143a );
 a1096a <=( a57130a  and  a57117a );
 a1097a <=( a57104a  and  a57091a );
 a1098a <=( a57078a  and  a57065a );
 a1099a <=( a57052a  and  a57039a );
 a1100a <=( a57026a  and  a57013a );
 a1101a <=( a57000a  and  a56987a );
 a1102a <=( a56974a  and  a56961a );
 a1103a <=( a56948a  and  a56935a );
 a1104a <=( a56922a  and  a56909a );
 a1105a <=( a56896a  and  a56883a );
 a1106a <=( a56870a  and  a56857a );
 a1107a <=( a56844a  and  a56831a );
 a1108a <=( a56818a  and  a56805a );
 a1109a <=( a56792a  and  a56779a );
 a1110a <=( a56766a  and  a56753a );
 a1111a <=( a56740a  and  a56727a );
 a1112a <=( a56714a  and  a56701a );
 a1113a <=( a56688a  and  a56675a );
 a1114a <=( a56662a  and  a56649a );
 a1115a <=( a56636a  and  a56623a );
 a1116a <=( a56610a  and  a56597a );
 a1117a <=( a56584a  and  a56571a );
 a1118a <=( a56558a  and  a56545a );
 a1119a <=( a56532a  and  a56519a );
 a1120a <=( a56506a  and  a56493a );
 a1121a <=( a56480a  and  a56467a );
 a1122a <=( a56454a  and  a56441a );
 a1123a <=( a56428a  and  a56415a );
 a1124a <=( a56402a  and  a56389a );
 a1125a <=( a56376a  and  a56363a );
 a1126a <=( a56350a  and  a56337a );
 a1127a <=( a56324a  and  a56311a );
 a1128a <=( a56298a  and  a56285a );
 a1129a <=( a56272a  and  a56259a );
 a1130a <=( a56246a  and  a56233a );
 a1131a <=( a56220a  and  a56207a );
 a1132a <=( a56194a  and  a56181a );
 a1133a <=( a56168a  and  a56155a );
 a1134a <=( a56142a  and  a56129a );
 a1135a <=( a56116a  and  a56103a );
 a1136a <=( a56090a  and  a56077a );
 a1137a <=( a56064a  and  a56051a );
 a1138a <=( a56038a  and  a56025a );
 a1139a <=( a56012a  and  a55999a );
 a1140a <=( a55986a  and  a55973a );
 a1141a <=( a55960a  and  a55947a );
 a1142a <=( a55934a  and  a55921a );
 a1143a <=( a55908a  and  a55895a );
 a1144a <=( a55882a  and  a55869a );
 a1145a <=( a55856a  and  a55843a );
 a1146a <=( a55830a  and  a55817a );
 a1147a <=( a55804a  and  a55791a );
 a1148a <=( a55778a  and  a55765a );
 a1149a <=( a55752a  and  a55739a );
 a1150a <=( a55726a  and  a55713a );
 a1151a <=( a55700a  and  a55687a );
 a1152a <=( a55674a  and  a55661a );
 a1153a <=( a55648a  and  a55635a );
 a1154a <=( a55622a  and  a55609a );
 a1155a <=( a55596a  and  a55583a );
 a1156a <=( a55570a  and  a55557a );
 a1157a <=( a55544a  and  a55531a );
 a1158a <=( a55518a  and  a55505a );
 a1159a <=( a55492a  and  a55479a );
 a1160a <=( a55466a  and  a55453a );
 a1161a <=( a55440a  and  a55427a );
 a1162a <=( a55414a  and  a55401a );
 a1163a <=( a55388a  and  a55375a );
 a1164a <=( a55362a  and  a55349a );
 a1165a <=( a55336a  and  a55323a );
 a1166a <=( a55310a  and  a55297a );
 a1167a <=( a55284a  and  a55271a );
 a1168a <=( a55258a  and  a55245a );
 a1169a <=( a55232a  and  a55219a );
 a1170a <=( a55206a  and  a55193a );
 a1171a <=( a55180a  and  a55167a );
 a1172a <=( a55154a  and  a55141a );
 a1173a <=( a55128a  and  a55115a );
 a1174a <=( a55102a  and  a55089a );
 a1175a <=( a55076a  and  a55063a );
 a1176a <=( a55050a  and  a55037a );
 a1177a <=( a55024a  and  a55011a );
 a1178a <=( a54998a  and  a54985a );
 a1179a <=( a54972a  and  a54959a );
 a1180a <=( a54946a  and  a54933a );
 a1181a <=( a54920a  and  a54907a );
 a1182a <=( a54894a  and  a54881a );
 a1183a <=( a54868a  and  a54855a );
 a1184a <=( a54842a  and  a54829a );
 a1185a <=( a54816a  and  a54803a );
 a1186a <=( a54790a  and  a54777a );
 a1187a <=( a54764a  and  a54751a );
 a1188a <=( a54738a  and  a54725a );
 a1189a <=( a54712a  and  a54699a );
 a1190a <=( a54686a  and  a54673a );
 a1191a <=( a54660a  and  a54647a );
 a1192a <=( a54634a  and  a54621a );
 a1193a <=( a54608a  and  a54595a );
 a1194a <=( a54582a  and  a54569a );
 a1195a <=( a54556a  and  a54543a );
 a1196a <=( a54530a  and  a54517a );
 a1197a <=( a54504a  and  a54491a );
 a1198a <=( a54478a  and  a54465a );
 a1199a <=( a54452a  and  a54439a );
 a1200a <=( a54426a  and  a54413a );
 a1201a <=( a54400a  and  a54387a );
 a1202a <=( a54374a  and  a54361a );
 a1203a <=( a54348a  and  a54335a );
 a1204a <=( a54322a  and  a54309a );
 a1205a <=( a54296a  and  a54283a );
 a1206a <=( a54270a  and  a54257a );
 a1207a <=( a54244a  and  a54231a );
 a1208a <=( a54218a  and  a54205a );
 a1209a <=( a54192a  and  a54179a );
 a1210a <=( a54166a  and  a54153a );
 a1211a <=( a54140a  and  a54127a );
 a1212a <=( a54114a  and  a54101a );
 a1213a <=( a54088a  and  a54075a );
 a1214a <=( a54062a  and  a54049a );
 a1215a <=( a54036a  and  a54023a );
 a1216a <=( a54010a  and  a53997a );
 a1217a <=( a53984a  and  a53971a );
 a1218a <=( a53958a  and  a53945a );
 a1219a <=( a53932a  and  a53919a );
 a1220a <=( a53906a  and  a53893a );
 a1221a <=( a53880a  and  a53867a );
 a1222a <=( a53854a  and  a53841a );
 a1223a <=( a53828a  and  a53815a );
 a1224a <=( a53802a  and  a53789a );
 a1225a <=( a53776a  and  a53763a );
 a1226a <=( a53750a  and  a53737a );
 a1227a <=( a53724a  and  a53711a );
 a1228a <=( a53698a  and  a53685a );
 a1229a <=( a53672a  and  a53659a );
 a1230a <=( a53646a  and  a53633a );
 a1231a <=( a53620a  and  a53607a );
 a1232a <=( a53594a  and  a53581a );
 a1233a <=( a53568a  and  a53555a );
 a1234a <=( a53542a  and  a53529a );
 a1235a <=( a53516a  and  a53503a );
 a1236a <=( a53490a  and  a53477a );
 a1237a <=( a53464a  and  a53451a );
 a1238a <=( a53438a  and  a53425a );
 a1239a <=( a53412a  and  a53399a );
 a1240a <=( a53386a  and  a53373a );
 a1241a <=( a53360a  and  a53347a );
 a1242a <=( a53334a  and  a53321a );
 a1243a <=( a53308a  and  a53295a );
 a1244a <=( a53282a  and  a53269a );
 a1245a <=( a53256a  and  a53243a );
 a1246a <=( a53230a  and  a53217a );
 a1247a <=( a53204a  and  a53191a );
 a1248a <=( a53178a  and  a53165a );
 a1249a <=( a53152a  and  a53139a );
 a1250a <=( a53126a  and  a53113a );
 a1251a <=( a53100a  and  a53087a );
 a1252a <=( a53074a  and  a53061a );
 a1253a <=( a53048a  and  a53035a );
 a1254a <=( a53022a  and  a53009a );
 a1255a <=( a52996a  and  a52983a );
 a1256a <=( a52970a  and  a52957a );
 a1257a <=( a52944a  and  a52931a );
 a1258a <=( a52918a  and  a52905a );
 a1259a <=( a52892a  and  a52879a );
 a1260a <=( a52866a  and  a52853a );
 a1261a <=( a52840a  and  a52827a );
 a1262a <=( a52814a  and  a52801a );
 a1263a <=( a52788a  and  a52775a );
 a1264a <=( a52762a  and  a52749a );
 a1265a <=( a52736a  and  a52723a );
 a1266a <=( a52710a  and  a52697a );
 a1267a <=( a52684a  and  a52671a );
 a1268a <=( a52658a  and  a52645a );
 a1269a <=( a52632a  and  a52619a );
 a1270a <=( a52606a  and  a52593a );
 a1271a <=( a52580a  and  a52567a );
 a1272a <=( a52554a  and  a52541a );
 a1273a <=( a52528a  and  a52515a );
 a1274a <=( a52502a  and  a52489a );
 a1275a <=( a52476a  and  a52463a );
 a1276a <=( a52450a  and  a52437a );
 a1277a <=( a52424a  and  a52411a );
 a1278a <=( a52398a  and  a52385a );
 a1279a <=( a52372a  and  a52359a );
 a1280a <=( a52346a  and  a52333a );
 a1281a <=( a52320a  and  a52307a );
 a1282a <=( a52294a  and  a52281a );
 a1283a <=( a52268a  and  a52255a );
 a1284a <=( a52242a  and  a52229a );
 a1285a <=( a52216a  and  a52203a );
 a1286a <=( a52190a  and  a52177a );
 a1287a <=( a52164a  and  a52151a );
 a1288a <=( a52138a  and  a52125a );
 a1289a <=( a52112a  and  a52099a );
 a1290a <=( a52086a  and  a52073a );
 a1291a <=( a52060a  and  a52047a );
 a1292a <=( a52034a  and  a52021a );
 a1293a <=( a52008a  and  a51995a );
 a1294a <=( a51982a  and  a51969a );
 a1295a <=( a51956a  and  a51943a );
 a1296a <=( a51930a  and  a51917a );
 a1297a <=( a51904a  and  a51891a );
 a1298a <=( a51878a  and  a51865a );
 a1299a <=( a51852a  and  a51839a );
 a1300a <=( a51826a  and  a51813a );
 a1301a <=( a51800a  and  a51787a );
 a1302a <=( a51774a  and  a51761a );
 a1303a <=( a51748a  and  a51735a );
 a1304a <=( a51722a  and  a51709a );
 a1305a <=( a51696a  and  a51683a );
 a1306a <=( a51670a  and  a51657a );
 a1307a <=( a51644a  and  a51631a );
 a1308a <=( a51618a  and  a51605a );
 a1309a <=( a51592a  and  a51579a );
 a1310a <=( a51566a  and  a51553a );
 a1311a <=( a51540a  and  a51527a );
 a1312a <=( a51514a  and  a51501a );
 a1313a <=( a51488a  and  a51475a );
 a1314a <=( a51462a  and  a51449a );
 a1315a <=( a51436a  and  a51423a );
 a1316a <=( a51410a  and  a51397a );
 a1317a <=( a51384a  and  a51371a );
 a1318a <=( a51358a  and  a51345a );
 a1319a <=( a51332a  and  a51319a );
 a1320a <=( a51306a  and  a51293a );
 a1321a <=( a51280a  and  a51267a );
 a1322a <=( a51254a  and  a51241a );
 a1323a <=( a51228a  and  a51215a );
 a1324a <=( a51202a  and  a51189a );
 a1325a <=( a51176a  and  a51163a );
 a1326a <=( a51150a  and  a51137a );
 a1327a <=( a51124a  and  a51111a );
 a1328a <=( a51098a  and  a51085a );
 a1329a <=( a51072a  and  a51059a );
 a1330a <=( a51046a  and  a51033a );
 a1331a <=( a51020a  and  a51007a );
 a1332a <=( a50994a  and  a50981a );
 a1333a <=( a50968a  and  a50955a );
 a1334a <=( a50942a  and  a50929a );
 a1335a <=( a50916a  and  a50903a );
 a1336a <=( a50890a  and  a50877a );
 a1337a <=( a50864a  and  a50851a );
 a1338a <=( a50838a  and  a50825a );
 a1339a <=( a50812a  and  a50799a );
 a1340a <=( a50786a  and  a50773a );
 a1341a <=( a50760a  and  a50747a );
 a1342a <=( a50734a  and  a50721a );
 a1343a <=( a50708a  and  a50695a );
 a1344a <=( a50682a  and  a50669a );
 a1345a <=( a50656a  and  a50643a );
 a1346a <=( a50630a  and  a50617a );
 a1347a <=( a50604a  and  a50591a );
 a1348a <=( a50578a  and  a50565a );
 a1349a <=( a50552a  and  a50539a );
 a1350a <=( a50526a  and  a50513a );
 a1351a <=( a50500a  and  a50487a );
 a1352a <=( a50474a  and  a50461a );
 a1353a <=( a50448a  and  a50435a );
 a1354a <=( a50422a  and  a50409a );
 a1355a <=( a50396a  and  a50383a );
 a1356a <=( a50370a  and  a50357a );
 a1357a <=( a50344a  and  a50331a );
 a1358a <=( a50318a  and  a50305a );
 a1359a <=( a50292a  and  a50279a );
 a1360a <=( a50266a  and  a50253a );
 a1361a <=( a50240a  and  a50227a );
 a1362a <=( a50214a  and  a50201a );
 a1363a <=( a50188a  and  a50175a );
 a1364a <=( a50162a  and  a50149a );
 a1365a <=( a50136a  and  a50123a );
 a1366a <=( a50110a  and  a50097a );
 a1367a <=( a50084a  and  a50071a );
 a1368a <=( a50058a  and  a50045a );
 a1369a <=( a50032a  and  a50019a );
 a1370a <=( a50006a  and  a49993a );
 a1371a <=( a49980a  and  a49967a );
 a1372a <=( a49954a  and  a49941a );
 a1373a <=( a49928a  and  a49915a );
 a1374a <=( a49902a  and  a49889a );
 a1375a <=( a49876a  and  a49863a );
 a1376a <=( a49850a  and  a49837a );
 a1377a <=( a49824a  and  a49811a );
 a1378a <=( a49798a  and  a49785a );
 a1379a <=( a49772a  and  a49759a );
 a1380a <=( a49746a  and  a49733a );
 a1381a <=( a49720a  and  a49707a );
 a1382a <=( a49694a  and  a49681a );
 a1383a <=( a49668a  and  a49655a );
 a1384a <=( a49642a  and  a49629a );
 a1385a <=( a49616a  and  a49603a );
 a1386a <=( a49590a  and  a49577a );
 a1387a <=( a49564a  and  a49551a );
 a1388a <=( a49538a  and  a49525a );
 a1389a <=( a49512a  and  a49499a );
 a1390a <=( a49486a  and  a49473a );
 a1391a <=( a49460a  and  a49447a );
 a1392a <=( a49434a  and  a49421a );
 a1393a <=( a49408a  and  a49395a );
 a1394a <=( a49382a  and  a49369a );
 a1395a <=( a49356a  and  a49343a );
 a1396a <=( a49330a  and  a49317a );
 a1397a <=( a49304a  and  a49291a );
 a1398a <=( a49278a  and  a49265a );
 a1399a <=( a49252a  and  a49239a );
 a1400a <=( a49226a  and  a49213a );
 a1401a <=( a49200a  and  a49187a );
 a1402a <=( a49174a  and  a49161a );
 a1403a <=( a49148a  and  a49135a );
 a1404a <=( a49122a  and  a49109a );
 a1405a <=( a49096a  and  a49083a );
 a1406a <=( a49070a  and  a49057a );
 a1407a <=( a49044a  and  a49031a );
 a1408a <=( a49018a  and  a49005a );
 a1409a <=( a48992a  and  a48979a );
 a1410a <=( a48966a  and  a48953a );
 a1411a <=( a48940a  and  a48927a );
 a1412a <=( a48914a  and  a48901a );
 a1413a <=( a48888a  and  a48875a );
 a1414a <=( a48862a  and  a48849a );
 a1415a <=( a48836a  and  a48823a );
 a1416a <=( a48810a  and  a48797a );
 a1417a <=( a48784a  and  a48771a );
 a1418a <=( a48758a  and  a48745a );
 a1419a <=( a48732a  and  a48719a );
 a1420a <=( a48706a  and  a48693a );
 a1421a <=( a48680a  and  a48667a );
 a1422a <=( a48654a  and  a48641a );
 a1423a <=( a48628a  and  a48615a );
 a1424a <=( a48602a  and  a48589a );
 a1425a <=( a48576a  and  a48563a );
 a1426a <=( a48550a  and  a48537a );
 a1427a <=( a48524a  and  a48511a );
 a1428a <=( a48498a  and  a48485a );
 a1429a <=( a48472a  and  a48459a );
 a1430a <=( a48446a  and  a48433a );
 a1431a <=( a48420a  and  a48407a );
 a1432a <=( a48394a  and  a48381a );
 a1433a <=( a48368a  and  a48355a );
 a1434a <=( a48342a  and  a48329a );
 a1435a <=( a48316a  and  a48303a );
 a1436a <=( a48290a  and  a48277a );
 a1437a <=( a48264a  and  a48251a );
 a1438a <=( a48238a  and  a48225a );
 a1439a <=( a48212a  and  a48199a );
 a1440a <=( a48186a  and  a48173a );
 a1441a <=( a48160a  and  a48147a );
 a1442a <=( a48134a  and  a48121a );
 a1443a <=( a48108a  and  a48095a );
 a1444a <=( a48082a  and  a48069a );
 a1445a <=( a48056a  and  a48043a );
 a1446a <=( a48030a  and  a48017a );
 a1447a <=( a48004a  and  a47991a );
 a1448a <=( a47978a  and  a47965a );
 a1449a <=( a47952a  and  a47939a );
 a1450a <=( a47926a  and  a47913a );
 a1451a <=( a47900a  and  a47887a );
 a1452a <=( a47874a  and  a47861a );
 a1453a <=( a47848a  and  a47835a );
 a1454a <=( a47822a  and  a47809a );
 a1455a <=( a47796a  and  a47783a );
 a1456a <=( a47770a  and  a47757a );
 a1457a <=( a47744a  and  a47731a );
 a1458a <=( a47718a  and  a47705a );
 a1459a <=( a47692a  and  a47679a );
 a1460a <=( a47666a  and  a47653a );
 a1461a <=( a47640a  and  a47627a );
 a1462a <=( a47614a  and  a47601a );
 a1463a <=( a47588a  and  a47575a );
 a1464a <=( a47562a  and  a47549a );
 a1465a <=( a47536a  and  a47523a );
 a1466a <=( a47510a  and  a47497a );
 a1467a <=( a47484a  and  a47471a );
 a1468a <=( a47458a  and  a47445a );
 a1469a <=( a47432a  and  a47419a );
 a1470a <=( a47406a  and  a47393a );
 a1471a <=( a47380a  and  a47367a );
 a1472a <=( a47354a  and  a47341a );
 a1473a <=( a47328a  and  a47315a );
 a1474a <=( a47302a  and  a47289a );
 a1475a <=( a47276a  and  a47263a );
 a1476a <=( a47250a  and  a47237a );
 a1477a <=( a47224a  and  a47211a );
 a1478a <=( a47198a  and  a47185a );
 a1479a <=( a47172a  and  a47159a );
 a1480a <=( a47146a  and  a47133a );
 a1481a <=( a47120a  and  a47107a );
 a1482a <=( a47094a  and  a47081a );
 a1483a <=( a47068a  and  a47055a );
 a1484a <=( a47042a  and  a47029a );
 a1485a <=( a47016a  and  a47003a );
 a1486a <=( a46990a  and  a46977a );
 a1487a <=( a46964a  and  a46951a );
 a1488a <=( a46938a  and  a46925a );
 a1489a <=( a46912a  and  a46899a );
 a1490a <=( a46886a  and  a46873a );
 a1491a <=( a46860a  and  a46847a );
 a1492a <=( a46834a  and  a46821a );
 a1493a <=( a46808a  and  a46795a );
 a1494a <=( a46782a  and  a46769a );
 a1495a <=( a46756a  and  a46743a );
 a1496a <=( a46730a  and  a46717a );
 a1497a <=( a46704a  and  a46691a );
 a1498a <=( a46678a  and  a46665a );
 a1499a <=( a46652a  and  a46639a );
 a1500a <=( a46626a  and  a46613a );
 a1501a <=( a46600a  and  a46587a );
 a1502a <=( a46574a  and  a46561a );
 a1503a <=( a46548a  and  a46535a );
 a1504a <=( a46522a  and  a46509a );
 a1505a <=( a46496a  and  a46483a );
 a1506a <=( a46470a  and  a46457a );
 a1507a <=( a46444a  and  a46431a );
 a1508a <=( a46418a  and  a46405a );
 a1509a <=( a46392a  and  a46379a );
 a1510a <=( a46366a  and  a46353a );
 a1511a <=( a46340a  and  a46327a );
 a1512a <=( a46314a  and  a46301a );
 a1513a <=( a46288a  and  a46275a );
 a1514a <=( a46262a  and  a46249a );
 a1515a <=( a46236a  and  a46223a );
 a1516a <=( a46210a  and  a46197a );
 a1517a <=( a46184a  and  a46171a );
 a1518a <=( a46158a  and  a46145a );
 a1519a <=( a46132a  and  a46119a );
 a1520a <=( a46106a  and  a46093a );
 a1521a <=( a46080a  and  a46067a );
 a1522a <=( a46054a  and  a46041a );
 a1523a <=( a46028a  and  a46015a );
 a1524a <=( a46002a  and  a45989a );
 a1525a <=( a45976a  and  a45963a );
 a1526a <=( a45950a  and  a45937a );
 a1527a <=( a45924a  and  a45911a );
 a1528a <=( a45898a  and  a45885a );
 a1529a <=( a45872a  and  a45859a );
 a1530a <=( a45846a  and  a45833a );
 a1531a <=( a45820a  and  a45807a );
 a1532a <=( a45794a  and  a45781a );
 a1533a <=( a45768a  and  a45755a );
 a1534a <=( a45742a  and  a45729a );
 a1535a <=( a45716a  and  a45703a );
 a1536a <=( a45690a  and  a45677a );
 a1537a <=( a45664a  and  a45651a );
 a1538a <=( a45638a  and  a45625a );
 a1539a <=( a45612a  and  a45599a );
 a1540a <=( a45586a  and  a45573a );
 a1541a <=( a45560a  and  a45547a );
 a1542a <=( a45534a  and  a45521a );
 a1543a <=( a45508a  and  a45495a );
 a1544a <=( a45482a  and  a45469a );
 a1545a <=( a45456a  and  a45443a );
 a1546a <=( a45430a  and  a45417a );
 a1547a <=( a45404a  and  a45391a );
 a1548a <=( a45378a  and  a45365a );
 a1549a <=( a45352a  and  a45339a );
 a1550a <=( a45326a  and  a45313a );
 a1551a <=( a45300a  and  a45287a );
 a1552a <=( a45274a  and  a45261a );
 a1553a <=( a45248a  and  a45235a );
 a1554a <=( a45222a  and  a45209a );
 a1555a <=( a45196a  and  a45183a );
 a1556a <=( a45170a  and  a45157a );
 a1557a <=( a45144a  and  a45131a );
 a1558a <=( a45118a  and  a45105a );
 a1559a <=( a45092a  and  a45079a );
 a1560a <=( a45066a  and  a45053a );
 a1561a <=( a45040a  and  a45027a );
 a1562a <=( a45014a  and  a45001a );
 a1563a <=( a44988a  and  a44975a );
 a1564a <=( a44962a  and  a44949a );
 a1565a <=( a44936a  and  a44923a );
 a1566a <=( a44910a  and  a44897a );
 a1567a <=( a44884a  and  a44871a );
 a1568a <=( a44858a  and  a44845a );
 a1569a <=( a44832a  and  a44819a );
 a1570a <=( a44806a  and  a44793a );
 a1571a <=( a44780a  and  a44767a );
 a1572a <=( a44754a  and  a44741a );
 a1573a <=( a44728a  and  a44715a );
 a1574a <=( a44702a  and  a44689a );
 a1575a <=( a44676a  and  a44663a );
 a1576a <=( a44650a  and  a44637a );
 a1577a <=( a44624a  and  a44611a );
 a1578a <=( a44598a  and  a44585a );
 a1579a <=( a44572a  and  a44559a );
 a1580a <=( a44546a  and  a44533a );
 a1581a <=( a44520a  and  a44507a );
 a1582a <=( a44494a  and  a44481a );
 a1583a <=( a44468a  and  a44455a );
 a1584a <=( a44442a  and  a44429a );
 a1585a <=( a44416a  and  a44403a );
 a1586a <=( a44390a  and  a44377a );
 a1587a <=( a44364a  and  a44351a );
 a1588a <=( a44338a  and  a44325a );
 a1589a <=( a44312a  and  a44299a );
 a1590a <=( a44286a  and  a44273a );
 a1591a <=( a44260a  and  a44247a );
 a1592a <=( a44234a  and  a44221a );
 a1593a <=( a44208a  and  a44195a );
 a1594a <=( a44182a  and  a44169a );
 a1595a <=( a44156a  and  a44143a );
 a1596a <=( a44130a  and  a44117a );
 a1597a <=( a44104a  and  a44091a );
 a1598a <=( a44078a  and  a44065a );
 a1599a <=( a44052a  and  a44039a );
 a1600a <=( a44026a  and  a44013a );
 a1601a <=( a44000a  and  a43987a );
 a1602a <=( a43974a  and  a43961a );
 a1603a <=( a43948a  and  a43935a );
 a1604a <=( a43922a  and  a43909a );
 a1605a <=( a43896a  and  a43883a );
 a1606a <=( a43870a  and  a43857a );
 a1607a <=( a43844a  and  a43831a );
 a1608a <=( a43818a  and  a43805a );
 a1609a <=( a43792a  and  a43779a );
 a1610a <=( a43766a  and  a43753a );
 a1611a <=( a43740a  and  a43727a );
 a1612a <=( a43714a  and  a43701a );
 a1613a <=( a43688a  and  a43675a );
 a1614a <=( a43662a  and  a43649a );
 a1615a <=( a43636a  and  a43623a );
 a1616a <=( a43610a  and  a43597a );
 a1617a <=( a43584a  and  a43571a );
 a1618a <=( a43558a  and  a43545a );
 a1619a <=( a43532a  and  a43519a );
 a1620a <=( a43506a  and  a43493a );
 a1621a <=( a43480a  and  a43467a );
 a1622a <=( a43454a  and  a43441a );
 a1623a <=( a43428a  and  a43415a );
 a1624a <=( a43402a  and  a43389a );
 a1625a <=( a43376a  and  a43363a );
 a1626a <=( a43350a  and  a43337a );
 a1627a <=( a43324a  and  a43311a );
 a1628a <=( a43298a  and  a43285a );
 a1629a <=( a43272a  and  a43259a );
 a1630a <=( a43246a  and  a43233a );
 a1631a <=( a43220a  and  a43207a );
 a1632a <=( a43194a  and  a43181a );
 a1633a <=( a43168a  and  a43155a );
 a1634a <=( a43142a  and  a43129a );
 a1635a <=( a43116a  and  a43103a );
 a1636a <=( a43090a  and  a43077a );
 a1637a <=( a43064a  and  a43051a );
 a1638a <=( a43038a  and  a43025a );
 a1639a <=( a43012a  and  a42999a );
 a1640a <=( a42986a  and  a42973a );
 a1641a <=( a42960a  and  a42947a );
 a1642a <=( a42934a  and  a42921a );
 a1643a <=( a42908a  and  a42895a );
 a1644a <=( a42882a  and  a42869a );
 a1645a <=( a42856a  and  a42843a );
 a1646a <=( a42830a  and  a42817a );
 a1647a <=( a42804a  and  a42791a );
 a1648a <=( a42778a  and  a42765a );
 a1649a <=( a42752a  and  a42739a );
 a1650a <=( a42726a  and  a42713a );
 a1651a <=( a42700a  and  a42687a );
 a1652a <=( a42674a  and  a42661a );
 a1653a <=( a42648a  and  a42635a );
 a1654a <=( a42622a  and  a42609a );
 a1655a <=( a42596a  and  a42583a );
 a1656a <=( a42570a  and  a42557a );
 a1657a <=( a42544a  and  a42531a );
 a1658a <=( a42518a  and  a42505a );
 a1659a <=( a42492a  and  a42479a );
 a1660a <=( a42468a  and  a42455a );
 a1661a <=( a42444a  and  a42431a );
 a1662a <=( a42420a  and  a42407a );
 a1663a <=( a42396a  and  a42383a );
 a1664a <=( a42372a  and  a42359a );
 a1665a <=( a42348a  and  a42335a );
 a1666a <=( a42324a  and  a42311a );
 a1667a <=( a42300a  and  a42287a );
 a1668a <=( a42276a  and  a42263a );
 a1669a <=( a42252a  and  a42239a );
 a1670a <=( a42228a  and  a42215a );
 a1671a <=( a42204a  and  a42191a );
 a1672a <=( a42180a  and  a42167a );
 a1673a <=( a42156a  and  a42143a );
 a1674a <=( a42132a  and  a42119a );
 a1675a <=( a42108a  and  a42095a );
 a1676a <=( a42084a  and  a42071a );
 a1677a <=( a42060a  and  a42047a );
 a1678a <=( a42036a  and  a42023a );
 a1679a <=( a42012a  and  a41999a );
 a1680a <=( a41988a  and  a41975a );
 a1681a <=( a41964a  and  a41951a );
 a1682a <=( a41940a  and  a41927a );
 a1683a <=( a41916a  and  a41903a );
 a1684a <=( a41892a  and  a41879a );
 a1685a <=( a41868a  and  a41855a );
 a1686a <=( a41844a  and  a41831a );
 a1687a <=( a41820a  and  a41807a );
 a1688a <=( a41796a  and  a41783a );
 a1689a <=( a41772a  and  a41759a );
 a1690a <=( a41748a  and  a41735a );
 a1691a <=( a41724a  and  a41711a );
 a1692a <=( a41700a  and  a41687a );
 a1693a <=( a41676a  and  a41663a );
 a1694a <=( a41652a  and  a41639a );
 a1695a <=( a41628a  and  a41615a );
 a1696a <=( a41604a  and  a41591a );
 a1697a <=( a41580a  and  a41567a );
 a1698a <=( a41556a  and  a41543a );
 a1699a <=( a41532a  and  a41519a );
 a1700a <=( a41508a  and  a41495a );
 a1701a <=( a41484a  and  a41471a );
 a1702a <=( a41460a  and  a41447a );
 a1703a <=( a41436a  and  a41423a );
 a1704a <=( a41412a  and  a41399a );
 a1705a <=( a41388a  and  a41375a );
 a1706a <=( a41364a  and  a41351a );
 a1707a <=( a41340a  and  a41327a );
 a1708a <=( a41316a  and  a41303a );
 a1709a <=( a41292a  and  a41279a );
 a1710a <=( a41268a  and  a41255a );
 a1711a <=( a41244a  and  a41231a );
 a1712a <=( a41220a  and  a41207a );
 a1713a <=( a41196a  and  a41183a );
 a1714a <=( a41172a  and  a41159a );
 a1715a <=( a41148a  and  a41135a );
 a1716a <=( a41124a  and  a41111a );
 a1717a <=( a41100a  and  a41087a );
 a1718a <=( a41076a  and  a41063a );
 a1719a <=( a41052a  and  a41039a );
 a1720a <=( a41028a  and  a41015a );
 a1721a <=( a41004a  and  a40991a );
 a1722a <=( a40980a  and  a40967a );
 a1723a <=( a40956a  and  a40943a );
 a1724a <=( a40932a  and  a40919a );
 a1725a <=( a40908a  and  a40895a );
 a1726a <=( a40884a  and  a40871a );
 a1727a <=( a40860a  and  a40847a );
 a1728a <=( a40836a  and  a40823a );
 a1729a <=( a40812a  and  a40799a );
 a1730a <=( a40788a  and  a40775a );
 a1731a <=( a40764a  and  a40751a );
 a1732a <=( a40740a  and  a40727a );
 a1733a <=( a40716a  and  a40703a );
 a1734a <=( a40692a  and  a40679a );
 a1735a <=( a40668a  and  a40655a );
 a1736a <=( a40644a  and  a40631a );
 a1737a <=( a40620a  and  a40607a );
 a1738a <=( a40596a  and  a40583a );
 a1739a <=( a40572a  and  a40559a );
 a1740a <=( a40548a  and  a40535a );
 a1741a <=( a40524a  and  a40511a );
 a1742a <=( a40500a  and  a40487a );
 a1743a <=( a40476a  and  a40463a );
 a1744a <=( a40452a  and  a40439a );
 a1745a <=( a40428a  and  a40415a );
 a1746a <=( a40404a  and  a40391a );
 a1747a <=( a40380a  and  a40367a );
 a1748a <=( a40356a  and  a40343a );
 a1749a <=( a40332a  and  a40319a );
 a1750a <=( a40308a  and  a40295a );
 a1751a <=( a40284a  and  a40271a );
 a1752a <=( a40260a  and  a40247a );
 a1753a <=( a40236a  and  a40223a );
 a1754a <=( a40212a  and  a40199a );
 a1755a <=( a40188a  and  a40175a );
 a1756a <=( a40164a  and  a40151a );
 a1757a <=( a40140a  and  a40127a );
 a1758a <=( a40116a  and  a40103a );
 a1759a <=( a40092a  and  a40079a );
 a1760a <=( a40068a  and  a40055a );
 a1761a <=( a40044a  and  a40031a );
 a1762a <=( a40020a  and  a40007a );
 a1763a <=( a39996a  and  a39983a );
 a1764a <=( a39972a  and  a39959a );
 a1765a <=( a39948a  and  a39935a );
 a1766a <=( a39924a  and  a39911a );
 a1767a <=( a39900a  and  a39887a );
 a1768a <=( a39876a  and  a39863a );
 a1769a <=( a39852a  and  a39839a );
 a1770a <=( a39828a  and  a39815a );
 a1771a <=( a39804a  and  a39791a );
 a1772a <=( a39780a  and  a39767a );
 a1773a <=( a39756a  and  a39743a );
 a1774a <=( a39732a  and  a39719a );
 a1775a <=( a39708a  and  a39695a );
 a1776a <=( a39684a  and  a39671a );
 a1777a <=( a39660a  and  a39647a );
 a1778a <=( a39636a  and  a39623a );
 a1779a <=( a39612a  and  a39599a );
 a1780a <=( a39588a  and  a39575a );
 a1781a <=( a39564a  and  a39551a );
 a1782a <=( a39540a  and  a39527a );
 a1783a <=( a39516a  and  a39503a );
 a1784a <=( a39492a  and  a39479a );
 a1785a <=( a39468a  and  a39455a );
 a1786a <=( a39444a  and  a39431a );
 a1787a <=( a39420a  and  a39407a );
 a1788a <=( a39396a  and  a39383a );
 a1789a <=( a39372a  and  a39359a );
 a1790a <=( a39348a  and  a39335a );
 a1791a <=( a39324a  and  a39311a );
 a1792a <=( a39300a  and  a39287a );
 a1793a <=( a39276a  and  a39263a );
 a1794a <=( a39252a  and  a39239a );
 a1795a <=( a39228a  and  a39215a );
 a1796a <=( a39204a  and  a39191a );
 a1797a <=( a39180a  and  a39167a );
 a1798a <=( a39156a  and  a39143a );
 a1799a <=( a39132a  and  a39119a );
 a1800a <=( a39108a  and  a39095a );
 a1801a <=( a39084a  and  a39071a );
 a1802a <=( a39060a  and  a39047a );
 a1803a <=( a39036a  and  a39023a );
 a1804a <=( a39012a  and  a38999a );
 a1805a <=( a38988a  and  a38975a );
 a1806a <=( a38964a  and  a38951a );
 a1807a <=( a38940a  and  a38927a );
 a1808a <=( a38916a  and  a38903a );
 a1809a <=( a38892a  and  a38879a );
 a1810a <=( a38868a  and  a38855a );
 a1811a <=( a38844a  and  a38831a );
 a1812a <=( a38820a  and  a38807a );
 a1813a <=( a38796a  and  a38783a );
 a1814a <=( a38772a  and  a38759a );
 a1815a <=( a38748a  and  a38735a );
 a1816a <=( a38724a  and  a38711a );
 a1817a <=( a38700a  and  a38687a );
 a1818a <=( a38676a  and  a38663a );
 a1819a <=( a38652a  and  a38639a );
 a1820a <=( a38628a  and  a38615a );
 a1821a <=( a38604a  and  a38591a );
 a1822a <=( a38580a  and  a38567a );
 a1823a <=( a38556a  and  a38543a );
 a1824a <=( a38532a  and  a38519a );
 a1825a <=( a38508a  and  a38495a );
 a1826a <=( a38484a  and  a38471a );
 a1827a <=( a38460a  and  a38447a );
 a1828a <=( a38436a  and  a38423a );
 a1829a <=( a38412a  and  a38399a );
 a1830a <=( a38388a  and  a38375a );
 a1831a <=( a38364a  and  a38351a );
 a1832a <=( a38340a  and  a38327a );
 a1833a <=( a38316a  and  a38303a );
 a1834a <=( a38292a  and  a38279a );
 a1835a <=( a38268a  and  a38255a );
 a1836a <=( a38244a  and  a38231a );
 a1837a <=( a38220a  and  a38207a );
 a1838a <=( a38196a  and  a38183a );
 a1839a <=( a38172a  and  a38159a );
 a1840a <=( a38148a  and  a38135a );
 a1841a <=( a38124a  and  a38111a );
 a1842a <=( a38100a  and  a38087a );
 a1843a <=( a38076a  and  a38063a );
 a1844a <=( a38052a  and  a38039a );
 a1845a <=( a38028a  and  a38015a );
 a1846a <=( a38004a  and  a37991a );
 a1847a <=( a37980a  and  a37967a );
 a1848a <=( a37956a  and  a37943a );
 a1849a <=( a37932a  and  a37919a );
 a1850a <=( a37908a  and  a37895a );
 a1851a <=( a37884a  and  a37871a );
 a1852a <=( a37860a  and  a37847a );
 a1853a <=( a37836a  and  a37823a );
 a1854a <=( a37812a  and  a37799a );
 a1855a <=( a37788a  and  a37775a );
 a1856a <=( a37764a  and  a37751a );
 a1857a <=( a37740a  and  a37727a );
 a1858a <=( a37716a  and  a37703a );
 a1859a <=( a37692a  and  a37679a );
 a1860a <=( a37668a  and  a37655a );
 a1861a <=( a37644a  and  a37631a );
 a1862a <=( a37620a  and  a37607a );
 a1863a <=( a37596a  and  a37583a );
 a1864a <=( a37572a  and  a37559a );
 a1865a <=( a37548a  and  a37535a );
 a1866a <=( a37524a  and  a37511a );
 a1867a <=( a37500a  and  a37487a );
 a1868a <=( a37476a  and  a37463a );
 a1869a <=( a37452a  and  a37439a );
 a1870a <=( a37428a  and  a37415a );
 a1871a <=( a37404a  and  a37391a );
 a1872a <=( a37380a  and  a37367a );
 a1873a <=( a37356a  and  a37343a );
 a1874a <=( a37332a  and  a37319a );
 a1875a <=( a37308a  and  a37295a );
 a1876a <=( a37284a  and  a37271a );
 a1877a <=( a37260a  and  a37247a );
 a1878a <=( a37236a  and  a37223a );
 a1879a <=( a37212a  and  a37199a );
 a1880a <=( a37188a  and  a37175a );
 a1881a <=( a37164a  and  a37151a );
 a1882a <=( a37140a  and  a37127a );
 a1883a <=( a37116a  and  a37103a );
 a1884a <=( a37092a  and  a37079a );
 a1885a <=( a37068a  and  a37055a );
 a1886a <=( a37044a  and  a37031a );
 a1887a <=( a37020a  and  a37007a );
 a1888a <=( a36996a  and  a36983a );
 a1889a <=( a36972a  and  a36959a );
 a1890a <=( a36948a  and  a36935a );
 a1891a <=( a36924a  and  a36911a );
 a1892a <=( a36900a  and  a36887a );
 a1893a <=( a36876a  and  a36863a );
 a1894a <=( a36852a  and  a36839a );
 a1895a <=( a36828a  and  a36815a );
 a1896a <=( a36804a  and  a36791a );
 a1897a <=( a36780a  and  a36767a );
 a1898a <=( a36756a  and  a36743a );
 a1899a <=( a36732a  and  a36719a );
 a1900a <=( a36708a  and  a36695a );
 a1901a <=( a36684a  and  a36671a );
 a1902a <=( a36660a  and  a36647a );
 a1903a <=( a36636a  and  a36623a );
 a1904a <=( a36612a  and  a36599a );
 a1905a <=( a36588a  and  a36575a );
 a1906a <=( a36564a  and  a36551a );
 a1907a <=( a36540a  and  a36527a );
 a1908a <=( a36516a  and  a36503a );
 a1909a <=( a36492a  and  a36479a );
 a1910a <=( a36468a  and  a36455a );
 a1911a <=( a36444a  and  a36431a );
 a1912a <=( a36420a  and  a36407a );
 a1913a <=( a36396a  and  a36383a );
 a1914a <=( a36372a  and  a36359a );
 a1915a <=( a36348a  and  a36335a );
 a1916a <=( a36324a  and  a36311a );
 a1917a <=( a36300a  and  a36287a );
 a1918a <=( a36276a  and  a36263a );
 a1919a <=( a36252a  and  a36239a );
 a1920a <=( a36228a  and  a36215a );
 a1921a <=( a36204a  and  a36191a );
 a1922a <=( a36180a  and  a36167a );
 a1923a <=( a36156a  and  a36143a );
 a1924a <=( a36132a  and  a36119a );
 a1925a <=( a36108a  and  a36095a );
 a1926a <=( a36084a  and  a36071a );
 a1927a <=( a36060a  and  a36047a );
 a1928a <=( a36036a  and  a36023a );
 a1929a <=( a36012a  and  a35999a );
 a1930a <=( a35988a  and  a35975a );
 a1931a <=( a35964a  and  a35951a );
 a1932a <=( a35940a  and  a35927a );
 a1933a <=( a35916a  and  a35903a );
 a1934a <=( a35892a  and  a35879a );
 a1935a <=( a35868a  and  a35855a );
 a1936a <=( a35844a  and  a35831a );
 a1937a <=( a35820a  and  a35807a );
 a1938a <=( a35796a  and  a35783a );
 a1939a <=( a35772a  and  a35759a );
 a1940a <=( a35748a  and  a35735a );
 a1941a <=( a35724a  and  a35711a );
 a1942a <=( a35700a  and  a35687a );
 a1943a <=( a35676a  and  a35663a );
 a1944a <=( a35652a  and  a35639a );
 a1945a <=( a35628a  and  a35615a );
 a1946a <=( a35604a  and  a35591a );
 a1947a <=( a35580a  and  a35567a );
 a1948a <=( a35556a  and  a35543a );
 a1949a <=( a35532a  and  a35519a );
 a1950a <=( a35508a  and  a35495a );
 a1951a <=( a35484a  and  a35471a );
 a1952a <=( a35460a  and  a35447a );
 a1953a <=( a35436a  and  a35423a );
 a1954a <=( a35412a  and  a35399a );
 a1955a <=( a35388a  and  a35375a );
 a1956a <=( a35364a  and  a35351a );
 a1957a <=( a35340a  and  a35327a );
 a1958a <=( a35316a  and  a35303a );
 a1959a <=( a35292a  and  a35279a );
 a1960a <=( a35268a  and  a35255a );
 a1961a <=( a35244a  and  a35231a );
 a1962a <=( a35220a  and  a35207a );
 a1963a <=( a35196a  and  a35183a );
 a1964a <=( a35172a  and  a35159a );
 a1965a <=( a35148a  and  a35135a );
 a1966a <=( a35124a  and  a35111a );
 a1967a <=( a35100a  and  a35087a );
 a1968a <=( a35076a  and  a35063a );
 a1969a <=( a35052a  and  a35039a );
 a1970a <=( a35028a  and  a35015a );
 a1971a <=( a35004a  and  a34991a );
 a1972a <=( a34980a  and  a34967a );
 a1973a <=( a34956a  and  a34943a );
 a1974a <=( a34932a  and  a34919a );
 a1975a <=( a34908a  and  a34895a );
 a1976a <=( a34884a  and  a34871a );
 a1977a <=( a34860a  and  a34847a );
 a1978a <=( a34836a  and  a34823a );
 a1979a <=( a34812a  and  a34799a );
 a1980a <=( a34788a  and  a34775a );
 a1981a <=( a34764a  and  a34751a );
 a1982a <=( a34740a  and  a34727a );
 a1983a <=( a34716a  and  a34703a );
 a1984a <=( a34692a  and  a34679a );
 a1985a <=( a34668a  and  a34655a );
 a1986a <=( a34644a  and  a34631a );
 a1987a <=( a34620a  and  a34607a );
 a1988a <=( a34596a  and  a34583a );
 a1989a <=( a34572a  and  a34559a );
 a1990a <=( a34548a  and  a34535a );
 a1991a <=( a34524a  and  a34511a );
 a1992a <=( a34500a  and  a34487a );
 a1993a <=( a34476a  and  a34463a );
 a1994a <=( a34452a  and  a34439a );
 a1995a <=( a34428a  and  a34415a );
 a1996a <=( a34404a  and  a34391a );
 a1997a <=( a34380a  and  a34367a );
 a1998a <=( a34356a  and  a34343a );
 a1999a <=( a34332a  and  a34319a );
 a2000a <=( a34308a  and  a34295a );
 a2001a <=( a34284a  and  a34271a );
 a2002a <=( a34260a  and  a34247a );
 a2003a <=( a34236a  and  a34223a );
 a2004a <=( a34212a  and  a34199a );
 a2005a <=( a34188a  and  a34175a );
 a2006a <=( a34164a  and  a34151a );
 a2007a <=( a34140a  and  a34127a );
 a2008a <=( a34116a  and  a34103a );
 a2009a <=( a34092a  and  a34079a );
 a2010a <=( a34068a  and  a34055a );
 a2011a <=( a34044a  and  a34031a );
 a2012a <=( a34020a  and  a34007a );
 a2013a <=( a33996a  and  a33983a );
 a2014a <=( a33972a  and  a33959a );
 a2015a <=( a33948a  and  a33935a );
 a2016a <=( a33924a  and  a33911a );
 a2017a <=( a33900a  and  a33887a );
 a2018a <=( a33876a  and  a33863a );
 a2019a <=( a33852a  and  a33839a );
 a2020a <=( a33828a  and  a33815a );
 a2021a <=( a33804a  and  a33791a );
 a2022a <=( a33780a  and  a33767a );
 a2023a <=( a33756a  and  a33743a );
 a2024a <=( a33732a  and  a33719a );
 a2025a <=( a33708a  and  a33695a );
 a2026a <=( a33684a  and  a33671a );
 a2027a <=( a33660a  and  a33647a );
 a2028a <=( a33636a  and  a33623a );
 a2029a <=( a33612a  and  a33599a );
 a2030a <=( a33588a  and  a33575a );
 a2031a <=( a33564a  and  a33551a );
 a2032a <=( a33540a  and  a33527a );
 a2033a <=( a33516a  and  a33503a );
 a2034a <=( a33492a  and  a33479a );
 a2035a <=( a33468a  and  a33455a );
 a2036a <=( a33444a  and  a33431a );
 a2037a <=( a33420a  and  a33407a );
 a2038a <=( a33396a  and  a33383a );
 a2039a <=( a33372a  and  a33359a );
 a2040a <=( a33348a  and  a33335a );
 a2041a <=( a33324a  and  a33311a );
 a2042a <=( a33300a  and  a33287a );
 a2043a <=( a33276a  and  a33263a );
 a2044a <=( a33252a  and  a33239a );
 a2045a <=( a33228a  and  a33215a );
 a2046a <=( a33204a  and  a33191a );
 a2047a <=( a33180a  and  a33167a );
 a2048a <=( a33156a  and  a33143a );
 a2049a <=( a33132a  and  a33119a );
 a2050a <=( a33108a  and  a33095a );
 a2051a <=( a33084a  and  a33071a );
 a2052a <=( a33060a  and  a33047a );
 a2053a <=( a33036a  and  a33023a );
 a2054a <=( a33012a  and  a32999a );
 a2055a <=( a32988a  and  a32975a );
 a2056a <=( a32964a  and  a32951a );
 a2057a <=( a32940a  and  a32927a );
 a2058a <=( a32916a  and  a32903a );
 a2059a <=( a32892a  and  a32879a );
 a2060a <=( a32868a  and  a32855a );
 a2061a <=( a32844a  and  a32831a );
 a2062a <=( a32820a  and  a32807a );
 a2063a <=( a32796a  and  a32783a );
 a2064a <=( a32772a  and  a32759a );
 a2065a <=( a32748a  and  a32735a );
 a2066a <=( a32724a  and  a32711a );
 a2067a <=( a32700a  and  a32687a );
 a2068a <=( a32676a  and  a32663a );
 a2069a <=( a32652a  and  a32639a );
 a2070a <=( a32628a  and  a32615a );
 a2071a <=( a32604a  and  a32591a );
 a2072a <=( a32580a  and  a32567a );
 a2073a <=( a32556a  and  a32543a );
 a2074a <=( a32532a  and  a32519a );
 a2075a <=( a32508a  and  a32495a );
 a2076a <=( a32484a  and  a32471a );
 a2077a <=( a32460a  and  a32447a );
 a2078a <=( a32436a  and  a32423a );
 a2079a <=( a32412a  and  a32399a );
 a2080a <=( a32388a  and  a32375a );
 a2081a <=( a32364a  and  a32351a );
 a2082a <=( a32340a  and  a32327a );
 a2083a <=( a32316a  and  a32303a );
 a2084a <=( a32292a  and  a32279a );
 a2085a <=( a32268a  and  a32255a );
 a2086a <=( a32244a  and  a32231a );
 a2087a <=( a32220a  and  a32207a );
 a2088a <=( a32196a  and  a32183a );
 a2089a <=( a32172a  and  a32159a );
 a2090a <=( a32148a  and  a32135a );
 a2091a <=( a32124a  and  a32111a );
 a2092a <=( a32100a  and  a32087a );
 a2093a <=( a32076a  and  a32063a );
 a2094a <=( a32052a  and  a32039a );
 a2095a <=( a32028a  and  a32015a );
 a2096a <=( a32004a  and  a31991a );
 a2097a <=( a31980a  and  a31967a );
 a2098a <=( a31956a  and  a31943a );
 a2099a <=( a31932a  and  a31919a );
 a2100a <=( a31908a  and  a31895a );
 a2101a <=( a31884a  and  a31871a );
 a2102a <=( a31860a  and  a31847a );
 a2103a <=( a31836a  and  a31823a );
 a2104a <=( a31812a  and  a31799a );
 a2105a <=( a31788a  and  a31775a );
 a2106a <=( a31764a  and  a31751a );
 a2107a <=( a31740a  and  a31727a );
 a2108a <=( a31716a  and  a31703a );
 a2109a <=( a31692a  and  a31679a );
 a2110a <=( a31668a  and  a31655a );
 a2111a <=( a31644a  and  a31631a );
 a2112a <=( a31620a  and  a31607a );
 a2113a <=( a31596a  and  a31583a );
 a2114a <=( a31572a  and  a31559a );
 a2115a <=( a31548a  and  a31535a );
 a2116a <=( a31524a  and  a31511a );
 a2117a <=( a31500a  and  a31487a );
 a2118a <=( a31476a  and  a31463a );
 a2119a <=( a31452a  and  a31439a );
 a2120a <=( a31428a  and  a31415a );
 a2121a <=( a31404a  and  a31391a );
 a2122a <=( a31380a  and  a31367a );
 a2123a <=( a31356a  and  a31343a );
 a2124a <=( a31332a  and  a31319a );
 a2125a <=( a31308a  and  a31295a );
 a2126a <=( a31284a  and  a31271a );
 a2127a <=( a31260a  and  a31247a );
 a2128a <=( a31236a  and  a31223a );
 a2129a <=( a31212a  and  a31199a );
 a2130a <=( a31188a  and  a31175a );
 a2131a <=( a31164a  and  a31151a );
 a2132a <=( a31140a  and  a31127a );
 a2133a <=( a31116a  and  a31103a );
 a2134a <=( a31092a  and  a31079a );
 a2135a <=( a31068a  and  a31055a );
 a2136a <=( a31044a  and  a31031a );
 a2137a <=( a31020a  and  a31007a );
 a2138a <=( a30996a  and  a30983a );
 a2139a <=( a30972a  and  a30959a );
 a2140a <=( a30948a  and  a30935a );
 a2141a <=( a30924a  and  a30911a );
 a2142a <=( a30900a  and  a30887a );
 a2143a <=( a30876a  and  a30863a );
 a2144a <=( a30852a  and  a30839a );
 a2145a <=( a30828a  and  a30815a );
 a2146a <=( a30804a  and  a30791a );
 a2147a <=( a30780a  and  a30767a );
 a2148a <=( a30756a  and  a30743a );
 a2149a <=( a30732a  and  a30719a );
 a2150a <=( a30708a  and  a30695a );
 a2151a <=( a30684a  and  a30671a );
 a2152a <=( a30660a  and  a30647a );
 a2153a <=( a30636a  and  a30623a );
 a2154a <=( a30612a  and  a30599a );
 a2155a <=( a30588a  and  a30575a );
 a2156a <=( a30564a  and  a30551a );
 a2157a <=( a30540a  and  a30527a );
 a2158a <=( a30516a  and  a30503a );
 a2159a <=( a30492a  and  a30479a );
 a2160a <=( a30468a  and  a30455a );
 a2161a <=( a30444a  and  a30431a );
 a2162a <=( a30420a  and  a30407a );
 a2163a <=( a30396a  and  a30383a );
 a2164a <=( a30372a  and  a30359a );
 a2165a <=( a30348a  and  a30335a );
 a2166a <=( a30324a  and  a30311a );
 a2167a <=( a30300a  and  a30287a );
 a2168a <=( a30276a  and  a30263a );
 a2169a <=( a30252a  and  a30239a );
 a2170a <=( a30228a  and  a30215a );
 a2171a <=( a30204a  and  a30191a );
 a2172a <=( a30180a  and  a30167a );
 a2173a <=( a30156a  and  a30143a );
 a2174a <=( a30132a  and  a30119a );
 a2175a <=( a30108a  and  a30095a );
 a2176a <=( a30084a  and  a30071a );
 a2177a <=( a30060a  and  a30047a );
 a2178a <=( a30036a  and  a30023a );
 a2179a <=( a30012a  and  a29999a );
 a2180a <=( a29988a  and  a29975a );
 a2181a <=( a29964a  and  a29951a );
 a2182a <=( a29940a  and  a29927a );
 a2183a <=( a29916a  and  a29903a );
 a2184a <=( a29892a  and  a29879a );
 a2185a <=( a29868a  and  a29855a );
 a2186a <=( a29844a  and  a29831a );
 a2187a <=( a29820a  and  a29807a );
 a2188a <=( a29796a  and  a29783a );
 a2189a <=( a29772a  and  a29759a );
 a2190a <=( a29748a  and  a29735a );
 a2191a <=( a29724a  and  a29711a );
 a2192a <=( a29700a  and  a29687a );
 a2193a <=( a29676a  and  a29663a );
 a2194a <=( a29652a  and  a29639a );
 a2195a <=( a29628a  and  a29615a );
 a2196a <=( a29604a  and  a29591a );
 a2197a <=( a29580a  and  a29567a );
 a2198a <=( a29556a  and  a29543a );
 a2199a <=( a29532a  and  a29519a );
 a2200a <=( a29508a  and  a29495a );
 a2201a <=( a29484a  and  a29473a );
 a2202a <=( a29462a  and  a29451a );
 a2203a <=( a29440a  and  a29429a );
 a2204a <=( a29418a  and  a29407a );
 a2205a <=( a29396a  and  a29385a );
 a2206a <=( a29374a  and  a29363a );
 a2207a <=( a29352a  and  a29341a );
 a2208a <=( a29330a  and  a29319a );
 a2209a <=( a29308a  and  a29297a );
 a2210a <=( a29286a  and  a29275a );
 a2211a <=( a29264a  and  a29253a );
 a2212a <=( a29242a  and  a29231a );
 a2213a <=( a29220a  and  a29209a );
 a2214a <=( a29198a  and  a29187a );
 a2215a <=( a29176a  and  a29165a );
 a2216a <=( a29154a  and  a29143a );
 a2217a <=( a29132a  and  a29121a );
 a2218a <=( a29110a  and  a29099a );
 a2219a <=( a29088a  and  a29077a );
 a2220a <=( a29066a  and  a29055a );
 a2221a <=( a29044a  and  a29033a );
 a2222a <=( a29022a  and  a29011a );
 a2223a <=( a29000a  and  a28989a );
 a2224a <=( a28978a  and  a28967a );
 a2225a <=( a28956a  and  a28945a );
 a2226a <=( a28934a  and  a28923a );
 a2227a <=( a28912a  and  a28901a );
 a2228a <=( a28890a  and  a28879a );
 a2229a <=( a28868a  and  a28857a );
 a2230a <=( a28846a  and  a28835a );
 a2231a <=( a28824a  and  a28813a );
 a2232a <=( a28802a  and  a28791a );
 a2233a <=( a28780a  and  a28769a );
 a2234a <=( a28758a  and  a28747a );
 a2235a <=( a28736a  and  a28725a );
 a2236a <=( a28714a  and  a28703a );
 a2237a <=( a28692a  and  a28681a );
 a2238a <=( a28670a  and  a28659a );
 a2239a <=( a28648a  and  a28637a );
 a2240a <=( a28626a  and  a28615a );
 a2241a <=( a28604a  and  a28593a );
 a2242a <=( a28582a  and  a28571a );
 a2243a <=( a28560a  and  a28549a );
 a2244a <=( a28538a  and  a28527a );
 a2245a <=( a28516a  and  a28505a );
 a2246a <=( a28494a  and  a28483a );
 a2247a <=( a28472a  and  a28461a );
 a2248a <=( a28450a  and  a28439a );
 a2249a <=( a28428a  and  a28417a );
 a2250a <=( a28406a  and  a28395a );
 a2251a <=( a28384a  and  a28373a );
 a2252a <=( a28362a  and  a28351a );
 a2253a <=( a28340a  and  a28329a );
 a2254a <=( a28318a  and  a28307a );
 a2255a <=( a28296a  and  a28285a );
 a2256a <=( a28274a  and  a28263a );
 a2257a <=( a28252a  and  a28241a );
 a2258a <=( a28230a  and  a28219a );
 a2259a <=( a28208a  and  a28197a );
 a2260a <=( a28186a  and  a28175a );
 a2261a <=( a28164a  and  a28153a );
 a2262a <=( a28142a  and  a28131a );
 a2263a <=( a28120a  and  a28109a );
 a2264a <=( a28098a  and  a28087a );
 a2265a <=( a28076a  and  a28065a );
 a2266a <=( a28054a  and  a28043a );
 a2267a <=( a28032a  and  a28021a );
 a2268a <=( a28010a  and  a27999a );
 a2269a <=( a27988a  and  a27977a );
 a2270a <=( a27966a  and  a27955a );
 a2271a <=( a27944a  and  a27933a );
 a2272a <=( a27922a  and  a27911a );
 a2273a <=( a27900a  and  a27889a );
 a2274a <=( a27878a  and  a27867a );
 a2275a <=( a27856a  and  a27845a );
 a2276a <=( a27834a  and  a27823a );
 a2277a <=( a27812a  and  a27801a );
 a2278a <=( a27790a  and  a27779a );
 a2279a <=( a27768a  and  a27757a );
 a2280a <=( a27746a  and  a27735a );
 a2281a <=( a27724a  and  a27713a );
 a2282a <=( a27702a  and  a27691a );
 a2283a <=( a27680a  and  a27669a );
 a2284a <=( a27658a  and  a27647a );
 a2285a <=( a27636a  and  a27625a );
 a2286a <=( a27614a  and  a27603a );
 a2287a <=( a27592a  and  a27581a );
 a2288a <=( a27570a  and  a27559a );
 a2289a <=( a27548a  and  a27537a );
 a2290a <=( a27526a  and  a27515a );
 a2291a <=( a27504a  and  a27493a );
 a2292a <=( a27482a  and  a27471a );
 a2293a <=( a27460a  and  a27449a );
 a2294a <=( a27438a  and  a27427a );
 a2295a <=( a27416a  and  a27405a );
 a2296a <=( a27394a  and  a27383a );
 a2297a <=( a27372a  and  a27361a );
 a2298a <=( a27350a  and  a27339a );
 a2299a <=( a27328a  and  a27317a );
 a2300a <=( a27306a  and  a27295a );
 a2301a <=( a27284a  and  a27273a );
 a2302a <=( a27262a  and  a27251a );
 a2303a <=( a27240a  and  a27229a );
 a2304a <=( a27218a  and  a27207a );
 a2305a <=( a27196a  and  a27185a );
 a2306a <=( a27174a  and  a27163a );
 a2307a <=( a27152a  and  a27141a );
 a2308a <=( a27130a  and  a27119a );
 a2309a <=( a27108a  and  a27097a );
 a2310a <=( a27086a  and  a27075a );
 a2311a <=( a27064a  and  a27053a );
 a2312a <=( a27042a  and  a27031a );
 a2313a <=( a27020a  and  a27009a );
 a2314a <=( a26998a  and  a26987a );
 a2315a <=( a26976a  and  a26965a );
 a2316a <=( a26954a  and  a26943a );
 a2317a <=( a26932a  and  a26921a );
 a2318a <=( a26910a  and  a26899a );
 a2319a <=( a26888a  and  a26877a );
 a2320a <=( a26866a  and  a26855a );
 a2321a <=( a26844a  and  a26833a );
 a2322a <=( a26822a  and  a26811a );
 a2323a <=( a26800a  and  a26789a );
 a2324a <=( a26778a  and  a26767a );
 a2325a <=( a26756a  and  a26745a );
 a2326a <=( a26734a  and  a26723a );
 a2327a <=( a26712a  and  a26701a );
 a2328a <=( a26690a  and  a26679a );
 a2329a <=( a26668a  and  a26657a );
 a2330a <=( a26646a  and  a26635a );
 a2331a <=( a26624a  and  a26613a );
 a2332a <=( a26602a  and  a26591a );
 a2333a <=( a26580a  and  a26569a );
 a2334a <=( a26558a  and  a26547a );
 a2335a <=( a26536a  and  a26525a );
 a2336a <=( a26514a  and  a26503a );
 a2337a <=( a26492a  and  a26481a );
 a2338a <=( a26470a  and  a26459a );
 a2339a <=( a26448a  and  a26437a );
 a2340a <=( a26426a  and  a26415a );
 a2341a <=( a26404a  and  a26393a );
 a2342a <=( a26382a  and  a26371a );
 a2343a <=( a26360a  and  a26349a );
 a2344a <=( a26338a  and  a26327a );
 a2345a <=( a26316a  and  a26305a );
 a2346a <=( a26294a  and  a26283a );
 a2347a <=( a26272a  and  a26261a );
 a2348a <=( a26250a  and  a26239a );
 a2349a <=( a26228a  and  a26217a );
 a2350a <=( a26206a  and  a26195a );
 a2351a <=( a26184a  and  a26173a );
 a2352a <=( a26162a  and  a26151a );
 a2353a <=( a26140a  and  a26129a );
 a2354a <=( a26118a  and  a26107a );
 a2355a <=( a26096a  and  a26085a );
 a2356a <=( a26074a  and  a26063a );
 a2357a <=( a26052a  and  a26041a );
 a2358a <=( a26030a  and  a26019a );
 a2359a <=( a26008a  and  a25997a );
 a2360a <=( a25986a  and  a25975a );
 a2361a <=( a25964a  and  a25953a );
 a2362a <=( a25942a  and  a25931a );
 a2363a <=( a25920a  and  a25909a );
 a2364a <=( a25898a  and  a25887a );
 a2365a <=( a25876a  and  a25865a );
 a2366a <=( a25854a  and  a25843a );
 a2367a <=( a25832a  and  a25821a );
 a2368a <=( a25810a  and  a25799a );
 a2369a <=( a25788a  and  a25777a );
 a2370a <=( a25766a  and  a25755a );
 a2371a <=( a25744a  and  a25733a );
 a2372a <=( a25722a  and  a25711a );
 a2373a <=( a25700a  and  a25689a );
 a2374a <=( a25678a  and  a25667a );
 a2375a <=( a25656a  and  a25645a );
 a2376a <=( a25634a  and  a25623a );
 a2377a <=( a25612a  and  a25601a );
 a2378a <=( a25590a  and  a25579a );
 a2379a <=( a25568a  and  a25557a );
 a2380a <=( a25546a  and  a25535a );
 a2381a <=( a25524a  and  a25513a );
 a2382a <=( a25502a  and  a25491a );
 a2383a <=( a25480a  and  a25469a );
 a2384a <=( a25458a  and  a25447a );
 a2385a <=( a25436a  and  a25425a );
 a2386a <=( a25414a  and  a25403a );
 a2387a <=( a25392a  and  a25381a );
 a2388a <=( a25370a  and  a25359a );
 a2389a <=( a25348a  and  a25337a );
 a2390a <=( a25326a  and  a25315a );
 a2391a <=( a25304a  and  a25293a );
 a2392a <=( a25282a  and  a25271a );
 a2393a <=( a25260a  and  a25249a );
 a2394a <=( a25238a  and  a25227a );
 a2395a <=( a25216a  and  a25205a );
 a2396a <=( a25194a  and  a25183a );
 a2397a <=( a25172a  and  a25161a );
 a2398a <=( a25150a  and  a25139a );
 a2399a <=( a25128a  and  a25117a );
 a2400a <=( a25106a  and  a25095a );
 a2401a <=( a25084a  and  a25073a );
 a2402a <=( a25062a  and  a25051a );
 a2403a <=( a25040a  and  a25029a );
 a2404a <=( a25018a  and  a25007a );
 a2405a <=( a24996a  and  a24985a );
 a2406a <=( a24974a  and  a24963a );
 a2407a <=( a24952a  and  a24941a );
 a2408a <=( a24930a  and  a24919a );
 a2409a <=( a24908a  and  a24897a );
 a2410a <=( a24886a  and  a24875a );
 a2411a <=( a24864a  and  a24853a );
 a2412a <=( a24842a  and  a24831a );
 a2413a <=( a24820a  and  a24809a );
 a2414a <=( a24798a  and  a24787a );
 a2415a <=( a24776a  and  a24765a );
 a2416a <=( a24754a  and  a24743a );
 a2417a <=( a24732a  and  a24721a );
 a2418a <=( a24710a  and  a24699a );
 a2419a <=( a24688a  and  a24677a );
 a2420a <=( a24666a  and  a24655a );
 a2421a <=( a24644a  and  a24633a );
 a2422a <=( a24622a  and  a24611a );
 a2423a <=( a24600a  and  a24589a );
 a2424a <=( a24578a  and  a24567a );
 a2425a <=( a24556a  and  a24545a );
 a2426a <=( a24534a  and  a24523a );
 a2427a <=( a24512a  and  a24501a );
 a2428a <=( a24490a  and  a24479a );
 a2429a <=( a24468a  and  a24457a );
 a2430a <=( a24446a  and  a24435a );
 a2431a <=( a24424a  and  a24413a );
 a2432a <=( a24402a  and  a24391a );
 a2433a <=( a24380a  and  a24369a );
 a2434a <=( a24358a  and  a24347a );
 a2435a <=( a24336a  and  a24325a );
 a2436a <=( a24314a  and  a24303a );
 a2437a <=( a24292a  and  a24281a );
 a2438a <=( a24270a  and  a24259a );
 a2439a <=( a24248a  and  a24237a );
 a2440a <=( a24226a  and  a24215a );
 a2441a <=( a24204a  and  a24193a );
 a2442a <=( a24182a  and  a24171a );
 a2443a <=( a24160a  and  a24149a );
 a2444a <=( a24138a  and  a24127a );
 a2445a <=( a24116a  and  a24105a );
 a2446a <=( a24094a  and  a24083a );
 a2447a <=( a24072a  and  a24061a );
 a2448a <=( a24050a  and  a24039a );
 a2449a <=( a24028a  and  a24017a );
 a2450a <=( a24006a  and  a23995a );
 a2451a <=( a23984a  and  a23973a );
 a2452a <=( a23962a  and  a23951a );
 a2453a <=( a23940a  and  a23929a );
 a2454a <=( a23918a  and  a23907a );
 a2455a <=( a23896a  and  a23885a );
 a2456a <=( a23874a  and  a23863a );
 a2457a <=( a23852a  and  a23841a );
 a2458a <=( a23830a  and  a23819a );
 a2459a <=( a23808a  and  a23797a );
 a2460a <=( a23786a  and  a23775a );
 a2461a <=( a23764a  and  a23753a );
 a2462a <=( a23742a  and  a23731a );
 a2463a <=( a23720a  and  a23709a );
 a2464a <=( a23698a  and  a23687a );
 a2465a <=( a23676a  and  a23665a );
 a2466a <=( a23654a  and  a23643a );
 a2467a <=( a23632a  and  a23621a );
 a2468a <=( a23610a  and  a23599a );
 a2469a <=( a23588a  and  a23577a );
 a2470a <=( a23566a  and  a23555a );
 a2471a <=( a23544a  and  a23533a );
 a2472a <=( a23522a  and  a23511a );
 a2473a <=( a23500a  and  a23489a );
 a2474a <=( a23478a  and  a23467a );
 a2475a <=( a23456a  and  a23445a );
 a2476a <=( a23434a  and  a23423a );
 a2477a <=( a23412a  and  a23401a );
 a2478a <=( a23390a  and  a23379a );
 a2479a <=( a23368a  and  a23357a );
 a2480a <=( a23346a  and  a23335a );
 a2481a <=( a23324a  and  a23313a );
 a2482a <=( a23302a  and  a23291a );
 a2483a <=( a23280a  and  a23269a );
 a2484a <=( a23258a  and  a23247a );
 a2485a <=( a23236a  and  a23225a );
 a2486a <=( a23214a  and  a23203a );
 a2487a <=( a23192a  and  a23181a );
 a2488a <=( a23170a  and  a23159a );
 a2489a <=( a23148a  and  a23137a );
 a2490a <=( a23126a  and  a23115a );
 a2491a <=( a23104a  and  a23093a );
 a2492a <=( a23082a  and  a23071a );
 a2493a <=( a23060a  and  a23049a );
 a2494a <=( a23038a  and  a23027a );
 a2495a <=( a23016a  and  a23005a );
 a2496a <=( a22994a  and  a22983a );
 a2497a <=( a22972a  and  a22961a );
 a2498a <=( a22950a  and  a22939a );
 a2499a <=( a22928a  and  a22917a );
 a2500a <=( a22906a  and  a22895a );
 a2501a <=( a22884a  and  a22873a );
 a2502a <=( a22862a  and  a22851a );
 a2503a <=( a22840a  and  a22829a );
 a2504a <=( a22818a  and  a22807a );
 a2505a <=( a22796a  and  a22785a );
 a2506a <=( a22774a  and  a22763a );
 a2507a <=( a22752a  and  a22741a );
 a2508a <=( a22730a  and  a22719a );
 a2509a <=( a22708a  and  a22697a );
 a2510a <=( a22686a  and  a22675a );
 a2511a <=( a22664a  and  a22653a );
 a2512a <=( a22642a  and  a22631a );
 a2513a <=( a22620a  and  a22609a );
 a2514a <=( a22598a  and  a22587a );
 a2515a <=( a22576a  and  a22565a );
 a2516a <=( a22554a  and  a22543a );
 a2517a <=( a22532a  and  a22521a );
 a2518a <=( a22510a  and  a22499a );
 a2519a <=( a22488a  and  a22477a );
 a2520a <=( a22466a  and  a22455a );
 a2521a <=( a22444a  and  a22433a );
 a2522a <=( a22422a  and  a22411a );
 a2523a <=( a22400a  and  a22389a );
 a2524a <=( a22378a  and  a22367a );
 a2525a <=( a22356a  and  a22345a );
 a2526a <=( a22334a  and  a22323a );
 a2527a <=( a22312a  and  a22301a );
 a2528a <=( a22290a  and  a22279a );
 a2529a <=( a22268a  and  a22257a );
 a2530a <=( a22246a  and  a22235a );
 a2531a <=( a22224a  and  a22213a );
 a2532a <=( a22202a  and  a22191a );
 a2533a <=( a22180a  and  a22169a );
 a2534a <=( a22158a  and  a22147a );
 a2535a <=( a22136a  and  a22125a );
 a2536a <=( a22114a  and  a22103a );
 a2537a <=( a22092a  and  a22081a );
 a2538a <=( a22070a  and  a22059a );
 a2539a <=( a22048a  and  a22037a );
 a2540a <=( a22026a  and  a22015a );
 a2541a <=( a22004a  and  a21993a );
 a2542a <=( a21982a  and  a21971a );
 a2543a <=( a21960a  and  a21949a );
 a2544a <=( a21938a  and  a21927a );
 a2545a <=( a21916a  and  a21905a );
 a2546a <=( a21894a  and  a21883a );
 a2547a <=( a21872a  and  a21861a );
 a2548a <=( a21850a  and  a21839a );
 a2549a <=( a21828a  and  a21817a );
 a2550a <=( a21806a  and  a21795a );
 a2551a <=( a21784a  and  a21773a );
 a2552a <=( a21762a  and  a21751a );
 a2553a <=( a21740a  and  a21729a );
 a2554a <=( a21718a  and  a21707a );
 a2555a <=( a21696a  and  a21685a );
 a2556a <=( a21674a  and  a21663a );
 a2557a <=( a21652a  and  a21641a );
 a2558a <=( a21630a  and  a21619a );
 a2559a <=( a21608a  and  a21597a );
 a2560a <=( a21586a  and  a21575a );
 a2561a <=( a21564a  and  a21553a );
 a2562a <=( a21542a  and  a21531a );
 a2563a <=( a21520a  and  a21509a );
 a2564a <=( a21498a  and  a21487a );
 a2565a <=( a21476a  and  a21465a );
 a2566a <=( a21454a  and  a21443a );
 a2567a <=( a21432a  and  a21421a );
 a2568a <=( a21410a  and  a21399a );
 a2569a <=( a21388a  and  a21377a );
 a2570a <=( a21366a  and  a21355a );
 a2571a <=( a21344a  and  a21333a );
 a2572a <=( a21322a  and  a21311a );
 a2573a <=( a21300a  and  a21289a );
 a2574a <=( a21278a  and  a21267a );
 a2575a <=( a21256a  and  a21245a );
 a2576a <=( a21234a  and  a21223a );
 a2577a <=( a21212a  and  a21201a );
 a2578a <=( a21190a  and  a21179a );
 a2579a <=( a21168a  and  a21157a );
 a2580a <=( a21146a  and  a21135a );
 a2581a <=( a21124a  and  a21113a );
 a2582a <=( a21102a  and  a21091a );
 a2583a <=( a21080a  and  a21069a );
 a2584a <=( a21058a  and  a21047a );
 a2585a <=( a21036a  and  a21025a );
 a2586a <=( a21014a  and  a21003a );
 a2587a <=( a20992a  and  a20981a );
 a2588a <=( a20970a  and  a20959a );
 a2589a <=( a20948a  and  a20937a );
 a2590a <=( a20926a  and  a20915a );
 a2591a <=( a20904a  and  a20893a );
 a2592a <=( a20882a  and  a20871a );
 a2593a <=( a20860a  and  a20849a );
 a2594a <=( a20838a  and  a20827a );
 a2595a <=( a20816a  and  a20805a );
 a2596a <=( a20794a  and  a20783a );
 a2597a <=( a20772a  and  a20761a );
 a2598a <=( a20750a  and  a20739a );
 a2599a <=( a20728a  and  a20717a );
 a2600a <=( a20706a  and  a20695a );
 a2601a <=( a20684a  and  a20673a );
 a2602a <=( a20662a  and  a20651a );
 a2603a <=( a20640a  and  a20629a );
 a2604a <=( a20618a  and  a20607a );
 a2605a <=( a20596a  and  a20585a );
 a2606a <=( a20574a  and  a20563a );
 a2607a <=( a20552a  and  a20541a );
 a2608a <=( a20530a  and  a20519a );
 a2609a <=( a20508a  and  a20497a );
 a2610a <=( a20486a  and  a20475a );
 a2611a <=( a20464a  and  a20453a );
 a2612a <=( a20442a  and  a20431a );
 a2613a <=( a20420a  and  a20409a );
 a2614a <=( a20398a  and  a20387a );
 a2615a <=( a20376a  and  a20365a );
 a2616a <=( a20354a  and  a20343a );
 a2617a <=( a20332a  and  a20321a );
 a2618a <=( a20310a  and  a20299a );
 a2619a <=( a20288a  and  a20277a );
 a2620a <=( a20266a  and  a20255a );
 a2621a <=( a20244a  and  a20233a );
 a2622a <=( a20222a  and  a20211a );
 a2623a <=( a20200a  and  a20189a );
 a2624a <=( a20178a  and  a20167a );
 a2625a <=( a20156a  and  a20145a );
 a2626a <=( a20134a  and  a20123a );
 a2627a <=( a20112a  and  a20101a );
 a2628a <=( a20090a  and  a20079a );
 a2629a <=( a20068a  and  a20057a );
 a2630a <=( a20046a  and  a20035a );
 a2631a <=( a20024a  and  a20013a );
 a2632a <=( a20002a  and  a19991a );
 a2633a <=( a19980a  and  a19969a );
 a2634a <=( a19958a  and  a19947a );
 a2635a <=( a19936a  and  a19925a );
 a2636a <=( a19914a  and  a19903a );
 a2637a <=( a19892a  and  a19881a );
 a2638a <=( a19870a  and  a19859a );
 a2639a <=( a19848a  and  a19837a );
 a2640a <=( a19826a  and  a19815a );
 a2641a <=( a19804a  and  a19793a );
 a2642a <=( a19782a  and  a19771a );
 a2643a <=( a19760a  and  a19749a );
 a2644a <=( a19738a  and  a19727a );
 a2645a <=( a19716a  and  a19705a );
 a2646a <=( a19694a  and  a19683a );
 a2647a <=( a19672a  and  a19661a );
 a2648a <=( a19650a  and  a19639a );
 a2649a <=( a19628a  and  a19617a );
 a2650a <=( a19606a  and  a19595a );
 a2651a <=( a19584a  and  a19573a );
 a2652a <=( a19562a  and  a19551a );
 a2653a <=( a19540a  and  a19529a );
 a2654a <=( a19518a  and  a19507a );
 a2655a <=( a19496a  and  a19485a );
 a2656a <=( a19474a  and  a19463a );
 a2657a <=( a19452a  and  a19441a );
 a2658a <=( a19430a  and  a19419a );
 a2659a <=( a19408a  and  a19397a );
 a2660a <=( a19386a  and  a19375a );
 a2661a <=( a19364a  and  a19353a );
 a2662a <=( a19342a  and  a19331a );
 a2663a <=( a19320a  and  a19309a );
 a2664a <=( a19298a  and  a19287a );
 a2665a <=( a19276a  and  a19265a );
 a2666a <=( a19254a  and  a19243a );
 a2667a <=( a19232a  and  a19221a );
 a2668a <=( a19210a  and  a19199a );
 a2669a <=( a19188a  and  a19177a );
 a2670a <=( a19166a  and  a19155a );
 a2671a <=( a19144a  and  a19133a );
 a2672a <=( a19122a  and  a19111a );
 a2673a <=( a19100a  and  a19089a );
 a2674a <=( a19078a  and  a19067a );
 a2675a <=( a19056a  and  a19045a );
 a2676a <=( a19034a  and  a19023a );
 a2677a <=( a19012a  and  a19001a );
 a2678a <=( a18990a  and  a18979a );
 a2679a <=( a18968a  and  a18957a );
 a2680a <=( a18946a  and  a18935a );
 a2681a <=( a18924a  and  a18913a );
 a2682a <=( a18902a  and  a18891a );
 a2683a <=( a18880a  and  a18869a );
 a2684a <=( a18858a  and  a18847a );
 a2685a <=( a18836a  and  a18825a );
 a2686a <=( a18814a  and  a18803a );
 a2687a <=( a18792a  and  a18781a );
 a2688a <=( a18770a  and  a18759a );
 a2689a <=( a18748a  and  a18737a );
 a2690a <=( a18726a  and  a18715a );
 a2691a <=( a18704a  and  a18693a );
 a2692a <=( a18682a  and  a18671a );
 a2693a <=( a18660a  and  a18649a );
 a2694a <=( a18638a  and  a18627a );
 a2695a <=( a18616a  and  a18605a );
 a2696a <=( a18594a  and  a18583a );
 a2697a <=( a18572a  and  a18561a );
 a2698a <=( a18550a  and  a18539a );
 a2699a <=( a18528a  and  a18517a );
 a2700a <=( a18506a  and  a18495a );
 a2701a <=( a18484a  and  a18473a );
 a2702a <=( a18462a  and  a18451a );
 a2703a <=( a18440a  and  a18429a );
 a2704a <=( a18418a  and  a18407a );
 a2705a <=( a18396a  and  a18385a );
 a2706a <=( a18374a  and  a18363a );
 a2707a <=( a18352a  and  a18341a );
 a2708a <=( a18330a  and  a18319a );
 a2709a <=( a18308a  and  a18297a );
 a2710a <=( a18286a  and  a18275a );
 a2711a <=( a18264a  and  a18253a );
 a2712a <=( a18242a  and  a18231a );
 a2713a <=( a18220a  and  a18209a );
 a2714a <=( a18198a  and  a18187a );
 a2715a <=( a18176a  and  a18165a );
 a2716a <=( a18154a  and  a18143a );
 a2717a <=( a18132a  and  a18121a );
 a2718a <=( a18110a  and  a18099a );
 a2719a <=( a18088a  and  a18077a );
 a2720a <=( a18066a  and  a18055a );
 a2721a <=( a18044a  and  a18033a );
 a2722a <=( a18022a  and  a18011a );
 a2723a <=( a18000a  and  a17989a );
 a2724a <=( a17978a  and  a17967a );
 a2725a <=( a17956a  and  a17945a );
 a2726a <=( a17934a  and  a17923a );
 a2727a <=( a17912a  and  a17901a );
 a2728a <=( a17890a  and  a17879a );
 a2729a <=( a17868a  and  a17857a );
 a2730a <=( a17846a  and  a17835a );
 a2731a <=( a17824a  and  a17813a );
 a2732a <=( a17802a  and  a17791a );
 a2733a <=( a17780a  and  a17769a );
 a2734a <=( a17758a  and  a17747a );
 a2735a <=( a17736a  and  a17725a );
 a2736a <=( a17714a  and  a17703a );
 a2737a <=( a17692a  and  a17681a );
 a2738a <=( a17670a  and  a17659a );
 a2739a <=( a17648a  and  a17637a );
 a2740a <=( a17626a  and  a17615a );
 a2741a <=( a17604a  and  a17593a );
 a2742a <=( a17582a  and  a17571a );
 a2743a <=( a17560a  and  a17549a );
 a2744a <=( a17538a  and  a17527a );
 a2745a <=( a17516a  and  a17505a );
 a2746a <=( a17494a  and  a17483a );
 a2747a <=( a17472a  and  a17461a );
 a2748a <=( a17450a  and  a17439a );
 a2749a <=( a17428a  and  a17417a );
 a2750a <=( a17408a  and  a17397a );
 a2751a <=( a17388a  and  a17377a );
 a2752a <=( a17368a  and  a17357a );
 a2753a <=( a17348a  and  a17337a );
 a2754a <=( a17328a  and  a17317a );
 a2755a <=( a17308a  and  a17297a );
 a2756a <=( a17288a  and  a17277a );
 a2757a <=( a17268a  and  a17257a );
 a2758a <=( a17248a  and  a17237a );
 a2759a <=( a17228a  and  a17217a );
 a2760a <=( a17208a  and  a17197a );
 a2761a <=( a17188a  and  a17177a );
 a2762a <=( a17168a  and  a17157a );
 a2763a <=( a17148a  and  a17137a );
 a2764a <=( a17128a  and  a17117a );
 a2765a <=( a17108a  and  a17097a );
 a2766a <=( a17088a  and  a17077a );
 a2767a <=( a17068a  and  a17057a );
 a2768a <=( a17048a  and  a17037a );
 a2769a <=( a17028a  and  a17017a );
 a2770a <=( a17008a  and  a16997a );
 a2771a <=( a16988a  and  a16977a );
 a2772a <=( a16968a  and  a16957a );
 a2773a <=( a16948a  and  a16937a );
 a2774a <=( a16928a  and  a16917a );
 a2775a <=( a16908a  and  a16897a );
 a2776a <=( a16888a  and  a16877a );
 a2777a <=( a16868a  and  a16857a );
 a2778a <=( a16848a  and  a16837a );
 a2779a <=( a16828a  and  a16817a );
 a2780a <=( a16808a  and  a16797a );
 a2781a <=( a16788a  and  a16777a );
 a2782a <=( a16768a  and  a16757a );
 a2783a <=( a16748a  and  a16737a );
 a2784a <=( a16728a  and  a16717a );
 a2785a <=( a16708a  and  a16697a );
 a2786a <=( a16688a  and  a16677a );
 a2787a <=( a16668a  and  a16657a );
 a2788a <=( a16648a  and  a16637a );
 a2789a <=( a16628a  and  a16617a );
 a2790a <=( a16608a  and  a16597a );
 a2791a <=( a16588a  and  a16577a );
 a2792a <=( a16568a  and  a16557a );
 a2793a <=( a16548a  and  a16537a );
 a2794a <=( a16528a  and  a16517a );
 a2795a <=( a16508a  and  a16497a );
 a2796a <=( a16488a  and  a16477a );
 a2797a <=( a16468a  and  a16457a );
 a2798a <=( a16448a  and  a16437a );
 a2799a <=( a16428a  and  a16417a );
 a2800a <=( a16408a  and  a16397a );
 a2801a <=( a16388a  and  a16377a );
 a2802a <=( a16368a  and  a16357a );
 a2803a <=( a16348a  and  a16337a );
 a2804a <=( a16328a  and  a16317a );
 a2805a <=( a16308a  and  a16297a );
 a2806a <=( a16288a  and  a16277a );
 a2807a <=( a16268a  and  a16257a );
 a2808a <=( a16248a  and  a16237a );
 a2809a <=( a16228a  and  a16217a );
 a2810a <=( a16208a  and  a16197a );
 a2811a <=( a16188a  and  a16177a );
 a2812a <=( a16168a  and  a16157a );
 a2813a <=( a16148a  and  a16137a );
 a2814a <=( a16128a  and  a16117a );
 a2815a <=( a16108a  and  a16097a );
 a2816a <=( a16088a  and  a16077a );
 a2817a <=( a16068a  and  a16057a );
 a2818a <=( a16048a  and  a16037a );
 a2819a <=( a16028a  and  a16017a );
 a2820a <=( a16008a  and  a15997a );
 a2821a <=( a15988a  and  a15977a );
 a2822a <=( a15968a  and  a15957a );
 a2823a <=( a15948a  and  a15937a );
 a2824a <=( a15928a  and  a15917a );
 a2825a <=( a15908a  and  a15897a );
 a2826a <=( a15888a  and  a15877a );
 a2827a <=( a15868a  and  a15857a );
 a2828a <=( a15848a  and  a15837a );
 a2829a <=( a15828a  and  a15817a );
 a2830a <=( a15808a  and  a15797a );
 a2831a <=( a15788a  and  a15777a );
 a2832a <=( a15768a  and  a15757a );
 a2833a <=( a15748a  and  a15737a );
 a2834a <=( a15728a  and  a15717a );
 a2835a <=( a15708a  and  a15697a );
 a2836a <=( a15688a  and  a15677a );
 a2837a <=( a15668a  and  a15657a );
 a2838a <=( a15648a  and  a15637a );
 a2839a <=( a15628a  and  a15617a );
 a2840a <=( a15608a  and  a15597a );
 a2841a <=( a15588a  and  a15577a );
 a2842a <=( a15568a  and  a15557a );
 a2843a <=( a15548a  and  a15537a );
 a2844a <=( a15528a  and  a15517a );
 a2845a <=( a15508a  and  a15497a );
 a2846a <=( a15488a  and  a15477a );
 a2847a <=( a15468a  and  a15457a );
 a2848a <=( a15448a  and  a15437a );
 a2849a <=( a15428a  and  a15417a );
 a2850a <=( a15408a  and  a15397a );
 a2851a <=( a15388a  and  a15377a );
 a2852a <=( a15368a  and  a15357a );
 a2853a <=( a15348a  and  a15337a );
 a2854a <=( a15328a  and  a15317a );
 a2855a <=( a15308a  and  a15297a );
 a2856a <=( a15288a  and  a15277a );
 a2857a <=( a15268a  and  a15257a );
 a2858a <=( a15248a  and  a15237a );
 a2859a <=( a15228a  and  a15217a );
 a2860a <=( a15208a  and  a15197a );
 a2861a <=( a15188a  and  a15177a );
 a2862a <=( a15168a  and  a15157a );
 a2863a <=( a15148a  and  a15137a );
 a2864a <=( a15128a  and  a15117a );
 a2865a <=( a15108a  and  a15097a );
 a2866a <=( a15088a  and  a15077a );
 a2867a <=( a15068a  and  a15057a );
 a2868a <=( a15048a  and  a15037a );
 a2869a <=( a15028a  and  a15017a );
 a2870a <=( a15008a  and  a14997a );
 a2871a <=( a14988a  and  a14977a );
 a2872a <=( a14968a  and  a14957a );
 a2873a <=( a14948a  and  a14937a );
 a2874a <=( a14928a  and  a14917a );
 a2875a <=( a14908a  and  a14897a );
 a2876a <=( a14888a  and  a14877a );
 a2877a <=( a14868a  and  a14857a );
 a2878a <=( a14848a  and  a14837a );
 a2879a <=( a14828a  and  a14817a );
 a2880a <=( a14808a  and  a14797a );
 a2881a <=( a14788a  and  a14777a );
 a2882a <=( a14768a  and  a14757a );
 a2883a <=( a14748a  and  a14737a );
 a2884a <=( a14728a  and  a14717a );
 a2885a <=( a14708a  and  a14697a );
 a2886a <=( a14688a  and  a14677a );
 a2887a <=( a14668a  and  a14657a );
 a2888a <=( a14648a  and  a14637a );
 a2889a <=( a14628a  and  a14617a );
 a2890a <=( a14608a  and  a14597a );
 a2891a <=( a14588a  and  a14577a );
 a2892a <=( a14568a  and  a14557a );
 a2893a <=( a14548a  and  a14537a );
 a2894a <=( a14528a  and  a14517a );
 a2895a <=( a14508a  and  a14497a );
 a2896a <=( a14488a  and  a14477a );
 a2897a <=( a14468a  and  a14457a );
 a2898a <=( a14448a  and  a14437a );
 a2899a <=( a14428a  and  a14417a );
 a2900a <=( a14408a  and  a14397a );
 a2901a <=( a14388a  and  a14377a );
 a2902a <=( a14368a  and  a14357a );
 a2903a <=( a14348a  and  a14337a );
 a2904a <=( a14328a  and  a14317a );
 a2905a <=( a14308a  and  a14297a );
 a2906a <=( a14288a  and  a14277a );
 a2907a <=( a14268a  and  a14257a );
 a2908a <=( a14248a  and  a14237a );
 a2909a <=( a14228a  and  a14217a );
 a2910a <=( a14208a  and  a14197a );
 a2911a <=( a14188a  and  a14177a );
 a2912a <=( a14168a  and  a14157a );
 a2913a <=( a14148a  and  a14137a );
 a2914a <=( a14128a  and  a14117a );
 a2915a <=( a14108a  and  a14097a );
 a2916a <=( a14088a  and  a14077a );
 a2917a <=( a14068a  and  a14057a );
 a2918a <=( a14048a  and  a14037a );
 a2919a <=( a14028a  and  a14017a );
 a2920a <=( a14008a  and  a13997a );
 a2921a <=( a13988a  and  a13977a );
 a2922a <=( a13968a  and  a13957a );
 a2923a <=( a13948a  and  a13937a );
 a2924a <=( a13928a  and  a13917a );
 a2925a <=( a13908a  and  a13897a );
 a2926a <=( a13888a  and  a13877a );
 a2927a <=( a13868a  and  a13857a );
 a2928a <=( a13848a  and  a13837a );
 a2929a <=( a13828a  and  a13817a );
 a2930a <=( a13808a  and  a13797a );
 a2931a <=( a13788a  and  a13777a );
 a2932a <=( a13768a  and  a13757a );
 a2933a <=( a13748a  and  a13737a );
 a2934a <=( a13728a  and  a13717a );
 a2935a <=( a13708a  and  a13697a );
 a2936a <=( a13688a  and  a13677a );
 a2937a <=( a13668a  and  a13657a );
 a2938a <=( a13648a  and  a13637a );
 a2939a <=( a13628a  and  a13619a );
 a2940a <=( a13610a  and  a13601a );
 a2941a <=( a13592a  and  a13583a );
 a2942a <=( a13574a  and  a13565a );
 a2943a <=( a13556a  and  a13547a );
 a2944a <=( a13538a  and  a13529a );
 a2945a <=( a13520a  and  a13511a );
 a2946a <=( a13502a  and  a13493a );
 a2947a <=( a13484a  and  a13475a );
 a2948a <=( a13466a  and  a13457a );
 a2949a <=( a13448a  and  a13439a );
 a2950a <=( a13430a  and  a13421a );
 a2951a <=( a13412a  and  a13403a );
 a2952a <=( a13394a  and  a13385a );
 a2953a <=( a13376a  and  a13367a );
 a2954a <=( a13358a  and  a13349a );
 a2955a <=( a13340a  and  a13331a );
 a2956a <=( a13322a  and  a13313a );
 a2957a <=( a13304a  and  a13295a );
 a2958a <=( a13286a  and  a13277a );
 a2959a <=( a13268a  and  a13259a );
 a2960a <=( a13250a  and  a13241a );
 a2961a <=( a13232a  and  a13223a );
 a2962a <=( a13214a  and  a13205a );
 a2963a <=( a13196a  and  a13187a );
 a2964a <=( a13178a  and  a13169a );
 a2965a <=( a13160a  and  a13151a );
 a2966a <=( a13142a  and  a13133a );
 a2967a <=( a13124a  and  a13115a );
 a2968a <=( a13106a  and  a13097a );
 a2969a <=( a13088a  and  a13079a );
 a2970a <=( a13070a  and  a13061a );
 a2971a <=( a13052a  and  a13043a );
 a2972a <=( a13034a  and  a13025a );
 a2973a <=( a13016a  and  a13007a );
 a2974a <=( a12998a  and  a12989a );
 a2975a <=( a12980a  and  a12971a );
 a2976a <=( a12962a  and  a12953a );
 a2977a <=( a12944a  and  a12935a );
 a2978a <=( a12926a  and  a12917a );
 a2979a <=( a12908a  and  a12899a );
 a2980a <=( a12890a  and  a12881a );
 a2981a <=( a12872a  and  a12863a );
 a2982a <=( a12854a  and  a12845a );
 a2983a <=( a12836a  and  a12827a );
 a2984a <=( a12818a  and  a12809a );
 a2985a <=( a12800a  and  a12791a );
 a2986a <=( a12782a  and  a12773a );
 a2987a <=( a12764a  and  a12755a );
 a2988a <=( a12746a  and  a12737a );
 a2989a <=( a12728a  and  a12719a );
 a2990a <=( a12710a  and  a12701a );
 a2991a <=( a12692a  and  a12683a );
 a2992a <=( a12674a  and  a12665a );
 a2993a <=( a12656a  and  a12647a );
 a2994a <=( a12638a  and  a12629a );
 a2995a <=( a12620a  and  a12611a );
 a2996a <=( a12602a  and  a12593a );
 a2997a <=( a12584a  and  a12575a );
 a2998a <=( a12566a  and  a12557a );
 a2999a <=( a12548a  and  a12539a );
 a3000a <=( a12530a  and  a12521a );
 a3001a <=( a12512a  and  a12503a );
 a3002a <=( a12494a  and  a12485a );
 a3003a <=( a12476a  and  a12467a );
 a3004a <=( a12458a  and  a12449a );
 a3005a <=( a12440a  and  a12431a );
 a3006a <=( a12422a  and  a12413a );
 a3007a <=( a12404a  and  a12395a );
 a3008a <=( a12386a  and  a12377a );
 a3009a <=( a12368a  and  a12359a );
 a3010a <=( a12350a  and  a12341a );
 a3011a <=( a12332a  and  a12323a );
 a3012a <=( a12314a  and  a12305a );
 a3013a <=( a12296a  and  a12287a );
 a3014a <=( a12278a  and  a12269a );
 a3015a <=( a12260a  and  a12251a );
 a3016a <=( a12242a  and  a12233a );
 a3017a <=( a12224a  and  a12215a );
 a3018a <=( a12206a  and  a12197a );
 a3019a <=( a12188a  and  a12179a );
 a3020a <=( a12170a  and  a12161a );
 a3021a <=( a12152a  and  a12143a );
 a3022a <=( a12134a  and  a12125a );
 a3023a <=( a12116a  and  a12107a );
 a3024a <=( a12098a  and  a12089a );
 a3025a <=( a12080a  and  a12071a );
 a3026a <=( a12062a  and  a12053a );
 a3027a <=( a12044a  and  a12035a );
 a3028a <=( a12026a  and  a12017a );
 a3029a <=( a12008a  and  a11999a );
 a3030a <=( a11990a  and  a11981a );
 a3031a <=( a11972a  and  a11963a );
 a3032a <=( a11954a  and  a11945a );
 a3033a <=( a11936a  and  a11927a );
 a3034a <=( a11918a  and  a11909a );
 a3035a <=( a11900a  and  a11891a );
 a3036a <=( a11882a  and  a11873a );
 a3037a <=( a11864a  and  a11855a );
 a3038a <=( a11846a  and  a11837a );
 a3039a <=( a11828a  and  a11819a );
 a3040a <=( a11810a  and  a11801a );
 a3041a <=( a11792a  and  a11783a );
 a3042a <=( a11774a  and  a11765a );
 a3043a <=( a11756a  and  a11747a );
 a3044a <=( a11738a  and  a11729a );
 a3045a <=( a11720a  and  a11711a );
 a3046a <=( a11702a  and  a11693a );
 a3047a <=( a11684a  and  a11675a );
 a3048a <=( a11666a  and  a11657a );
 a3049a <=( a11648a  and  a11639a );
 a3050a <=( a11630a  and  a11621a );
 a3051a <=( a11612a  and  a11603a );
 a3052a <=( a11594a  and  a11585a );
 a3053a <=( a11576a  and  a11567a );
 a3054a <=( a11558a  and  a11549a );
 a3055a <=( a11540a  and  a11531a );
 a3056a <=( a11522a  and  a11513a );
 a3057a <=( a11504a  and  a11495a );
 a3058a <=( a11486a  and  a11477a );
 a3059a <=( a11468a  and  a11459a );
 a3060a <=( a11450a  and  a11441a );
 a3061a <=( a11432a  and  a11423a );
 a3062a <=( a11414a  and  a11405a );
 a3063a <=( a11396a  and  a11387a );
 a3064a <=( a11378a  and  a11369a );
 a3065a <=( a11360a  and  a11351a );
 a3066a <=( a11342a  and  a11333a );
 a3067a <=( a11324a  and  a11315a );
 a3068a <=( a11306a  and  a11297a );
 a3069a <=( a11288a  and  a11279a );
 a3070a <=( a11270a  and  a11261a );
 a3071a <=( a11252a  and  a11243a );
 a3072a <=( a11234a  and  a11225a );
 a3073a <=( a11216a  and  a11207a );
 a3074a <=( a11198a  and  a11189a );
 a3075a <=( a11180a  and  a11171a );
 a3076a <=( a11162a  and  a11153a );
 a3077a <=( a11144a  and  a11135a );
 a3078a <=( a11126a  and  a11117a );
 a3079a <=( a11108a  and  a11099a );
 a3080a <=( a11090a  and  a11081a );
 a3081a <=( a11072a  and  a11063a );
 a3082a <=( a11054a  and  a11045a );
 a3083a <=( a11036a  and  a11027a );
 a3084a <=( a11018a  and  a11009a );
 a3085a <=( a11000a  and  a10991a );
 a3086a <=( a10982a  and  a10973a );
 a3087a <=( a10964a  and  a10955a );
 a3088a <=( a10946a  and  a10937a );
 a3089a <=( a10928a  and  a10919a );
 a3090a <=( a10910a  and  a10901a );
 a3091a <=( a10892a  and  a10883a );
 a3092a <=( a10874a  and  a10865a );
 a3093a <=( a10856a  and  a10847a );
 a3094a <=( a10838a  and  a10829a );
 a3095a <=( a10820a  and  a10811a );
 a3096a <=( a10802a  and  a10793a );
 a3097a <=( a10784a  and  a10775a );
 a3098a <=( a10766a  and  a10757a );
 a3099a <=( a10748a  and  a10739a );
 a3100a <=( a10730a  and  a10721a );
 a3101a <=( a10712a  and  a10703a );
 a3102a <=( a10694a  and  a10685a );
 a3103a <=( a10676a  and  a10667a );
 a3104a <=( a10658a  and  a10649a );
 a3105a <=( a10640a  and  a10631a );
 a3106a <=( a10622a  and  a10613a );
 a3107a <=( a10604a  and  a10595a );
 a3108a <=( a10586a  and  a10577a );
 a3109a <=( a10568a  and  a10559a );
 a3110a <=( a10550a  and  a10541a );
 a3111a <=( a10532a  and  a10523a );
 a3112a <=( a10514a  and  a10505a );
 a3113a <=( a10496a  and  a10487a );
 a3114a <=( a10478a  and  a10469a );
 a3115a <=( a10460a  and  a10451a );
 a3116a <=( a10442a  and  a10433a );
 a3117a <=( a10424a  and  a10415a );
 a3118a <=( a10406a  and  a10397a );
 a3119a <=( a10388a  and  a10379a );
 a3120a <=( a10370a  and  a10361a );
 a3121a <=( a10352a  and  a10343a );
 a3122a <=( a10334a  and  a10325a );
 a3123a <=( a10316a  and  a10307a );
 a3124a <=( a10298a  and  a10289a );
 a3125a <=( a10280a  and  a10271a );
 a3126a <=( a10262a  and  a10253a );
 a3127a <=( a10244a  and  a10235a );
 a3128a <=( a10226a  and  a10217a );
 a3129a <=( a10208a  and  a10199a );
 a3130a <=( a10192a  and  a10183a );
 a3131a <=( a10176a  and  a10167a );
 a3132a <=( a10160a  and  a10151a );
 a3133a <=( a10144a  and  a10135a );
 a3134a <=( a10128a  and  a10119a );
 a3135a <=( a10112a  and  a10103a );
 a3136a <=( a10096a  and  a10087a );
 a3137a <=( a10080a  and  a10071a );
 a3138a <=( a10064a  and  a10055a );
 a3139a <=( a10048a  and  a10039a );
 a3140a <=( a10032a  and  a10023a );
 a3141a <=( a10016a  and  a10007a );
 a3142a <=( a10000a  and  a9991a );
 a3143a <=( a9984a  and  a9975a );
 a3144a <=( a9968a  and  a9959a );
 a3145a <=( a9952a  and  a9943a );
 a3146a <=( a9936a  and  a9927a );
 a3147a <=( a9920a  and  a9911a );
 a3148a <=( a9904a  and  a9895a );
 a3149a <=( a9888a  and  a9879a );
 a3150a <=( a9872a  and  a9863a );
 a3151a <=( a9856a  and  a9849a );
 a3152a <=( a9842a  and  a9835a );
 a3153a <=( a9828a  and  a9821a );
 a3154a <=( a9814a  and  a9807a );
 a3155a <=( a9800a  and  a9793a );
 a3156a <=( a9786a  and  a9779a );
 a3157a <=( a9772a  and  a9765a );
 a3158a <=( a9758a  and  a9751a );
 a3159a <=( a9744a  and  a9737a );
 a3160a <=( a9730a  and  a9723a );
 a3161a <=( a9716a  and  a9709a );
 a3162a <=( a9702a  and  a9695a );
 a3163a <=( a9688a  and  a9681a );
 a3164a <=( a9674a  and  a9667a );
 a3165a <=( a9660a  and  a9653a );
 a3166a <=( a9646a  and  a9639a );
 a3167a <=( a9632a  and  a9625a );
 a3168a <=( a9618a  and  a9611a );
 a3169a <=( a9604a  and  a9597a );
 a3170a <=( a9590a  and  a9583a );
 a3171a <=( a9576a  and  a9569a );
 a3172a <=( a9562a  and  a9555a );
 a3173a <=( a9548a  and  a9541a );
 a3174a <=( a9534a  and  a9527a );
 a3178a <=( a3172a ) or ( a3173a );
 a3179a <=( a3174a ) or ( a3178a );
 a3183a <=( a3169a ) or ( a3170a );
 a3184a <=( a3171a ) or ( a3183a );
 a3185a <=( a3184a ) or ( a3179a );
 a3189a <=( a3166a ) or ( a3167a );
 a3190a <=( a3168a ) or ( a3189a );
 a3194a <=( a3163a ) or ( a3164a );
 a3195a <=( a3165a ) or ( a3194a );
 a3196a <=( a3195a ) or ( a3190a );
 a3197a <=( a3196a ) or ( a3185a );
 a3201a <=( a3160a ) or ( a3161a );
 a3202a <=( a3162a ) or ( a3201a );
 a3206a <=( a3157a ) or ( a3158a );
 a3207a <=( a3159a ) or ( a3206a );
 a3208a <=( a3207a ) or ( a3202a );
 a3212a <=( a3154a ) or ( a3155a );
 a3213a <=( a3156a ) or ( a3212a );
 a3217a <=( a3151a ) or ( a3152a );
 a3218a <=( a3153a ) or ( a3217a );
 a3219a <=( a3218a ) or ( a3213a );
 a3220a <=( a3219a ) or ( a3208a );
 a3221a <=( a3220a ) or ( a3197a );
 a3225a <=( a3148a ) or ( a3149a );
 a3226a <=( a3150a ) or ( a3225a );
 a3230a <=( a3145a ) or ( a3146a );
 a3231a <=( a3147a ) or ( a3230a );
 a3232a <=( a3231a ) or ( a3226a );
 a3236a <=( a3142a ) or ( a3143a );
 a3237a <=( a3144a ) or ( a3236a );
 a3241a <=( a3139a ) or ( a3140a );
 a3242a <=( a3141a ) or ( a3241a );
 a3243a <=( a3242a ) or ( a3237a );
 a3244a <=( a3243a ) or ( a3232a );
 a3248a <=( a3136a ) or ( a3137a );
 a3249a <=( a3138a ) or ( a3248a );
 a3253a <=( a3133a ) or ( a3134a );
 a3254a <=( a3135a ) or ( a3253a );
 a3255a <=( a3254a ) or ( a3249a );
 a3259a <=( a3130a ) or ( a3131a );
 a3260a <=( a3132a ) or ( a3259a );
 a3263a <=( a3128a ) or ( a3129a );
 a3266a <=( a3126a ) or ( a3127a );
 a3267a <=( a3266a ) or ( a3263a );
 a3268a <=( a3267a ) or ( a3260a );
 a3269a <=( a3268a ) or ( a3255a );
 a3270a <=( a3269a ) or ( a3244a );
 a3271a <=( a3270a ) or ( a3221a );
 a3275a <=( a3123a ) or ( a3124a );
 a3276a <=( a3125a ) or ( a3275a );
 a3280a <=( a3120a ) or ( a3121a );
 a3281a <=( a3122a ) or ( a3280a );
 a3282a <=( a3281a ) or ( a3276a );
 a3286a <=( a3117a ) or ( a3118a );
 a3287a <=( a3119a ) or ( a3286a );
 a3291a <=( a3114a ) or ( a3115a );
 a3292a <=( a3116a ) or ( a3291a );
 a3293a <=( a3292a ) or ( a3287a );
 a3294a <=( a3293a ) or ( a3282a );
 a3298a <=( a3111a ) or ( a3112a );
 a3299a <=( a3113a ) or ( a3298a );
 a3303a <=( a3108a ) or ( a3109a );
 a3304a <=( a3110a ) or ( a3303a );
 a3305a <=( a3304a ) or ( a3299a );
 a3309a <=( a3105a ) or ( a3106a );
 a3310a <=( a3107a ) or ( a3309a );
 a3313a <=( a3103a ) or ( a3104a );
 a3316a <=( a3101a ) or ( a3102a );
 a3317a <=( a3316a ) or ( a3313a );
 a3318a <=( a3317a ) or ( a3310a );
 a3319a <=( a3318a ) or ( a3305a );
 a3320a <=( a3319a ) or ( a3294a );
 a3324a <=( a3098a ) or ( a3099a );
 a3325a <=( a3100a ) or ( a3324a );
 a3329a <=( a3095a ) or ( a3096a );
 a3330a <=( a3097a ) or ( a3329a );
 a3331a <=( a3330a ) or ( a3325a );
 a3335a <=( a3092a ) or ( a3093a );
 a3336a <=( a3094a ) or ( a3335a );
 a3340a <=( a3089a ) or ( a3090a );
 a3341a <=( a3091a ) or ( a3340a );
 a3342a <=( a3341a ) or ( a3336a );
 a3343a <=( a3342a ) or ( a3331a );
 a3347a <=( a3086a ) or ( a3087a );
 a3348a <=( a3088a ) or ( a3347a );
 a3352a <=( a3083a ) or ( a3084a );
 a3353a <=( a3085a ) or ( a3352a );
 a3354a <=( a3353a ) or ( a3348a );
 a3358a <=( a3080a ) or ( a3081a );
 a3359a <=( a3082a ) or ( a3358a );
 a3362a <=( a3078a ) or ( a3079a );
 a3365a <=( a3076a ) or ( a3077a );
 a3366a <=( a3365a ) or ( a3362a );
 a3367a <=( a3366a ) or ( a3359a );
 a3368a <=( a3367a ) or ( a3354a );
 a3369a <=( a3368a ) or ( a3343a );
 a3370a <=( a3369a ) or ( a3320a );
 a3371a <=( a3370a ) or ( a3271a );
 a3375a <=( a3073a ) or ( a3074a );
 a3376a <=( a3075a ) or ( a3375a );
 a3380a <=( a3070a ) or ( a3071a );
 a3381a <=( a3072a ) or ( a3380a );
 a3382a <=( a3381a ) or ( a3376a );
 a3386a <=( a3067a ) or ( a3068a );
 a3387a <=( a3069a ) or ( a3386a );
 a3391a <=( a3064a ) or ( a3065a );
 a3392a <=( a3066a ) or ( a3391a );
 a3393a <=( a3392a ) or ( a3387a );
 a3394a <=( a3393a ) or ( a3382a );
 a3398a <=( a3061a ) or ( a3062a );
 a3399a <=( a3063a ) or ( a3398a );
 a3403a <=( a3058a ) or ( a3059a );
 a3404a <=( a3060a ) or ( a3403a );
 a3405a <=( a3404a ) or ( a3399a );
 a3409a <=( a3055a ) or ( a3056a );
 a3410a <=( a3057a ) or ( a3409a );
 a3414a <=( a3052a ) or ( a3053a );
 a3415a <=( a3054a ) or ( a3414a );
 a3416a <=( a3415a ) or ( a3410a );
 a3417a <=( a3416a ) or ( a3405a );
 a3418a <=( a3417a ) or ( a3394a );
 a3422a <=( a3049a ) or ( a3050a );
 a3423a <=( a3051a ) or ( a3422a );
 a3427a <=( a3046a ) or ( a3047a );
 a3428a <=( a3048a ) or ( a3427a );
 a3429a <=( a3428a ) or ( a3423a );
 a3433a <=( a3043a ) or ( a3044a );
 a3434a <=( a3045a ) or ( a3433a );
 a3438a <=( a3040a ) or ( a3041a );
 a3439a <=( a3042a ) or ( a3438a );
 a3440a <=( a3439a ) or ( a3434a );
 a3441a <=( a3440a ) or ( a3429a );
 a3445a <=( a3037a ) or ( a3038a );
 a3446a <=( a3039a ) or ( a3445a );
 a3450a <=( a3034a ) or ( a3035a );
 a3451a <=( a3036a ) or ( a3450a );
 a3452a <=( a3451a ) or ( a3446a );
 a3456a <=( a3031a ) or ( a3032a );
 a3457a <=( a3033a ) or ( a3456a );
 a3460a <=( a3029a ) or ( a3030a );
 a3463a <=( a3027a ) or ( a3028a );
 a3464a <=( a3463a ) or ( a3460a );
 a3465a <=( a3464a ) or ( a3457a );
 a3466a <=( a3465a ) or ( a3452a );
 a3467a <=( a3466a ) or ( a3441a );
 a3468a <=( a3467a ) or ( a3418a );
 a3472a <=( a3024a ) or ( a3025a );
 a3473a <=( a3026a ) or ( a3472a );
 a3477a <=( a3021a ) or ( a3022a );
 a3478a <=( a3023a ) or ( a3477a );
 a3479a <=( a3478a ) or ( a3473a );
 a3483a <=( a3018a ) or ( a3019a );
 a3484a <=( a3020a ) or ( a3483a );
 a3488a <=( a3015a ) or ( a3016a );
 a3489a <=( a3017a ) or ( a3488a );
 a3490a <=( a3489a ) or ( a3484a );
 a3491a <=( a3490a ) or ( a3479a );
 a3495a <=( a3012a ) or ( a3013a );
 a3496a <=( a3014a ) or ( a3495a );
 a3500a <=( a3009a ) or ( a3010a );
 a3501a <=( a3011a ) or ( a3500a );
 a3502a <=( a3501a ) or ( a3496a );
 a3506a <=( a3006a ) or ( a3007a );
 a3507a <=( a3008a ) or ( a3506a );
 a3510a <=( a3004a ) or ( a3005a );
 a3513a <=( a3002a ) or ( a3003a );
 a3514a <=( a3513a ) or ( a3510a );
 a3515a <=( a3514a ) or ( a3507a );
 a3516a <=( a3515a ) or ( a3502a );
 a3517a <=( a3516a ) or ( a3491a );
 a3521a <=( a2999a ) or ( a3000a );
 a3522a <=( a3001a ) or ( a3521a );
 a3526a <=( a2996a ) or ( a2997a );
 a3527a <=( a2998a ) or ( a3526a );
 a3528a <=( a3527a ) or ( a3522a );
 a3532a <=( a2993a ) or ( a2994a );
 a3533a <=( a2995a ) or ( a3532a );
 a3537a <=( a2990a ) or ( a2991a );
 a3538a <=( a2992a ) or ( a3537a );
 a3539a <=( a3538a ) or ( a3533a );
 a3540a <=( a3539a ) or ( a3528a );
 a3544a <=( a2987a ) or ( a2988a );
 a3545a <=( a2989a ) or ( a3544a );
 a3549a <=( a2984a ) or ( a2985a );
 a3550a <=( a2986a ) or ( a3549a );
 a3551a <=( a3550a ) or ( a3545a );
 a3555a <=( a2981a ) or ( a2982a );
 a3556a <=( a2983a ) or ( a3555a );
 a3559a <=( a2979a ) or ( a2980a );
 a3562a <=( a2977a ) or ( a2978a );
 a3563a <=( a3562a ) or ( a3559a );
 a3564a <=( a3563a ) or ( a3556a );
 a3565a <=( a3564a ) or ( a3551a );
 a3566a <=( a3565a ) or ( a3540a );
 a3567a <=( a3566a ) or ( a3517a );
 a3568a <=( a3567a ) or ( a3468a );
 a3569a <=( a3568a ) or ( a3371a );
 a3573a <=( a2974a ) or ( a2975a );
 a3574a <=( a2976a ) or ( a3573a );
 a3578a <=( a2971a ) or ( a2972a );
 a3579a <=( a2973a ) or ( a3578a );
 a3580a <=( a3579a ) or ( a3574a );
 a3584a <=( a2968a ) or ( a2969a );
 a3585a <=( a2970a ) or ( a3584a );
 a3589a <=( a2965a ) or ( a2966a );
 a3590a <=( a2967a ) or ( a3589a );
 a3591a <=( a3590a ) or ( a3585a );
 a3592a <=( a3591a ) or ( a3580a );
 a3596a <=( a2962a ) or ( a2963a );
 a3597a <=( a2964a ) or ( a3596a );
 a3601a <=( a2959a ) or ( a2960a );
 a3602a <=( a2961a ) or ( a3601a );
 a3603a <=( a3602a ) or ( a3597a );
 a3607a <=( a2956a ) or ( a2957a );
 a3608a <=( a2958a ) or ( a3607a );
 a3612a <=( a2953a ) or ( a2954a );
 a3613a <=( a2955a ) or ( a3612a );
 a3614a <=( a3613a ) or ( a3608a );
 a3615a <=( a3614a ) or ( a3603a );
 a3616a <=( a3615a ) or ( a3592a );
 a3620a <=( a2950a ) or ( a2951a );
 a3621a <=( a2952a ) or ( a3620a );
 a3625a <=( a2947a ) or ( a2948a );
 a3626a <=( a2949a ) or ( a3625a );
 a3627a <=( a3626a ) or ( a3621a );
 a3631a <=( a2944a ) or ( a2945a );
 a3632a <=( a2946a ) or ( a3631a );
 a3636a <=( a2941a ) or ( a2942a );
 a3637a <=( a2943a ) or ( a3636a );
 a3638a <=( a3637a ) or ( a3632a );
 a3639a <=( a3638a ) or ( a3627a );
 a3643a <=( a2938a ) or ( a2939a );
 a3644a <=( a2940a ) or ( a3643a );
 a3648a <=( a2935a ) or ( a2936a );
 a3649a <=( a2937a ) or ( a3648a );
 a3650a <=( a3649a ) or ( a3644a );
 a3654a <=( a2932a ) or ( a2933a );
 a3655a <=( a2934a ) or ( a3654a );
 a3658a <=( a2930a ) or ( a2931a );
 a3661a <=( a2928a ) or ( a2929a );
 a3662a <=( a3661a ) or ( a3658a );
 a3663a <=( a3662a ) or ( a3655a );
 a3664a <=( a3663a ) or ( a3650a );
 a3665a <=( a3664a ) or ( a3639a );
 a3666a <=( a3665a ) or ( a3616a );
 a3670a <=( a2925a ) or ( a2926a );
 a3671a <=( a2927a ) or ( a3670a );
 a3675a <=( a2922a ) or ( a2923a );
 a3676a <=( a2924a ) or ( a3675a );
 a3677a <=( a3676a ) or ( a3671a );
 a3681a <=( a2919a ) or ( a2920a );
 a3682a <=( a2921a ) or ( a3681a );
 a3686a <=( a2916a ) or ( a2917a );
 a3687a <=( a2918a ) or ( a3686a );
 a3688a <=( a3687a ) or ( a3682a );
 a3689a <=( a3688a ) or ( a3677a );
 a3693a <=( a2913a ) or ( a2914a );
 a3694a <=( a2915a ) or ( a3693a );
 a3698a <=( a2910a ) or ( a2911a );
 a3699a <=( a2912a ) or ( a3698a );
 a3700a <=( a3699a ) or ( a3694a );
 a3704a <=( a2907a ) or ( a2908a );
 a3705a <=( a2909a ) or ( a3704a );
 a3708a <=( a2905a ) or ( a2906a );
 a3711a <=( a2903a ) or ( a2904a );
 a3712a <=( a3711a ) or ( a3708a );
 a3713a <=( a3712a ) or ( a3705a );
 a3714a <=( a3713a ) or ( a3700a );
 a3715a <=( a3714a ) or ( a3689a );
 a3719a <=( a2900a ) or ( a2901a );
 a3720a <=( a2902a ) or ( a3719a );
 a3724a <=( a2897a ) or ( a2898a );
 a3725a <=( a2899a ) or ( a3724a );
 a3726a <=( a3725a ) or ( a3720a );
 a3730a <=( a2894a ) or ( a2895a );
 a3731a <=( a2896a ) or ( a3730a );
 a3735a <=( a2891a ) or ( a2892a );
 a3736a <=( a2893a ) or ( a3735a );
 a3737a <=( a3736a ) or ( a3731a );
 a3738a <=( a3737a ) or ( a3726a );
 a3742a <=( a2888a ) or ( a2889a );
 a3743a <=( a2890a ) or ( a3742a );
 a3747a <=( a2885a ) or ( a2886a );
 a3748a <=( a2887a ) or ( a3747a );
 a3749a <=( a3748a ) or ( a3743a );
 a3753a <=( a2882a ) or ( a2883a );
 a3754a <=( a2884a ) or ( a3753a );
 a3757a <=( a2880a ) or ( a2881a );
 a3760a <=( a2878a ) or ( a2879a );
 a3761a <=( a3760a ) or ( a3757a );
 a3762a <=( a3761a ) or ( a3754a );
 a3763a <=( a3762a ) or ( a3749a );
 a3764a <=( a3763a ) or ( a3738a );
 a3765a <=( a3764a ) or ( a3715a );
 a3766a <=( a3765a ) or ( a3666a );
 a3770a <=( a2875a ) or ( a2876a );
 a3771a <=( a2877a ) or ( a3770a );
 a3775a <=( a2872a ) or ( a2873a );
 a3776a <=( a2874a ) or ( a3775a );
 a3777a <=( a3776a ) or ( a3771a );
 a3781a <=( a2869a ) or ( a2870a );
 a3782a <=( a2871a ) or ( a3781a );
 a3786a <=( a2866a ) or ( a2867a );
 a3787a <=( a2868a ) or ( a3786a );
 a3788a <=( a3787a ) or ( a3782a );
 a3789a <=( a3788a ) or ( a3777a );
 a3793a <=( a2863a ) or ( a2864a );
 a3794a <=( a2865a ) or ( a3793a );
 a3798a <=( a2860a ) or ( a2861a );
 a3799a <=( a2862a ) or ( a3798a );
 a3800a <=( a3799a ) or ( a3794a );
 a3804a <=( a2857a ) or ( a2858a );
 a3805a <=( a2859a ) or ( a3804a );
 a3809a <=( a2854a ) or ( a2855a );
 a3810a <=( a2856a ) or ( a3809a );
 a3811a <=( a3810a ) or ( a3805a );
 a3812a <=( a3811a ) or ( a3800a );
 a3813a <=( a3812a ) or ( a3789a );
 a3817a <=( a2851a ) or ( a2852a );
 a3818a <=( a2853a ) or ( a3817a );
 a3822a <=( a2848a ) or ( a2849a );
 a3823a <=( a2850a ) or ( a3822a );
 a3824a <=( a3823a ) or ( a3818a );
 a3828a <=( a2845a ) or ( a2846a );
 a3829a <=( a2847a ) or ( a3828a );
 a3833a <=( a2842a ) or ( a2843a );
 a3834a <=( a2844a ) or ( a3833a );
 a3835a <=( a3834a ) or ( a3829a );
 a3836a <=( a3835a ) or ( a3824a );
 a3840a <=( a2839a ) or ( a2840a );
 a3841a <=( a2841a ) or ( a3840a );
 a3845a <=( a2836a ) or ( a2837a );
 a3846a <=( a2838a ) or ( a3845a );
 a3847a <=( a3846a ) or ( a3841a );
 a3851a <=( a2833a ) or ( a2834a );
 a3852a <=( a2835a ) or ( a3851a );
 a3855a <=( a2831a ) or ( a2832a );
 a3858a <=( a2829a ) or ( a2830a );
 a3859a <=( a3858a ) or ( a3855a );
 a3860a <=( a3859a ) or ( a3852a );
 a3861a <=( a3860a ) or ( a3847a );
 a3862a <=( a3861a ) or ( a3836a );
 a3863a <=( a3862a ) or ( a3813a );
 a3867a <=( a2826a ) or ( a2827a );
 a3868a <=( a2828a ) or ( a3867a );
 a3872a <=( a2823a ) or ( a2824a );
 a3873a <=( a2825a ) or ( a3872a );
 a3874a <=( a3873a ) or ( a3868a );
 a3878a <=( a2820a ) or ( a2821a );
 a3879a <=( a2822a ) or ( a3878a );
 a3883a <=( a2817a ) or ( a2818a );
 a3884a <=( a2819a ) or ( a3883a );
 a3885a <=( a3884a ) or ( a3879a );
 a3886a <=( a3885a ) or ( a3874a );
 a3890a <=( a2814a ) or ( a2815a );
 a3891a <=( a2816a ) or ( a3890a );
 a3895a <=( a2811a ) or ( a2812a );
 a3896a <=( a2813a ) or ( a3895a );
 a3897a <=( a3896a ) or ( a3891a );
 a3901a <=( a2808a ) or ( a2809a );
 a3902a <=( a2810a ) or ( a3901a );
 a3905a <=( a2806a ) or ( a2807a );
 a3908a <=( a2804a ) or ( a2805a );
 a3909a <=( a3908a ) or ( a3905a );
 a3910a <=( a3909a ) or ( a3902a );
 a3911a <=( a3910a ) or ( a3897a );
 a3912a <=( a3911a ) or ( a3886a );
 a3916a <=( a2801a ) or ( a2802a );
 a3917a <=( a2803a ) or ( a3916a );
 a3921a <=( a2798a ) or ( a2799a );
 a3922a <=( a2800a ) or ( a3921a );
 a3923a <=( a3922a ) or ( a3917a );
 a3927a <=( a2795a ) or ( a2796a );
 a3928a <=( a2797a ) or ( a3927a );
 a3932a <=( a2792a ) or ( a2793a );
 a3933a <=( a2794a ) or ( a3932a );
 a3934a <=( a3933a ) or ( a3928a );
 a3935a <=( a3934a ) or ( a3923a );
 a3939a <=( a2789a ) or ( a2790a );
 a3940a <=( a2791a ) or ( a3939a );
 a3944a <=( a2786a ) or ( a2787a );
 a3945a <=( a2788a ) or ( a3944a );
 a3946a <=( a3945a ) or ( a3940a );
 a3950a <=( a2783a ) or ( a2784a );
 a3951a <=( a2785a ) or ( a3950a );
 a3954a <=( a2781a ) or ( a2782a );
 a3957a <=( a2779a ) or ( a2780a );
 a3958a <=( a3957a ) or ( a3954a );
 a3959a <=( a3958a ) or ( a3951a );
 a3960a <=( a3959a ) or ( a3946a );
 a3961a <=( a3960a ) or ( a3935a );
 a3962a <=( a3961a ) or ( a3912a );
 a3963a <=( a3962a ) or ( a3863a );
 a3964a <=( a3963a ) or ( a3766a );
 a3965a <=( a3964a ) or ( a3569a );
 a3969a <=( a2776a ) or ( a2777a );
 a3970a <=( a2778a ) or ( a3969a );
 a3974a <=( a2773a ) or ( a2774a );
 a3975a <=( a2775a ) or ( a3974a );
 a3976a <=( a3975a ) or ( a3970a );
 a3980a <=( a2770a ) or ( a2771a );
 a3981a <=( a2772a ) or ( a3980a );
 a3985a <=( a2767a ) or ( a2768a );
 a3986a <=( a2769a ) or ( a3985a );
 a3987a <=( a3986a ) or ( a3981a );
 a3988a <=( a3987a ) or ( a3976a );
 a3992a <=( a2764a ) or ( a2765a );
 a3993a <=( a2766a ) or ( a3992a );
 a3997a <=( a2761a ) or ( a2762a );
 a3998a <=( a2763a ) or ( a3997a );
 a3999a <=( a3998a ) or ( a3993a );
 a4003a <=( a2758a ) or ( a2759a );
 a4004a <=( a2760a ) or ( a4003a );
 a4008a <=( a2755a ) or ( a2756a );
 a4009a <=( a2757a ) or ( a4008a );
 a4010a <=( a4009a ) or ( a4004a );
 a4011a <=( a4010a ) or ( a3999a );
 a4012a <=( a4011a ) or ( a3988a );
 a4016a <=( a2752a ) or ( a2753a );
 a4017a <=( a2754a ) or ( a4016a );
 a4021a <=( a2749a ) or ( a2750a );
 a4022a <=( a2751a ) or ( a4021a );
 a4023a <=( a4022a ) or ( a4017a );
 a4027a <=( a2746a ) or ( a2747a );
 a4028a <=( a2748a ) or ( a4027a );
 a4032a <=( a2743a ) or ( a2744a );
 a4033a <=( a2745a ) or ( a4032a );
 a4034a <=( a4033a ) or ( a4028a );
 a4035a <=( a4034a ) or ( a4023a );
 a4039a <=( a2740a ) or ( a2741a );
 a4040a <=( a2742a ) or ( a4039a );
 a4044a <=( a2737a ) or ( a2738a );
 a4045a <=( a2739a ) or ( a4044a );
 a4046a <=( a4045a ) or ( a4040a );
 a4050a <=( a2734a ) or ( a2735a );
 a4051a <=( a2736a ) or ( a4050a );
 a4054a <=( a2732a ) or ( a2733a );
 a4057a <=( a2730a ) or ( a2731a );
 a4058a <=( a4057a ) or ( a4054a );
 a4059a <=( a4058a ) or ( a4051a );
 a4060a <=( a4059a ) or ( a4046a );
 a4061a <=( a4060a ) or ( a4035a );
 a4062a <=( a4061a ) or ( a4012a );
 a4066a <=( a2727a ) or ( a2728a );
 a4067a <=( a2729a ) or ( a4066a );
 a4071a <=( a2724a ) or ( a2725a );
 a4072a <=( a2726a ) or ( a4071a );
 a4073a <=( a4072a ) or ( a4067a );
 a4077a <=( a2721a ) or ( a2722a );
 a4078a <=( a2723a ) or ( a4077a );
 a4082a <=( a2718a ) or ( a2719a );
 a4083a <=( a2720a ) or ( a4082a );
 a4084a <=( a4083a ) or ( a4078a );
 a4085a <=( a4084a ) or ( a4073a );
 a4089a <=( a2715a ) or ( a2716a );
 a4090a <=( a2717a ) or ( a4089a );
 a4094a <=( a2712a ) or ( a2713a );
 a4095a <=( a2714a ) or ( a4094a );
 a4096a <=( a4095a ) or ( a4090a );
 a4100a <=( a2709a ) or ( a2710a );
 a4101a <=( a2711a ) or ( a4100a );
 a4104a <=( a2707a ) or ( a2708a );
 a4107a <=( a2705a ) or ( a2706a );
 a4108a <=( a4107a ) or ( a4104a );
 a4109a <=( a4108a ) or ( a4101a );
 a4110a <=( a4109a ) or ( a4096a );
 a4111a <=( a4110a ) or ( a4085a );
 a4115a <=( a2702a ) or ( a2703a );
 a4116a <=( a2704a ) or ( a4115a );
 a4120a <=( a2699a ) or ( a2700a );
 a4121a <=( a2701a ) or ( a4120a );
 a4122a <=( a4121a ) or ( a4116a );
 a4126a <=( a2696a ) or ( a2697a );
 a4127a <=( a2698a ) or ( a4126a );
 a4131a <=( a2693a ) or ( a2694a );
 a4132a <=( a2695a ) or ( a4131a );
 a4133a <=( a4132a ) or ( a4127a );
 a4134a <=( a4133a ) or ( a4122a );
 a4138a <=( a2690a ) or ( a2691a );
 a4139a <=( a2692a ) or ( a4138a );
 a4143a <=( a2687a ) or ( a2688a );
 a4144a <=( a2689a ) or ( a4143a );
 a4145a <=( a4144a ) or ( a4139a );
 a4149a <=( a2684a ) or ( a2685a );
 a4150a <=( a2686a ) or ( a4149a );
 a4153a <=( a2682a ) or ( a2683a );
 a4156a <=( a2680a ) or ( a2681a );
 a4157a <=( a4156a ) or ( a4153a );
 a4158a <=( a4157a ) or ( a4150a );
 a4159a <=( a4158a ) or ( a4145a );
 a4160a <=( a4159a ) or ( a4134a );
 a4161a <=( a4160a ) or ( a4111a );
 a4162a <=( a4161a ) or ( a4062a );
 a4166a <=( a2677a ) or ( a2678a );
 a4167a <=( a2679a ) or ( a4166a );
 a4171a <=( a2674a ) or ( a2675a );
 a4172a <=( a2676a ) or ( a4171a );
 a4173a <=( a4172a ) or ( a4167a );
 a4177a <=( a2671a ) or ( a2672a );
 a4178a <=( a2673a ) or ( a4177a );
 a4182a <=( a2668a ) or ( a2669a );
 a4183a <=( a2670a ) or ( a4182a );
 a4184a <=( a4183a ) or ( a4178a );
 a4185a <=( a4184a ) or ( a4173a );
 a4189a <=( a2665a ) or ( a2666a );
 a4190a <=( a2667a ) or ( a4189a );
 a4194a <=( a2662a ) or ( a2663a );
 a4195a <=( a2664a ) or ( a4194a );
 a4196a <=( a4195a ) or ( a4190a );
 a4200a <=( a2659a ) or ( a2660a );
 a4201a <=( a2661a ) or ( a4200a );
 a4205a <=( a2656a ) or ( a2657a );
 a4206a <=( a2658a ) or ( a4205a );
 a4207a <=( a4206a ) or ( a4201a );
 a4208a <=( a4207a ) or ( a4196a );
 a4209a <=( a4208a ) or ( a4185a );
 a4213a <=( a2653a ) or ( a2654a );
 a4214a <=( a2655a ) or ( a4213a );
 a4218a <=( a2650a ) or ( a2651a );
 a4219a <=( a2652a ) or ( a4218a );
 a4220a <=( a4219a ) or ( a4214a );
 a4224a <=( a2647a ) or ( a2648a );
 a4225a <=( a2649a ) or ( a4224a );
 a4229a <=( a2644a ) or ( a2645a );
 a4230a <=( a2646a ) or ( a4229a );
 a4231a <=( a4230a ) or ( a4225a );
 a4232a <=( a4231a ) or ( a4220a );
 a4236a <=( a2641a ) or ( a2642a );
 a4237a <=( a2643a ) or ( a4236a );
 a4241a <=( a2638a ) or ( a2639a );
 a4242a <=( a2640a ) or ( a4241a );
 a4243a <=( a4242a ) or ( a4237a );
 a4247a <=( a2635a ) or ( a2636a );
 a4248a <=( a2637a ) or ( a4247a );
 a4251a <=( a2633a ) or ( a2634a );
 a4254a <=( a2631a ) or ( a2632a );
 a4255a <=( a4254a ) or ( a4251a );
 a4256a <=( a4255a ) or ( a4248a );
 a4257a <=( a4256a ) or ( a4243a );
 a4258a <=( a4257a ) or ( a4232a );
 a4259a <=( a4258a ) or ( a4209a );
 a4263a <=( a2628a ) or ( a2629a );
 a4264a <=( a2630a ) or ( a4263a );
 a4268a <=( a2625a ) or ( a2626a );
 a4269a <=( a2627a ) or ( a4268a );
 a4270a <=( a4269a ) or ( a4264a );
 a4274a <=( a2622a ) or ( a2623a );
 a4275a <=( a2624a ) or ( a4274a );
 a4279a <=( a2619a ) or ( a2620a );
 a4280a <=( a2621a ) or ( a4279a );
 a4281a <=( a4280a ) or ( a4275a );
 a4282a <=( a4281a ) or ( a4270a );
 a4286a <=( a2616a ) or ( a2617a );
 a4287a <=( a2618a ) or ( a4286a );
 a4291a <=( a2613a ) or ( a2614a );
 a4292a <=( a2615a ) or ( a4291a );
 a4293a <=( a4292a ) or ( a4287a );
 a4297a <=( a2610a ) or ( a2611a );
 a4298a <=( a2612a ) or ( a4297a );
 a4301a <=( a2608a ) or ( a2609a );
 a4304a <=( a2606a ) or ( a2607a );
 a4305a <=( a4304a ) or ( a4301a );
 a4306a <=( a4305a ) or ( a4298a );
 a4307a <=( a4306a ) or ( a4293a );
 a4308a <=( a4307a ) or ( a4282a );
 a4312a <=( a2603a ) or ( a2604a );
 a4313a <=( a2605a ) or ( a4312a );
 a4317a <=( a2600a ) or ( a2601a );
 a4318a <=( a2602a ) or ( a4317a );
 a4319a <=( a4318a ) or ( a4313a );
 a4323a <=( a2597a ) or ( a2598a );
 a4324a <=( a2599a ) or ( a4323a );
 a4328a <=( a2594a ) or ( a2595a );
 a4329a <=( a2596a ) or ( a4328a );
 a4330a <=( a4329a ) or ( a4324a );
 a4331a <=( a4330a ) or ( a4319a );
 a4335a <=( a2591a ) or ( a2592a );
 a4336a <=( a2593a ) or ( a4335a );
 a4340a <=( a2588a ) or ( a2589a );
 a4341a <=( a2590a ) or ( a4340a );
 a4342a <=( a4341a ) or ( a4336a );
 a4346a <=( a2585a ) or ( a2586a );
 a4347a <=( a2587a ) or ( a4346a );
 a4350a <=( a2583a ) or ( a2584a );
 a4353a <=( a2581a ) or ( a2582a );
 a4354a <=( a4353a ) or ( a4350a );
 a4355a <=( a4354a ) or ( a4347a );
 a4356a <=( a4355a ) or ( a4342a );
 a4357a <=( a4356a ) or ( a4331a );
 a4358a <=( a4357a ) or ( a4308a );
 a4359a <=( a4358a ) or ( a4259a );
 a4360a <=( a4359a ) or ( a4162a );
 a4364a <=( a2578a ) or ( a2579a );
 a4365a <=( a2580a ) or ( a4364a );
 a4369a <=( a2575a ) or ( a2576a );
 a4370a <=( a2577a ) or ( a4369a );
 a4371a <=( a4370a ) or ( a4365a );
 a4375a <=( a2572a ) or ( a2573a );
 a4376a <=( a2574a ) or ( a4375a );
 a4380a <=( a2569a ) or ( a2570a );
 a4381a <=( a2571a ) or ( a4380a );
 a4382a <=( a4381a ) or ( a4376a );
 a4383a <=( a4382a ) or ( a4371a );
 a4387a <=( a2566a ) or ( a2567a );
 a4388a <=( a2568a ) or ( a4387a );
 a4392a <=( a2563a ) or ( a2564a );
 a4393a <=( a2565a ) or ( a4392a );
 a4394a <=( a4393a ) or ( a4388a );
 a4398a <=( a2560a ) or ( a2561a );
 a4399a <=( a2562a ) or ( a4398a );
 a4403a <=( a2557a ) or ( a2558a );
 a4404a <=( a2559a ) or ( a4403a );
 a4405a <=( a4404a ) or ( a4399a );
 a4406a <=( a4405a ) or ( a4394a );
 a4407a <=( a4406a ) or ( a4383a );
 a4411a <=( a2554a ) or ( a2555a );
 a4412a <=( a2556a ) or ( a4411a );
 a4416a <=( a2551a ) or ( a2552a );
 a4417a <=( a2553a ) or ( a4416a );
 a4418a <=( a4417a ) or ( a4412a );
 a4422a <=( a2548a ) or ( a2549a );
 a4423a <=( a2550a ) or ( a4422a );
 a4427a <=( a2545a ) or ( a2546a );
 a4428a <=( a2547a ) or ( a4427a );
 a4429a <=( a4428a ) or ( a4423a );
 a4430a <=( a4429a ) or ( a4418a );
 a4434a <=( a2542a ) or ( a2543a );
 a4435a <=( a2544a ) or ( a4434a );
 a4439a <=( a2539a ) or ( a2540a );
 a4440a <=( a2541a ) or ( a4439a );
 a4441a <=( a4440a ) or ( a4435a );
 a4445a <=( a2536a ) or ( a2537a );
 a4446a <=( a2538a ) or ( a4445a );
 a4449a <=( a2534a ) or ( a2535a );
 a4452a <=( a2532a ) or ( a2533a );
 a4453a <=( a4452a ) or ( a4449a );
 a4454a <=( a4453a ) or ( a4446a );
 a4455a <=( a4454a ) or ( a4441a );
 a4456a <=( a4455a ) or ( a4430a );
 a4457a <=( a4456a ) or ( a4407a );
 a4461a <=( a2529a ) or ( a2530a );
 a4462a <=( a2531a ) or ( a4461a );
 a4466a <=( a2526a ) or ( a2527a );
 a4467a <=( a2528a ) or ( a4466a );
 a4468a <=( a4467a ) or ( a4462a );
 a4472a <=( a2523a ) or ( a2524a );
 a4473a <=( a2525a ) or ( a4472a );
 a4477a <=( a2520a ) or ( a2521a );
 a4478a <=( a2522a ) or ( a4477a );
 a4479a <=( a4478a ) or ( a4473a );
 a4480a <=( a4479a ) or ( a4468a );
 a4484a <=( a2517a ) or ( a2518a );
 a4485a <=( a2519a ) or ( a4484a );
 a4489a <=( a2514a ) or ( a2515a );
 a4490a <=( a2516a ) or ( a4489a );
 a4491a <=( a4490a ) or ( a4485a );
 a4495a <=( a2511a ) or ( a2512a );
 a4496a <=( a2513a ) or ( a4495a );
 a4499a <=( a2509a ) or ( a2510a );
 a4502a <=( a2507a ) or ( a2508a );
 a4503a <=( a4502a ) or ( a4499a );
 a4504a <=( a4503a ) or ( a4496a );
 a4505a <=( a4504a ) or ( a4491a );
 a4506a <=( a4505a ) or ( a4480a );
 a4510a <=( a2504a ) or ( a2505a );
 a4511a <=( a2506a ) or ( a4510a );
 a4515a <=( a2501a ) or ( a2502a );
 a4516a <=( a2503a ) or ( a4515a );
 a4517a <=( a4516a ) or ( a4511a );
 a4521a <=( a2498a ) or ( a2499a );
 a4522a <=( a2500a ) or ( a4521a );
 a4526a <=( a2495a ) or ( a2496a );
 a4527a <=( a2497a ) or ( a4526a );
 a4528a <=( a4527a ) or ( a4522a );
 a4529a <=( a4528a ) or ( a4517a );
 a4533a <=( a2492a ) or ( a2493a );
 a4534a <=( a2494a ) or ( a4533a );
 a4538a <=( a2489a ) or ( a2490a );
 a4539a <=( a2491a ) or ( a4538a );
 a4540a <=( a4539a ) or ( a4534a );
 a4544a <=( a2486a ) or ( a2487a );
 a4545a <=( a2488a ) or ( a4544a );
 a4548a <=( a2484a ) or ( a2485a );
 a4551a <=( a2482a ) or ( a2483a );
 a4552a <=( a4551a ) or ( a4548a );
 a4553a <=( a4552a ) or ( a4545a );
 a4554a <=( a4553a ) or ( a4540a );
 a4555a <=( a4554a ) or ( a4529a );
 a4556a <=( a4555a ) or ( a4506a );
 a4557a <=( a4556a ) or ( a4457a );
 a4561a <=( a2479a ) or ( a2480a );
 a4562a <=( a2481a ) or ( a4561a );
 a4566a <=( a2476a ) or ( a2477a );
 a4567a <=( a2478a ) or ( a4566a );
 a4568a <=( a4567a ) or ( a4562a );
 a4572a <=( a2473a ) or ( a2474a );
 a4573a <=( a2475a ) or ( a4572a );
 a4577a <=( a2470a ) or ( a2471a );
 a4578a <=( a2472a ) or ( a4577a );
 a4579a <=( a4578a ) or ( a4573a );
 a4580a <=( a4579a ) or ( a4568a );
 a4584a <=( a2467a ) or ( a2468a );
 a4585a <=( a2469a ) or ( a4584a );
 a4589a <=( a2464a ) or ( a2465a );
 a4590a <=( a2466a ) or ( a4589a );
 a4591a <=( a4590a ) or ( a4585a );
 a4595a <=( a2461a ) or ( a2462a );
 a4596a <=( a2463a ) or ( a4595a );
 a4599a <=( a2459a ) or ( a2460a );
 a4602a <=( a2457a ) or ( a2458a );
 a4603a <=( a4602a ) or ( a4599a );
 a4604a <=( a4603a ) or ( a4596a );
 a4605a <=( a4604a ) or ( a4591a );
 a4606a <=( a4605a ) or ( a4580a );
 a4610a <=( a2454a ) or ( a2455a );
 a4611a <=( a2456a ) or ( a4610a );
 a4615a <=( a2451a ) or ( a2452a );
 a4616a <=( a2453a ) or ( a4615a );
 a4617a <=( a4616a ) or ( a4611a );
 a4621a <=( a2448a ) or ( a2449a );
 a4622a <=( a2450a ) or ( a4621a );
 a4626a <=( a2445a ) or ( a2446a );
 a4627a <=( a2447a ) or ( a4626a );
 a4628a <=( a4627a ) or ( a4622a );
 a4629a <=( a4628a ) or ( a4617a );
 a4633a <=( a2442a ) or ( a2443a );
 a4634a <=( a2444a ) or ( a4633a );
 a4638a <=( a2439a ) or ( a2440a );
 a4639a <=( a2441a ) or ( a4638a );
 a4640a <=( a4639a ) or ( a4634a );
 a4644a <=( a2436a ) or ( a2437a );
 a4645a <=( a2438a ) or ( a4644a );
 a4648a <=( a2434a ) or ( a2435a );
 a4651a <=( a2432a ) or ( a2433a );
 a4652a <=( a4651a ) or ( a4648a );
 a4653a <=( a4652a ) or ( a4645a );
 a4654a <=( a4653a ) or ( a4640a );
 a4655a <=( a4654a ) or ( a4629a );
 a4656a <=( a4655a ) or ( a4606a );
 a4660a <=( a2429a ) or ( a2430a );
 a4661a <=( a2431a ) or ( a4660a );
 a4665a <=( a2426a ) or ( a2427a );
 a4666a <=( a2428a ) or ( a4665a );
 a4667a <=( a4666a ) or ( a4661a );
 a4671a <=( a2423a ) or ( a2424a );
 a4672a <=( a2425a ) or ( a4671a );
 a4676a <=( a2420a ) or ( a2421a );
 a4677a <=( a2422a ) or ( a4676a );
 a4678a <=( a4677a ) or ( a4672a );
 a4679a <=( a4678a ) or ( a4667a );
 a4683a <=( a2417a ) or ( a2418a );
 a4684a <=( a2419a ) or ( a4683a );
 a4688a <=( a2414a ) or ( a2415a );
 a4689a <=( a2416a ) or ( a4688a );
 a4690a <=( a4689a ) or ( a4684a );
 a4694a <=( a2411a ) or ( a2412a );
 a4695a <=( a2413a ) or ( a4694a );
 a4698a <=( a2409a ) or ( a2410a );
 a4701a <=( a2407a ) or ( a2408a );
 a4702a <=( a4701a ) or ( a4698a );
 a4703a <=( a4702a ) or ( a4695a );
 a4704a <=( a4703a ) or ( a4690a );
 a4705a <=( a4704a ) or ( a4679a );
 a4709a <=( a2404a ) or ( a2405a );
 a4710a <=( a2406a ) or ( a4709a );
 a4714a <=( a2401a ) or ( a2402a );
 a4715a <=( a2403a ) or ( a4714a );
 a4716a <=( a4715a ) or ( a4710a );
 a4720a <=( a2398a ) or ( a2399a );
 a4721a <=( a2400a ) or ( a4720a );
 a4725a <=( a2395a ) or ( a2396a );
 a4726a <=( a2397a ) or ( a4725a );
 a4727a <=( a4726a ) or ( a4721a );
 a4728a <=( a4727a ) or ( a4716a );
 a4732a <=( a2392a ) or ( a2393a );
 a4733a <=( a2394a ) or ( a4732a );
 a4737a <=( a2389a ) or ( a2390a );
 a4738a <=( a2391a ) or ( a4737a );
 a4739a <=( a4738a ) or ( a4733a );
 a4743a <=( a2386a ) or ( a2387a );
 a4744a <=( a2388a ) or ( a4743a );
 a4747a <=( a2384a ) or ( a2385a );
 a4750a <=( a2382a ) or ( a2383a );
 a4751a <=( a4750a ) or ( a4747a );
 a4752a <=( a4751a ) or ( a4744a );
 a4753a <=( a4752a ) or ( a4739a );
 a4754a <=( a4753a ) or ( a4728a );
 a4755a <=( a4754a ) or ( a4705a );
 a4756a <=( a4755a ) or ( a4656a );
 a4757a <=( a4756a ) or ( a4557a );
 a4758a <=( a4757a ) or ( a4360a );
 a4759a <=( a4758a ) or ( a3965a );
 a4763a <=( a2379a ) or ( a2380a );
 a4764a <=( a2381a ) or ( a4763a );
 a4768a <=( a2376a ) or ( a2377a );
 a4769a <=( a2378a ) or ( a4768a );
 a4770a <=( a4769a ) or ( a4764a );
 a4774a <=( a2373a ) or ( a2374a );
 a4775a <=( a2375a ) or ( a4774a );
 a4779a <=( a2370a ) or ( a2371a );
 a4780a <=( a2372a ) or ( a4779a );
 a4781a <=( a4780a ) or ( a4775a );
 a4782a <=( a4781a ) or ( a4770a );
 a4786a <=( a2367a ) or ( a2368a );
 a4787a <=( a2369a ) or ( a4786a );
 a4791a <=( a2364a ) or ( a2365a );
 a4792a <=( a2366a ) or ( a4791a );
 a4793a <=( a4792a ) or ( a4787a );
 a4797a <=( a2361a ) or ( a2362a );
 a4798a <=( a2363a ) or ( a4797a );
 a4802a <=( a2358a ) or ( a2359a );
 a4803a <=( a2360a ) or ( a4802a );
 a4804a <=( a4803a ) or ( a4798a );
 a4805a <=( a4804a ) or ( a4793a );
 a4806a <=( a4805a ) or ( a4782a );
 a4810a <=( a2355a ) or ( a2356a );
 a4811a <=( a2357a ) or ( a4810a );
 a4815a <=( a2352a ) or ( a2353a );
 a4816a <=( a2354a ) or ( a4815a );
 a4817a <=( a4816a ) or ( a4811a );
 a4821a <=( a2349a ) or ( a2350a );
 a4822a <=( a2351a ) or ( a4821a );
 a4826a <=( a2346a ) or ( a2347a );
 a4827a <=( a2348a ) or ( a4826a );
 a4828a <=( a4827a ) or ( a4822a );
 a4829a <=( a4828a ) or ( a4817a );
 a4833a <=( a2343a ) or ( a2344a );
 a4834a <=( a2345a ) or ( a4833a );
 a4838a <=( a2340a ) or ( a2341a );
 a4839a <=( a2342a ) or ( a4838a );
 a4840a <=( a4839a ) or ( a4834a );
 a4844a <=( a2337a ) or ( a2338a );
 a4845a <=( a2339a ) or ( a4844a );
 a4848a <=( a2335a ) or ( a2336a );
 a4851a <=( a2333a ) or ( a2334a );
 a4852a <=( a4851a ) or ( a4848a );
 a4853a <=( a4852a ) or ( a4845a );
 a4854a <=( a4853a ) or ( a4840a );
 a4855a <=( a4854a ) or ( a4829a );
 a4856a <=( a4855a ) or ( a4806a );
 a4860a <=( a2330a ) or ( a2331a );
 a4861a <=( a2332a ) or ( a4860a );
 a4865a <=( a2327a ) or ( a2328a );
 a4866a <=( a2329a ) or ( a4865a );
 a4867a <=( a4866a ) or ( a4861a );
 a4871a <=( a2324a ) or ( a2325a );
 a4872a <=( a2326a ) or ( a4871a );
 a4876a <=( a2321a ) or ( a2322a );
 a4877a <=( a2323a ) or ( a4876a );
 a4878a <=( a4877a ) or ( a4872a );
 a4879a <=( a4878a ) or ( a4867a );
 a4883a <=( a2318a ) or ( a2319a );
 a4884a <=( a2320a ) or ( a4883a );
 a4888a <=( a2315a ) or ( a2316a );
 a4889a <=( a2317a ) or ( a4888a );
 a4890a <=( a4889a ) or ( a4884a );
 a4894a <=( a2312a ) or ( a2313a );
 a4895a <=( a2314a ) or ( a4894a );
 a4898a <=( a2310a ) or ( a2311a );
 a4901a <=( a2308a ) or ( a2309a );
 a4902a <=( a4901a ) or ( a4898a );
 a4903a <=( a4902a ) or ( a4895a );
 a4904a <=( a4903a ) or ( a4890a );
 a4905a <=( a4904a ) or ( a4879a );
 a4909a <=( a2305a ) or ( a2306a );
 a4910a <=( a2307a ) or ( a4909a );
 a4914a <=( a2302a ) or ( a2303a );
 a4915a <=( a2304a ) or ( a4914a );
 a4916a <=( a4915a ) or ( a4910a );
 a4920a <=( a2299a ) or ( a2300a );
 a4921a <=( a2301a ) or ( a4920a );
 a4925a <=( a2296a ) or ( a2297a );
 a4926a <=( a2298a ) or ( a4925a );
 a4927a <=( a4926a ) or ( a4921a );
 a4928a <=( a4927a ) or ( a4916a );
 a4932a <=( a2293a ) or ( a2294a );
 a4933a <=( a2295a ) or ( a4932a );
 a4937a <=( a2290a ) or ( a2291a );
 a4938a <=( a2292a ) or ( a4937a );
 a4939a <=( a4938a ) or ( a4933a );
 a4943a <=( a2287a ) or ( a2288a );
 a4944a <=( a2289a ) or ( a4943a );
 a4947a <=( a2285a ) or ( a2286a );
 a4950a <=( a2283a ) or ( a2284a );
 a4951a <=( a4950a ) or ( a4947a );
 a4952a <=( a4951a ) or ( a4944a );
 a4953a <=( a4952a ) or ( a4939a );
 a4954a <=( a4953a ) or ( a4928a );
 a4955a <=( a4954a ) or ( a4905a );
 a4956a <=( a4955a ) or ( a4856a );
 a4960a <=( a2280a ) or ( a2281a );
 a4961a <=( a2282a ) or ( a4960a );
 a4965a <=( a2277a ) or ( a2278a );
 a4966a <=( a2279a ) or ( a4965a );
 a4967a <=( a4966a ) or ( a4961a );
 a4971a <=( a2274a ) or ( a2275a );
 a4972a <=( a2276a ) or ( a4971a );
 a4976a <=( a2271a ) or ( a2272a );
 a4977a <=( a2273a ) or ( a4976a );
 a4978a <=( a4977a ) or ( a4972a );
 a4979a <=( a4978a ) or ( a4967a );
 a4983a <=( a2268a ) or ( a2269a );
 a4984a <=( a2270a ) or ( a4983a );
 a4988a <=( a2265a ) or ( a2266a );
 a4989a <=( a2267a ) or ( a4988a );
 a4990a <=( a4989a ) or ( a4984a );
 a4994a <=( a2262a ) or ( a2263a );
 a4995a <=( a2264a ) or ( a4994a );
 a4999a <=( a2259a ) or ( a2260a );
 a5000a <=( a2261a ) or ( a4999a );
 a5001a <=( a5000a ) or ( a4995a );
 a5002a <=( a5001a ) or ( a4990a );
 a5003a <=( a5002a ) or ( a4979a );
 a5007a <=( a2256a ) or ( a2257a );
 a5008a <=( a2258a ) or ( a5007a );
 a5012a <=( a2253a ) or ( a2254a );
 a5013a <=( a2255a ) or ( a5012a );
 a5014a <=( a5013a ) or ( a5008a );
 a5018a <=( a2250a ) or ( a2251a );
 a5019a <=( a2252a ) or ( a5018a );
 a5023a <=( a2247a ) or ( a2248a );
 a5024a <=( a2249a ) or ( a5023a );
 a5025a <=( a5024a ) or ( a5019a );
 a5026a <=( a5025a ) or ( a5014a );
 a5030a <=( a2244a ) or ( a2245a );
 a5031a <=( a2246a ) or ( a5030a );
 a5035a <=( a2241a ) or ( a2242a );
 a5036a <=( a2243a ) or ( a5035a );
 a5037a <=( a5036a ) or ( a5031a );
 a5041a <=( a2238a ) or ( a2239a );
 a5042a <=( a2240a ) or ( a5041a );
 a5045a <=( a2236a ) or ( a2237a );
 a5048a <=( a2234a ) or ( a2235a );
 a5049a <=( a5048a ) or ( a5045a );
 a5050a <=( a5049a ) or ( a5042a );
 a5051a <=( a5050a ) or ( a5037a );
 a5052a <=( a5051a ) or ( a5026a );
 a5053a <=( a5052a ) or ( a5003a );
 a5057a <=( a2231a ) or ( a2232a );
 a5058a <=( a2233a ) or ( a5057a );
 a5062a <=( a2228a ) or ( a2229a );
 a5063a <=( a2230a ) or ( a5062a );
 a5064a <=( a5063a ) or ( a5058a );
 a5068a <=( a2225a ) or ( a2226a );
 a5069a <=( a2227a ) or ( a5068a );
 a5073a <=( a2222a ) or ( a2223a );
 a5074a <=( a2224a ) or ( a5073a );
 a5075a <=( a5074a ) or ( a5069a );
 a5076a <=( a5075a ) or ( a5064a );
 a5080a <=( a2219a ) or ( a2220a );
 a5081a <=( a2221a ) or ( a5080a );
 a5085a <=( a2216a ) or ( a2217a );
 a5086a <=( a2218a ) or ( a5085a );
 a5087a <=( a5086a ) or ( a5081a );
 a5091a <=( a2213a ) or ( a2214a );
 a5092a <=( a2215a ) or ( a5091a );
 a5095a <=( a2211a ) or ( a2212a );
 a5098a <=( a2209a ) or ( a2210a );
 a5099a <=( a5098a ) or ( a5095a );
 a5100a <=( a5099a ) or ( a5092a );
 a5101a <=( a5100a ) or ( a5087a );
 a5102a <=( a5101a ) or ( a5076a );
 a5106a <=( a2206a ) or ( a2207a );
 a5107a <=( a2208a ) or ( a5106a );
 a5111a <=( a2203a ) or ( a2204a );
 a5112a <=( a2205a ) or ( a5111a );
 a5113a <=( a5112a ) or ( a5107a );
 a5117a <=( a2200a ) or ( a2201a );
 a5118a <=( a2202a ) or ( a5117a );
 a5122a <=( a2197a ) or ( a2198a );
 a5123a <=( a2199a ) or ( a5122a );
 a5124a <=( a5123a ) or ( a5118a );
 a5125a <=( a5124a ) or ( a5113a );
 a5129a <=( a2194a ) or ( a2195a );
 a5130a <=( a2196a ) or ( a5129a );
 a5134a <=( a2191a ) or ( a2192a );
 a5135a <=( a2193a ) or ( a5134a );
 a5136a <=( a5135a ) or ( a5130a );
 a5140a <=( a2188a ) or ( a2189a );
 a5141a <=( a2190a ) or ( a5140a );
 a5144a <=( a2186a ) or ( a2187a );
 a5147a <=( a2184a ) or ( a2185a );
 a5148a <=( a5147a ) or ( a5144a );
 a5149a <=( a5148a ) or ( a5141a );
 a5150a <=( a5149a ) or ( a5136a );
 a5151a <=( a5150a ) or ( a5125a );
 a5152a <=( a5151a ) or ( a5102a );
 a5153a <=( a5152a ) or ( a5053a );
 a5154a <=( a5153a ) or ( a4956a );
 a5158a <=( a2181a ) or ( a2182a );
 a5159a <=( a2183a ) or ( a5158a );
 a5163a <=( a2178a ) or ( a2179a );
 a5164a <=( a2180a ) or ( a5163a );
 a5165a <=( a5164a ) or ( a5159a );
 a5169a <=( a2175a ) or ( a2176a );
 a5170a <=( a2177a ) or ( a5169a );
 a5174a <=( a2172a ) or ( a2173a );
 a5175a <=( a2174a ) or ( a5174a );
 a5176a <=( a5175a ) or ( a5170a );
 a5177a <=( a5176a ) or ( a5165a );
 a5181a <=( a2169a ) or ( a2170a );
 a5182a <=( a2171a ) or ( a5181a );
 a5186a <=( a2166a ) or ( a2167a );
 a5187a <=( a2168a ) or ( a5186a );
 a5188a <=( a5187a ) or ( a5182a );
 a5192a <=( a2163a ) or ( a2164a );
 a5193a <=( a2165a ) or ( a5192a );
 a5197a <=( a2160a ) or ( a2161a );
 a5198a <=( a2162a ) or ( a5197a );
 a5199a <=( a5198a ) or ( a5193a );
 a5200a <=( a5199a ) or ( a5188a );
 a5201a <=( a5200a ) or ( a5177a );
 a5205a <=( a2157a ) or ( a2158a );
 a5206a <=( a2159a ) or ( a5205a );
 a5210a <=( a2154a ) or ( a2155a );
 a5211a <=( a2156a ) or ( a5210a );
 a5212a <=( a5211a ) or ( a5206a );
 a5216a <=( a2151a ) or ( a2152a );
 a5217a <=( a2153a ) or ( a5216a );
 a5221a <=( a2148a ) or ( a2149a );
 a5222a <=( a2150a ) or ( a5221a );
 a5223a <=( a5222a ) or ( a5217a );
 a5224a <=( a5223a ) or ( a5212a );
 a5228a <=( a2145a ) or ( a2146a );
 a5229a <=( a2147a ) or ( a5228a );
 a5233a <=( a2142a ) or ( a2143a );
 a5234a <=( a2144a ) or ( a5233a );
 a5235a <=( a5234a ) or ( a5229a );
 a5239a <=( a2139a ) or ( a2140a );
 a5240a <=( a2141a ) or ( a5239a );
 a5243a <=( a2137a ) or ( a2138a );
 a5246a <=( a2135a ) or ( a2136a );
 a5247a <=( a5246a ) or ( a5243a );
 a5248a <=( a5247a ) or ( a5240a );
 a5249a <=( a5248a ) or ( a5235a );
 a5250a <=( a5249a ) or ( a5224a );
 a5251a <=( a5250a ) or ( a5201a );
 a5255a <=( a2132a ) or ( a2133a );
 a5256a <=( a2134a ) or ( a5255a );
 a5260a <=( a2129a ) or ( a2130a );
 a5261a <=( a2131a ) or ( a5260a );
 a5262a <=( a5261a ) or ( a5256a );
 a5266a <=( a2126a ) or ( a2127a );
 a5267a <=( a2128a ) or ( a5266a );
 a5271a <=( a2123a ) or ( a2124a );
 a5272a <=( a2125a ) or ( a5271a );
 a5273a <=( a5272a ) or ( a5267a );
 a5274a <=( a5273a ) or ( a5262a );
 a5278a <=( a2120a ) or ( a2121a );
 a5279a <=( a2122a ) or ( a5278a );
 a5283a <=( a2117a ) or ( a2118a );
 a5284a <=( a2119a ) or ( a5283a );
 a5285a <=( a5284a ) or ( a5279a );
 a5289a <=( a2114a ) or ( a2115a );
 a5290a <=( a2116a ) or ( a5289a );
 a5293a <=( a2112a ) or ( a2113a );
 a5296a <=( a2110a ) or ( a2111a );
 a5297a <=( a5296a ) or ( a5293a );
 a5298a <=( a5297a ) or ( a5290a );
 a5299a <=( a5298a ) or ( a5285a );
 a5300a <=( a5299a ) or ( a5274a );
 a5304a <=( a2107a ) or ( a2108a );
 a5305a <=( a2109a ) or ( a5304a );
 a5309a <=( a2104a ) or ( a2105a );
 a5310a <=( a2106a ) or ( a5309a );
 a5311a <=( a5310a ) or ( a5305a );
 a5315a <=( a2101a ) or ( a2102a );
 a5316a <=( a2103a ) or ( a5315a );
 a5320a <=( a2098a ) or ( a2099a );
 a5321a <=( a2100a ) or ( a5320a );
 a5322a <=( a5321a ) or ( a5316a );
 a5323a <=( a5322a ) or ( a5311a );
 a5327a <=( a2095a ) or ( a2096a );
 a5328a <=( a2097a ) or ( a5327a );
 a5332a <=( a2092a ) or ( a2093a );
 a5333a <=( a2094a ) or ( a5332a );
 a5334a <=( a5333a ) or ( a5328a );
 a5338a <=( a2089a ) or ( a2090a );
 a5339a <=( a2091a ) or ( a5338a );
 a5342a <=( a2087a ) or ( a2088a );
 a5345a <=( a2085a ) or ( a2086a );
 a5346a <=( a5345a ) or ( a5342a );
 a5347a <=( a5346a ) or ( a5339a );
 a5348a <=( a5347a ) or ( a5334a );
 a5349a <=( a5348a ) or ( a5323a );
 a5350a <=( a5349a ) or ( a5300a );
 a5351a <=( a5350a ) or ( a5251a );
 a5355a <=( a2082a ) or ( a2083a );
 a5356a <=( a2084a ) or ( a5355a );
 a5360a <=( a2079a ) or ( a2080a );
 a5361a <=( a2081a ) or ( a5360a );
 a5362a <=( a5361a ) or ( a5356a );
 a5366a <=( a2076a ) or ( a2077a );
 a5367a <=( a2078a ) or ( a5366a );
 a5371a <=( a2073a ) or ( a2074a );
 a5372a <=( a2075a ) or ( a5371a );
 a5373a <=( a5372a ) or ( a5367a );
 a5374a <=( a5373a ) or ( a5362a );
 a5378a <=( a2070a ) or ( a2071a );
 a5379a <=( a2072a ) or ( a5378a );
 a5383a <=( a2067a ) or ( a2068a );
 a5384a <=( a2069a ) or ( a5383a );
 a5385a <=( a5384a ) or ( a5379a );
 a5389a <=( a2064a ) or ( a2065a );
 a5390a <=( a2066a ) or ( a5389a );
 a5393a <=( a2062a ) or ( a2063a );
 a5396a <=( a2060a ) or ( a2061a );
 a5397a <=( a5396a ) or ( a5393a );
 a5398a <=( a5397a ) or ( a5390a );
 a5399a <=( a5398a ) or ( a5385a );
 a5400a <=( a5399a ) or ( a5374a );
 a5404a <=( a2057a ) or ( a2058a );
 a5405a <=( a2059a ) or ( a5404a );
 a5409a <=( a2054a ) or ( a2055a );
 a5410a <=( a2056a ) or ( a5409a );
 a5411a <=( a5410a ) or ( a5405a );
 a5415a <=( a2051a ) or ( a2052a );
 a5416a <=( a2053a ) or ( a5415a );
 a5420a <=( a2048a ) or ( a2049a );
 a5421a <=( a2050a ) or ( a5420a );
 a5422a <=( a5421a ) or ( a5416a );
 a5423a <=( a5422a ) or ( a5411a );
 a5427a <=( a2045a ) or ( a2046a );
 a5428a <=( a2047a ) or ( a5427a );
 a5432a <=( a2042a ) or ( a2043a );
 a5433a <=( a2044a ) or ( a5432a );
 a5434a <=( a5433a ) or ( a5428a );
 a5438a <=( a2039a ) or ( a2040a );
 a5439a <=( a2041a ) or ( a5438a );
 a5442a <=( a2037a ) or ( a2038a );
 a5445a <=( a2035a ) or ( a2036a );
 a5446a <=( a5445a ) or ( a5442a );
 a5447a <=( a5446a ) or ( a5439a );
 a5448a <=( a5447a ) or ( a5434a );
 a5449a <=( a5448a ) or ( a5423a );
 a5450a <=( a5449a ) or ( a5400a );
 a5454a <=( a2032a ) or ( a2033a );
 a5455a <=( a2034a ) or ( a5454a );
 a5459a <=( a2029a ) or ( a2030a );
 a5460a <=( a2031a ) or ( a5459a );
 a5461a <=( a5460a ) or ( a5455a );
 a5465a <=( a2026a ) or ( a2027a );
 a5466a <=( a2028a ) or ( a5465a );
 a5470a <=( a2023a ) or ( a2024a );
 a5471a <=( a2025a ) or ( a5470a );
 a5472a <=( a5471a ) or ( a5466a );
 a5473a <=( a5472a ) or ( a5461a );
 a5477a <=( a2020a ) or ( a2021a );
 a5478a <=( a2022a ) or ( a5477a );
 a5482a <=( a2017a ) or ( a2018a );
 a5483a <=( a2019a ) or ( a5482a );
 a5484a <=( a5483a ) or ( a5478a );
 a5488a <=( a2014a ) or ( a2015a );
 a5489a <=( a2016a ) or ( a5488a );
 a5492a <=( a2012a ) or ( a2013a );
 a5495a <=( a2010a ) or ( a2011a );
 a5496a <=( a5495a ) or ( a5492a );
 a5497a <=( a5496a ) or ( a5489a );
 a5498a <=( a5497a ) or ( a5484a );
 a5499a <=( a5498a ) or ( a5473a );
 a5503a <=( a2007a ) or ( a2008a );
 a5504a <=( a2009a ) or ( a5503a );
 a5508a <=( a2004a ) or ( a2005a );
 a5509a <=( a2006a ) or ( a5508a );
 a5510a <=( a5509a ) or ( a5504a );
 a5514a <=( a2001a ) or ( a2002a );
 a5515a <=( a2003a ) or ( a5514a );
 a5519a <=( a1998a ) or ( a1999a );
 a5520a <=( a2000a ) or ( a5519a );
 a5521a <=( a5520a ) or ( a5515a );
 a5522a <=( a5521a ) or ( a5510a );
 a5526a <=( a1995a ) or ( a1996a );
 a5527a <=( a1997a ) or ( a5526a );
 a5531a <=( a1992a ) or ( a1993a );
 a5532a <=( a1994a ) or ( a5531a );
 a5533a <=( a5532a ) or ( a5527a );
 a5537a <=( a1989a ) or ( a1990a );
 a5538a <=( a1991a ) or ( a5537a );
 a5541a <=( a1987a ) or ( a1988a );
 a5544a <=( a1985a ) or ( a1986a );
 a5545a <=( a5544a ) or ( a5541a );
 a5546a <=( a5545a ) or ( a5538a );
 a5547a <=( a5546a ) or ( a5533a );
 a5548a <=( a5547a ) or ( a5522a );
 a5549a <=( a5548a ) or ( a5499a );
 a5550a <=( a5549a ) or ( a5450a );
 a5551a <=( a5550a ) or ( a5351a );
 a5552a <=( a5551a ) or ( a5154a );
 a5556a <=( a1982a ) or ( a1983a );
 a5557a <=( a1984a ) or ( a5556a );
 a5561a <=( a1979a ) or ( a1980a );
 a5562a <=( a1981a ) or ( a5561a );
 a5563a <=( a5562a ) or ( a5557a );
 a5567a <=( a1976a ) or ( a1977a );
 a5568a <=( a1978a ) or ( a5567a );
 a5572a <=( a1973a ) or ( a1974a );
 a5573a <=( a1975a ) or ( a5572a );
 a5574a <=( a5573a ) or ( a5568a );
 a5575a <=( a5574a ) or ( a5563a );
 a5579a <=( a1970a ) or ( a1971a );
 a5580a <=( a1972a ) or ( a5579a );
 a5584a <=( a1967a ) or ( a1968a );
 a5585a <=( a1969a ) or ( a5584a );
 a5586a <=( a5585a ) or ( a5580a );
 a5590a <=( a1964a ) or ( a1965a );
 a5591a <=( a1966a ) or ( a5590a );
 a5595a <=( a1961a ) or ( a1962a );
 a5596a <=( a1963a ) or ( a5595a );
 a5597a <=( a5596a ) or ( a5591a );
 a5598a <=( a5597a ) or ( a5586a );
 a5599a <=( a5598a ) or ( a5575a );
 a5603a <=( a1958a ) or ( a1959a );
 a5604a <=( a1960a ) or ( a5603a );
 a5608a <=( a1955a ) or ( a1956a );
 a5609a <=( a1957a ) or ( a5608a );
 a5610a <=( a5609a ) or ( a5604a );
 a5614a <=( a1952a ) or ( a1953a );
 a5615a <=( a1954a ) or ( a5614a );
 a5619a <=( a1949a ) or ( a1950a );
 a5620a <=( a1951a ) or ( a5619a );
 a5621a <=( a5620a ) or ( a5615a );
 a5622a <=( a5621a ) or ( a5610a );
 a5626a <=( a1946a ) or ( a1947a );
 a5627a <=( a1948a ) or ( a5626a );
 a5631a <=( a1943a ) or ( a1944a );
 a5632a <=( a1945a ) or ( a5631a );
 a5633a <=( a5632a ) or ( a5627a );
 a5637a <=( a1940a ) or ( a1941a );
 a5638a <=( a1942a ) or ( a5637a );
 a5641a <=( a1938a ) or ( a1939a );
 a5644a <=( a1936a ) or ( a1937a );
 a5645a <=( a5644a ) or ( a5641a );
 a5646a <=( a5645a ) or ( a5638a );
 a5647a <=( a5646a ) or ( a5633a );
 a5648a <=( a5647a ) or ( a5622a );
 a5649a <=( a5648a ) or ( a5599a );
 a5653a <=( a1933a ) or ( a1934a );
 a5654a <=( a1935a ) or ( a5653a );
 a5658a <=( a1930a ) or ( a1931a );
 a5659a <=( a1932a ) or ( a5658a );
 a5660a <=( a5659a ) or ( a5654a );
 a5664a <=( a1927a ) or ( a1928a );
 a5665a <=( a1929a ) or ( a5664a );
 a5669a <=( a1924a ) or ( a1925a );
 a5670a <=( a1926a ) or ( a5669a );
 a5671a <=( a5670a ) or ( a5665a );
 a5672a <=( a5671a ) or ( a5660a );
 a5676a <=( a1921a ) or ( a1922a );
 a5677a <=( a1923a ) or ( a5676a );
 a5681a <=( a1918a ) or ( a1919a );
 a5682a <=( a1920a ) or ( a5681a );
 a5683a <=( a5682a ) or ( a5677a );
 a5687a <=( a1915a ) or ( a1916a );
 a5688a <=( a1917a ) or ( a5687a );
 a5691a <=( a1913a ) or ( a1914a );
 a5694a <=( a1911a ) or ( a1912a );
 a5695a <=( a5694a ) or ( a5691a );
 a5696a <=( a5695a ) or ( a5688a );
 a5697a <=( a5696a ) or ( a5683a );
 a5698a <=( a5697a ) or ( a5672a );
 a5702a <=( a1908a ) or ( a1909a );
 a5703a <=( a1910a ) or ( a5702a );
 a5707a <=( a1905a ) or ( a1906a );
 a5708a <=( a1907a ) or ( a5707a );
 a5709a <=( a5708a ) or ( a5703a );
 a5713a <=( a1902a ) or ( a1903a );
 a5714a <=( a1904a ) or ( a5713a );
 a5718a <=( a1899a ) or ( a1900a );
 a5719a <=( a1901a ) or ( a5718a );
 a5720a <=( a5719a ) or ( a5714a );
 a5721a <=( a5720a ) or ( a5709a );
 a5725a <=( a1896a ) or ( a1897a );
 a5726a <=( a1898a ) or ( a5725a );
 a5730a <=( a1893a ) or ( a1894a );
 a5731a <=( a1895a ) or ( a5730a );
 a5732a <=( a5731a ) or ( a5726a );
 a5736a <=( a1890a ) or ( a1891a );
 a5737a <=( a1892a ) or ( a5736a );
 a5740a <=( a1888a ) or ( a1889a );
 a5743a <=( a1886a ) or ( a1887a );
 a5744a <=( a5743a ) or ( a5740a );
 a5745a <=( a5744a ) or ( a5737a );
 a5746a <=( a5745a ) or ( a5732a );
 a5747a <=( a5746a ) or ( a5721a );
 a5748a <=( a5747a ) or ( a5698a );
 a5749a <=( a5748a ) or ( a5649a );
 a5753a <=( a1883a ) or ( a1884a );
 a5754a <=( a1885a ) or ( a5753a );
 a5758a <=( a1880a ) or ( a1881a );
 a5759a <=( a1882a ) or ( a5758a );
 a5760a <=( a5759a ) or ( a5754a );
 a5764a <=( a1877a ) or ( a1878a );
 a5765a <=( a1879a ) or ( a5764a );
 a5769a <=( a1874a ) or ( a1875a );
 a5770a <=( a1876a ) or ( a5769a );
 a5771a <=( a5770a ) or ( a5765a );
 a5772a <=( a5771a ) or ( a5760a );
 a5776a <=( a1871a ) or ( a1872a );
 a5777a <=( a1873a ) or ( a5776a );
 a5781a <=( a1868a ) or ( a1869a );
 a5782a <=( a1870a ) or ( a5781a );
 a5783a <=( a5782a ) or ( a5777a );
 a5787a <=( a1865a ) or ( a1866a );
 a5788a <=( a1867a ) or ( a5787a );
 a5792a <=( a1862a ) or ( a1863a );
 a5793a <=( a1864a ) or ( a5792a );
 a5794a <=( a5793a ) or ( a5788a );
 a5795a <=( a5794a ) or ( a5783a );
 a5796a <=( a5795a ) or ( a5772a );
 a5800a <=( a1859a ) or ( a1860a );
 a5801a <=( a1861a ) or ( a5800a );
 a5805a <=( a1856a ) or ( a1857a );
 a5806a <=( a1858a ) or ( a5805a );
 a5807a <=( a5806a ) or ( a5801a );
 a5811a <=( a1853a ) or ( a1854a );
 a5812a <=( a1855a ) or ( a5811a );
 a5816a <=( a1850a ) or ( a1851a );
 a5817a <=( a1852a ) or ( a5816a );
 a5818a <=( a5817a ) or ( a5812a );
 a5819a <=( a5818a ) or ( a5807a );
 a5823a <=( a1847a ) or ( a1848a );
 a5824a <=( a1849a ) or ( a5823a );
 a5828a <=( a1844a ) or ( a1845a );
 a5829a <=( a1846a ) or ( a5828a );
 a5830a <=( a5829a ) or ( a5824a );
 a5834a <=( a1841a ) or ( a1842a );
 a5835a <=( a1843a ) or ( a5834a );
 a5838a <=( a1839a ) or ( a1840a );
 a5841a <=( a1837a ) or ( a1838a );
 a5842a <=( a5841a ) or ( a5838a );
 a5843a <=( a5842a ) or ( a5835a );
 a5844a <=( a5843a ) or ( a5830a );
 a5845a <=( a5844a ) or ( a5819a );
 a5846a <=( a5845a ) or ( a5796a );
 a5850a <=( a1834a ) or ( a1835a );
 a5851a <=( a1836a ) or ( a5850a );
 a5855a <=( a1831a ) or ( a1832a );
 a5856a <=( a1833a ) or ( a5855a );
 a5857a <=( a5856a ) or ( a5851a );
 a5861a <=( a1828a ) or ( a1829a );
 a5862a <=( a1830a ) or ( a5861a );
 a5866a <=( a1825a ) or ( a1826a );
 a5867a <=( a1827a ) or ( a5866a );
 a5868a <=( a5867a ) or ( a5862a );
 a5869a <=( a5868a ) or ( a5857a );
 a5873a <=( a1822a ) or ( a1823a );
 a5874a <=( a1824a ) or ( a5873a );
 a5878a <=( a1819a ) or ( a1820a );
 a5879a <=( a1821a ) or ( a5878a );
 a5880a <=( a5879a ) or ( a5874a );
 a5884a <=( a1816a ) or ( a1817a );
 a5885a <=( a1818a ) or ( a5884a );
 a5888a <=( a1814a ) or ( a1815a );
 a5891a <=( a1812a ) or ( a1813a );
 a5892a <=( a5891a ) or ( a5888a );
 a5893a <=( a5892a ) or ( a5885a );
 a5894a <=( a5893a ) or ( a5880a );
 a5895a <=( a5894a ) or ( a5869a );
 a5899a <=( a1809a ) or ( a1810a );
 a5900a <=( a1811a ) or ( a5899a );
 a5904a <=( a1806a ) or ( a1807a );
 a5905a <=( a1808a ) or ( a5904a );
 a5906a <=( a5905a ) or ( a5900a );
 a5910a <=( a1803a ) or ( a1804a );
 a5911a <=( a1805a ) or ( a5910a );
 a5915a <=( a1800a ) or ( a1801a );
 a5916a <=( a1802a ) or ( a5915a );
 a5917a <=( a5916a ) or ( a5911a );
 a5918a <=( a5917a ) or ( a5906a );
 a5922a <=( a1797a ) or ( a1798a );
 a5923a <=( a1799a ) or ( a5922a );
 a5927a <=( a1794a ) or ( a1795a );
 a5928a <=( a1796a ) or ( a5927a );
 a5929a <=( a5928a ) or ( a5923a );
 a5933a <=( a1791a ) or ( a1792a );
 a5934a <=( a1793a ) or ( a5933a );
 a5937a <=( a1789a ) or ( a1790a );
 a5940a <=( a1787a ) or ( a1788a );
 a5941a <=( a5940a ) or ( a5937a );
 a5942a <=( a5941a ) or ( a5934a );
 a5943a <=( a5942a ) or ( a5929a );
 a5944a <=( a5943a ) or ( a5918a );
 a5945a <=( a5944a ) or ( a5895a );
 a5946a <=( a5945a ) or ( a5846a );
 a5947a <=( a5946a ) or ( a5749a );
 a5951a <=( a1784a ) or ( a1785a );
 a5952a <=( a1786a ) or ( a5951a );
 a5956a <=( a1781a ) or ( a1782a );
 a5957a <=( a1783a ) or ( a5956a );
 a5958a <=( a5957a ) or ( a5952a );
 a5962a <=( a1778a ) or ( a1779a );
 a5963a <=( a1780a ) or ( a5962a );
 a5967a <=( a1775a ) or ( a1776a );
 a5968a <=( a1777a ) or ( a5967a );
 a5969a <=( a5968a ) or ( a5963a );
 a5970a <=( a5969a ) or ( a5958a );
 a5974a <=( a1772a ) or ( a1773a );
 a5975a <=( a1774a ) or ( a5974a );
 a5979a <=( a1769a ) or ( a1770a );
 a5980a <=( a1771a ) or ( a5979a );
 a5981a <=( a5980a ) or ( a5975a );
 a5985a <=( a1766a ) or ( a1767a );
 a5986a <=( a1768a ) or ( a5985a );
 a5990a <=( a1763a ) or ( a1764a );
 a5991a <=( a1765a ) or ( a5990a );
 a5992a <=( a5991a ) or ( a5986a );
 a5993a <=( a5992a ) or ( a5981a );
 a5994a <=( a5993a ) or ( a5970a );
 a5998a <=( a1760a ) or ( a1761a );
 a5999a <=( a1762a ) or ( a5998a );
 a6003a <=( a1757a ) or ( a1758a );
 a6004a <=( a1759a ) or ( a6003a );
 a6005a <=( a6004a ) or ( a5999a );
 a6009a <=( a1754a ) or ( a1755a );
 a6010a <=( a1756a ) or ( a6009a );
 a6014a <=( a1751a ) or ( a1752a );
 a6015a <=( a1753a ) or ( a6014a );
 a6016a <=( a6015a ) or ( a6010a );
 a6017a <=( a6016a ) or ( a6005a );
 a6021a <=( a1748a ) or ( a1749a );
 a6022a <=( a1750a ) or ( a6021a );
 a6026a <=( a1745a ) or ( a1746a );
 a6027a <=( a1747a ) or ( a6026a );
 a6028a <=( a6027a ) or ( a6022a );
 a6032a <=( a1742a ) or ( a1743a );
 a6033a <=( a1744a ) or ( a6032a );
 a6036a <=( a1740a ) or ( a1741a );
 a6039a <=( a1738a ) or ( a1739a );
 a6040a <=( a6039a ) or ( a6036a );
 a6041a <=( a6040a ) or ( a6033a );
 a6042a <=( a6041a ) or ( a6028a );
 a6043a <=( a6042a ) or ( a6017a );
 a6044a <=( a6043a ) or ( a5994a );
 a6048a <=( a1735a ) or ( a1736a );
 a6049a <=( a1737a ) or ( a6048a );
 a6053a <=( a1732a ) or ( a1733a );
 a6054a <=( a1734a ) or ( a6053a );
 a6055a <=( a6054a ) or ( a6049a );
 a6059a <=( a1729a ) or ( a1730a );
 a6060a <=( a1731a ) or ( a6059a );
 a6064a <=( a1726a ) or ( a1727a );
 a6065a <=( a1728a ) or ( a6064a );
 a6066a <=( a6065a ) or ( a6060a );
 a6067a <=( a6066a ) or ( a6055a );
 a6071a <=( a1723a ) or ( a1724a );
 a6072a <=( a1725a ) or ( a6071a );
 a6076a <=( a1720a ) or ( a1721a );
 a6077a <=( a1722a ) or ( a6076a );
 a6078a <=( a6077a ) or ( a6072a );
 a6082a <=( a1717a ) or ( a1718a );
 a6083a <=( a1719a ) or ( a6082a );
 a6086a <=( a1715a ) or ( a1716a );
 a6089a <=( a1713a ) or ( a1714a );
 a6090a <=( a6089a ) or ( a6086a );
 a6091a <=( a6090a ) or ( a6083a );
 a6092a <=( a6091a ) or ( a6078a );
 a6093a <=( a6092a ) or ( a6067a );
 a6097a <=( a1710a ) or ( a1711a );
 a6098a <=( a1712a ) or ( a6097a );
 a6102a <=( a1707a ) or ( a1708a );
 a6103a <=( a1709a ) or ( a6102a );
 a6104a <=( a6103a ) or ( a6098a );
 a6108a <=( a1704a ) or ( a1705a );
 a6109a <=( a1706a ) or ( a6108a );
 a6113a <=( a1701a ) or ( a1702a );
 a6114a <=( a1703a ) or ( a6113a );
 a6115a <=( a6114a ) or ( a6109a );
 a6116a <=( a6115a ) or ( a6104a );
 a6120a <=( a1698a ) or ( a1699a );
 a6121a <=( a1700a ) or ( a6120a );
 a6125a <=( a1695a ) or ( a1696a );
 a6126a <=( a1697a ) or ( a6125a );
 a6127a <=( a6126a ) or ( a6121a );
 a6131a <=( a1692a ) or ( a1693a );
 a6132a <=( a1694a ) or ( a6131a );
 a6135a <=( a1690a ) or ( a1691a );
 a6138a <=( a1688a ) or ( a1689a );
 a6139a <=( a6138a ) or ( a6135a );
 a6140a <=( a6139a ) or ( a6132a );
 a6141a <=( a6140a ) or ( a6127a );
 a6142a <=( a6141a ) or ( a6116a );
 a6143a <=( a6142a ) or ( a6093a );
 a6144a <=( a6143a ) or ( a6044a );
 a6148a <=( a1685a ) or ( a1686a );
 a6149a <=( a1687a ) or ( a6148a );
 a6153a <=( a1682a ) or ( a1683a );
 a6154a <=( a1684a ) or ( a6153a );
 a6155a <=( a6154a ) or ( a6149a );
 a6159a <=( a1679a ) or ( a1680a );
 a6160a <=( a1681a ) or ( a6159a );
 a6164a <=( a1676a ) or ( a1677a );
 a6165a <=( a1678a ) or ( a6164a );
 a6166a <=( a6165a ) or ( a6160a );
 a6167a <=( a6166a ) or ( a6155a );
 a6171a <=( a1673a ) or ( a1674a );
 a6172a <=( a1675a ) or ( a6171a );
 a6176a <=( a1670a ) or ( a1671a );
 a6177a <=( a1672a ) or ( a6176a );
 a6178a <=( a6177a ) or ( a6172a );
 a6182a <=( a1667a ) or ( a1668a );
 a6183a <=( a1669a ) or ( a6182a );
 a6186a <=( a1665a ) or ( a1666a );
 a6189a <=( a1663a ) or ( a1664a );
 a6190a <=( a6189a ) or ( a6186a );
 a6191a <=( a6190a ) or ( a6183a );
 a6192a <=( a6191a ) or ( a6178a );
 a6193a <=( a6192a ) or ( a6167a );
 a6197a <=( a1660a ) or ( a1661a );
 a6198a <=( a1662a ) or ( a6197a );
 a6202a <=( a1657a ) or ( a1658a );
 a6203a <=( a1659a ) or ( a6202a );
 a6204a <=( a6203a ) or ( a6198a );
 a6208a <=( a1654a ) or ( a1655a );
 a6209a <=( a1656a ) or ( a6208a );
 a6213a <=( a1651a ) or ( a1652a );
 a6214a <=( a1653a ) or ( a6213a );
 a6215a <=( a6214a ) or ( a6209a );
 a6216a <=( a6215a ) or ( a6204a );
 a6220a <=( a1648a ) or ( a1649a );
 a6221a <=( a1650a ) or ( a6220a );
 a6225a <=( a1645a ) or ( a1646a );
 a6226a <=( a1647a ) or ( a6225a );
 a6227a <=( a6226a ) or ( a6221a );
 a6231a <=( a1642a ) or ( a1643a );
 a6232a <=( a1644a ) or ( a6231a );
 a6235a <=( a1640a ) or ( a1641a );
 a6238a <=( a1638a ) or ( a1639a );
 a6239a <=( a6238a ) or ( a6235a );
 a6240a <=( a6239a ) or ( a6232a );
 a6241a <=( a6240a ) or ( a6227a );
 a6242a <=( a6241a ) or ( a6216a );
 a6243a <=( a6242a ) or ( a6193a );
 a6247a <=( a1635a ) or ( a1636a );
 a6248a <=( a1637a ) or ( a6247a );
 a6252a <=( a1632a ) or ( a1633a );
 a6253a <=( a1634a ) or ( a6252a );
 a6254a <=( a6253a ) or ( a6248a );
 a6258a <=( a1629a ) or ( a1630a );
 a6259a <=( a1631a ) or ( a6258a );
 a6263a <=( a1626a ) or ( a1627a );
 a6264a <=( a1628a ) or ( a6263a );
 a6265a <=( a6264a ) or ( a6259a );
 a6266a <=( a6265a ) or ( a6254a );
 a6270a <=( a1623a ) or ( a1624a );
 a6271a <=( a1625a ) or ( a6270a );
 a6275a <=( a1620a ) or ( a1621a );
 a6276a <=( a1622a ) or ( a6275a );
 a6277a <=( a6276a ) or ( a6271a );
 a6281a <=( a1617a ) or ( a1618a );
 a6282a <=( a1619a ) or ( a6281a );
 a6285a <=( a1615a ) or ( a1616a );
 a6288a <=( a1613a ) or ( a1614a );
 a6289a <=( a6288a ) or ( a6285a );
 a6290a <=( a6289a ) or ( a6282a );
 a6291a <=( a6290a ) or ( a6277a );
 a6292a <=( a6291a ) or ( a6266a );
 a6296a <=( a1610a ) or ( a1611a );
 a6297a <=( a1612a ) or ( a6296a );
 a6301a <=( a1607a ) or ( a1608a );
 a6302a <=( a1609a ) or ( a6301a );
 a6303a <=( a6302a ) or ( a6297a );
 a6307a <=( a1604a ) or ( a1605a );
 a6308a <=( a1606a ) or ( a6307a );
 a6312a <=( a1601a ) or ( a1602a );
 a6313a <=( a1603a ) or ( a6312a );
 a6314a <=( a6313a ) or ( a6308a );
 a6315a <=( a6314a ) or ( a6303a );
 a6319a <=( a1598a ) or ( a1599a );
 a6320a <=( a1600a ) or ( a6319a );
 a6324a <=( a1595a ) or ( a1596a );
 a6325a <=( a1597a ) or ( a6324a );
 a6326a <=( a6325a ) or ( a6320a );
 a6330a <=( a1592a ) or ( a1593a );
 a6331a <=( a1594a ) or ( a6330a );
 a6334a <=( a1590a ) or ( a1591a );
 a6337a <=( a1588a ) or ( a1589a );
 a6338a <=( a6337a ) or ( a6334a );
 a6339a <=( a6338a ) or ( a6331a );
 a6340a <=( a6339a ) or ( a6326a );
 a6341a <=( a6340a ) or ( a6315a );
 a6342a <=( a6341a ) or ( a6292a );
 a6343a <=( a6342a ) or ( a6243a );
 a6344a <=( a6343a ) or ( a6144a );
 a6345a <=( a6344a ) or ( a5947a );
 a6346a <=( a6345a ) or ( a5552a );
 a6347a <=( a6346a ) or ( a4759a );
 a6351a <=( a1585a ) or ( a1586a );
 a6352a <=( a1587a ) or ( a6351a );
 a6356a <=( a1582a ) or ( a1583a );
 a6357a <=( a1584a ) or ( a6356a );
 a6358a <=( a6357a ) or ( a6352a );
 a6362a <=( a1579a ) or ( a1580a );
 a6363a <=( a1581a ) or ( a6362a );
 a6367a <=( a1576a ) or ( a1577a );
 a6368a <=( a1578a ) or ( a6367a );
 a6369a <=( a6368a ) or ( a6363a );
 a6370a <=( a6369a ) or ( a6358a );
 a6374a <=( a1573a ) or ( a1574a );
 a6375a <=( a1575a ) or ( a6374a );
 a6379a <=( a1570a ) or ( a1571a );
 a6380a <=( a1572a ) or ( a6379a );
 a6381a <=( a6380a ) or ( a6375a );
 a6385a <=( a1567a ) or ( a1568a );
 a6386a <=( a1569a ) or ( a6385a );
 a6390a <=( a1564a ) or ( a1565a );
 a6391a <=( a1566a ) or ( a6390a );
 a6392a <=( a6391a ) or ( a6386a );
 a6393a <=( a6392a ) or ( a6381a );
 a6394a <=( a6393a ) or ( a6370a );
 a6398a <=( a1561a ) or ( a1562a );
 a6399a <=( a1563a ) or ( a6398a );
 a6403a <=( a1558a ) or ( a1559a );
 a6404a <=( a1560a ) or ( a6403a );
 a6405a <=( a6404a ) or ( a6399a );
 a6409a <=( a1555a ) or ( a1556a );
 a6410a <=( a1557a ) or ( a6409a );
 a6414a <=( a1552a ) or ( a1553a );
 a6415a <=( a1554a ) or ( a6414a );
 a6416a <=( a6415a ) or ( a6410a );
 a6417a <=( a6416a ) or ( a6405a );
 a6421a <=( a1549a ) or ( a1550a );
 a6422a <=( a1551a ) or ( a6421a );
 a6426a <=( a1546a ) or ( a1547a );
 a6427a <=( a1548a ) or ( a6426a );
 a6428a <=( a6427a ) or ( a6422a );
 a6432a <=( a1543a ) or ( a1544a );
 a6433a <=( a1545a ) or ( a6432a );
 a6436a <=( a1541a ) or ( a1542a );
 a6439a <=( a1539a ) or ( a1540a );
 a6440a <=( a6439a ) or ( a6436a );
 a6441a <=( a6440a ) or ( a6433a );
 a6442a <=( a6441a ) or ( a6428a );
 a6443a <=( a6442a ) or ( a6417a );
 a6444a <=( a6443a ) or ( a6394a );
 a6448a <=( a1536a ) or ( a1537a );
 a6449a <=( a1538a ) or ( a6448a );
 a6453a <=( a1533a ) or ( a1534a );
 a6454a <=( a1535a ) or ( a6453a );
 a6455a <=( a6454a ) or ( a6449a );
 a6459a <=( a1530a ) or ( a1531a );
 a6460a <=( a1532a ) or ( a6459a );
 a6464a <=( a1527a ) or ( a1528a );
 a6465a <=( a1529a ) or ( a6464a );
 a6466a <=( a6465a ) or ( a6460a );
 a6467a <=( a6466a ) or ( a6455a );
 a6471a <=( a1524a ) or ( a1525a );
 a6472a <=( a1526a ) or ( a6471a );
 a6476a <=( a1521a ) or ( a1522a );
 a6477a <=( a1523a ) or ( a6476a );
 a6478a <=( a6477a ) or ( a6472a );
 a6482a <=( a1518a ) or ( a1519a );
 a6483a <=( a1520a ) or ( a6482a );
 a6486a <=( a1516a ) or ( a1517a );
 a6489a <=( a1514a ) or ( a1515a );
 a6490a <=( a6489a ) or ( a6486a );
 a6491a <=( a6490a ) or ( a6483a );
 a6492a <=( a6491a ) or ( a6478a );
 a6493a <=( a6492a ) or ( a6467a );
 a6497a <=( a1511a ) or ( a1512a );
 a6498a <=( a1513a ) or ( a6497a );
 a6502a <=( a1508a ) or ( a1509a );
 a6503a <=( a1510a ) or ( a6502a );
 a6504a <=( a6503a ) or ( a6498a );
 a6508a <=( a1505a ) or ( a1506a );
 a6509a <=( a1507a ) or ( a6508a );
 a6513a <=( a1502a ) or ( a1503a );
 a6514a <=( a1504a ) or ( a6513a );
 a6515a <=( a6514a ) or ( a6509a );
 a6516a <=( a6515a ) or ( a6504a );
 a6520a <=( a1499a ) or ( a1500a );
 a6521a <=( a1501a ) or ( a6520a );
 a6525a <=( a1496a ) or ( a1497a );
 a6526a <=( a1498a ) or ( a6525a );
 a6527a <=( a6526a ) or ( a6521a );
 a6531a <=( a1493a ) or ( a1494a );
 a6532a <=( a1495a ) or ( a6531a );
 a6535a <=( a1491a ) or ( a1492a );
 a6538a <=( a1489a ) or ( a1490a );
 a6539a <=( a6538a ) or ( a6535a );
 a6540a <=( a6539a ) or ( a6532a );
 a6541a <=( a6540a ) or ( a6527a );
 a6542a <=( a6541a ) or ( a6516a );
 a6543a <=( a6542a ) or ( a6493a );
 a6544a <=( a6543a ) or ( a6444a );
 a6548a <=( a1486a ) or ( a1487a );
 a6549a <=( a1488a ) or ( a6548a );
 a6553a <=( a1483a ) or ( a1484a );
 a6554a <=( a1485a ) or ( a6553a );
 a6555a <=( a6554a ) or ( a6549a );
 a6559a <=( a1480a ) or ( a1481a );
 a6560a <=( a1482a ) or ( a6559a );
 a6564a <=( a1477a ) or ( a1478a );
 a6565a <=( a1479a ) or ( a6564a );
 a6566a <=( a6565a ) or ( a6560a );
 a6567a <=( a6566a ) or ( a6555a );
 a6571a <=( a1474a ) or ( a1475a );
 a6572a <=( a1476a ) or ( a6571a );
 a6576a <=( a1471a ) or ( a1472a );
 a6577a <=( a1473a ) or ( a6576a );
 a6578a <=( a6577a ) or ( a6572a );
 a6582a <=( a1468a ) or ( a1469a );
 a6583a <=( a1470a ) or ( a6582a );
 a6587a <=( a1465a ) or ( a1466a );
 a6588a <=( a1467a ) or ( a6587a );
 a6589a <=( a6588a ) or ( a6583a );
 a6590a <=( a6589a ) or ( a6578a );
 a6591a <=( a6590a ) or ( a6567a );
 a6595a <=( a1462a ) or ( a1463a );
 a6596a <=( a1464a ) or ( a6595a );
 a6600a <=( a1459a ) or ( a1460a );
 a6601a <=( a1461a ) or ( a6600a );
 a6602a <=( a6601a ) or ( a6596a );
 a6606a <=( a1456a ) or ( a1457a );
 a6607a <=( a1458a ) or ( a6606a );
 a6611a <=( a1453a ) or ( a1454a );
 a6612a <=( a1455a ) or ( a6611a );
 a6613a <=( a6612a ) or ( a6607a );
 a6614a <=( a6613a ) or ( a6602a );
 a6618a <=( a1450a ) or ( a1451a );
 a6619a <=( a1452a ) or ( a6618a );
 a6623a <=( a1447a ) or ( a1448a );
 a6624a <=( a1449a ) or ( a6623a );
 a6625a <=( a6624a ) or ( a6619a );
 a6629a <=( a1444a ) or ( a1445a );
 a6630a <=( a1446a ) or ( a6629a );
 a6633a <=( a1442a ) or ( a1443a );
 a6636a <=( a1440a ) or ( a1441a );
 a6637a <=( a6636a ) or ( a6633a );
 a6638a <=( a6637a ) or ( a6630a );
 a6639a <=( a6638a ) or ( a6625a );
 a6640a <=( a6639a ) or ( a6614a );
 a6641a <=( a6640a ) or ( a6591a );
 a6645a <=( a1437a ) or ( a1438a );
 a6646a <=( a1439a ) or ( a6645a );
 a6650a <=( a1434a ) or ( a1435a );
 a6651a <=( a1436a ) or ( a6650a );
 a6652a <=( a6651a ) or ( a6646a );
 a6656a <=( a1431a ) or ( a1432a );
 a6657a <=( a1433a ) or ( a6656a );
 a6661a <=( a1428a ) or ( a1429a );
 a6662a <=( a1430a ) or ( a6661a );
 a6663a <=( a6662a ) or ( a6657a );
 a6664a <=( a6663a ) or ( a6652a );
 a6668a <=( a1425a ) or ( a1426a );
 a6669a <=( a1427a ) or ( a6668a );
 a6673a <=( a1422a ) or ( a1423a );
 a6674a <=( a1424a ) or ( a6673a );
 a6675a <=( a6674a ) or ( a6669a );
 a6679a <=( a1419a ) or ( a1420a );
 a6680a <=( a1421a ) or ( a6679a );
 a6683a <=( a1417a ) or ( a1418a );
 a6686a <=( a1415a ) or ( a1416a );
 a6687a <=( a6686a ) or ( a6683a );
 a6688a <=( a6687a ) or ( a6680a );
 a6689a <=( a6688a ) or ( a6675a );
 a6690a <=( a6689a ) or ( a6664a );
 a6694a <=( a1412a ) or ( a1413a );
 a6695a <=( a1414a ) or ( a6694a );
 a6699a <=( a1409a ) or ( a1410a );
 a6700a <=( a1411a ) or ( a6699a );
 a6701a <=( a6700a ) or ( a6695a );
 a6705a <=( a1406a ) or ( a1407a );
 a6706a <=( a1408a ) or ( a6705a );
 a6710a <=( a1403a ) or ( a1404a );
 a6711a <=( a1405a ) or ( a6710a );
 a6712a <=( a6711a ) or ( a6706a );
 a6713a <=( a6712a ) or ( a6701a );
 a6717a <=( a1400a ) or ( a1401a );
 a6718a <=( a1402a ) or ( a6717a );
 a6722a <=( a1397a ) or ( a1398a );
 a6723a <=( a1399a ) or ( a6722a );
 a6724a <=( a6723a ) or ( a6718a );
 a6728a <=( a1394a ) or ( a1395a );
 a6729a <=( a1396a ) or ( a6728a );
 a6732a <=( a1392a ) or ( a1393a );
 a6735a <=( a1390a ) or ( a1391a );
 a6736a <=( a6735a ) or ( a6732a );
 a6737a <=( a6736a ) or ( a6729a );
 a6738a <=( a6737a ) or ( a6724a );
 a6739a <=( a6738a ) or ( a6713a );
 a6740a <=( a6739a ) or ( a6690a );
 a6741a <=( a6740a ) or ( a6641a );
 a6742a <=( a6741a ) or ( a6544a );
 a6746a <=( a1387a ) or ( a1388a );
 a6747a <=( a1389a ) or ( a6746a );
 a6751a <=( a1384a ) or ( a1385a );
 a6752a <=( a1386a ) or ( a6751a );
 a6753a <=( a6752a ) or ( a6747a );
 a6757a <=( a1381a ) or ( a1382a );
 a6758a <=( a1383a ) or ( a6757a );
 a6762a <=( a1378a ) or ( a1379a );
 a6763a <=( a1380a ) or ( a6762a );
 a6764a <=( a6763a ) or ( a6758a );
 a6765a <=( a6764a ) or ( a6753a );
 a6769a <=( a1375a ) or ( a1376a );
 a6770a <=( a1377a ) or ( a6769a );
 a6774a <=( a1372a ) or ( a1373a );
 a6775a <=( a1374a ) or ( a6774a );
 a6776a <=( a6775a ) or ( a6770a );
 a6780a <=( a1369a ) or ( a1370a );
 a6781a <=( a1371a ) or ( a6780a );
 a6785a <=( a1366a ) or ( a1367a );
 a6786a <=( a1368a ) or ( a6785a );
 a6787a <=( a6786a ) or ( a6781a );
 a6788a <=( a6787a ) or ( a6776a );
 a6789a <=( a6788a ) or ( a6765a );
 a6793a <=( a1363a ) or ( a1364a );
 a6794a <=( a1365a ) or ( a6793a );
 a6798a <=( a1360a ) or ( a1361a );
 a6799a <=( a1362a ) or ( a6798a );
 a6800a <=( a6799a ) or ( a6794a );
 a6804a <=( a1357a ) or ( a1358a );
 a6805a <=( a1359a ) or ( a6804a );
 a6809a <=( a1354a ) or ( a1355a );
 a6810a <=( a1356a ) or ( a6809a );
 a6811a <=( a6810a ) or ( a6805a );
 a6812a <=( a6811a ) or ( a6800a );
 a6816a <=( a1351a ) or ( a1352a );
 a6817a <=( a1353a ) or ( a6816a );
 a6821a <=( a1348a ) or ( a1349a );
 a6822a <=( a1350a ) or ( a6821a );
 a6823a <=( a6822a ) or ( a6817a );
 a6827a <=( a1345a ) or ( a1346a );
 a6828a <=( a1347a ) or ( a6827a );
 a6831a <=( a1343a ) or ( a1344a );
 a6834a <=( a1341a ) or ( a1342a );
 a6835a <=( a6834a ) or ( a6831a );
 a6836a <=( a6835a ) or ( a6828a );
 a6837a <=( a6836a ) or ( a6823a );
 a6838a <=( a6837a ) or ( a6812a );
 a6839a <=( a6838a ) or ( a6789a );
 a6843a <=( a1338a ) or ( a1339a );
 a6844a <=( a1340a ) or ( a6843a );
 a6848a <=( a1335a ) or ( a1336a );
 a6849a <=( a1337a ) or ( a6848a );
 a6850a <=( a6849a ) or ( a6844a );
 a6854a <=( a1332a ) or ( a1333a );
 a6855a <=( a1334a ) or ( a6854a );
 a6859a <=( a1329a ) or ( a1330a );
 a6860a <=( a1331a ) or ( a6859a );
 a6861a <=( a6860a ) or ( a6855a );
 a6862a <=( a6861a ) or ( a6850a );
 a6866a <=( a1326a ) or ( a1327a );
 a6867a <=( a1328a ) or ( a6866a );
 a6871a <=( a1323a ) or ( a1324a );
 a6872a <=( a1325a ) or ( a6871a );
 a6873a <=( a6872a ) or ( a6867a );
 a6877a <=( a1320a ) or ( a1321a );
 a6878a <=( a1322a ) or ( a6877a );
 a6881a <=( a1318a ) or ( a1319a );
 a6884a <=( a1316a ) or ( a1317a );
 a6885a <=( a6884a ) or ( a6881a );
 a6886a <=( a6885a ) or ( a6878a );
 a6887a <=( a6886a ) or ( a6873a );
 a6888a <=( a6887a ) or ( a6862a );
 a6892a <=( a1313a ) or ( a1314a );
 a6893a <=( a1315a ) or ( a6892a );
 a6897a <=( a1310a ) or ( a1311a );
 a6898a <=( a1312a ) or ( a6897a );
 a6899a <=( a6898a ) or ( a6893a );
 a6903a <=( a1307a ) or ( a1308a );
 a6904a <=( a1309a ) or ( a6903a );
 a6908a <=( a1304a ) or ( a1305a );
 a6909a <=( a1306a ) or ( a6908a );
 a6910a <=( a6909a ) or ( a6904a );
 a6911a <=( a6910a ) or ( a6899a );
 a6915a <=( a1301a ) or ( a1302a );
 a6916a <=( a1303a ) or ( a6915a );
 a6920a <=( a1298a ) or ( a1299a );
 a6921a <=( a1300a ) or ( a6920a );
 a6922a <=( a6921a ) or ( a6916a );
 a6926a <=( a1295a ) or ( a1296a );
 a6927a <=( a1297a ) or ( a6926a );
 a6930a <=( a1293a ) or ( a1294a );
 a6933a <=( a1291a ) or ( a1292a );
 a6934a <=( a6933a ) or ( a6930a );
 a6935a <=( a6934a ) or ( a6927a );
 a6936a <=( a6935a ) or ( a6922a );
 a6937a <=( a6936a ) or ( a6911a );
 a6938a <=( a6937a ) or ( a6888a );
 a6939a <=( a6938a ) or ( a6839a );
 a6943a <=( a1288a ) or ( a1289a );
 a6944a <=( a1290a ) or ( a6943a );
 a6948a <=( a1285a ) or ( a1286a );
 a6949a <=( a1287a ) or ( a6948a );
 a6950a <=( a6949a ) or ( a6944a );
 a6954a <=( a1282a ) or ( a1283a );
 a6955a <=( a1284a ) or ( a6954a );
 a6959a <=( a1279a ) or ( a1280a );
 a6960a <=( a1281a ) or ( a6959a );
 a6961a <=( a6960a ) or ( a6955a );
 a6962a <=( a6961a ) or ( a6950a );
 a6966a <=( a1276a ) or ( a1277a );
 a6967a <=( a1278a ) or ( a6966a );
 a6971a <=( a1273a ) or ( a1274a );
 a6972a <=( a1275a ) or ( a6971a );
 a6973a <=( a6972a ) or ( a6967a );
 a6977a <=( a1270a ) or ( a1271a );
 a6978a <=( a1272a ) or ( a6977a );
 a6982a <=( a1267a ) or ( a1268a );
 a6983a <=( a1269a ) or ( a6982a );
 a6984a <=( a6983a ) or ( a6978a );
 a6985a <=( a6984a ) or ( a6973a );
 a6986a <=( a6985a ) or ( a6962a );
 a6990a <=( a1264a ) or ( a1265a );
 a6991a <=( a1266a ) or ( a6990a );
 a6995a <=( a1261a ) or ( a1262a );
 a6996a <=( a1263a ) or ( a6995a );
 a6997a <=( a6996a ) or ( a6991a );
 a7001a <=( a1258a ) or ( a1259a );
 a7002a <=( a1260a ) or ( a7001a );
 a7006a <=( a1255a ) or ( a1256a );
 a7007a <=( a1257a ) or ( a7006a );
 a7008a <=( a7007a ) or ( a7002a );
 a7009a <=( a7008a ) or ( a6997a );
 a7013a <=( a1252a ) or ( a1253a );
 a7014a <=( a1254a ) or ( a7013a );
 a7018a <=( a1249a ) or ( a1250a );
 a7019a <=( a1251a ) or ( a7018a );
 a7020a <=( a7019a ) or ( a7014a );
 a7024a <=( a1246a ) or ( a1247a );
 a7025a <=( a1248a ) or ( a7024a );
 a7028a <=( a1244a ) or ( a1245a );
 a7031a <=( a1242a ) or ( a1243a );
 a7032a <=( a7031a ) or ( a7028a );
 a7033a <=( a7032a ) or ( a7025a );
 a7034a <=( a7033a ) or ( a7020a );
 a7035a <=( a7034a ) or ( a7009a );
 a7036a <=( a7035a ) or ( a6986a );
 a7040a <=( a1239a ) or ( a1240a );
 a7041a <=( a1241a ) or ( a7040a );
 a7045a <=( a1236a ) or ( a1237a );
 a7046a <=( a1238a ) or ( a7045a );
 a7047a <=( a7046a ) or ( a7041a );
 a7051a <=( a1233a ) or ( a1234a );
 a7052a <=( a1235a ) or ( a7051a );
 a7056a <=( a1230a ) or ( a1231a );
 a7057a <=( a1232a ) or ( a7056a );
 a7058a <=( a7057a ) or ( a7052a );
 a7059a <=( a7058a ) or ( a7047a );
 a7063a <=( a1227a ) or ( a1228a );
 a7064a <=( a1229a ) or ( a7063a );
 a7068a <=( a1224a ) or ( a1225a );
 a7069a <=( a1226a ) or ( a7068a );
 a7070a <=( a7069a ) or ( a7064a );
 a7074a <=( a1221a ) or ( a1222a );
 a7075a <=( a1223a ) or ( a7074a );
 a7078a <=( a1219a ) or ( a1220a );
 a7081a <=( a1217a ) or ( a1218a );
 a7082a <=( a7081a ) or ( a7078a );
 a7083a <=( a7082a ) or ( a7075a );
 a7084a <=( a7083a ) or ( a7070a );
 a7085a <=( a7084a ) or ( a7059a );
 a7089a <=( a1214a ) or ( a1215a );
 a7090a <=( a1216a ) or ( a7089a );
 a7094a <=( a1211a ) or ( a1212a );
 a7095a <=( a1213a ) or ( a7094a );
 a7096a <=( a7095a ) or ( a7090a );
 a7100a <=( a1208a ) or ( a1209a );
 a7101a <=( a1210a ) or ( a7100a );
 a7105a <=( a1205a ) or ( a1206a );
 a7106a <=( a1207a ) or ( a7105a );
 a7107a <=( a7106a ) or ( a7101a );
 a7108a <=( a7107a ) or ( a7096a );
 a7112a <=( a1202a ) or ( a1203a );
 a7113a <=( a1204a ) or ( a7112a );
 a7117a <=( a1199a ) or ( a1200a );
 a7118a <=( a1201a ) or ( a7117a );
 a7119a <=( a7118a ) or ( a7113a );
 a7123a <=( a1196a ) or ( a1197a );
 a7124a <=( a1198a ) or ( a7123a );
 a7127a <=( a1194a ) or ( a1195a );
 a7130a <=( a1192a ) or ( a1193a );
 a7131a <=( a7130a ) or ( a7127a );
 a7132a <=( a7131a ) or ( a7124a );
 a7133a <=( a7132a ) or ( a7119a );
 a7134a <=( a7133a ) or ( a7108a );
 a7135a <=( a7134a ) or ( a7085a );
 a7136a <=( a7135a ) or ( a7036a );
 a7137a <=( a7136a ) or ( a6939a );
 a7138a <=( a7137a ) or ( a6742a );
 a7142a <=( a1189a ) or ( a1190a );
 a7143a <=( a1191a ) or ( a7142a );
 a7147a <=( a1186a ) or ( a1187a );
 a7148a <=( a1188a ) or ( a7147a );
 a7149a <=( a7148a ) or ( a7143a );
 a7153a <=( a1183a ) or ( a1184a );
 a7154a <=( a1185a ) or ( a7153a );
 a7158a <=( a1180a ) or ( a1181a );
 a7159a <=( a1182a ) or ( a7158a );
 a7160a <=( a7159a ) or ( a7154a );
 a7161a <=( a7160a ) or ( a7149a );
 a7165a <=( a1177a ) or ( a1178a );
 a7166a <=( a1179a ) or ( a7165a );
 a7170a <=( a1174a ) or ( a1175a );
 a7171a <=( a1176a ) or ( a7170a );
 a7172a <=( a7171a ) or ( a7166a );
 a7176a <=( a1171a ) or ( a1172a );
 a7177a <=( a1173a ) or ( a7176a );
 a7181a <=( a1168a ) or ( a1169a );
 a7182a <=( a1170a ) or ( a7181a );
 a7183a <=( a7182a ) or ( a7177a );
 a7184a <=( a7183a ) or ( a7172a );
 a7185a <=( a7184a ) or ( a7161a );
 a7189a <=( a1165a ) or ( a1166a );
 a7190a <=( a1167a ) or ( a7189a );
 a7194a <=( a1162a ) or ( a1163a );
 a7195a <=( a1164a ) or ( a7194a );
 a7196a <=( a7195a ) or ( a7190a );
 a7200a <=( a1159a ) or ( a1160a );
 a7201a <=( a1161a ) or ( a7200a );
 a7205a <=( a1156a ) or ( a1157a );
 a7206a <=( a1158a ) or ( a7205a );
 a7207a <=( a7206a ) or ( a7201a );
 a7208a <=( a7207a ) or ( a7196a );
 a7212a <=( a1153a ) or ( a1154a );
 a7213a <=( a1155a ) or ( a7212a );
 a7217a <=( a1150a ) or ( a1151a );
 a7218a <=( a1152a ) or ( a7217a );
 a7219a <=( a7218a ) or ( a7213a );
 a7223a <=( a1147a ) or ( a1148a );
 a7224a <=( a1149a ) or ( a7223a );
 a7227a <=( a1145a ) or ( a1146a );
 a7230a <=( a1143a ) or ( a1144a );
 a7231a <=( a7230a ) or ( a7227a );
 a7232a <=( a7231a ) or ( a7224a );
 a7233a <=( a7232a ) or ( a7219a );
 a7234a <=( a7233a ) or ( a7208a );
 a7235a <=( a7234a ) or ( a7185a );
 a7239a <=( a1140a ) or ( a1141a );
 a7240a <=( a1142a ) or ( a7239a );
 a7244a <=( a1137a ) or ( a1138a );
 a7245a <=( a1139a ) or ( a7244a );
 a7246a <=( a7245a ) or ( a7240a );
 a7250a <=( a1134a ) or ( a1135a );
 a7251a <=( a1136a ) or ( a7250a );
 a7255a <=( a1131a ) or ( a1132a );
 a7256a <=( a1133a ) or ( a7255a );
 a7257a <=( a7256a ) or ( a7251a );
 a7258a <=( a7257a ) or ( a7246a );
 a7262a <=( a1128a ) or ( a1129a );
 a7263a <=( a1130a ) or ( a7262a );
 a7267a <=( a1125a ) or ( a1126a );
 a7268a <=( a1127a ) or ( a7267a );
 a7269a <=( a7268a ) or ( a7263a );
 a7273a <=( a1122a ) or ( a1123a );
 a7274a <=( a1124a ) or ( a7273a );
 a7277a <=( a1120a ) or ( a1121a );
 a7280a <=( a1118a ) or ( a1119a );
 a7281a <=( a7280a ) or ( a7277a );
 a7282a <=( a7281a ) or ( a7274a );
 a7283a <=( a7282a ) or ( a7269a );
 a7284a <=( a7283a ) or ( a7258a );
 a7288a <=( a1115a ) or ( a1116a );
 a7289a <=( a1117a ) or ( a7288a );
 a7293a <=( a1112a ) or ( a1113a );
 a7294a <=( a1114a ) or ( a7293a );
 a7295a <=( a7294a ) or ( a7289a );
 a7299a <=( a1109a ) or ( a1110a );
 a7300a <=( a1111a ) or ( a7299a );
 a7304a <=( a1106a ) or ( a1107a );
 a7305a <=( a1108a ) or ( a7304a );
 a7306a <=( a7305a ) or ( a7300a );
 a7307a <=( a7306a ) or ( a7295a );
 a7311a <=( a1103a ) or ( a1104a );
 a7312a <=( a1105a ) or ( a7311a );
 a7316a <=( a1100a ) or ( a1101a );
 a7317a <=( a1102a ) or ( a7316a );
 a7318a <=( a7317a ) or ( a7312a );
 a7322a <=( a1097a ) or ( a1098a );
 a7323a <=( a1099a ) or ( a7322a );
 a7326a <=( a1095a ) or ( a1096a );
 a7329a <=( a1093a ) or ( a1094a );
 a7330a <=( a7329a ) or ( a7326a );
 a7331a <=( a7330a ) or ( a7323a );
 a7332a <=( a7331a ) or ( a7318a );
 a7333a <=( a7332a ) or ( a7307a );
 a7334a <=( a7333a ) or ( a7284a );
 a7335a <=( a7334a ) or ( a7235a );
 a7339a <=( a1090a ) or ( a1091a );
 a7340a <=( a1092a ) or ( a7339a );
 a7344a <=( a1087a ) or ( a1088a );
 a7345a <=( a1089a ) or ( a7344a );
 a7346a <=( a7345a ) or ( a7340a );
 a7350a <=( a1084a ) or ( a1085a );
 a7351a <=( a1086a ) or ( a7350a );
 a7355a <=( a1081a ) or ( a1082a );
 a7356a <=( a1083a ) or ( a7355a );
 a7357a <=( a7356a ) or ( a7351a );
 a7358a <=( a7357a ) or ( a7346a );
 a7362a <=( a1078a ) or ( a1079a );
 a7363a <=( a1080a ) or ( a7362a );
 a7367a <=( a1075a ) or ( a1076a );
 a7368a <=( a1077a ) or ( a7367a );
 a7369a <=( a7368a ) or ( a7363a );
 a7373a <=( a1072a ) or ( a1073a );
 a7374a <=( a1074a ) or ( a7373a );
 a7378a <=( a1069a ) or ( a1070a );
 a7379a <=( a1071a ) or ( a7378a );
 a7380a <=( a7379a ) or ( a7374a );
 a7381a <=( a7380a ) or ( a7369a );
 a7382a <=( a7381a ) or ( a7358a );
 a7386a <=( a1066a ) or ( a1067a );
 a7387a <=( a1068a ) or ( a7386a );
 a7391a <=( a1063a ) or ( a1064a );
 a7392a <=( a1065a ) or ( a7391a );
 a7393a <=( a7392a ) or ( a7387a );
 a7397a <=( a1060a ) or ( a1061a );
 a7398a <=( a1062a ) or ( a7397a );
 a7402a <=( a1057a ) or ( a1058a );
 a7403a <=( a1059a ) or ( a7402a );
 a7404a <=( a7403a ) or ( a7398a );
 a7405a <=( a7404a ) or ( a7393a );
 a7409a <=( a1054a ) or ( a1055a );
 a7410a <=( a1056a ) or ( a7409a );
 a7414a <=( a1051a ) or ( a1052a );
 a7415a <=( a1053a ) or ( a7414a );
 a7416a <=( a7415a ) or ( a7410a );
 a7420a <=( a1048a ) or ( a1049a );
 a7421a <=( a1050a ) or ( a7420a );
 a7424a <=( a1046a ) or ( a1047a );
 a7427a <=( a1044a ) or ( a1045a );
 a7428a <=( a7427a ) or ( a7424a );
 a7429a <=( a7428a ) or ( a7421a );
 a7430a <=( a7429a ) or ( a7416a );
 a7431a <=( a7430a ) or ( a7405a );
 a7432a <=( a7431a ) or ( a7382a );
 a7436a <=( a1041a ) or ( a1042a );
 a7437a <=( a1043a ) or ( a7436a );
 a7441a <=( a1038a ) or ( a1039a );
 a7442a <=( a1040a ) or ( a7441a );
 a7443a <=( a7442a ) or ( a7437a );
 a7447a <=( a1035a ) or ( a1036a );
 a7448a <=( a1037a ) or ( a7447a );
 a7452a <=( a1032a ) or ( a1033a );
 a7453a <=( a1034a ) or ( a7452a );
 a7454a <=( a7453a ) or ( a7448a );
 a7455a <=( a7454a ) or ( a7443a );
 a7459a <=( a1029a ) or ( a1030a );
 a7460a <=( a1031a ) or ( a7459a );
 a7464a <=( a1026a ) or ( a1027a );
 a7465a <=( a1028a ) or ( a7464a );
 a7466a <=( a7465a ) or ( a7460a );
 a7470a <=( a1023a ) or ( a1024a );
 a7471a <=( a1025a ) or ( a7470a );
 a7474a <=( a1021a ) or ( a1022a );
 a7477a <=( a1019a ) or ( a1020a );
 a7478a <=( a7477a ) or ( a7474a );
 a7479a <=( a7478a ) or ( a7471a );
 a7480a <=( a7479a ) or ( a7466a );
 a7481a <=( a7480a ) or ( a7455a );
 a7485a <=( a1016a ) or ( a1017a );
 a7486a <=( a1018a ) or ( a7485a );
 a7490a <=( a1013a ) or ( a1014a );
 a7491a <=( a1015a ) or ( a7490a );
 a7492a <=( a7491a ) or ( a7486a );
 a7496a <=( a1010a ) or ( a1011a );
 a7497a <=( a1012a ) or ( a7496a );
 a7501a <=( a1007a ) or ( a1008a );
 a7502a <=( a1009a ) or ( a7501a );
 a7503a <=( a7502a ) or ( a7497a );
 a7504a <=( a7503a ) or ( a7492a );
 a7508a <=( a1004a ) or ( a1005a );
 a7509a <=( a1006a ) or ( a7508a );
 a7513a <=( a1001a ) or ( a1002a );
 a7514a <=( a1003a ) or ( a7513a );
 a7515a <=( a7514a ) or ( a7509a );
 a7519a <=( a998a ) or ( a999a );
 a7520a <=( a1000a ) or ( a7519a );
 a7523a <=( a996a ) or ( a997a );
 a7526a <=( a994a ) or ( a995a );
 a7527a <=( a7526a ) or ( a7523a );
 a7528a <=( a7527a ) or ( a7520a );
 a7529a <=( a7528a ) or ( a7515a );
 a7530a <=( a7529a ) or ( a7504a );
 a7531a <=( a7530a ) or ( a7481a );
 a7532a <=( a7531a ) or ( a7432a );
 a7533a <=( a7532a ) or ( a7335a );
 a7537a <=( a991a ) or ( a992a );
 a7538a <=( a993a ) or ( a7537a );
 a7542a <=( a988a ) or ( a989a );
 a7543a <=( a990a ) or ( a7542a );
 a7544a <=( a7543a ) or ( a7538a );
 a7548a <=( a985a ) or ( a986a );
 a7549a <=( a987a ) or ( a7548a );
 a7553a <=( a982a ) or ( a983a );
 a7554a <=( a984a ) or ( a7553a );
 a7555a <=( a7554a ) or ( a7549a );
 a7556a <=( a7555a ) or ( a7544a );
 a7560a <=( a979a ) or ( a980a );
 a7561a <=( a981a ) or ( a7560a );
 a7565a <=( a976a ) or ( a977a );
 a7566a <=( a978a ) or ( a7565a );
 a7567a <=( a7566a ) or ( a7561a );
 a7571a <=( a973a ) or ( a974a );
 a7572a <=( a975a ) or ( a7571a );
 a7576a <=( a970a ) or ( a971a );
 a7577a <=( a972a ) or ( a7576a );
 a7578a <=( a7577a ) or ( a7572a );
 a7579a <=( a7578a ) or ( a7567a );
 a7580a <=( a7579a ) or ( a7556a );
 a7584a <=( a967a ) or ( a968a );
 a7585a <=( a969a ) or ( a7584a );
 a7589a <=( a964a ) or ( a965a );
 a7590a <=( a966a ) or ( a7589a );
 a7591a <=( a7590a ) or ( a7585a );
 a7595a <=( a961a ) or ( a962a );
 a7596a <=( a963a ) or ( a7595a );
 a7600a <=( a958a ) or ( a959a );
 a7601a <=( a960a ) or ( a7600a );
 a7602a <=( a7601a ) or ( a7596a );
 a7603a <=( a7602a ) or ( a7591a );
 a7607a <=( a955a ) or ( a956a );
 a7608a <=( a957a ) or ( a7607a );
 a7612a <=( a952a ) or ( a953a );
 a7613a <=( a954a ) or ( a7612a );
 a7614a <=( a7613a ) or ( a7608a );
 a7618a <=( a949a ) or ( a950a );
 a7619a <=( a951a ) or ( a7618a );
 a7622a <=( a947a ) or ( a948a );
 a7625a <=( a945a ) or ( a946a );
 a7626a <=( a7625a ) or ( a7622a );
 a7627a <=( a7626a ) or ( a7619a );
 a7628a <=( a7627a ) or ( a7614a );
 a7629a <=( a7628a ) or ( a7603a );
 a7630a <=( a7629a ) or ( a7580a );
 a7634a <=( a942a ) or ( a943a );
 a7635a <=( a944a ) or ( a7634a );
 a7639a <=( a939a ) or ( a940a );
 a7640a <=( a941a ) or ( a7639a );
 a7641a <=( a7640a ) or ( a7635a );
 a7645a <=( a936a ) or ( a937a );
 a7646a <=( a938a ) or ( a7645a );
 a7650a <=( a933a ) or ( a934a );
 a7651a <=( a935a ) or ( a7650a );
 a7652a <=( a7651a ) or ( a7646a );
 a7653a <=( a7652a ) or ( a7641a );
 a7657a <=( a930a ) or ( a931a );
 a7658a <=( a932a ) or ( a7657a );
 a7662a <=( a927a ) or ( a928a );
 a7663a <=( a929a ) or ( a7662a );
 a7664a <=( a7663a ) or ( a7658a );
 a7668a <=( a924a ) or ( a925a );
 a7669a <=( a926a ) or ( a7668a );
 a7672a <=( a922a ) or ( a923a );
 a7675a <=( a920a ) or ( a921a );
 a7676a <=( a7675a ) or ( a7672a );
 a7677a <=( a7676a ) or ( a7669a );
 a7678a <=( a7677a ) or ( a7664a );
 a7679a <=( a7678a ) or ( a7653a );
 a7683a <=( a917a ) or ( a918a );
 a7684a <=( a919a ) or ( a7683a );
 a7688a <=( a914a ) or ( a915a );
 a7689a <=( a916a ) or ( a7688a );
 a7690a <=( a7689a ) or ( a7684a );
 a7694a <=( a911a ) or ( a912a );
 a7695a <=( a913a ) or ( a7694a );
 a7699a <=( a908a ) or ( a909a );
 a7700a <=( a910a ) or ( a7699a );
 a7701a <=( a7700a ) or ( a7695a );
 a7702a <=( a7701a ) or ( a7690a );
 a7706a <=( a905a ) or ( a906a );
 a7707a <=( a907a ) or ( a7706a );
 a7711a <=( a902a ) or ( a903a );
 a7712a <=( a904a ) or ( a7711a );
 a7713a <=( a7712a ) or ( a7707a );
 a7717a <=( a899a ) or ( a900a );
 a7718a <=( a901a ) or ( a7717a );
 a7721a <=( a897a ) or ( a898a );
 a7724a <=( a895a ) or ( a896a );
 a7725a <=( a7724a ) or ( a7721a );
 a7726a <=( a7725a ) or ( a7718a );
 a7727a <=( a7726a ) or ( a7713a );
 a7728a <=( a7727a ) or ( a7702a );
 a7729a <=( a7728a ) or ( a7679a );
 a7730a <=( a7729a ) or ( a7630a );
 a7734a <=( a892a ) or ( a893a );
 a7735a <=( a894a ) or ( a7734a );
 a7739a <=( a889a ) or ( a890a );
 a7740a <=( a891a ) or ( a7739a );
 a7741a <=( a7740a ) or ( a7735a );
 a7745a <=( a886a ) or ( a887a );
 a7746a <=( a888a ) or ( a7745a );
 a7750a <=( a883a ) or ( a884a );
 a7751a <=( a885a ) or ( a7750a );
 a7752a <=( a7751a ) or ( a7746a );
 a7753a <=( a7752a ) or ( a7741a );
 a7757a <=( a880a ) or ( a881a );
 a7758a <=( a882a ) or ( a7757a );
 a7762a <=( a877a ) or ( a878a );
 a7763a <=( a879a ) or ( a7762a );
 a7764a <=( a7763a ) or ( a7758a );
 a7768a <=( a874a ) or ( a875a );
 a7769a <=( a876a ) or ( a7768a );
 a7772a <=( a872a ) or ( a873a );
 a7775a <=( a870a ) or ( a871a );
 a7776a <=( a7775a ) or ( a7772a );
 a7777a <=( a7776a ) or ( a7769a );
 a7778a <=( a7777a ) or ( a7764a );
 a7779a <=( a7778a ) or ( a7753a );
 a7783a <=( a867a ) or ( a868a );
 a7784a <=( a869a ) or ( a7783a );
 a7788a <=( a864a ) or ( a865a );
 a7789a <=( a866a ) or ( a7788a );
 a7790a <=( a7789a ) or ( a7784a );
 a7794a <=( a861a ) or ( a862a );
 a7795a <=( a863a ) or ( a7794a );
 a7799a <=( a858a ) or ( a859a );
 a7800a <=( a860a ) or ( a7799a );
 a7801a <=( a7800a ) or ( a7795a );
 a7802a <=( a7801a ) or ( a7790a );
 a7806a <=( a855a ) or ( a856a );
 a7807a <=( a857a ) or ( a7806a );
 a7811a <=( a852a ) or ( a853a );
 a7812a <=( a854a ) or ( a7811a );
 a7813a <=( a7812a ) or ( a7807a );
 a7817a <=( a849a ) or ( a850a );
 a7818a <=( a851a ) or ( a7817a );
 a7821a <=( a847a ) or ( a848a );
 a7824a <=( a845a ) or ( a846a );
 a7825a <=( a7824a ) or ( a7821a );
 a7826a <=( a7825a ) or ( a7818a );
 a7827a <=( a7826a ) or ( a7813a );
 a7828a <=( a7827a ) or ( a7802a );
 a7829a <=( a7828a ) or ( a7779a );
 a7833a <=( a842a ) or ( a843a );
 a7834a <=( a844a ) or ( a7833a );
 a7838a <=( a839a ) or ( a840a );
 a7839a <=( a841a ) or ( a7838a );
 a7840a <=( a7839a ) or ( a7834a );
 a7844a <=( a836a ) or ( a837a );
 a7845a <=( a838a ) or ( a7844a );
 a7849a <=( a833a ) or ( a834a );
 a7850a <=( a835a ) or ( a7849a );
 a7851a <=( a7850a ) or ( a7845a );
 a7852a <=( a7851a ) or ( a7840a );
 a7856a <=( a830a ) or ( a831a );
 a7857a <=( a832a ) or ( a7856a );
 a7861a <=( a827a ) or ( a828a );
 a7862a <=( a829a ) or ( a7861a );
 a7863a <=( a7862a ) or ( a7857a );
 a7867a <=( a824a ) or ( a825a );
 a7868a <=( a826a ) or ( a7867a );
 a7871a <=( a822a ) or ( a823a );
 a7874a <=( a820a ) or ( a821a );
 a7875a <=( a7874a ) or ( a7871a );
 a7876a <=( a7875a ) or ( a7868a );
 a7877a <=( a7876a ) or ( a7863a );
 a7878a <=( a7877a ) or ( a7852a );
 a7882a <=( a817a ) or ( a818a );
 a7883a <=( a819a ) or ( a7882a );
 a7887a <=( a814a ) or ( a815a );
 a7888a <=( a816a ) or ( a7887a );
 a7889a <=( a7888a ) or ( a7883a );
 a7893a <=( a811a ) or ( a812a );
 a7894a <=( a813a ) or ( a7893a );
 a7898a <=( a808a ) or ( a809a );
 a7899a <=( a810a ) or ( a7898a );
 a7900a <=( a7899a ) or ( a7894a );
 a7901a <=( a7900a ) or ( a7889a );
 a7905a <=( a805a ) or ( a806a );
 a7906a <=( a807a ) or ( a7905a );
 a7910a <=( a802a ) or ( a803a );
 a7911a <=( a804a ) or ( a7910a );
 a7912a <=( a7911a ) or ( a7906a );
 a7916a <=( a799a ) or ( a800a );
 a7917a <=( a801a ) or ( a7916a );
 a7920a <=( a797a ) or ( a798a );
 a7923a <=( a795a ) or ( a796a );
 a7924a <=( a7923a ) or ( a7920a );
 a7925a <=( a7924a ) or ( a7917a );
 a7926a <=( a7925a ) or ( a7912a );
 a7927a <=( a7926a ) or ( a7901a );
 a7928a <=( a7927a ) or ( a7878a );
 a7929a <=( a7928a ) or ( a7829a );
 a7930a <=( a7929a ) or ( a7730a );
 a7931a <=( a7930a ) or ( a7533a );
 a7932a <=( a7931a ) or ( a7138a );
 a7936a <=( a792a ) or ( a793a );
 a7937a <=( a794a ) or ( a7936a );
 a7941a <=( a789a ) or ( a790a );
 a7942a <=( a791a ) or ( a7941a );
 a7943a <=( a7942a ) or ( a7937a );
 a7947a <=( a786a ) or ( a787a );
 a7948a <=( a788a ) or ( a7947a );
 a7952a <=( a783a ) or ( a784a );
 a7953a <=( a785a ) or ( a7952a );
 a7954a <=( a7953a ) or ( a7948a );
 a7955a <=( a7954a ) or ( a7943a );
 a7959a <=( a780a ) or ( a781a );
 a7960a <=( a782a ) or ( a7959a );
 a7964a <=( a777a ) or ( a778a );
 a7965a <=( a779a ) or ( a7964a );
 a7966a <=( a7965a ) or ( a7960a );
 a7970a <=( a774a ) or ( a775a );
 a7971a <=( a776a ) or ( a7970a );
 a7975a <=( a771a ) or ( a772a );
 a7976a <=( a773a ) or ( a7975a );
 a7977a <=( a7976a ) or ( a7971a );
 a7978a <=( a7977a ) or ( a7966a );
 a7979a <=( a7978a ) or ( a7955a );
 a7983a <=( a768a ) or ( a769a );
 a7984a <=( a770a ) or ( a7983a );
 a7988a <=( a765a ) or ( a766a );
 a7989a <=( a767a ) or ( a7988a );
 a7990a <=( a7989a ) or ( a7984a );
 a7994a <=( a762a ) or ( a763a );
 a7995a <=( a764a ) or ( a7994a );
 a7999a <=( a759a ) or ( a760a );
 a8000a <=( a761a ) or ( a7999a );
 a8001a <=( a8000a ) or ( a7995a );
 a8002a <=( a8001a ) or ( a7990a );
 a8006a <=( a756a ) or ( a757a );
 a8007a <=( a758a ) or ( a8006a );
 a8011a <=( a753a ) or ( a754a );
 a8012a <=( a755a ) or ( a8011a );
 a8013a <=( a8012a ) or ( a8007a );
 a8017a <=( a750a ) or ( a751a );
 a8018a <=( a752a ) or ( a8017a );
 a8021a <=( a748a ) or ( a749a );
 a8024a <=( a746a ) or ( a747a );
 a8025a <=( a8024a ) or ( a8021a );
 a8026a <=( a8025a ) or ( a8018a );
 a8027a <=( a8026a ) or ( a8013a );
 a8028a <=( a8027a ) or ( a8002a );
 a8029a <=( a8028a ) or ( a7979a );
 a8033a <=( a743a ) or ( a744a );
 a8034a <=( a745a ) or ( a8033a );
 a8038a <=( a740a ) or ( a741a );
 a8039a <=( a742a ) or ( a8038a );
 a8040a <=( a8039a ) or ( a8034a );
 a8044a <=( a737a ) or ( a738a );
 a8045a <=( a739a ) or ( a8044a );
 a8049a <=( a734a ) or ( a735a );
 a8050a <=( a736a ) or ( a8049a );
 a8051a <=( a8050a ) or ( a8045a );
 a8052a <=( a8051a ) or ( a8040a );
 a8056a <=( a731a ) or ( a732a );
 a8057a <=( a733a ) or ( a8056a );
 a8061a <=( a728a ) or ( a729a );
 a8062a <=( a730a ) or ( a8061a );
 a8063a <=( a8062a ) or ( a8057a );
 a8067a <=( a725a ) or ( a726a );
 a8068a <=( a727a ) or ( a8067a );
 a8071a <=( a723a ) or ( a724a );
 a8074a <=( a721a ) or ( a722a );
 a8075a <=( a8074a ) or ( a8071a );
 a8076a <=( a8075a ) or ( a8068a );
 a8077a <=( a8076a ) or ( a8063a );
 a8078a <=( a8077a ) or ( a8052a );
 a8082a <=( a718a ) or ( a719a );
 a8083a <=( a720a ) or ( a8082a );
 a8087a <=( a715a ) or ( a716a );
 a8088a <=( a717a ) or ( a8087a );
 a8089a <=( a8088a ) or ( a8083a );
 a8093a <=( a712a ) or ( a713a );
 a8094a <=( a714a ) or ( a8093a );
 a8098a <=( a709a ) or ( a710a );
 a8099a <=( a711a ) or ( a8098a );
 a8100a <=( a8099a ) or ( a8094a );
 a8101a <=( a8100a ) or ( a8089a );
 a8105a <=( a706a ) or ( a707a );
 a8106a <=( a708a ) or ( a8105a );
 a8110a <=( a703a ) or ( a704a );
 a8111a <=( a705a ) or ( a8110a );
 a8112a <=( a8111a ) or ( a8106a );
 a8116a <=( a700a ) or ( a701a );
 a8117a <=( a702a ) or ( a8116a );
 a8120a <=( a698a ) or ( a699a );
 a8123a <=( a696a ) or ( a697a );
 a8124a <=( a8123a ) or ( a8120a );
 a8125a <=( a8124a ) or ( a8117a );
 a8126a <=( a8125a ) or ( a8112a );
 a8127a <=( a8126a ) or ( a8101a );
 a8128a <=( a8127a ) or ( a8078a );
 a8129a <=( a8128a ) or ( a8029a );
 a8133a <=( a693a ) or ( a694a );
 a8134a <=( a695a ) or ( a8133a );
 a8138a <=( a690a ) or ( a691a );
 a8139a <=( a692a ) or ( a8138a );
 a8140a <=( a8139a ) or ( a8134a );
 a8144a <=( a687a ) or ( a688a );
 a8145a <=( a689a ) or ( a8144a );
 a8149a <=( a684a ) or ( a685a );
 a8150a <=( a686a ) or ( a8149a );
 a8151a <=( a8150a ) or ( a8145a );
 a8152a <=( a8151a ) or ( a8140a );
 a8156a <=( a681a ) or ( a682a );
 a8157a <=( a683a ) or ( a8156a );
 a8161a <=( a678a ) or ( a679a );
 a8162a <=( a680a ) or ( a8161a );
 a8163a <=( a8162a ) or ( a8157a );
 a8167a <=( a675a ) or ( a676a );
 a8168a <=( a677a ) or ( a8167a );
 a8172a <=( a672a ) or ( a673a );
 a8173a <=( a674a ) or ( a8172a );
 a8174a <=( a8173a ) or ( a8168a );
 a8175a <=( a8174a ) or ( a8163a );
 a8176a <=( a8175a ) or ( a8152a );
 a8180a <=( a669a ) or ( a670a );
 a8181a <=( a671a ) or ( a8180a );
 a8185a <=( a666a ) or ( a667a );
 a8186a <=( a668a ) or ( a8185a );
 a8187a <=( a8186a ) or ( a8181a );
 a8191a <=( a663a ) or ( a664a );
 a8192a <=( a665a ) or ( a8191a );
 a8196a <=( a660a ) or ( a661a );
 a8197a <=( a662a ) or ( a8196a );
 a8198a <=( a8197a ) or ( a8192a );
 a8199a <=( a8198a ) or ( a8187a );
 a8203a <=( a657a ) or ( a658a );
 a8204a <=( a659a ) or ( a8203a );
 a8208a <=( a654a ) or ( a655a );
 a8209a <=( a656a ) or ( a8208a );
 a8210a <=( a8209a ) or ( a8204a );
 a8214a <=( a651a ) or ( a652a );
 a8215a <=( a653a ) or ( a8214a );
 a8218a <=( a649a ) or ( a650a );
 a8221a <=( a647a ) or ( a648a );
 a8222a <=( a8221a ) or ( a8218a );
 a8223a <=( a8222a ) or ( a8215a );
 a8224a <=( a8223a ) or ( a8210a );
 a8225a <=( a8224a ) or ( a8199a );
 a8226a <=( a8225a ) or ( a8176a );
 a8230a <=( a644a ) or ( a645a );
 a8231a <=( a646a ) or ( a8230a );
 a8235a <=( a641a ) or ( a642a );
 a8236a <=( a643a ) or ( a8235a );
 a8237a <=( a8236a ) or ( a8231a );
 a8241a <=( a638a ) or ( a639a );
 a8242a <=( a640a ) or ( a8241a );
 a8246a <=( a635a ) or ( a636a );
 a8247a <=( a637a ) or ( a8246a );
 a8248a <=( a8247a ) or ( a8242a );
 a8249a <=( a8248a ) or ( a8237a );
 a8253a <=( a632a ) or ( a633a );
 a8254a <=( a634a ) or ( a8253a );
 a8258a <=( a629a ) or ( a630a );
 a8259a <=( a631a ) or ( a8258a );
 a8260a <=( a8259a ) or ( a8254a );
 a8264a <=( a626a ) or ( a627a );
 a8265a <=( a628a ) or ( a8264a );
 a8268a <=( a624a ) or ( a625a );
 a8271a <=( a622a ) or ( a623a );
 a8272a <=( a8271a ) or ( a8268a );
 a8273a <=( a8272a ) or ( a8265a );
 a8274a <=( a8273a ) or ( a8260a );
 a8275a <=( a8274a ) or ( a8249a );
 a8279a <=( a619a ) or ( a620a );
 a8280a <=( a621a ) or ( a8279a );
 a8284a <=( a616a ) or ( a617a );
 a8285a <=( a618a ) or ( a8284a );
 a8286a <=( a8285a ) or ( a8280a );
 a8290a <=( a613a ) or ( a614a );
 a8291a <=( a615a ) or ( a8290a );
 a8295a <=( a610a ) or ( a611a );
 a8296a <=( a612a ) or ( a8295a );
 a8297a <=( a8296a ) or ( a8291a );
 a8298a <=( a8297a ) or ( a8286a );
 a8302a <=( a607a ) or ( a608a );
 a8303a <=( a609a ) or ( a8302a );
 a8307a <=( a604a ) or ( a605a );
 a8308a <=( a606a ) or ( a8307a );
 a8309a <=( a8308a ) or ( a8303a );
 a8313a <=( a601a ) or ( a602a );
 a8314a <=( a603a ) or ( a8313a );
 a8317a <=( a599a ) or ( a600a );
 a8320a <=( a597a ) or ( a598a );
 a8321a <=( a8320a ) or ( a8317a );
 a8322a <=( a8321a ) or ( a8314a );
 a8323a <=( a8322a ) or ( a8309a );
 a8324a <=( a8323a ) or ( a8298a );
 a8325a <=( a8324a ) or ( a8275a );
 a8326a <=( a8325a ) or ( a8226a );
 a8327a <=( a8326a ) or ( a8129a );
 a8331a <=( a594a ) or ( a595a );
 a8332a <=( a596a ) or ( a8331a );
 a8336a <=( a591a ) or ( a592a );
 a8337a <=( a593a ) or ( a8336a );
 a8338a <=( a8337a ) or ( a8332a );
 a8342a <=( a588a ) or ( a589a );
 a8343a <=( a590a ) or ( a8342a );
 a8347a <=( a585a ) or ( a586a );
 a8348a <=( a587a ) or ( a8347a );
 a8349a <=( a8348a ) or ( a8343a );
 a8350a <=( a8349a ) or ( a8338a );
 a8354a <=( a582a ) or ( a583a );
 a8355a <=( a584a ) or ( a8354a );
 a8359a <=( a579a ) or ( a580a );
 a8360a <=( a581a ) or ( a8359a );
 a8361a <=( a8360a ) or ( a8355a );
 a8365a <=( a576a ) or ( a577a );
 a8366a <=( a578a ) or ( a8365a );
 a8370a <=( a573a ) or ( a574a );
 a8371a <=( a575a ) or ( a8370a );
 a8372a <=( a8371a ) or ( a8366a );
 a8373a <=( a8372a ) or ( a8361a );
 a8374a <=( a8373a ) or ( a8350a );
 a8378a <=( a570a ) or ( a571a );
 a8379a <=( a572a ) or ( a8378a );
 a8383a <=( a567a ) or ( a568a );
 a8384a <=( a569a ) or ( a8383a );
 a8385a <=( a8384a ) or ( a8379a );
 a8389a <=( a564a ) or ( a565a );
 a8390a <=( a566a ) or ( a8389a );
 a8394a <=( a561a ) or ( a562a );
 a8395a <=( a563a ) or ( a8394a );
 a8396a <=( a8395a ) or ( a8390a );
 a8397a <=( a8396a ) or ( a8385a );
 a8401a <=( a558a ) or ( a559a );
 a8402a <=( a560a ) or ( a8401a );
 a8406a <=( a555a ) or ( a556a );
 a8407a <=( a557a ) or ( a8406a );
 a8408a <=( a8407a ) or ( a8402a );
 a8412a <=( a552a ) or ( a553a );
 a8413a <=( a554a ) or ( a8412a );
 a8416a <=( a550a ) or ( a551a );
 a8419a <=( a548a ) or ( a549a );
 a8420a <=( a8419a ) or ( a8416a );
 a8421a <=( a8420a ) or ( a8413a );
 a8422a <=( a8421a ) or ( a8408a );
 a8423a <=( a8422a ) or ( a8397a );
 a8424a <=( a8423a ) or ( a8374a );
 a8428a <=( a545a ) or ( a546a );
 a8429a <=( a547a ) or ( a8428a );
 a8433a <=( a542a ) or ( a543a );
 a8434a <=( a544a ) or ( a8433a );
 a8435a <=( a8434a ) or ( a8429a );
 a8439a <=( a539a ) or ( a540a );
 a8440a <=( a541a ) or ( a8439a );
 a8444a <=( a536a ) or ( a537a );
 a8445a <=( a538a ) or ( a8444a );
 a8446a <=( a8445a ) or ( a8440a );
 a8447a <=( a8446a ) or ( a8435a );
 a8451a <=( a533a ) or ( a534a );
 a8452a <=( a535a ) or ( a8451a );
 a8456a <=( a530a ) or ( a531a );
 a8457a <=( a532a ) or ( a8456a );
 a8458a <=( a8457a ) or ( a8452a );
 a8462a <=( a527a ) or ( a528a );
 a8463a <=( a529a ) or ( a8462a );
 a8466a <=( a525a ) or ( a526a );
 a8469a <=( a523a ) or ( a524a );
 a8470a <=( a8469a ) or ( a8466a );
 a8471a <=( a8470a ) or ( a8463a );
 a8472a <=( a8471a ) or ( a8458a );
 a8473a <=( a8472a ) or ( a8447a );
 a8477a <=( a520a ) or ( a521a );
 a8478a <=( a522a ) or ( a8477a );
 a8482a <=( a517a ) or ( a518a );
 a8483a <=( a519a ) or ( a8482a );
 a8484a <=( a8483a ) or ( a8478a );
 a8488a <=( a514a ) or ( a515a );
 a8489a <=( a516a ) or ( a8488a );
 a8493a <=( a511a ) or ( a512a );
 a8494a <=( a513a ) or ( a8493a );
 a8495a <=( a8494a ) or ( a8489a );
 a8496a <=( a8495a ) or ( a8484a );
 a8500a <=( a508a ) or ( a509a );
 a8501a <=( a510a ) or ( a8500a );
 a8505a <=( a505a ) or ( a506a );
 a8506a <=( a507a ) or ( a8505a );
 a8507a <=( a8506a ) or ( a8501a );
 a8511a <=( a502a ) or ( a503a );
 a8512a <=( a504a ) or ( a8511a );
 a8515a <=( a500a ) or ( a501a );
 a8518a <=( a498a ) or ( a499a );
 a8519a <=( a8518a ) or ( a8515a );
 a8520a <=( a8519a ) or ( a8512a );
 a8521a <=( a8520a ) or ( a8507a );
 a8522a <=( a8521a ) or ( a8496a );
 a8523a <=( a8522a ) or ( a8473a );
 a8524a <=( a8523a ) or ( a8424a );
 a8528a <=( a495a ) or ( a496a );
 a8529a <=( a497a ) or ( a8528a );
 a8533a <=( a492a ) or ( a493a );
 a8534a <=( a494a ) or ( a8533a );
 a8535a <=( a8534a ) or ( a8529a );
 a8539a <=( a489a ) or ( a490a );
 a8540a <=( a491a ) or ( a8539a );
 a8544a <=( a486a ) or ( a487a );
 a8545a <=( a488a ) or ( a8544a );
 a8546a <=( a8545a ) or ( a8540a );
 a8547a <=( a8546a ) or ( a8535a );
 a8551a <=( a483a ) or ( a484a );
 a8552a <=( a485a ) or ( a8551a );
 a8556a <=( a480a ) or ( a481a );
 a8557a <=( a482a ) or ( a8556a );
 a8558a <=( a8557a ) or ( a8552a );
 a8562a <=( a477a ) or ( a478a );
 a8563a <=( a479a ) or ( a8562a );
 a8566a <=( a475a ) or ( a476a );
 a8569a <=( a473a ) or ( a474a );
 a8570a <=( a8569a ) or ( a8566a );
 a8571a <=( a8570a ) or ( a8563a );
 a8572a <=( a8571a ) or ( a8558a );
 a8573a <=( a8572a ) or ( a8547a );
 a8577a <=( a470a ) or ( a471a );
 a8578a <=( a472a ) or ( a8577a );
 a8582a <=( a467a ) or ( a468a );
 a8583a <=( a469a ) or ( a8582a );
 a8584a <=( a8583a ) or ( a8578a );
 a8588a <=( a464a ) or ( a465a );
 a8589a <=( a466a ) or ( a8588a );
 a8593a <=( a461a ) or ( a462a );
 a8594a <=( a463a ) or ( a8593a );
 a8595a <=( a8594a ) or ( a8589a );
 a8596a <=( a8595a ) or ( a8584a );
 a8600a <=( a458a ) or ( a459a );
 a8601a <=( a460a ) or ( a8600a );
 a8605a <=( a455a ) or ( a456a );
 a8606a <=( a457a ) or ( a8605a );
 a8607a <=( a8606a ) or ( a8601a );
 a8611a <=( a452a ) or ( a453a );
 a8612a <=( a454a ) or ( a8611a );
 a8615a <=( a450a ) or ( a451a );
 a8618a <=( a448a ) or ( a449a );
 a8619a <=( a8618a ) or ( a8615a );
 a8620a <=( a8619a ) or ( a8612a );
 a8621a <=( a8620a ) or ( a8607a );
 a8622a <=( a8621a ) or ( a8596a );
 a8623a <=( a8622a ) or ( a8573a );
 a8627a <=( a445a ) or ( a446a );
 a8628a <=( a447a ) or ( a8627a );
 a8632a <=( a442a ) or ( a443a );
 a8633a <=( a444a ) or ( a8632a );
 a8634a <=( a8633a ) or ( a8628a );
 a8638a <=( a439a ) or ( a440a );
 a8639a <=( a441a ) or ( a8638a );
 a8643a <=( a436a ) or ( a437a );
 a8644a <=( a438a ) or ( a8643a );
 a8645a <=( a8644a ) or ( a8639a );
 a8646a <=( a8645a ) or ( a8634a );
 a8650a <=( a433a ) or ( a434a );
 a8651a <=( a435a ) or ( a8650a );
 a8655a <=( a430a ) or ( a431a );
 a8656a <=( a432a ) or ( a8655a );
 a8657a <=( a8656a ) or ( a8651a );
 a8661a <=( a427a ) or ( a428a );
 a8662a <=( a429a ) or ( a8661a );
 a8665a <=( a425a ) or ( a426a );
 a8668a <=( a423a ) or ( a424a );
 a8669a <=( a8668a ) or ( a8665a );
 a8670a <=( a8669a ) or ( a8662a );
 a8671a <=( a8670a ) or ( a8657a );
 a8672a <=( a8671a ) or ( a8646a );
 a8676a <=( a420a ) or ( a421a );
 a8677a <=( a422a ) or ( a8676a );
 a8681a <=( a417a ) or ( a418a );
 a8682a <=( a419a ) or ( a8681a );
 a8683a <=( a8682a ) or ( a8677a );
 a8687a <=( a414a ) or ( a415a );
 a8688a <=( a416a ) or ( a8687a );
 a8692a <=( a411a ) or ( a412a );
 a8693a <=( a413a ) or ( a8692a );
 a8694a <=( a8693a ) or ( a8688a );
 a8695a <=( a8694a ) or ( a8683a );
 a8699a <=( a408a ) or ( a409a );
 a8700a <=( a410a ) or ( a8699a );
 a8704a <=( a405a ) or ( a406a );
 a8705a <=( a407a ) or ( a8704a );
 a8706a <=( a8705a ) or ( a8700a );
 a8710a <=( a402a ) or ( a403a );
 a8711a <=( a404a ) or ( a8710a );
 a8714a <=( a400a ) or ( a401a );
 a8717a <=( a398a ) or ( a399a );
 a8718a <=( a8717a ) or ( a8714a );
 a8719a <=( a8718a ) or ( a8711a );
 a8720a <=( a8719a ) or ( a8706a );
 a8721a <=( a8720a ) or ( a8695a );
 a8722a <=( a8721a ) or ( a8672a );
 a8723a <=( a8722a ) or ( a8623a );
 a8724a <=( a8723a ) or ( a8524a );
 a8725a <=( a8724a ) or ( a8327a );
 a8729a <=( a395a ) or ( a396a );
 a8730a <=( a397a ) or ( a8729a );
 a8734a <=( a392a ) or ( a393a );
 a8735a <=( a394a ) or ( a8734a );
 a8736a <=( a8735a ) or ( a8730a );
 a8740a <=( a389a ) or ( a390a );
 a8741a <=( a391a ) or ( a8740a );
 a8745a <=( a386a ) or ( a387a );
 a8746a <=( a388a ) or ( a8745a );
 a8747a <=( a8746a ) or ( a8741a );
 a8748a <=( a8747a ) or ( a8736a );
 a8752a <=( a383a ) or ( a384a );
 a8753a <=( a385a ) or ( a8752a );
 a8757a <=( a380a ) or ( a381a );
 a8758a <=( a382a ) or ( a8757a );
 a8759a <=( a8758a ) or ( a8753a );
 a8763a <=( a377a ) or ( a378a );
 a8764a <=( a379a ) or ( a8763a );
 a8768a <=( a374a ) or ( a375a );
 a8769a <=( a376a ) or ( a8768a );
 a8770a <=( a8769a ) or ( a8764a );
 a8771a <=( a8770a ) or ( a8759a );
 a8772a <=( a8771a ) or ( a8748a );
 a8776a <=( a371a ) or ( a372a );
 a8777a <=( a373a ) or ( a8776a );
 a8781a <=( a368a ) or ( a369a );
 a8782a <=( a370a ) or ( a8781a );
 a8783a <=( a8782a ) or ( a8777a );
 a8787a <=( a365a ) or ( a366a );
 a8788a <=( a367a ) or ( a8787a );
 a8792a <=( a362a ) or ( a363a );
 a8793a <=( a364a ) or ( a8792a );
 a8794a <=( a8793a ) or ( a8788a );
 a8795a <=( a8794a ) or ( a8783a );
 a8799a <=( a359a ) or ( a360a );
 a8800a <=( a361a ) or ( a8799a );
 a8804a <=( a356a ) or ( a357a );
 a8805a <=( a358a ) or ( a8804a );
 a8806a <=( a8805a ) or ( a8800a );
 a8810a <=( a353a ) or ( a354a );
 a8811a <=( a355a ) or ( a8810a );
 a8814a <=( a351a ) or ( a352a );
 a8817a <=( a349a ) or ( a350a );
 a8818a <=( a8817a ) or ( a8814a );
 a8819a <=( a8818a ) or ( a8811a );
 a8820a <=( a8819a ) or ( a8806a );
 a8821a <=( a8820a ) or ( a8795a );
 a8822a <=( a8821a ) or ( a8772a );
 a8826a <=( a346a ) or ( a347a );
 a8827a <=( a348a ) or ( a8826a );
 a8831a <=( a343a ) or ( a344a );
 a8832a <=( a345a ) or ( a8831a );
 a8833a <=( a8832a ) or ( a8827a );
 a8837a <=( a340a ) or ( a341a );
 a8838a <=( a342a ) or ( a8837a );
 a8842a <=( a337a ) or ( a338a );
 a8843a <=( a339a ) or ( a8842a );
 a8844a <=( a8843a ) or ( a8838a );
 a8845a <=( a8844a ) or ( a8833a );
 a8849a <=( a334a ) or ( a335a );
 a8850a <=( a336a ) or ( a8849a );
 a8854a <=( a331a ) or ( a332a );
 a8855a <=( a333a ) or ( a8854a );
 a8856a <=( a8855a ) or ( a8850a );
 a8860a <=( a328a ) or ( a329a );
 a8861a <=( a330a ) or ( a8860a );
 a8864a <=( a326a ) or ( a327a );
 a8867a <=( a324a ) or ( a325a );
 a8868a <=( a8867a ) or ( a8864a );
 a8869a <=( a8868a ) or ( a8861a );
 a8870a <=( a8869a ) or ( a8856a );
 a8871a <=( a8870a ) or ( a8845a );
 a8875a <=( a321a ) or ( a322a );
 a8876a <=( a323a ) or ( a8875a );
 a8880a <=( a318a ) or ( a319a );
 a8881a <=( a320a ) or ( a8880a );
 a8882a <=( a8881a ) or ( a8876a );
 a8886a <=( a315a ) or ( a316a );
 a8887a <=( a317a ) or ( a8886a );
 a8891a <=( a312a ) or ( a313a );
 a8892a <=( a314a ) or ( a8891a );
 a8893a <=( a8892a ) or ( a8887a );
 a8894a <=( a8893a ) or ( a8882a );
 a8898a <=( a309a ) or ( a310a );
 a8899a <=( a311a ) or ( a8898a );
 a8903a <=( a306a ) or ( a307a );
 a8904a <=( a308a ) or ( a8903a );
 a8905a <=( a8904a ) or ( a8899a );
 a8909a <=( a303a ) or ( a304a );
 a8910a <=( a305a ) or ( a8909a );
 a8913a <=( a301a ) or ( a302a );
 a8916a <=( a299a ) or ( a300a );
 a8917a <=( a8916a ) or ( a8913a );
 a8918a <=( a8917a ) or ( a8910a );
 a8919a <=( a8918a ) or ( a8905a );
 a8920a <=( a8919a ) or ( a8894a );
 a8921a <=( a8920a ) or ( a8871a );
 a8922a <=( a8921a ) or ( a8822a );
 a8926a <=( a296a ) or ( a297a );
 a8927a <=( a298a ) or ( a8926a );
 a8931a <=( a293a ) or ( a294a );
 a8932a <=( a295a ) or ( a8931a );
 a8933a <=( a8932a ) or ( a8927a );
 a8937a <=( a290a ) or ( a291a );
 a8938a <=( a292a ) or ( a8937a );
 a8942a <=( a287a ) or ( a288a );
 a8943a <=( a289a ) or ( a8942a );
 a8944a <=( a8943a ) or ( a8938a );
 a8945a <=( a8944a ) or ( a8933a );
 a8949a <=( a284a ) or ( a285a );
 a8950a <=( a286a ) or ( a8949a );
 a8954a <=( a281a ) or ( a282a );
 a8955a <=( a283a ) or ( a8954a );
 a8956a <=( a8955a ) or ( a8950a );
 a8960a <=( a278a ) or ( a279a );
 a8961a <=( a280a ) or ( a8960a );
 a8965a <=( a275a ) or ( a276a );
 a8966a <=( a277a ) or ( a8965a );
 a8967a <=( a8966a ) or ( a8961a );
 a8968a <=( a8967a ) or ( a8956a );
 a8969a <=( a8968a ) or ( a8945a );
 a8973a <=( a272a ) or ( a273a );
 a8974a <=( a274a ) or ( a8973a );
 a8978a <=( a269a ) or ( a270a );
 a8979a <=( a271a ) or ( a8978a );
 a8980a <=( a8979a ) or ( a8974a );
 a8984a <=( a266a ) or ( a267a );
 a8985a <=( a268a ) or ( a8984a );
 a8989a <=( a263a ) or ( a264a );
 a8990a <=( a265a ) or ( a8989a );
 a8991a <=( a8990a ) or ( a8985a );
 a8992a <=( a8991a ) or ( a8980a );
 a8996a <=( a260a ) or ( a261a );
 a8997a <=( a262a ) or ( a8996a );
 a9001a <=( a257a ) or ( a258a );
 a9002a <=( a259a ) or ( a9001a );
 a9003a <=( a9002a ) or ( a8997a );
 a9007a <=( a254a ) or ( a255a );
 a9008a <=( a256a ) or ( a9007a );
 a9011a <=( a252a ) or ( a253a );
 a9014a <=( a250a ) or ( a251a );
 a9015a <=( a9014a ) or ( a9011a );
 a9016a <=( a9015a ) or ( a9008a );
 a9017a <=( a9016a ) or ( a9003a );
 a9018a <=( a9017a ) or ( a8992a );
 a9019a <=( a9018a ) or ( a8969a );
 a9023a <=( a247a ) or ( a248a );
 a9024a <=( a249a ) or ( a9023a );
 a9028a <=( a244a ) or ( a245a );
 a9029a <=( a246a ) or ( a9028a );
 a9030a <=( a9029a ) or ( a9024a );
 a9034a <=( a241a ) or ( a242a );
 a9035a <=( a243a ) or ( a9034a );
 a9039a <=( a238a ) or ( a239a );
 a9040a <=( a240a ) or ( a9039a );
 a9041a <=( a9040a ) or ( a9035a );
 a9042a <=( a9041a ) or ( a9030a );
 a9046a <=( a235a ) or ( a236a );
 a9047a <=( a237a ) or ( a9046a );
 a9051a <=( a232a ) or ( a233a );
 a9052a <=( a234a ) or ( a9051a );
 a9053a <=( a9052a ) or ( a9047a );
 a9057a <=( a229a ) or ( a230a );
 a9058a <=( a231a ) or ( a9057a );
 a9061a <=( a227a ) or ( a228a );
 a9064a <=( a225a ) or ( a226a );
 a9065a <=( a9064a ) or ( a9061a );
 a9066a <=( a9065a ) or ( a9058a );
 a9067a <=( a9066a ) or ( a9053a );
 a9068a <=( a9067a ) or ( a9042a );
 a9072a <=( a222a ) or ( a223a );
 a9073a <=( a224a ) or ( a9072a );
 a9077a <=( a219a ) or ( a220a );
 a9078a <=( a221a ) or ( a9077a );
 a9079a <=( a9078a ) or ( a9073a );
 a9083a <=( a216a ) or ( a217a );
 a9084a <=( a218a ) or ( a9083a );
 a9088a <=( a213a ) or ( a214a );
 a9089a <=( a215a ) or ( a9088a );
 a9090a <=( a9089a ) or ( a9084a );
 a9091a <=( a9090a ) or ( a9079a );
 a9095a <=( a210a ) or ( a211a );
 a9096a <=( a212a ) or ( a9095a );
 a9100a <=( a207a ) or ( a208a );
 a9101a <=( a209a ) or ( a9100a );
 a9102a <=( a9101a ) or ( a9096a );
 a9106a <=( a204a ) or ( a205a );
 a9107a <=( a206a ) or ( a9106a );
 a9110a <=( a202a ) or ( a203a );
 a9113a <=( a200a ) or ( a201a );
 a9114a <=( a9113a ) or ( a9110a );
 a9115a <=( a9114a ) or ( a9107a );
 a9116a <=( a9115a ) or ( a9102a );
 a9117a <=( a9116a ) or ( a9091a );
 a9118a <=( a9117a ) or ( a9068a );
 a9119a <=( a9118a ) or ( a9019a );
 a9120a <=( a9119a ) or ( a8922a );
 a9124a <=( a197a ) or ( a198a );
 a9125a <=( a199a ) or ( a9124a );
 a9129a <=( a194a ) or ( a195a );
 a9130a <=( a196a ) or ( a9129a );
 a9131a <=( a9130a ) or ( a9125a );
 a9135a <=( a191a ) or ( a192a );
 a9136a <=( a193a ) or ( a9135a );
 a9140a <=( a188a ) or ( a189a );
 a9141a <=( a190a ) or ( a9140a );
 a9142a <=( a9141a ) or ( a9136a );
 a9143a <=( a9142a ) or ( a9131a );
 a9147a <=( a185a ) or ( a186a );
 a9148a <=( a187a ) or ( a9147a );
 a9152a <=( a182a ) or ( a183a );
 a9153a <=( a184a ) or ( a9152a );
 a9154a <=( a9153a ) or ( a9148a );
 a9158a <=( a179a ) or ( a180a );
 a9159a <=( a181a ) or ( a9158a );
 a9163a <=( a176a ) or ( a177a );
 a9164a <=( a178a ) or ( a9163a );
 a9165a <=( a9164a ) or ( a9159a );
 a9166a <=( a9165a ) or ( a9154a );
 a9167a <=( a9166a ) or ( a9143a );
 a9171a <=( a173a ) or ( a174a );
 a9172a <=( a175a ) or ( a9171a );
 a9176a <=( a170a ) or ( a171a );
 a9177a <=( a172a ) or ( a9176a );
 a9178a <=( a9177a ) or ( a9172a );
 a9182a <=( a167a ) or ( a168a );
 a9183a <=( a169a ) or ( a9182a );
 a9187a <=( a164a ) or ( a165a );
 a9188a <=( a166a ) or ( a9187a );
 a9189a <=( a9188a ) or ( a9183a );
 a9190a <=( a9189a ) or ( a9178a );
 a9194a <=( a161a ) or ( a162a );
 a9195a <=( a163a ) or ( a9194a );
 a9199a <=( a158a ) or ( a159a );
 a9200a <=( a160a ) or ( a9199a );
 a9201a <=( a9200a ) or ( a9195a );
 a9205a <=( a155a ) or ( a156a );
 a9206a <=( a157a ) or ( a9205a );
 a9209a <=( a153a ) or ( a154a );
 a9212a <=( a151a ) or ( a152a );
 a9213a <=( a9212a ) or ( a9209a );
 a9214a <=( a9213a ) or ( a9206a );
 a9215a <=( a9214a ) or ( a9201a );
 a9216a <=( a9215a ) or ( a9190a );
 a9217a <=( a9216a ) or ( a9167a );
 a9221a <=( a148a ) or ( a149a );
 a9222a <=( a150a ) or ( a9221a );
 a9226a <=( a145a ) or ( a146a );
 a9227a <=( a147a ) or ( a9226a );
 a9228a <=( a9227a ) or ( a9222a );
 a9232a <=( a142a ) or ( a143a );
 a9233a <=( a144a ) or ( a9232a );
 a9237a <=( a139a ) or ( a140a );
 a9238a <=( a141a ) or ( a9237a );
 a9239a <=( a9238a ) or ( a9233a );
 a9240a <=( a9239a ) or ( a9228a );
 a9244a <=( a136a ) or ( a137a );
 a9245a <=( a138a ) or ( a9244a );
 a9249a <=( a133a ) or ( a134a );
 a9250a <=( a135a ) or ( a9249a );
 a9251a <=( a9250a ) or ( a9245a );
 a9255a <=( a130a ) or ( a131a );
 a9256a <=( a132a ) or ( a9255a );
 a9259a <=( a128a ) or ( a129a );
 a9262a <=( a126a ) or ( a127a );
 a9263a <=( a9262a ) or ( a9259a );
 a9264a <=( a9263a ) or ( a9256a );
 a9265a <=( a9264a ) or ( a9251a );
 a9266a <=( a9265a ) or ( a9240a );
 a9270a <=( a123a ) or ( a124a );
 a9271a <=( a125a ) or ( a9270a );
 a9275a <=( a120a ) or ( a121a );
 a9276a <=( a122a ) or ( a9275a );
 a9277a <=( a9276a ) or ( a9271a );
 a9281a <=( a117a ) or ( a118a );
 a9282a <=( a119a ) or ( a9281a );
 a9286a <=( a114a ) or ( a115a );
 a9287a <=( a116a ) or ( a9286a );
 a9288a <=( a9287a ) or ( a9282a );
 a9289a <=( a9288a ) or ( a9277a );
 a9293a <=( a111a ) or ( a112a );
 a9294a <=( a113a ) or ( a9293a );
 a9298a <=( a108a ) or ( a109a );
 a9299a <=( a110a ) or ( a9298a );
 a9300a <=( a9299a ) or ( a9294a );
 a9304a <=( a105a ) or ( a106a );
 a9305a <=( a107a ) or ( a9304a );
 a9308a <=( a103a ) or ( a104a );
 a9311a <=( a101a ) or ( a102a );
 a9312a <=( a9311a ) or ( a9308a );
 a9313a <=( a9312a ) or ( a9305a );
 a9314a <=( a9313a ) or ( a9300a );
 a9315a <=( a9314a ) or ( a9289a );
 a9316a <=( a9315a ) or ( a9266a );
 a9317a <=( a9316a ) or ( a9217a );
 a9321a <=( a98a ) or ( a99a );
 a9322a <=( a100a ) or ( a9321a );
 a9326a <=( a95a ) or ( a96a );
 a9327a <=( a97a ) or ( a9326a );
 a9328a <=( a9327a ) or ( a9322a );
 a9332a <=( a92a ) or ( a93a );
 a9333a <=( a94a ) or ( a9332a );
 a9337a <=( a89a ) or ( a90a );
 a9338a <=( a91a ) or ( a9337a );
 a9339a <=( a9338a ) or ( a9333a );
 a9340a <=( a9339a ) or ( a9328a );
 a9344a <=( a86a ) or ( a87a );
 a9345a <=( a88a ) or ( a9344a );
 a9349a <=( a83a ) or ( a84a );
 a9350a <=( a85a ) or ( a9349a );
 a9351a <=( a9350a ) or ( a9345a );
 a9355a <=( a80a ) or ( a81a );
 a9356a <=( a82a ) or ( a9355a );
 a9359a <=( a78a ) or ( a79a );
 a9362a <=( a76a ) or ( a77a );
 a9363a <=( a9362a ) or ( a9359a );
 a9364a <=( a9363a ) or ( a9356a );
 a9365a <=( a9364a ) or ( a9351a );
 a9366a <=( a9365a ) or ( a9340a );
 a9370a <=( a73a ) or ( a74a );
 a9371a <=( a75a ) or ( a9370a );
 a9375a <=( a70a ) or ( a71a );
 a9376a <=( a72a ) or ( a9375a );
 a9377a <=( a9376a ) or ( a9371a );
 a9381a <=( a67a ) or ( a68a );
 a9382a <=( a69a ) or ( a9381a );
 a9386a <=( a64a ) or ( a65a );
 a9387a <=( a66a ) or ( a9386a );
 a9388a <=( a9387a ) or ( a9382a );
 a9389a <=( a9388a ) or ( a9377a );
 a9393a <=( a61a ) or ( a62a );
 a9394a <=( a63a ) or ( a9393a );
 a9398a <=( a58a ) or ( a59a );
 a9399a <=( a60a ) or ( a9398a );
 a9400a <=( a9399a ) or ( a9394a );
 a9404a <=( a55a ) or ( a56a );
 a9405a <=( a57a ) or ( a9404a );
 a9408a <=( a53a ) or ( a54a );
 a9411a <=( a51a ) or ( a52a );
 a9412a <=( a9411a ) or ( a9408a );
 a9413a <=( a9412a ) or ( a9405a );
 a9414a <=( a9413a ) or ( a9400a );
 a9415a <=( a9414a ) or ( a9389a );
 a9416a <=( a9415a ) or ( a9366a );
 a9420a <=( a48a ) or ( a49a );
 a9421a <=( a50a ) or ( a9420a );
 a9425a <=( a45a ) or ( a46a );
 a9426a <=( a47a ) or ( a9425a );
 a9427a <=( a9426a ) or ( a9421a );
 a9431a <=( a42a ) or ( a43a );
 a9432a <=( a44a ) or ( a9431a );
 a9436a <=( a39a ) or ( a40a );
 a9437a <=( a41a ) or ( a9436a );
 a9438a <=( a9437a ) or ( a9432a );
 a9439a <=( a9438a ) or ( a9427a );
 a9443a <=( a36a ) or ( a37a );
 a9444a <=( a38a ) or ( a9443a );
 a9448a <=( a33a ) or ( a34a );
 a9449a <=( a35a ) or ( a9448a );
 a9450a <=( a9449a ) or ( a9444a );
 a9454a <=( a30a ) or ( a31a );
 a9455a <=( a32a ) or ( a9454a );
 a9458a <=( a28a ) or ( a29a );
 a9461a <=( a26a ) or ( a27a );
 a9462a <=( a9461a ) or ( a9458a );
 a9463a <=( a9462a ) or ( a9455a );
 a9464a <=( a9463a ) or ( a9450a );
 a9465a <=( a9464a ) or ( a9439a );
 a9469a <=( a23a ) or ( a24a );
 a9470a <=( a25a ) or ( a9469a );
 a9474a <=( a20a ) or ( a21a );
 a9475a <=( a22a ) or ( a9474a );
 a9476a <=( a9475a ) or ( a9470a );
 a9480a <=( a17a ) or ( a18a );
 a9481a <=( a19a ) or ( a9480a );
 a9485a <=( a14a ) or ( a15a );
 a9486a <=( a16a ) or ( a9485a );
 a9487a <=( a9486a ) or ( a9481a );
 a9488a <=( a9487a ) or ( a9476a );
 a9492a <=( a11a ) or ( a12a );
 a9493a <=( a13a ) or ( a9492a );
 a9497a <=( a8a ) or ( a9a );
 a9498a <=( a10a ) or ( a9497a );
 a9499a <=( a9498a ) or ( a9493a );
 a9503a <=( a5a ) or ( a6a );
 a9504a <=( a7a ) or ( a9503a );
 a9507a <=( a3a ) or ( a4a );
 a9510a <=( a1a ) or ( a2a );
 a9511a <=( a9510a ) or ( a9507a );
 a9512a <=( a9511a ) or ( a9504a );
 a9513a <=( a9512a ) or ( a9499a );
 a9514a <=( a9513a ) or ( a9488a );
 a9515a <=( a9514a ) or ( a9465a );
 a9516a <=( a9515a ) or ( a9416a );
 a9517a <=( a9516a ) or ( a9317a );
 a9518a <=( a9517a ) or ( a9120a );
 a9519a <=( a9518a ) or ( a8725a );
 a9520a <=( a9519a ) or ( a7932a );
 a9523a <=( A166  and  A168 );
 a9526a <=( A200  and  A199 );
 a9527a <=( a9526a  and  a9523a );
 a9530a <=( A233  and  (not A232) );
 a9533a <=( (not A300)  and  (not A299) );
 a9534a <=( a9533a  and  a9530a );
 a9537a <=( A166  and  A168 );
 a9540a <=( A200  and  A199 );
 a9541a <=( a9540a  and  a9537a );
 a9544a <=( A233  and  (not A232) );
 a9547a <=( A299  and  A298 );
 a9548a <=( a9547a  and  a9544a );
 a9551a <=( A166  and  A168 );
 a9554a <=( A200  and  A199 );
 a9555a <=( a9554a  and  a9551a );
 a9558a <=( A233  and  (not A232) );
 a9561a <=( (not A299)  and  (not A298) );
 a9562a <=( a9561a  and  a9558a );
 a9565a <=( A166  and  A168 );
 a9568a <=( A200  and  A199 );
 a9569a <=( a9568a  and  a9565a );
 a9572a <=( A233  and  (not A232) );
 a9575a <=( A266  and  (not A265) );
 a9576a <=( a9575a  and  a9572a );
 a9579a <=( A166  and  A168 );
 a9582a <=( (not A201)  and  (not A200) );
 a9583a <=( a9582a  and  a9579a );
 a9586a <=( A233  and  (not A232) );
 a9589a <=( (not A300)  and  (not A299) );
 a9590a <=( a9589a  and  a9586a );
 a9593a <=( A166  and  A168 );
 a9596a <=( (not A201)  and  (not A200) );
 a9597a <=( a9596a  and  a9593a );
 a9600a <=( A233  and  (not A232) );
 a9603a <=( A299  and  A298 );
 a9604a <=( a9603a  and  a9600a );
 a9607a <=( A166  and  A168 );
 a9610a <=( (not A201)  and  (not A200) );
 a9611a <=( a9610a  and  a9607a );
 a9614a <=( A233  and  (not A232) );
 a9617a <=( (not A299)  and  (not A298) );
 a9618a <=( a9617a  and  a9614a );
 a9621a <=( A166  and  A168 );
 a9624a <=( (not A201)  and  (not A200) );
 a9625a <=( a9624a  and  a9621a );
 a9628a <=( A233  and  (not A232) );
 a9631a <=( A266  and  (not A265) );
 a9632a <=( a9631a  and  a9628a );
 a9635a <=( A166  and  A168 );
 a9638a <=( (not A200)  and  (not A199) );
 a9639a <=( a9638a  and  a9635a );
 a9642a <=( A233  and  (not A232) );
 a9645a <=( (not A300)  and  (not A299) );
 a9646a <=( a9645a  and  a9642a );
 a9649a <=( A166  and  A168 );
 a9652a <=( (not A200)  and  (not A199) );
 a9653a <=( a9652a  and  a9649a );
 a9656a <=( A233  and  (not A232) );
 a9659a <=( A299  and  A298 );
 a9660a <=( a9659a  and  a9656a );
 a9663a <=( A166  and  A168 );
 a9666a <=( (not A200)  and  (not A199) );
 a9667a <=( a9666a  and  a9663a );
 a9670a <=( A233  and  (not A232) );
 a9673a <=( (not A299)  and  (not A298) );
 a9674a <=( a9673a  and  a9670a );
 a9677a <=( A166  and  A168 );
 a9680a <=( (not A200)  and  (not A199) );
 a9681a <=( a9680a  and  a9677a );
 a9684a <=( A233  and  (not A232) );
 a9687a <=( A266  and  (not A265) );
 a9688a <=( a9687a  and  a9684a );
 a9691a <=( A167  and  A168 );
 a9694a <=( A200  and  A199 );
 a9695a <=( a9694a  and  a9691a );
 a9698a <=( A233  and  (not A232) );
 a9701a <=( (not A300)  and  (not A299) );
 a9702a <=( a9701a  and  a9698a );
 a9705a <=( A167  and  A168 );
 a9708a <=( A200  and  A199 );
 a9709a <=( a9708a  and  a9705a );
 a9712a <=( A233  and  (not A232) );
 a9715a <=( A299  and  A298 );
 a9716a <=( a9715a  and  a9712a );
 a9719a <=( A167  and  A168 );
 a9722a <=( A200  and  A199 );
 a9723a <=( a9722a  and  a9719a );
 a9726a <=( A233  and  (not A232) );
 a9729a <=( (not A299)  and  (not A298) );
 a9730a <=( a9729a  and  a9726a );
 a9733a <=( A167  and  A168 );
 a9736a <=( A200  and  A199 );
 a9737a <=( a9736a  and  a9733a );
 a9740a <=( A233  and  (not A232) );
 a9743a <=( A266  and  (not A265) );
 a9744a <=( a9743a  and  a9740a );
 a9747a <=( A167  and  A168 );
 a9750a <=( (not A201)  and  (not A200) );
 a9751a <=( a9750a  and  a9747a );
 a9754a <=( A233  and  (not A232) );
 a9757a <=( (not A300)  and  (not A299) );
 a9758a <=( a9757a  and  a9754a );
 a9761a <=( A167  and  A168 );
 a9764a <=( (not A201)  and  (not A200) );
 a9765a <=( a9764a  and  a9761a );
 a9768a <=( A233  and  (not A232) );
 a9771a <=( A299  and  A298 );
 a9772a <=( a9771a  and  a9768a );
 a9775a <=( A167  and  A168 );
 a9778a <=( (not A201)  and  (not A200) );
 a9779a <=( a9778a  and  a9775a );
 a9782a <=( A233  and  (not A232) );
 a9785a <=( (not A299)  and  (not A298) );
 a9786a <=( a9785a  and  a9782a );
 a9789a <=( A167  and  A168 );
 a9792a <=( (not A201)  and  (not A200) );
 a9793a <=( a9792a  and  a9789a );
 a9796a <=( A233  and  (not A232) );
 a9799a <=( A266  and  (not A265) );
 a9800a <=( a9799a  and  a9796a );
 a9803a <=( A167  and  A168 );
 a9806a <=( (not A200)  and  (not A199) );
 a9807a <=( a9806a  and  a9803a );
 a9810a <=( A233  and  (not A232) );
 a9813a <=( (not A300)  and  (not A299) );
 a9814a <=( a9813a  and  a9810a );
 a9817a <=( A167  and  A168 );
 a9820a <=( (not A200)  and  (not A199) );
 a9821a <=( a9820a  and  a9817a );
 a9824a <=( A233  and  (not A232) );
 a9827a <=( A299  and  A298 );
 a9828a <=( a9827a  and  a9824a );
 a9831a <=( A167  and  A168 );
 a9834a <=( (not A200)  and  (not A199) );
 a9835a <=( a9834a  and  a9831a );
 a9838a <=( A233  and  (not A232) );
 a9841a <=( (not A299)  and  (not A298) );
 a9842a <=( a9841a  and  a9838a );
 a9845a <=( A167  and  A168 );
 a9848a <=( (not A200)  and  (not A199) );
 a9849a <=( a9848a  and  a9845a );
 a9852a <=( A233  and  (not A232) );
 a9855a <=( A266  and  (not A265) );
 a9856a <=( a9855a  and  a9852a );
 a9859a <=( A166  and  A168 );
 a9862a <=( A200  and  A199 );
 a9863a <=( a9862a  and  a9859a );
 a9866a <=( A233  and  (not A232) );
 a9870a <=( (not A302)  and  (not A301) );
 a9871a <=( (not A299)  and  a9870a );
 a9872a <=( a9871a  and  a9866a );
 a9875a <=( A166  and  A168 );
 a9878a <=( (not A202)  and  (not A200) );
 a9879a <=( a9878a  and  a9875a );
 a9882a <=( (not A232)  and  (not A203) );
 a9886a <=( (not A300)  and  (not A299) );
 a9887a <=( A233  and  a9886a );
 a9888a <=( a9887a  and  a9882a );
 a9891a <=( A166  and  A168 );
 a9894a <=( (not A202)  and  (not A200) );
 a9895a <=( a9894a  and  a9891a );
 a9898a <=( (not A232)  and  (not A203) );
 a9902a <=( A299  and  A298 );
 a9903a <=( A233  and  a9902a );
 a9904a <=( a9903a  and  a9898a );
 a9907a <=( A166  and  A168 );
 a9910a <=( (not A202)  and  (not A200) );
 a9911a <=( a9910a  and  a9907a );
 a9914a <=( (not A232)  and  (not A203) );
 a9918a <=( (not A299)  and  (not A298) );
 a9919a <=( A233  and  a9918a );
 a9920a <=( a9919a  and  a9914a );
 a9923a <=( A166  and  A168 );
 a9926a <=( (not A202)  and  (not A200) );
 a9927a <=( a9926a  and  a9923a );
 a9930a <=( (not A232)  and  (not A203) );
 a9934a <=( A266  and  (not A265) );
 a9935a <=( A233  and  a9934a );
 a9936a <=( a9935a  and  a9930a );
 a9939a <=( A166  and  A168 );
 a9942a <=( (not A201)  and  (not A200) );
 a9943a <=( a9942a  and  a9939a );
 a9946a <=( A233  and  (not A232) );
 a9950a <=( (not A302)  and  (not A301) );
 a9951a <=( (not A299)  and  a9950a );
 a9952a <=( a9951a  and  a9946a );
 a9955a <=( A166  and  A168 );
 a9958a <=( (not A200)  and  (not A199) );
 a9959a <=( a9958a  and  a9955a );
 a9962a <=( A233  and  (not A232) );
 a9966a <=( (not A302)  and  (not A301) );
 a9967a <=( (not A299)  and  a9966a );
 a9968a <=( a9967a  and  a9962a );
 a9971a <=( A167  and  A168 );
 a9974a <=( A200  and  A199 );
 a9975a <=( a9974a  and  a9971a );
 a9978a <=( A233  and  (not A232) );
 a9982a <=( (not A302)  and  (not A301) );
 a9983a <=( (not A299)  and  a9982a );
 a9984a <=( a9983a  and  a9978a );
 a9987a <=( A167  and  A168 );
 a9990a <=( (not A202)  and  (not A200) );
 a9991a <=( a9990a  and  a9987a );
 a9994a <=( (not A232)  and  (not A203) );
 a9998a <=( (not A300)  and  (not A299) );
 a9999a <=( A233  and  a9998a );
 a10000a <=( a9999a  and  a9994a );
 a10003a <=( A167  and  A168 );
 a10006a <=( (not A202)  and  (not A200) );
 a10007a <=( a10006a  and  a10003a );
 a10010a <=( (not A232)  and  (not A203) );
 a10014a <=( A299  and  A298 );
 a10015a <=( A233  and  a10014a );
 a10016a <=( a10015a  and  a10010a );
 a10019a <=( A167  and  A168 );
 a10022a <=( (not A202)  and  (not A200) );
 a10023a <=( a10022a  and  a10019a );
 a10026a <=( (not A232)  and  (not A203) );
 a10030a <=( (not A299)  and  (not A298) );
 a10031a <=( A233  and  a10030a );
 a10032a <=( a10031a  and  a10026a );
 a10035a <=( A167  and  A168 );
 a10038a <=( (not A202)  and  (not A200) );
 a10039a <=( a10038a  and  a10035a );
 a10042a <=( (not A232)  and  (not A203) );
 a10046a <=( A266  and  (not A265) );
 a10047a <=( A233  and  a10046a );
 a10048a <=( a10047a  and  a10042a );
 a10051a <=( A167  and  A168 );
 a10054a <=( (not A201)  and  (not A200) );
 a10055a <=( a10054a  and  a10051a );
 a10058a <=( A233  and  (not A232) );
 a10062a <=( (not A302)  and  (not A301) );
 a10063a <=( (not A299)  and  a10062a );
 a10064a <=( a10063a  and  a10058a );
 a10067a <=( A167  and  A168 );
 a10070a <=( (not A200)  and  (not A199) );
 a10071a <=( a10070a  and  a10067a );
 a10074a <=( A233  and  (not A232) );
 a10078a <=( (not A302)  and  (not A301) );
 a10079a <=( (not A299)  and  a10078a );
 a10080a <=( a10079a  and  a10074a );
 a10083a <=( (not A167)  and  A170 );
 a10086a <=( (not A199)  and  (not A166) );
 a10087a <=( a10086a  and  a10083a );
 a10090a <=( (not A232)  and  A200 );
 a10094a <=( (not A300)  and  (not A299) );
 a10095a <=( A233  and  a10094a );
 a10096a <=( a10095a  and  a10090a );
 a10099a <=( (not A167)  and  A170 );
 a10102a <=( (not A199)  and  (not A166) );
 a10103a <=( a10102a  and  a10099a );
 a10106a <=( (not A232)  and  A200 );
 a10110a <=( A299  and  A298 );
 a10111a <=( A233  and  a10110a );
 a10112a <=( a10111a  and  a10106a );
 a10115a <=( (not A167)  and  A170 );
 a10118a <=( (not A199)  and  (not A166) );
 a10119a <=( a10118a  and  a10115a );
 a10122a <=( (not A232)  and  A200 );
 a10126a <=( (not A299)  and  (not A298) );
 a10127a <=( A233  and  a10126a );
 a10128a <=( a10127a  and  a10122a );
 a10131a <=( (not A167)  and  A170 );
 a10134a <=( (not A199)  and  (not A166) );
 a10135a <=( a10134a  and  a10131a );
 a10138a <=( (not A232)  and  A200 );
 a10142a <=( A266  and  (not A265) );
 a10143a <=( A233  and  a10142a );
 a10144a <=( a10143a  and  a10138a );
 a10147a <=( (not A167)  and  (not A169) );
 a10150a <=( (not A199)  and  (not A166) );
 a10151a <=( a10150a  and  a10147a );
 a10154a <=( (not A232)  and  A200 );
 a10158a <=( (not A300)  and  (not A299) );
 a10159a <=( A233  and  a10158a );
 a10160a <=( a10159a  and  a10154a );
 a10163a <=( (not A167)  and  (not A169) );
 a10166a <=( (not A199)  and  (not A166) );
 a10167a <=( a10166a  and  a10163a );
 a10170a <=( (not A232)  and  A200 );
 a10174a <=( A299  and  A298 );
 a10175a <=( A233  and  a10174a );
 a10176a <=( a10175a  and  a10170a );
 a10179a <=( (not A167)  and  (not A169) );
 a10182a <=( (not A199)  and  (not A166) );
 a10183a <=( a10182a  and  a10179a );
 a10186a <=( (not A232)  and  A200 );
 a10190a <=( (not A299)  and  (not A298) );
 a10191a <=( A233  and  a10190a );
 a10192a <=( a10191a  and  a10186a );
 a10195a <=( (not A167)  and  (not A169) );
 a10198a <=( (not A199)  and  (not A166) );
 a10199a <=( a10198a  and  a10195a );
 a10202a <=( (not A232)  and  A200 );
 a10206a <=( A266  and  (not A265) );
 a10207a <=( A233  and  a10206a );
 a10208a <=( a10207a  and  a10202a );
 a10211a <=( A166  and  A168 );
 a10215a <=( A232  and  A200 );
 a10216a <=( A199  and  a10215a );
 a10217a <=( a10216a  and  a10211a );
 a10220a <=( A265  and  A233 );
 a10224a <=( A299  and  (not A298) );
 a10225a <=( (not A267)  and  a10224a );
 a10226a <=( a10225a  and  a10220a );
 a10229a <=( A166  and  A168 );
 a10233a <=( A232  and  A200 );
 a10234a <=( A199  and  a10233a );
 a10235a <=( a10234a  and  a10229a );
 a10238a <=( A265  and  A233 );
 a10242a <=( A299  and  (not A298) );
 a10243a <=( A266  and  a10242a );
 a10244a <=( a10243a  and  a10238a );
 a10247a <=( A166  and  A168 );
 a10251a <=( A232  and  A200 );
 a10252a <=( A199  and  a10251a );
 a10253a <=( a10252a  and  a10247a );
 a10256a <=( (not A265)  and  A233 );
 a10260a <=( A299  and  (not A298) );
 a10261a <=( (not A266)  and  a10260a );
 a10262a <=( a10261a  and  a10256a );
 a10265a <=( A166  and  A168 );
 a10269a <=( (not A232)  and  A200 );
 a10270a <=( A199  and  a10269a );
 a10271a <=( a10270a  and  a10265a );
 a10274a <=( A265  and  A233 );
 a10278a <=( A268  and  A267 );
 a10279a <=( (not A266)  and  a10278a );
 a10280a <=( a10279a  and  a10274a );
 a10283a <=( A166  and  A168 );
 a10287a <=( (not A232)  and  A200 );
 a10288a <=( A199  and  a10287a );
 a10289a <=( a10288a  and  a10283a );
 a10292a <=( A265  and  A233 );
 a10296a <=( A269  and  A267 );
 a10297a <=( (not A266)  and  a10296a );
 a10298a <=( a10297a  and  a10292a );
 a10301a <=( A166  and  A168 );
 a10305a <=( (not A233)  and  A200 );
 a10306a <=( A199  and  a10305a );
 a10307a <=( a10306a  and  a10301a );
 a10310a <=( A265  and  (not A234) );
 a10314a <=( A299  and  (not A298) );
 a10315a <=( A266  and  a10314a );
 a10316a <=( a10315a  and  a10310a );
 a10319a <=( A166  and  A168 );
 a10323a <=( (not A233)  and  A200 );
 a10324a <=( A199  and  a10323a );
 a10325a <=( a10324a  and  a10319a );
 a10328a <=( (not A266)  and  (not A234) );
 a10332a <=( A299  and  (not A298) );
 a10333a <=( (not A267)  and  a10332a );
 a10334a <=( a10333a  and  a10328a );
 a10337a <=( A166  and  A168 );
 a10341a <=( (not A233)  and  A200 );
 a10342a <=( A199  and  a10341a );
 a10343a <=( a10342a  and  a10337a );
 a10346a <=( (not A265)  and  (not A234) );
 a10350a <=( A299  and  (not A298) );
 a10351a <=( (not A266)  and  a10350a );
 a10352a <=( a10351a  and  a10346a );
 a10355a <=( A166  and  A168 );
 a10359a <=( A232  and  A200 );
 a10360a <=( A199  and  a10359a );
 a10361a <=( a10360a  and  a10355a );
 a10364a <=( A234  and  (not A233) );
 a10368a <=( (not A300)  and  A298 );
 a10369a <=( A235  and  a10368a );
 a10370a <=( a10369a  and  a10364a );
 a10373a <=( A166  and  A168 );
 a10377a <=( A232  and  A200 );
 a10378a <=( A199  and  a10377a );
 a10379a <=( a10378a  and  a10373a );
 a10382a <=( A234  and  (not A233) );
 a10386a <=( A299  and  A298 );
 a10387a <=( A235  and  a10386a );
 a10388a <=( a10387a  and  a10382a );
 a10391a <=( A166  and  A168 );
 a10395a <=( A232  and  A200 );
 a10396a <=( A199  and  a10395a );
 a10397a <=( a10396a  and  a10391a );
 a10400a <=( A234  and  (not A233) );
 a10404a <=( (not A299)  and  (not A298) );
 a10405a <=( A235  and  a10404a );
 a10406a <=( a10405a  and  a10400a );
 a10409a <=( A166  and  A168 );
 a10413a <=( A232  and  A200 );
 a10414a <=( A199  and  a10413a );
 a10415a <=( a10414a  and  a10409a );
 a10418a <=( A234  and  (not A233) );
 a10422a <=( A266  and  (not A265) );
 a10423a <=( A235  and  a10422a );
 a10424a <=( a10423a  and  a10418a );
 a10427a <=( A166  and  A168 );
 a10431a <=( A232  and  A200 );
 a10432a <=( A199  and  a10431a );
 a10433a <=( a10432a  and  a10427a );
 a10436a <=( A234  and  (not A233) );
 a10440a <=( (not A300)  and  A298 );
 a10441a <=( A236  and  a10440a );
 a10442a <=( a10441a  and  a10436a );
 a10445a <=( A166  and  A168 );
 a10449a <=( A232  and  A200 );
 a10450a <=( A199  and  a10449a );
 a10451a <=( a10450a  and  a10445a );
 a10454a <=( A234  and  (not A233) );
 a10458a <=( A299  and  A298 );
 a10459a <=( A236  and  a10458a );
 a10460a <=( a10459a  and  a10454a );
 a10463a <=( A166  and  A168 );
 a10467a <=( A232  and  A200 );
 a10468a <=( A199  and  a10467a );
 a10469a <=( a10468a  and  a10463a );
 a10472a <=( A234  and  (not A233) );
 a10476a <=( (not A299)  and  (not A298) );
 a10477a <=( A236  and  a10476a );
 a10478a <=( a10477a  and  a10472a );
 a10481a <=( A166  and  A168 );
 a10485a <=( A232  and  A200 );
 a10486a <=( A199  and  a10485a );
 a10487a <=( a10486a  and  a10481a );
 a10490a <=( A234  and  (not A233) );
 a10494a <=( A266  and  (not A265) );
 a10495a <=( A236  and  a10494a );
 a10496a <=( a10495a  and  a10490a );
 a10499a <=( A166  and  A168 );
 a10503a <=( (not A232)  and  A200 );
 a10504a <=( A199  and  a10503a );
 a10505a <=( a10504a  and  a10499a );
 a10508a <=( A265  and  (not A233) );
 a10512a <=( A299  and  (not A298) );
 a10513a <=( A266  and  a10512a );
 a10514a <=( a10513a  and  a10508a );
 a10517a <=( A166  and  A168 );
 a10521a <=( (not A232)  and  A200 );
 a10522a <=( A199  and  a10521a );
 a10523a <=( a10522a  and  a10517a );
 a10526a <=( (not A266)  and  (not A233) );
 a10530a <=( A299  and  (not A298) );
 a10531a <=( (not A267)  and  a10530a );
 a10532a <=( a10531a  and  a10526a );
 a10535a <=( A166  and  A168 );
 a10539a <=( (not A232)  and  A200 );
 a10540a <=( A199  and  a10539a );
 a10541a <=( a10540a  and  a10535a );
 a10544a <=( (not A265)  and  (not A233) );
 a10548a <=( A299  and  (not A298) );
 a10549a <=( (not A266)  and  a10548a );
 a10550a <=( a10549a  and  a10544a );
 a10553a <=( A166  and  A168 );
 a10557a <=( (not A203)  and  (not A202) );
 a10558a <=( (not A200)  and  a10557a );
 a10559a <=( a10558a  and  a10553a );
 a10562a <=( A233  and  (not A232) );
 a10566a <=( (not A302)  and  (not A301) );
 a10567a <=( (not A299)  and  a10566a );
 a10568a <=( a10567a  and  a10562a );
 a10571a <=( A166  and  A168 );
 a10575a <=( A232  and  (not A201) );
 a10576a <=( (not A200)  and  a10575a );
 a10577a <=( a10576a  and  a10571a );
 a10580a <=( A265  and  A233 );
 a10584a <=( A299  and  (not A298) );
 a10585a <=( (not A267)  and  a10584a );
 a10586a <=( a10585a  and  a10580a );
 a10589a <=( A166  and  A168 );
 a10593a <=( A232  and  (not A201) );
 a10594a <=( (not A200)  and  a10593a );
 a10595a <=( a10594a  and  a10589a );
 a10598a <=( A265  and  A233 );
 a10602a <=( A299  and  (not A298) );
 a10603a <=( A266  and  a10602a );
 a10604a <=( a10603a  and  a10598a );
 a10607a <=( A166  and  A168 );
 a10611a <=( A232  and  (not A201) );
 a10612a <=( (not A200)  and  a10611a );
 a10613a <=( a10612a  and  a10607a );
 a10616a <=( (not A265)  and  A233 );
 a10620a <=( A299  and  (not A298) );
 a10621a <=( (not A266)  and  a10620a );
 a10622a <=( a10621a  and  a10616a );
 a10625a <=( A166  and  A168 );
 a10629a <=( (not A232)  and  (not A201) );
 a10630a <=( (not A200)  and  a10629a );
 a10631a <=( a10630a  and  a10625a );
 a10634a <=( A265  and  A233 );
 a10638a <=( A268  and  A267 );
 a10639a <=( (not A266)  and  a10638a );
 a10640a <=( a10639a  and  a10634a );
 a10643a <=( A166  and  A168 );
 a10647a <=( (not A232)  and  (not A201) );
 a10648a <=( (not A200)  and  a10647a );
 a10649a <=( a10648a  and  a10643a );
 a10652a <=( A265  and  A233 );
 a10656a <=( A269  and  A267 );
 a10657a <=( (not A266)  and  a10656a );
 a10658a <=( a10657a  and  a10652a );
 a10661a <=( A166  and  A168 );
 a10665a <=( (not A233)  and  (not A201) );
 a10666a <=( (not A200)  and  a10665a );
 a10667a <=( a10666a  and  a10661a );
 a10670a <=( A265  and  (not A234) );
 a10674a <=( A299  and  (not A298) );
 a10675a <=( A266  and  a10674a );
 a10676a <=( a10675a  and  a10670a );
 a10679a <=( A166  and  A168 );
 a10683a <=( (not A233)  and  (not A201) );
 a10684a <=( (not A200)  and  a10683a );
 a10685a <=( a10684a  and  a10679a );
 a10688a <=( (not A266)  and  (not A234) );
 a10692a <=( A299  and  (not A298) );
 a10693a <=( (not A267)  and  a10692a );
 a10694a <=( a10693a  and  a10688a );
 a10697a <=( A166  and  A168 );
 a10701a <=( (not A233)  and  (not A201) );
 a10702a <=( (not A200)  and  a10701a );
 a10703a <=( a10702a  and  a10697a );
 a10706a <=( (not A265)  and  (not A234) );
 a10710a <=( A299  and  (not A298) );
 a10711a <=( (not A266)  and  a10710a );
 a10712a <=( a10711a  and  a10706a );
 a10715a <=( A166  and  A168 );
 a10719a <=( A232  and  (not A201) );
 a10720a <=( (not A200)  and  a10719a );
 a10721a <=( a10720a  and  a10715a );
 a10724a <=( A234  and  (not A233) );
 a10728a <=( (not A300)  and  A298 );
 a10729a <=( A235  and  a10728a );
 a10730a <=( a10729a  and  a10724a );
 a10733a <=( A166  and  A168 );
 a10737a <=( A232  and  (not A201) );
 a10738a <=( (not A200)  and  a10737a );
 a10739a <=( a10738a  and  a10733a );
 a10742a <=( A234  and  (not A233) );
 a10746a <=( A299  and  A298 );
 a10747a <=( A235  and  a10746a );
 a10748a <=( a10747a  and  a10742a );
 a10751a <=( A166  and  A168 );
 a10755a <=( A232  and  (not A201) );
 a10756a <=( (not A200)  and  a10755a );
 a10757a <=( a10756a  and  a10751a );
 a10760a <=( A234  and  (not A233) );
 a10764a <=( (not A299)  and  (not A298) );
 a10765a <=( A235  and  a10764a );
 a10766a <=( a10765a  and  a10760a );
 a10769a <=( A166  and  A168 );
 a10773a <=( A232  and  (not A201) );
 a10774a <=( (not A200)  and  a10773a );
 a10775a <=( a10774a  and  a10769a );
 a10778a <=( A234  and  (not A233) );
 a10782a <=( A266  and  (not A265) );
 a10783a <=( A235  and  a10782a );
 a10784a <=( a10783a  and  a10778a );
 a10787a <=( A166  and  A168 );
 a10791a <=( A232  and  (not A201) );
 a10792a <=( (not A200)  and  a10791a );
 a10793a <=( a10792a  and  a10787a );
 a10796a <=( A234  and  (not A233) );
 a10800a <=( (not A300)  and  A298 );
 a10801a <=( A236  and  a10800a );
 a10802a <=( a10801a  and  a10796a );
 a10805a <=( A166  and  A168 );
 a10809a <=( A232  and  (not A201) );
 a10810a <=( (not A200)  and  a10809a );
 a10811a <=( a10810a  and  a10805a );
 a10814a <=( A234  and  (not A233) );
 a10818a <=( A299  and  A298 );
 a10819a <=( A236  and  a10818a );
 a10820a <=( a10819a  and  a10814a );
 a10823a <=( A166  and  A168 );
 a10827a <=( A232  and  (not A201) );
 a10828a <=( (not A200)  and  a10827a );
 a10829a <=( a10828a  and  a10823a );
 a10832a <=( A234  and  (not A233) );
 a10836a <=( (not A299)  and  (not A298) );
 a10837a <=( A236  and  a10836a );
 a10838a <=( a10837a  and  a10832a );
 a10841a <=( A166  and  A168 );
 a10845a <=( A232  and  (not A201) );
 a10846a <=( (not A200)  and  a10845a );
 a10847a <=( a10846a  and  a10841a );
 a10850a <=( A234  and  (not A233) );
 a10854a <=( A266  and  (not A265) );
 a10855a <=( A236  and  a10854a );
 a10856a <=( a10855a  and  a10850a );
 a10859a <=( A166  and  A168 );
 a10863a <=( (not A232)  and  (not A201) );
 a10864a <=( (not A200)  and  a10863a );
 a10865a <=( a10864a  and  a10859a );
 a10868a <=( A265  and  (not A233) );
 a10872a <=( A299  and  (not A298) );
 a10873a <=( A266  and  a10872a );
 a10874a <=( a10873a  and  a10868a );
 a10877a <=( A166  and  A168 );
 a10881a <=( (not A232)  and  (not A201) );
 a10882a <=( (not A200)  and  a10881a );
 a10883a <=( a10882a  and  a10877a );
 a10886a <=( (not A266)  and  (not A233) );
 a10890a <=( A299  and  (not A298) );
 a10891a <=( (not A267)  and  a10890a );
 a10892a <=( a10891a  and  a10886a );
 a10895a <=( A166  and  A168 );
 a10899a <=( (not A232)  and  (not A201) );
 a10900a <=( (not A200)  and  a10899a );
 a10901a <=( a10900a  and  a10895a );
 a10904a <=( (not A265)  and  (not A233) );
 a10908a <=( A299  and  (not A298) );
 a10909a <=( (not A266)  and  a10908a );
 a10910a <=( a10909a  and  a10904a );
 a10913a <=( A166  and  A168 );
 a10917a <=( A232  and  (not A200) );
 a10918a <=( (not A199)  and  a10917a );
 a10919a <=( a10918a  and  a10913a );
 a10922a <=( A265  and  A233 );
 a10926a <=( A299  and  (not A298) );
 a10927a <=( (not A267)  and  a10926a );
 a10928a <=( a10927a  and  a10922a );
 a10931a <=( A166  and  A168 );
 a10935a <=( A232  and  (not A200) );
 a10936a <=( (not A199)  and  a10935a );
 a10937a <=( a10936a  and  a10931a );
 a10940a <=( A265  and  A233 );
 a10944a <=( A299  and  (not A298) );
 a10945a <=( A266  and  a10944a );
 a10946a <=( a10945a  and  a10940a );
 a10949a <=( A166  and  A168 );
 a10953a <=( A232  and  (not A200) );
 a10954a <=( (not A199)  and  a10953a );
 a10955a <=( a10954a  and  a10949a );
 a10958a <=( (not A265)  and  A233 );
 a10962a <=( A299  and  (not A298) );
 a10963a <=( (not A266)  and  a10962a );
 a10964a <=( a10963a  and  a10958a );
 a10967a <=( A166  and  A168 );
 a10971a <=( (not A232)  and  (not A200) );
 a10972a <=( (not A199)  and  a10971a );
 a10973a <=( a10972a  and  a10967a );
 a10976a <=( A265  and  A233 );
 a10980a <=( A268  and  A267 );
 a10981a <=( (not A266)  and  a10980a );
 a10982a <=( a10981a  and  a10976a );
 a10985a <=( A166  and  A168 );
 a10989a <=( (not A232)  and  (not A200) );
 a10990a <=( (not A199)  and  a10989a );
 a10991a <=( a10990a  and  a10985a );
 a10994a <=( A265  and  A233 );
 a10998a <=( A269  and  A267 );
 a10999a <=( (not A266)  and  a10998a );
 a11000a <=( a10999a  and  a10994a );
 a11003a <=( A166  and  A168 );
 a11007a <=( (not A233)  and  (not A200) );
 a11008a <=( (not A199)  and  a11007a );
 a11009a <=( a11008a  and  a11003a );
 a11012a <=( A265  and  (not A234) );
 a11016a <=( A299  and  (not A298) );
 a11017a <=( A266  and  a11016a );
 a11018a <=( a11017a  and  a11012a );
 a11021a <=( A166  and  A168 );
 a11025a <=( (not A233)  and  (not A200) );
 a11026a <=( (not A199)  and  a11025a );
 a11027a <=( a11026a  and  a11021a );
 a11030a <=( (not A266)  and  (not A234) );
 a11034a <=( A299  and  (not A298) );
 a11035a <=( (not A267)  and  a11034a );
 a11036a <=( a11035a  and  a11030a );
 a11039a <=( A166  and  A168 );
 a11043a <=( (not A233)  and  (not A200) );
 a11044a <=( (not A199)  and  a11043a );
 a11045a <=( a11044a  and  a11039a );
 a11048a <=( (not A265)  and  (not A234) );
 a11052a <=( A299  and  (not A298) );
 a11053a <=( (not A266)  and  a11052a );
 a11054a <=( a11053a  and  a11048a );
 a11057a <=( A166  and  A168 );
 a11061a <=( A232  and  (not A200) );
 a11062a <=( (not A199)  and  a11061a );
 a11063a <=( a11062a  and  a11057a );
 a11066a <=( A234  and  (not A233) );
 a11070a <=( (not A300)  and  A298 );
 a11071a <=( A235  and  a11070a );
 a11072a <=( a11071a  and  a11066a );
 a11075a <=( A166  and  A168 );
 a11079a <=( A232  and  (not A200) );
 a11080a <=( (not A199)  and  a11079a );
 a11081a <=( a11080a  and  a11075a );
 a11084a <=( A234  and  (not A233) );
 a11088a <=( A299  and  A298 );
 a11089a <=( A235  and  a11088a );
 a11090a <=( a11089a  and  a11084a );
 a11093a <=( A166  and  A168 );
 a11097a <=( A232  and  (not A200) );
 a11098a <=( (not A199)  and  a11097a );
 a11099a <=( a11098a  and  a11093a );
 a11102a <=( A234  and  (not A233) );
 a11106a <=( (not A299)  and  (not A298) );
 a11107a <=( A235  and  a11106a );
 a11108a <=( a11107a  and  a11102a );
 a11111a <=( A166  and  A168 );
 a11115a <=( A232  and  (not A200) );
 a11116a <=( (not A199)  and  a11115a );
 a11117a <=( a11116a  and  a11111a );
 a11120a <=( A234  and  (not A233) );
 a11124a <=( A266  and  (not A265) );
 a11125a <=( A235  and  a11124a );
 a11126a <=( a11125a  and  a11120a );
 a11129a <=( A166  and  A168 );
 a11133a <=( A232  and  (not A200) );
 a11134a <=( (not A199)  and  a11133a );
 a11135a <=( a11134a  and  a11129a );
 a11138a <=( A234  and  (not A233) );
 a11142a <=( (not A300)  and  A298 );
 a11143a <=( A236  and  a11142a );
 a11144a <=( a11143a  and  a11138a );
 a11147a <=( A166  and  A168 );
 a11151a <=( A232  and  (not A200) );
 a11152a <=( (not A199)  and  a11151a );
 a11153a <=( a11152a  and  a11147a );
 a11156a <=( A234  and  (not A233) );
 a11160a <=( A299  and  A298 );
 a11161a <=( A236  and  a11160a );
 a11162a <=( a11161a  and  a11156a );
 a11165a <=( A166  and  A168 );
 a11169a <=( A232  and  (not A200) );
 a11170a <=( (not A199)  and  a11169a );
 a11171a <=( a11170a  and  a11165a );
 a11174a <=( A234  and  (not A233) );
 a11178a <=( (not A299)  and  (not A298) );
 a11179a <=( A236  and  a11178a );
 a11180a <=( a11179a  and  a11174a );
 a11183a <=( A166  and  A168 );
 a11187a <=( A232  and  (not A200) );
 a11188a <=( (not A199)  and  a11187a );
 a11189a <=( a11188a  and  a11183a );
 a11192a <=( A234  and  (not A233) );
 a11196a <=( A266  and  (not A265) );
 a11197a <=( A236  and  a11196a );
 a11198a <=( a11197a  and  a11192a );
 a11201a <=( A166  and  A168 );
 a11205a <=( (not A232)  and  (not A200) );
 a11206a <=( (not A199)  and  a11205a );
 a11207a <=( a11206a  and  a11201a );
 a11210a <=( A265  and  (not A233) );
 a11214a <=( A299  and  (not A298) );
 a11215a <=( A266  and  a11214a );
 a11216a <=( a11215a  and  a11210a );
 a11219a <=( A166  and  A168 );
 a11223a <=( (not A232)  and  (not A200) );
 a11224a <=( (not A199)  and  a11223a );
 a11225a <=( a11224a  and  a11219a );
 a11228a <=( (not A266)  and  (not A233) );
 a11232a <=( A299  and  (not A298) );
 a11233a <=( (not A267)  and  a11232a );
 a11234a <=( a11233a  and  a11228a );
 a11237a <=( A166  and  A168 );
 a11241a <=( (not A232)  and  (not A200) );
 a11242a <=( (not A199)  and  a11241a );
 a11243a <=( a11242a  and  a11237a );
 a11246a <=( (not A265)  and  (not A233) );
 a11250a <=( A299  and  (not A298) );
 a11251a <=( (not A266)  and  a11250a );
 a11252a <=( a11251a  and  a11246a );
 a11255a <=( A167  and  A168 );
 a11259a <=( A232  and  A200 );
 a11260a <=( A199  and  a11259a );
 a11261a <=( a11260a  and  a11255a );
 a11264a <=( A265  and  A233 );
 a11268a <=( A299  and  (not A298) );
 a11269a <=( (not A267)  and  a11268a );
 a11270a <=( a11269a  and  a11264a );
 a11273a <=( A167  and  A168 );
 a11277a <=( A232  and  A200 );
 a11278a <=( A199  and  a11277a );
 a11279a <=( a11278a  and  a11273a );
 a11282a <=( A265  and  A233 );
 a11286a <=( A299  and  (not A298) );
 a11287a <=( A266  and  a11286a );
 a11288a <=( a11287a  and  a11282a );
 a11291a <=( A167  and  A168 );
 a11295a <=( A232  and  A200 );
 a11296a <=( A199  and  a11295a );
 a11297a <=( a11296a  and  a11291a );
 a11300a <=( (not A265)  and  A233 );
 a11304a <=( A299  and  (not A298) );
 a11305a <=( (not A266)  and  a11304a );
 a11306a <=( a11305a  and  a11300a );
 a11309a <=( A167  and  A168 );
 a11313a <=( (not A232)  and  A200 );
 a11314a <=( A199  and  a11313a );
 a11315a <=( a11314a  and  a11309a );
 a11318a <=( A265  and  A233 );
 a11322a <=( A268  and  A267 );
 a11323a <=( (not A266)  and  a11322a );
 a11324a <=( a11323a  and  a11318a );
 a11327a <=( A167  and  A168 );
 a11331a <=( (not A232)  and  A200 );
 a11332a <=( A199  and  a11331a );
 a11333a <=( a11332a  and  a11327a );
 a11336a <=( A265  and  A233 );
 a11340a <=( A269  and  A267 );
 a11341a <=( (not A266)  and  a11340a );
 a11342a <=( a11341a  and  a11336a );
 a11345a <=( A167  and  A168 );
 a11349a <=( (not A233)  and  A200 );
 a11350a <=( A199  and  a11349a );
 a11351a <=( a11350a  and  a11345a );
 a11354a <=( A265  and  (not A234) );
 a11358a <=( A299  and  (not A298) );
 a11359a <=( A266  and  a11358a );
 a11360a <=( a11359a  and  a11354a );
 a11363a <=( A167  and  A168 );
 a11367a <=( (not A233)  and  A200 );
 a11368a <=( A199  and  a11367a );
 a11369a <=( a11368a  and  a11363a );
 a11372a <=( (not A266)  and  (not A234) );
 a11376a <=( A299  and  (not A298) );
 a11377a <=( (not A267)  and  a11376a );
 a11378a <=( a11377a  and  a11372a );
 a11381a <=( A167  and  A168 );
 a11385a <=( (not A233)  and  A200 );
 a11386a <=( A199  and  a11385a );
 a11387a <=( a11386a  and  a11381a );
 a11390a <=( (not A265)  and  (not A234) );
 a11394a <=( A299  and  (not A298) );
 a11395a <=( (not A266)  and  a11394a );
 a11396a <=( a11395a  and  a11390a );
 a11399a <=( A167  and  A168 );
 a11403a <=( A232  and  A200 );
 a11404a <=( A199  and  a11403a );
 a11405a <=( a11404a  and  a11399a );
 a11408a <=( A234  and  (not A233) );
 a11412a <=( (not A300)  and  A298 );
 a11413a <=( A235  and  a11412a );
 a11414a <=( a11413a  and  a11408a );
 a11417a <=( A167  and  A168 );
 a11421a <=( A232  and  A200 );
 a11422a <=( A199  and  a11421a );
 a11423a <=( a11422a  and  a11417a );
 a11426a <=( A234  and  (not A233) );
 a11430a <=( A299  and  A298 );
 a11431a <=( A235  and  a11430a );
 a11432a <=( a11431a  and  a11426a );
 a11435a <=( A167  and  A168 );
 a11439a <=( A232  and  A200 );
 a11440a <=( A199  and  a11439a );
 a11441a <=( a11440a  and  a11435a );
 a11444a <=( A234  and  (not A233) );
 a11448a <=( (not A299)  and  (not A298) );
 a11449a <=( A235  and  a11448a );
 a11450a <=( a11449a  and  a11444a );
 a11453a <=( A167  and  A168 );
 a11457a <=( A232  and  A200 );
 a11458a <=( A199  and  a11457a );
 a11459a <=( a11458a  and  a11453a );
 a11462a <=( A234  and  (not A233) );
 a11466a <=( A266  and  (not A265) );
 a11467a <=( A235  and  a11466a );
 a11468a <=( a11467a  and  a11462a );
 a11471a <=( A167  and  A168 );
 a11475a <=( A232  and  A200 );
 a11476a <=( A199  and  a11475a );
 a11477a <=( a11476a  and  a11471a );
 a11480a <=( A234  and  (not A233) );
 a11484a <=( (not A300)  and  A298 );
 a11485a <=( A236  and  a11484a );
 a11486a <=( a11485a  and  a11480a );
 a11489a <=( A167  and  A168 );
 a11493a <=( A232  and  A200 );
 a11494a <=( A199  and  a11493a );
 a11495a <=( a11494a  and  a11489a );
 a11498a <=( A234  and  (not A233) );
 a11502a <=( A299  and  A298 );
 a11503a <=( A236  and  a11502a );
 a11504a <=( a11503a  and  a11498a );
 a11507a <=( A167  and  A168 );
 a11511a <=( A232  and  A200 );
 a11512a <=( A199  and  a11511a );
 a11513a <=( a11512a  and  a11507a );
 a11516a <=( A234  and  (not A233) );
 a11520a <=( (not A299)  and  (not A298) );
 a11521a <=( A236  and  a11520a );
 a11522a <=( a11521a  and  a11516a );
 a11525a <=( A167  and  A168 );
 a11529a <=( A232  and  A200 );
 a11530a <=( A199  and  a11529a );
 a11531a <=( a11530a  and  a11525a );
 a11534a <=( A234  and  (not A233) );
 a11538a <=( A266  and  (not A265) );
 a11539a <=( A236  and  a11538a );
 a11540a <=( a11539a  and  a11534a );
 a11543a <=( A167  and  A168 );
 a11547a <=( (not A232)  and  A200 );
 a11548a <=( A199  and  a11547a );
 a11549a <=( a11548a  and  a11543a );
 a11552a <=( A265  and  (not A233) );
 a11556a <=( A299  and  (not A298) );
 a11557a <=( A266  and  a11556a );
 a11558a <=( a11557a  and  a11552a );
 a11561a <=( A167  and  A168 );
 a11565a <=( (not A232)  and  A200 );
 a11566a <=( A199  and  a11565a );
 a11567a <=( a11566a  and  a11561a );
 a11570a <=( (not A266)  and  (not A233) );
 a11574a <=( A299  and  (not A298) );
 a11575a <=( (not A267)  and  a11574a );
 a11576a <=( a11575a  and  a11570a );
 a11579a <=( A167  and  A168 );
 a11583a <=( (not A232)  and  A200 );
 a11584a <=( A199  and  a11583a );
 a11585a <=( a11584a  and  a11579a );
 a11588a <=( (not A265)  and  (not A233) );
 a11592a <=( A299  and  (not A298) );
 a11593a <=( (not A266)  and  a11592a );
 a11594a <=( a11593a  and  a11588a );
 a11597a <=( A167  and  A168 );
 a11601a <=( (not A203)  and  (not A202) );
 a11602a <=( (not A200)  and  a11601a );
 a11603a <=( a11602a  and  a11597a );
 a11606a <=( A233  and  (not A232) );
 a11610a <=( (not A302)  and  (not A301) );
 a11611a <=( (not A299)  and  a11610a );
 a11612a <=( a11611a  and  a11606a );
 a11615a <=( A167  and  A168 );
 a11619a <=( A232  and  (not A201) );
 a11620a <=( (not A200)  and  a11619a );
 a11621a <=( a11620a  and  a11615a );
 a11624a <=( A265  and  A233 );
 a11628a <=( A299  and  (not A298) );
 a11629a <=( (not A267)  and  a11628a );
 a11630a <=( a11629a  and  a11624a );
 a11633a <=( A167  and  A168 );
 a11637a <=( A232  and  (not A201) );
 a11638a <=( (not A200)  and  a11637a );
 a11639a <=( a11638a  and  a11633a );
 a11642a <=( A265  and  A233 );
 a11646a <=( A299  and  (not A298) );
 a11647a <=( A266  and  a11646a );
 a11648a <=( a11647a  and  a11642a );
 a11651a <=( A167  and  A168 );
 a11655a <=( A232  and  (not A201) );
 a11656a <=( (not A200)  and  a11655a );
 a11657a <=( a11656a  and  a11651a );
 a11660a <=( (not A265)  and  A233 );
 a11664a <=( A299  and  (not A298) );
 a11665a <=( (not A266)  and  a11664a );
 a11666a <=( a11665a  and  a11660a );
 a11669a <=( A167  and  A168 );
 a11673a <=( (not A232)  and  (not A201) );
 a11674a <=( (not A200)  and  a11673a );
 a11675a <=( a11674a  and  a11669a );
 a11678a <=( A265  and  A233 );
 a11682a <=( A268  and  A267 );
 a11683a <=( (not A266)  and  a11682a );
 a11684a <=( a11683a  and  a11678a );
 a11687a <=( A167  and  A168 );
 a11691a <=( (not A232)  and  (not A201) );
 a11692a <=( (not A200)  and  a11691a );
 a11693a <=( a11692a  and  a11687a );
 a11696a <=( A265  and  A233 );
 a11700a <=( A269  and  A267 );
 a11701a <=( (not A266)  and  a11700a );
 a11702a <=( a11701a  and  a11696a );
 a11705a <=( A167  and  A168 );
 a11709a <=( (not A233)  and  (not A201) );
 a11710a <=( (not A200)  and  a11709a );
 a11711a <=( a11710a  and  a11705a );
 a11714a <=( A265  and  (not A234) );
 a11718a <=( A299  and  (not A298) );
 a11719a <=( A266  and  a11718a );
 a11720a <=( a11719a  and  a11714a );
 a11723a <=( A167  and  A168 );
 a11727a <=( (not A233)  and  (not A201) );
 a11728a <=( (not A200)  and  a11727a );
 a11729a <=( a11728a  and  a11723a );
 a11732a <=( (not A266)  and  (not A234) );
 a11736a <=( A299  and  (not A298) );
 a11737a <=( (not A267)  and  a11736a );
 a11738a <=( a11737a  and  a11732a );
 a11741a <=( A167  and  A168 );
 a11745a <=( (not A233)  and  (not A201) );
 a11746a <=( (not A200)  and  a11745a );
 a11747a <=( a11746a  and  a11741a );
 a11750a <=( (not A265)  and  (not A234) );
 a11754a <=( A299  and  (not A298) );
 a11755a <=( (not A266)  and  a11754a );
 a11756a <=( a11755a  and  a11750a );
 a11759a <=( A167  and  A168 );
 a11763a <=( A232  and  (not A201) );
 a11764a <=( (not A200)  and  a11763a );
 a11765a <=( a11764a  and  a11759a );
 a11768a <=( A234  and  (not A233) );
 a11772a <=( (not A300)  and  A298 );
 a11773a <=( A235  and  a11772a );
 a11774a <=( a11773a  and  a11768a );
 a11777a <=( A167  and  A168 );
 a11781a <=( A232  and  (not A201) );
 a11782a <=( (not A200)  and  a11781a );
 a11783a <=( a11782a  and  a11777a );
 a11786a <=( A234  and  (not A233) );
 a11790a <=( A299  and  A298 );
 a11791a <=( A235  and  a11790a );
 a11792a <=( a11791a  and  a11786a );
 a11795a <=( A167  and  A168 );
 a11799a <=( A232  and  (not A201) );
 a11800a <=( (not A200)  and  a11799a );
 a11801a <=( a11800a  and  a11795a );
 a11804a <=( A234  and  (not A233) );
 a11808a <=( (not A299)  and  (not A298) );
 a11809a <=( A235  and  a11808a );
 a11810a <=( a11809a  and  a11804a );
 a11813a <=( A167  and  A168 );
 a11817a <=( A232  and  (not A201) );
 a11818a <=( (not A200)  and  a11817a );
 a11819a <=( a11818a  and  a11813a );
 a11822a <=( A234  and  (not A233) );
 a11826a <=( A266  and  (not A265) );
 a11827a <=( A235  and  a11826a );
 a11828a <=( a11827a  and  a11822a );
 a11831a <=( A167  and  A168 );
 a11835a <=( A232  and  (not A201) );
 a11836a <=( (not A200)  and  a11835a );
 a11837a <=( a11836a  and  a11831a );
 a11840a <=( A234  and  (not A233) );
 a11844a <=( (not A300)  and  A298 );
 a11845a <=( A236  and  a11844a );
 a11846a <=( a11845a  and  a11840a );
 a11849a <=( A167  and  A168 );
 a11853a <=( A232  and  (not A201) );
 a11854a <=( (not A200)  and  a11853a );
 a11855a <=( a11854a  and  a11849a );
 a11858a <=( A234  and  (not A233) );
 a11862a <=( A299  and  A298 );
 a11863a <=( A236  and  a11862a );
 a11864a <=( a11863a  and  a11858a );
 a11867a <=( A167  and  A168 );
 a11871a <=( A232  and  (not A201) );
 a11872a <=( (not A200)  and  a11871a );
 a11873a <=( a11872a  and  a11867a );
 a11876a <=( A234  and  (not A233) );
 a11880a <=( (not A299)  and  (not A298) );
 a11881a <=( A236  and  a11880a );
 a11882a <=( a11881a  and  a11876a );
 a11885a <=( A167  and  A168 );
 a11889a <=( A232  and  (not A201) );
 a11890a <=( (not A200)  and  a11889a );
 a11891a <=( a11890a  and  a11885a );
 a11894a <=( A234  and  (not A233) );
 a11898a <=( A266  and  (not A265) );
 a11899a <=( A236  and  a11898a );
 a11900a <=( a11899a  and  a11894a );
 a11903a <=( A167  and  A168 );
 a11907a <=( (not A232)  and  (not A201) );
 a11908a <=( (not A200)  and  a11907a );
 a11909a <=( a11908a  and  a11903a );
 a11912a <=( A265  and  (not A233) );
 a11916a <=( A299  and  (not A298) );
 a11917a <=( A266  and  a11916a );
 a11918a <=( a11917a  and  a11912a );
 a11921a <=( A167  and  A168 );
 a11925a <=( (not A232)  and  (not A201) );
 a11926a <=( (not A200)  and  a11925a );
 a11927a <=( a11926a  and  a11921a );
 a11930a <=( (not A266)  and  (not A233) );
 a11934a <=( A299  and  (not A298) );
 a11935a <=( (not A267)  and  a11934a );
 a11936a <=( a11935a  and  a11930a );
 a11939a <=( A167  and  A168 );
 a11943a <=( (not A232)  and  (not A201) );
 a11944a <=( (not A200)  and  a11943a );
 a11945a <=( a11944a  and  a11939a );
 a11948a <=( (not A265)  and  (not A233) );
 a11952a <=( A299  and  (not A298) );
 a11953a <=( (not A266)  and  a11952a );
 a11954a <=( a11953a  and  a11948a );
 a11957a <=( A167  and  A168 );
 a11961a <=( A232  and  (not A200) );
 a11962a <=( (not A199)  and  a11961a );
 a11963a <=( a11962a  and  a11957a );
 a11966a <=( A265  and  A233 );
 a11970a <=( A299  and  (not A298) );
 a11971a <=( (not A267)  and  a11970a );
 a11972a <=( a11971a  and  a11966a );
 a11975a <=( A167  and  A168 );
 a11979a <=( A232  and  (not A200) );
 a11980a <=( (not A199)  and  a11979a );
 a11981a <=( a11980a  and  a11975a );
 a11984a <=( A265  and  A233 );
 a11988a <=( A299  and  (not A298) );
 a11989a <=( A266  and  a11988a );
 a11990a <=( a11989a  and  a11984a );
 a11993a <=( A167  and  A168 );
 a11997a <=( A232  and  (not A200) );
 a11998a <=( (not A199)  and  a11997a );
 a11999a <=( a11998a  and  a11993a );
 a12002a <=( (not A265)  and  A233 );
 a12006a <=( A299  and  (not A298) );
 a12007a <=( (not A266)  and  a12006a );
 a12008a <=( a12007a  and  a12002a );
 a12011a <=( A167  and  A168 );
 a12015a <=( (not A232)  and  (not A200) );
 a12016a <=( (not A199)  and  a12015a );
 a12017a <=( a12016a  and  a12011a );
 a12020a <=( A265  and  A233 );
 a12024a <=( A268  and  A267 );
 a12025a <=( (not A266)  and  a12024a );
 a12026a <=( a12025a  and  a12020a );
 a12029a <=( A167  and  A168 );
 a12033a <=( (not A232)  and  (not A200) );
 a12034a <=( (not A199)  and  a12033a );
 a12035a <=( a12034a  and  a12029a );
 a12038a <=( A265  and  A233 );
 a12042a <=( A269  and  A267 );
 a12043a <=( (not A266)  and  a12042a );
 a12044a <=( a12043a  and  a12038a );
 a12047a <=( A167  and  A168 );
 a12051a <=( (not A233)  and  (not A200) );
 a12052a <=( (not A199)  and  a12051a );
 a12053a <=( a12052a  and  a12047a );
 a12056a <=( A265  and  (not A234) );
 a12060a <=( A299  and  (not A298) );
 a12061a <=( A266  and  a12060a );
 a12062a <=( a12061a  and  a12056a );
 a12065a <=( A167  and  A168 );
 a12069a <=( (not A233)  and  (not A200) );
 a12070a <=( (not A199)  and  a12069a );
 a12071a <=( a12070a  and  a12065a );
 a12074a <=( (not A266)  and  (not A234) );
 a12078a <=( A299  and  (not A298) );
 a12079a <=( (not A267)  and  a12078a );
 a12080a <=( a12079a  and  a12074a );
 a12083a <=( A167  and  A168 );
 a12087a <=( (not A233)  and  (not A200) );
 a12088a <=( (not A199)  and  a12087a );
 a12089a <=( a12088a  and  a12083a );
 a12092a <=( (not A265)  and  (not A234) );
 a12096a <=( A299  and  (not A298) );
 a12097a <=( (not A266)  and  a12096a );
 a12098a <=( a12097a  and  a12092a );
 a12101a <=( A167  and  A168 );
 a12105a <=( A232  and  (not A200) );
 a12106a <=( (not A199)  and  a12105a );
 a12107a <=( a12106a  and  a12101a );
 a12110a <=( A234  and  (not A233) );
 a12114a <=( (not A300)  and  A298 );
 a12115a <=( A235  and  a12114a );
 a12116a <=( a12115a  and  a12110a );
 a12119a <=( A167  and  A168 );
 a12123a <=( A232  and  (not A200) );
 a12124a <=( (not A199)  and  a12123a );
 a12125a <=( a12124a  and  a12119a );
 a12128a <=( A234  and  (not A233) );
 a12132a <=( A299  and  A298 );
 a12133a <=( A235  and  a12132a );
 a12134a <=( a12133a  and  a12128a );
 a12137a <=( A167  and  A168 );
 a12141a <=( A232  and  (not A200) );
 a12142a <=( (not A199)  and  a12141a );
 a12143a <=( a12142a  and  a12137a );
 a12146a <=( A234  and  (not A233) );
 a12150a <=( (not A299)  and  (not A298) );
 a12151a <=( A235  and  a12150a );
 a12152a <=( a12151a  and  a12146a );
 a12155a <=( A167  and  A168 );
 a12159a <=( A232  and  (not A200) );
 a12160a <=( (not A199)  and  a12159a );
 a12161a <=( a12160a  and  a12155a );
 a12164a <=( A234  and  (not A233) );
 a12168a <=( A266  and  (not A265) );
 a12169a <=( A235  and  a12168a );
 a12170a <=( a12169a  and  a12164a );
 a12173a <=( A167  and  A168 );
 a12177a <=( A232  and  (not A200) );
 a12178a <=( (not A199)  and  a12177a );
 a12179a <=( a12178a  and  a12173a );
 a12182a <=( A234  and  (not A233) );
 a12186a <=( (not A300)  and  A298 );
 a12187a <=( A236  and  a12186a );
 a12188a <=( a12187a  and  a12182a );
 a12191a <=( A167  and  A168 );
 a12195a <=( A232  and  (not A200) );
 a12196a <=( (not A199)  and  a12195a );
 a12197a <=( a12196a  and  a12191a );
 a12200a <=( A234  and  (not A233) );
 a12204a <=( A299  and  A298 );
 a12205a <=( A236  and  a12204a );
 a12206a <=( a12205a  and  a12200a );
 a12209a <=( A167  and  A168 );
 a12213a <=( A232  and  (not A200) );
 a12214a <=( (not A199)  and  a12213a );
 a12215a <=( a12214a  and  a12209a );
 a12218a <=( A234  and  (not A233) );
 a12222a <=( (not A299)  and  (not A298) );
 a12223a <=( A236  and  a12222a );
 a12224a <=( a12223a  and  a12218a );
 a12227a <=( A167  and  A168 );
 a12231a <=( A232  and  (not A200) );
 a12232a <=( (not A199)  and  a12231a );
 a12233a <=( a12232a  and  a12227a );
 a12236a <=( A234  and  (not A233) );
 a12240a <=( A266  and  (not A265) );
 a12241a <=( A236  and  a12240a );
 a12242a <=( a12241a  and  a12236a );
 a12245a <=( A167  and  A168 );
 a12249a <=( (not A232)  and  (not A200) );
 a12250a <=( (not A199)  and  a12249a );
 a12251a <=( a12250a  and  a12245a );
 a12254a <=( A265  and  (not A233) );
 a12258a <=( A299  and  (not A298) );
 a12259a <=( A266  and  a12258a );
 a12260a <=( a12259a  and  a12254a );
 a12263a <=( A167  and  A168 );
 a12267a <=( (not A232)  and  (not A200) );
 a12268a <=( (not A199)  and  a12267a );
 a12269a <=( a12268a  and  a12263a );
 a12272a <=( (not A266)  and  (not A233) );
 a12276a <=( A299  and  (not A298) );
 a12277a <=( (not A267)  and  a12276a );
 a12278a <=( a12277a  and  a12272a );
 a12281a <=( A167  and  A168 );
 a12285a <=( (not A232)  and  (not A200) );
 a12286a <=( (not A199)  and  a12285a );
 a12287a <=( a12286a  and  a12281a );
 a12290a <=( (not A265)  and  (not A233) );
 a12294a <=( A299  and  (not A298) );
 a12295a <=( (not A266)  and  a12294a );
 a12296a <=( a12295a  and  a12290a );
 a12299a <=( (not A167)  and  A170 );
 a12303a <=( A200  and  (not A199) );
 a12304a <=( (not A166)  and  a12303a );
 a12305a <=( a12304a  and  a12299a );
 a12308a <=( A233  and  (not A232) );
 a12312a <=( (not A302)  and  (not A301) );
 a12313a <=( (not A299)  and  a12312a );
 a12314a <=( a12313a  and  a12308a );
 a12317a <=( (not A168)  and  A170 );
 a12321a <=( (not A199)  and  A166 );
 a12322a <=( A167  and  a12321a );
 a12323a <=( a12322a  and  a12317a );
 a12326a <=( (not A232)  and  A200 );
 a12330a <=( (not A300)  and  (not A299) );
 a12331a <=( A233  and  a12330a );
 a12332a <=( a12331a  and  a12326a );
 a12335a <=( (not A168)  and  A170 );
 a12339a <=( (not A199)  and  A166 );
 a12340a <=( A167  and  a12339a );
 a12341a <=( a12340a  and  a12335a );
 a12344a <=( (not A232)  and  A200 );
 a12348a <=( A299  and  A298 );
 a12349a <=( A233  and  a12348a );
 a12350a <=( a12349a  and  a12344a );
 a12353a <=( (not A168)  and  A170 );
 a12357a <=( (not A199)  and  A166 );
 a12358a <=( A167  and  a12357a );
 a12359a <=( a12358a  and  a12353a );
 a12362a <=( (not A232)  and  A200 );
 a12366a <=( (not A299)  and  (not A298) );
 a12367a <=( A233  and  a12366a );
 a12368a <=( a12367a  and  a12362a );
 a12371a <=( (not A168)  and  A170 );
 a12375a <=( (not A199)  and  A166 );
 a12376a <=( A167  and  a12375a );
 a12377a <=( a12376a  and  a12371a );
 a12380a <=( (not A232)  and  A200 );
 a12384a <=( A266  and  (not A265) );
 a12385a <=( A233  and  a12384a );
 a12386a <=( a12385a  and  a12380a );
 a12389a <=( (not A168)  and  (not A170) );
 a12393a <=( (not A199)  and  (not A166) );
 a12394a <=( A167  and  a12393a );
 a12395a <=( a12394a  and  a12389a );
 a12398a <=( (not A232)  and  A200 );
 a12402a <=( (not A300)  and  (not A299) );
 a12403a <=( A233  and  a12402a );
 a12404a <=( a12403a  and  a12398a );
 a12407a <=( (not A168)  and  (not A170) );
 a12411a <=( (not A199)  and  (not A166) );
 a12412a <=( A167  and  a12411a );
 a12413a <=( a12412a  and  a12407a );
 a12416a <=( (not A232)  and  A200 );
 a12420a <=( A299  and  A298 );
 a12421a <=( A233  and  a12420a );
 a12422a <=( a12421a  and  a12416a );
 a12425a <=( (not A168)  and  (not A170) );
 a12429a <=( (not A199)  and  (not A166) );
 a12430a <=( A167  and  a12429a );
 a12431a <=( a12430a  and  a12425a );
 a12434a <=( (not A232)  and  A200 );
 a12438a <=( (not A299)  and  (not A298) );
 a12439a <=( A233  and  a12438a );
 a12440a <=( a12439a  and  a12434a );
 a12443a <=( (not A168)  and  (not A170) );
 a12447a <=( (not A199)  and  (not A166) );
 a12448a <=( A167  and  a12447a );
 a12449a <=( a12448a  and  a12443a );
 a12452a <=( (not A232)  and  A200 );
 a12456a <=( A266  and  (not A265) );
 a12457a <=( A233  and  a12456a );
 a12458a <=( a12457a  and  a12452a );
 a12461a <=( (not A168)  and  (not A170) );
 a12465a <=( (not A199)  and  A166 );
 a12466a <=( (not A167)  and  a12465a );
 a12467a <=( a12466a  and  a12461a );
 a12470a <=( (not A232)  and  A200 );
 a12474a <=( (not A300)  and  (not A299) );
 a12475a <=( A233  and  a12474a );
 a12476a <=( a12475a  and  a12470a );
 a12479a <=( (not A168)  and  (not A170) );
 a12483a <=( (not A199)  and  A166 );
 a12484a <=( (not A167)  and  a12483a );
 a12485a <=( a12484a  and  a12479a );
 a12488a <=( (not A232)  and  A200 );
 a12492a <=( A299  and  A298 );
 a12493a <=( A233  and  a12492a );
 a12494a <=( a12493a  and  a12488a );
 a12497a <=( (not A168)  and  (not A170) );
 a12501a <=( (not A199)  and  A166 );
 a12502a <=( (not A167)  and  a12501a );
 a12503a <=( a12502a  and  a12497a );
 a12506a <=( (not A232)  and  A200 );
 a12510a <=( (not A299)  and  (not A298) );
 a12511a <=( A233  and  a12510a );
 a12512a <=( a12511a  and  a12506a );
 a12515a <=( (not A168)  and  (not A170) );
 a12519a <=( (not A199)  and  A166 );
 a12520a <=( (not A167)  and  a12519a );
 a12521a <=( a12520a  and  a12515a );
 a12524a <=( (not A232)  and  A200 );
 a12528a <=( A266  and  (not A265) );
 a12529a <=( A233  and  a12528a );
 a12530a <=( a12529a  and  a12524a );
 a12533a <=( (not A168)  and  A169 );
 a12537a <=( (not A199)  and  (not A166) );
 a12538a <=( A167  and  a12537a );
 a12539a <=( a12538a  and  a12533a );
 a12542a <=( (not A232)  and  A200 );
 a12546a <=( (not A300)  and  (not A299) );
 a12547a <=( A233  and  a12546a );
 a12548a <=( a12547a  and  a12542a );
 a12551a <=( (not A168)  and  A169 );
 a12555a <=( (not A199)  and  (not A166) );
 a12556a <=( A167  and  a12555a );
 a12557a <=( a12556a  and  a12551a );
 a12560a <=( (not A232)  and  A200 );
 a12564a <=( A299  and  A298 );
 a12565a <=( A233  and  a12564a );
 a12566a <=( a12565a  and  a12560a );
 a12569a <=( (not A168)  and  A169 );
 a12573a <=( (not A199)  and  (not A166) );
 a12574a <=( A167  and  a12573a );
 a12575a <=( a12574a  and  a12569a );
 a12578a <=( (not A232)  and  A200 );
 a12582a <=( (not A299)  and  (not A298) );
 a12583a <=( A233  and  a12582a );
 a12584a <=( a12583a  and  a12578a );
 a12587a <=( (not A168)  and  A169 );
 a12591a <=( (not A199)  and  (not A166) );
 a12592a <=( A167  and  a12591a );
 a12593a <=( a12592a  and  a12587a );
 a12596a <=( (not A232)  and  A200 );
 a12600a <=( A266  and  (not A265) );
 a12601a <=( A233  and  a12600a );
 a12602a <=( a12601a  and  a12596a );
 a12605a <=( (not A168)  and  A169 );
 a12609a <=( (not A199)  and  A166 );
 a12610a <=( (not A167)  and  a12609a );
 a12611a <=( a12610a  and  a12605a );
 a12614a <=( (not A232)  and  A200 );
 a12618a <=( (not A300)  and  (not A299) );
 a12619a <=( A233  and  a12618a );
 a12620a <=( a12619a  and  a12614a );
 a12623a <=( (not A168)  and  A169 );
 a12627a <=( (not A199)  and  A166 );
 a12628a <=( (not A167)  and  a12627a );
 a12629a <=( a12628a  and  a12623a );
 a12632a <=( (not A232)  and  A200 );
 a12636a <=( A299  and  A298 );
 a12637a <=( A233  and  a12636a );
 a12638a <=( a12637a  and  a12632a );
 a12641a <=( (not A168)  and  A169 );
 a12645a <=( (not A199)  and  A166 );
 a12646a <=( (not A167)  and  a12645a );
 a12647a <=( a12646a  and  a12641a );
 a12650a <=( (not A232)  and  A200 );
 a12654a <=( (not A299)  and  (not A298) );
 a12655a <=( A233  and  a12654a );
 a12656a <=( a12655a  and  a12650a );
 a12659a <=( (not A168)  and  A169 );
 a12663a <=( (not A199)  and  A166 );
 a12664a <=( (not A167)  and  a12663a );
 a12665a <=( a12664a  and  a12659a );
 a12668a <=( (not A232)  and  A200 );
 a12672a <=( A266  and  (not A265) );
 a12673a <=( A233  and  a12672a );
 a12674a <=( a12673a  and  a12668a );
 a12677a <=( A169  and  (not A170) );
 a12681a <=( A199  and  A166 );
 a12682a <=( A167  and  a12681a );
 a12683a <=( a12682a  and  a12677a );
 a12686a <=( (not A232)  and  A200 );
 a12690a <=( (not A300)  and  (not A299) );
 a12691a <=( A233  and  a12690a );
 a12692a <=( a12691a  and  a12686a );
 a12695a <=( A169  and  (not A170) );
 a12699a <=( A199  and  A166 );
 a12700a <=( A167  and  a12699a );
 a12701a <=( a12700a  and  a12695a );
 a12704a <=( (not A232)  and  A200 );
 a12708a <=( A299  and  A298 );
 a12709a <=( A233  and  a12708a );
 a12710a <=( a12709a  and  a12704a );
 a12713a <=( A169  and  (not A170) );
 a12717a <=( A199  and  A166 );
 a12718a <=( A167  and  a12717a );
 a12719a <=( a12718a  and  a12713a );
 a12722a <=( (not A232)  and  A200 );
 a12726a <=( (not A299)  and  (not A298) );
 a12727a <=( A233  and  a12726a );
 a12728a <=( a12727a  and  a12722a );
 a12731a <=( A169  and  (not A170) );
 a12735a <=( A199  and  A166 );
 a12736a <=( A167  and  a12735a );
 a12737a <=( a12736a  and  a12731a );
 a12740a <=( (not A232)  and  A200 );
 a12744a <=( A266  and  (not A265) );
 a12745a <=( A233  and  a12744a );
 a12746a <=( a12745a  and  a12740a );
 a12749a <=( A169  and  (not A170) );
 a12753a <=( (not A200)  and  A166 );
 a12754a <=( A167  and  a12753a );
 a12755a <=( a12754a  and  a12749a );
 a12758a <=( (not A232)  and  (not A201) );
 a12762a <=( (not A300)  and  (not A299) );
 a12763a <=( A233  and  a12762a );
 a12764a <=( a12763a  and  a12758a );
 a12767a <=( A169  and  (not A170) );
 a12771a <=( (not A200)  and  A166 );
 a12772a <=( A167  and  a12771a );
 a12773a <=( a12772a  and  a12767a );
 a12776a <=( (not A232)  and  (not A201) );
 a12780a <=( A299  and  A298 );
 a12781a <=( A233  and  a12780a );
 a12782a <=( a12781a  and  a12776a );
 a12785a <=( A169  and  (not A170) );
 a12789a <=( (not A200)  and  A166 );
 a12790a <=( A167  and  a12789a );
 a12791a <=( a12790a  and  a12785a );
 a12794a <=( (not A232)  and  (not A201) );
 a12798a <=( (not A299)  and  (not A298) );
 a12799a <=( A233  and  a12798a );
 a12800a <=( a12799a  and  a12794a );
 a12803a <=( A169  and  (not A170) );
 a12807a <=( (not A200)  and  A166 );
 a12808a <=( A167  and  a12807a );
 a12809a <=( a12808a  and  a12803a );
 a12812a <=( (not A232)  and  (not A201) );
 a12816a <=( A266  and  (not A265) );
 a12817a <=( A233  and  a12816a );
 a12818a <=( a12817a  and  a12812a );
 a12821a <=( A169  and  (not A170) );
 a12825a <=( (not A199)  and  A166 );
 a12826a <=( A167  and  a12825a );
 a12827a <=( a12826a  and  a12821a );
 a12830a <=( (not A232)  and  (not A200) );
 a12834a <=( (not A300)  and  (not A299) );
 a12835a <=( A233  and  a12834a );
 a12836a <=( a12835a  and  a12830a );
 a12839a <=( A169  and  (not A170) );
 a12843a <=( (not A199)  and  A166 );
 a12844a <=( A167  and  a12843a );
 a12845a <=( a12844a  and  a12839a );
 a12848a <=( (not A232)  and  (not A200) );
 a12852a <=( A299  and  A298 );
 a12853a <=( A233  and  a12852a );
 a12854a <=( a12853a  and  a12848a );
 a12857a <=( A169  and  (not A170) );
 a12861a <=( (not A199)  and  A166 );
 a12862a <=( A167  and  a12861a );
 a12863a <=( a12862a  and  a12857a );
 a12866a <=( (not A232)  and  (not A200) );
 a12870a <=( (not A299)  and  (not A298) );
 a12871a <=( A233  and  a12870a );
 a12872a <=( a12871a  and  a12866a );
 a12875a <=( A169  and  (not A170) );
 a12879a <=( (not A199)  and  A166 );
 a12880a <=( A167  and  a12879a );
 a12881a <=( a12880a  and  a12875a );
 a12884a <=( (not A232)  and  (not A200) );
 a12888a <=( A266  and  (not A265) );
 a12889a <=( A233  and  a12888a );
 a12890a <=( a12889a  and  a12884a );
 a12893a <=( A169  and  (not A170) );
 a12897a <=( A199  and  (not A166) );
 a12898a <=( (not A167)  and  a12897a );
 a12899a <=( a12898a  and  a12893a );
 a12902a <=( (not A232)  and  A200 );
 a12906a <=( (not A300)  and  (not A299) );
 a12907a <=( A233  and  a12906a );
 a12908a <=( a12907a  and  a12902a );
 a12911a <=( A169  and  (not A170) );
 a12915a <=( A199  and  (not A166) );
 a12916a <=( (not A167)  and  a12915a );
 a12917a <=( a12916a  and  a12911a );
 a12920a <=( (not A232)  and  A200 );
 a12924a <=( A299  and  A298 );
 a12925a <=( A233  and  a12924a );
 a12926a <=( a12925a  and  a12920a );
 a12929a <=( A169  and  (not A170) );
 a12933a <=( A199  and  (not A166) );
 a12934a <=( (not A167)  and  a12933a );
 a12935a <=( a12934a  and  a12929a );
 a12938a <=( (not A232)  and  A200 );
 a12942a <=( (not A299)  and  (not A298) );
 a12943a <=( A233  and  a12942a );
 a12944a <=( a12943a  and  a12938a );
 a12947a <=( A169  and  (not A170) );
 a12951a <=( A199  and  (not A166) );
 a12952a <=( (not A167)  and  a12951a );
 a12953a <=( a12952a  and  a12947a );
 a12956a <=( (not A232)  and  A200 );
 a12960a <=( A266  and  (not A265) );
 a12961a <=( A233  and  a12960a );
 a12962a <=( a12961a  and  a12956a );
 a12965a <=( A169  and  (not A170) );
 a12969a <=( (not A200)  and  (not A166) );
 a12970a <=( (not A167)  and  a12969a );
 a12971a <=( a12970a  and  a12965a );
 a12974a <=( (not A232)  and  (not A201) );
 a12978a <=( (not A300)  and  (not A299) );
 a12979a <=( A233  and  a12978a );
 a12980a <=( a12979a  and  a12974a );
 a12983a <=( A169  and  (not A170) );
 a12987a <=( (not A200)  and  (not A166) );
 a12988a <=( (not A167)  and  a12987a );
 a12989a <=( a12988a  and  a12983a );
 a12992a <=( (not A232)  and  (not A201) );
 a12996a <=( A299  and  A298 );
 a12997a <=( A233  and  a12996a );
 a12998a <=( a12997a  and  a12992a );
 a13001a <=( A169  and  (not A170) );
 a13005a <=( (not A200)  and  (not A166) );
 a13006a <=( (not A167)  and  a13005a );
 a13007a <=( a13006a  and  a13001a );
 a13010a <=( (not A232)  and  (not A201) );
 a13014a <=( (not A299)  and  (not A298) );
 a13015a <=( A233  and  a13014a );
 a13016a <=( a13015a  and  a13010a );
 a13019a <=( A169  and  (not A170) );
 a13023a <=( (not A200)  and  (not A166) );
 a13024a <=( (not A167)  and  a13023a );
 a13025a <=( a13024a  and  a13019a );
 a13028a <=( (not A232)  and  (not A201) );
 a13032a <=( A266  and  (not A265) );
 a13033a <=( A233  and  a13032a );
 a13034a <=( a13033a  and  a13028a );
 a13037a <=( A169  and  (not A170) );
 a13041a <=( (not A199)  and  (not A166) );
 a13042a <=( (not A167)  and  a13041a );
 a13043a <=( a13042a  and  a13037a );
 a13046a <=( (not A232)  and  (not A200) );
 a13050a <=( (not A300)  and  (not A299) );
 a13051a <=( A233  and  a13050a );
 a13052a <=( a13051a  and  a13046a );
 a13055a <=( A169  and  (not A170) );
 a13059a <=( (not A199)  and  (not A166) );
 a13060a <=( (not A167)  and  a13059a );
 a13061a <=( a13060a  and  a13055a );
 a13064a <=( (not A232)  and  (not A200) );
 a13068a <=( A299  and  A298 );
 a13069a <=( A233  and  a13068a );
 a13070a <=( a13069a  and  a13064a );
 a13073a <=( A169  and  (not A170) );
 a13077a <=( (not A199)  and  (not A166) );
 a13078a <=( (not A167)  and  a13077a );
 a13079a <=( a13078a  and  a13073a );
 a13082a <=( (not A232)  and  (not A200) );
 a13086a <=( (not A299)  and  (not A298) );
 a13087a <=( A233  and  a13086a );
 a13088a <=( a13087a  and  a13082a );
 a13091a <=( A169  and  (not A170) );
 a13095a <=( (not A199)  and  (not A166) );
 a13096a <=( (not A167)  and  a13095a );
 a13097a <=( a13096a  and  a13091a );
 a13100a <=( (not A232)  and  (not A200) );
 a13104a <=( A266  and  (not A265) );
 a13105a <=( A233  and  a13104a );
 a13106a <=( a13105a  and  a13100a );
 a13109a <=( (not A167)  and  (not A169) );
 a13113a <=( A200  and  (not A199) );
 a13114a <=( (not A166)  and  a13113a );
 a13115a <=( a13114a  and  a13109a );
 a13118a <=( A233  and  (not A232) );
 a13122a <=( (not A302)  and  (not A301) );
 a13123a <=( (not A299)  and  a13122a );
 a13124a <=( a13123a  and  a13118a );
 a13127a <=( (not A168)  and  (not A169) );
 a13131a <=( (not A199)  and  A166 );
 a13132a <=( A167  and  a13131a );
 a13133a <=( a13132a  and  a13127a );
 a13136a <=( (not A232)  and  A200 );
 a13140a <=( (not A300)  and  (not A299) );
 a13141a <=( A233  and  a13140a );
 a13142a <=( a13141a  and  a13136a );
 a13145a <=( (not A168)  and  (not A169) );
 a13149a <=( (not A199)  and  A166 );
 a13150a <=( A167  and  a13149a );
 a13151a <=( a13150a  and  a13145a );
 a13154a <=( (not A232)  and  A200 );
 a13158a <=( A299  and  A298 );
 a13159a <=( A233  and  a13158a );
 a13160a <=( a13159a  and  a13154a );
 a13163a <=( (not A168)  and  (not A169) );
 a13167a <=( (not A199)  and  A166 );
 a13168a <=( A167  and  a13167a );
 a13169a <=( a13168a  and  a13163a );
 a13172a <=( (not A232)  and  A200 );
 a13176a <=( (not A299)  and  (not A298) );
 a13177a <=( A233  and  a13176a );
 a13178a <=( a13177a  and  a13172a );
 a13181a <=( (not A168)  and  (not A169) );
 a13185a <=( (not A199)  and  A166 );
 a13186a <=( A167  and  a13185a );
 a13187a <=( a13186a  and  a13181a );
 a13190a <=( (not A232)  and  A200 );
 a13194a <=( A266  and  (not A265) );
 a13195a <=( A233  and  a13194a );
 a13196a <=( a13195a  and  a13190a );
 a13199a <=( (not A169)  and  A170 );
 a13203a <=( A199  and  (not A166) );
 a13204a <=( A167  and  a13203a );
 a13205a <=( a13204a  and  a13199a );
 a13208a <=( (not A232)  and  A200 );
 a13212a <=( (not A300)  and  (not A299) );
 a13213a <=( A233  and  a13212a );
 a13214a <=( a13213a  and  a13208a );
 a13217a <=( (not A169)  and  A170 );
 a13221a <=( A199  and  (not A166) );
 a13222a <=( A167  and  a13221a );
 a13223a <=( a13222a  and  a13217a );
 a13226a <=( (not A232)  and  A200 );
 a13230a <=( A299  and  A298 );
 a13231a <=( A233  and  a13230a );
 a13232a <=( a13231a  and  a13226a );
 a13235a <=( (not A169)  and  A170 );
 a13239a <=( A199  and  (not A166) );
 a13240a <=( A167  and  a13239a );
 a13241a <=( a13240a  and  a13235a );
 a13244a <=( (not A232)  and  A200 );
 a13248a <=( (not A299)  and  (not A298) );
 a13249a <=( A233  and  a13248a );
 a13250a <=( a13249a  and  a13244a );
 a13253a <=( (not A169)  and  A170 );
 a13257a <=( A199  and  (not A166) );
 a13258a <=( A167  and  a13257a );
 a13259a <=( a13258a  and  a13253a );
 a13262a <=( (not A232)  and  A200 );
 a13266a <=( A266  and  (not A265) );
 a13267a <=( A233  and  a13266a );
 a13268a <=( a13267a  and  a13262a );
 a13271a <=( (not A169)  and  A170 );
 a13275a <=( (not A200)  and  (not A166) );
 a13276a <=( A167  and  a13275a );
 a13277a <=( a13276a  and  a13271a );
 a13280a <=( (not A232)  and  (not A201) );
 a13284a <=( (not A300)  and  (not A299) );
 a13285a <=( A233  and  a13284a );
 a13286a <=( a13285a  and  a13280a );
 a13289a <=( (not A169)  and  A170 );
 a13293a <=( (not A200)  and  (not A166) );
 a13294a <=( A167  and  a13293a );
 a13295a <=( a13294a  and  a13289a );
 a13298a <=( (not A232)  and  (not A201) );
 a13302a <=( A299  and  A298 );
 a13303a <=( A233  and  a13302a );
 a13304a <=( a13303a  and  a13298a );
 a13307a <=( (not A169)  and  A170 );
 a13311a <=( (not A200)  and  (not A166) );
 a13312a <=( A167  and  a13311a );
 a13313a <=( a13312a  and  a13307a );
 a13316a <=( (not A232)  and  (not A201) );
 a13320a <=( (not A299)  and  (not A298) );
 a13321a <=( A233  and  a13320a );
 a13322a <=( a13321a  and  a13316a );
 a13325a <=( (not A169)  and  A170 );
 a13329a <=( (not A200)  and  (not A166) );
 a13330a <=( A167  and  a13329a );
 a13331a <=( a13330a  and  a13325a );
 a13334a <=( (not A232)  and  (not A201) );
 a13338a <=( A266  and  (not A265) );
 a13339a <=( A233  and  a13338a );
 a13340a <=( a13339a  and  a13334a );
 a13343a <=( (not A169)  and  A170 );
 a13347a <=( (not A199)  and  (not A166) );
 a13348a <=( A167  and  a13347a );
 a13349a <=( a13348a  and  a13343a );
 a13352a <=( (not A232)  and  (not A200) );
 a13356a <=( (not A300)  and  (not A299) );
 a13357a <=( A233  and  a13356a );
 a13358a <=( a13357a  and  a13352a );
 a13361a <=( (not A169)  and  A170 );
 a13365a <=( (not A199)  and  (not A166) );
 a13366a <=( A167  and  a13365a );
 a13367a <=( a13366a  and  a13361a );
 a13370a <=( (not A232)  and  (not A200) );
 a13374a <=( A299  and  A298 );
 a13375a <=( A233  and  a13374a );
 a13376a <=( a13375a  and  a13370a );
 a13379a <=( (not A169)  and  A170 );
 a13383a <=( (not A199)  and  (not A166) );
 a13384a <=( A167  and  a13383a );
 a13385a <=( a13384a  and  a13379a );
 a13388a <=( (not A232)  and  (not A200) );
 a13392a <=( (not A299)  and  (not A298) );
 a13393a <=( A233  and  a13392a );
 a13394a <=( a13393a  and  a13388a );
 a13397a <=( (not A169)  and  A170 );
 a13401a <=( (not A199)  and  (not A166) );
 a13402a <=( A167  and  a13401a );
 a13403a <=( a13402a  and  a13397a );
 a13406a <=( (not A232)  and  (not A200) );
 a13410a <=( A266  and  (not A265) );
 a13411a <=( A233  and  a13410a );
 a13412a <=( a13411a  and  a13406a );
 a13415a <=( (not A169)  and  A170 );
 a13419a <=( A199  and  A166 );
 a13420a <=( (not A167)  and  a13419a );
 a13421a <=( a13420a  and  a13415a );
 a13424a <=( (not A232)  and  A200 );
 a13428a <=( (not A300)  and  (not A299) );
 a13429a <=( A233  and  a13428a );
 a13430a <=( a13429a  and  a13424a );
 a13433a <=( (not A169)  and  A170 );
 a13437a <=( A199  and  A166 );
 a13438a <=( (not A167)  and  a13437a );
 a13439a <=( a13438a  and  a13433a );
 a13442a <=( (not A232)  and  A200 );
 a13446a <=( A299  and  A298 );
 a13447a <=( A233  and  a13446a );
 a13448a <=( a13447a  and  a13442a );
 a13451a <=( (not A169)  and  A170 );
 a13455a <=( A199  and  A166 );
 a13456a <=( (not A167)  and  a13455a );
 a13457a <=( a13456a  and  a13451a );
 a13460a <=( (not A232)  and  A200 );
 a13464a <=( (not A299)  and  (not A298) );
 a13465a <=( A233  and  a13464a );
 a13466a <=( a13465a  and  a13460a );
 a13469a <=( (not A169)  and  A170 );
 a13473a <=( A199  and  A166 );
 a13474a <=( (not A167)  and  a13473a );
 a13475a <=( a13474a  and  a13469a );
 a13478a <=( (not A232)  and  A200 );
 a13482a <=( A266  and  (not A265) );
 a13483a <=( A233  and  a13482a );
 a13484a <=( a13483a  and  a13478a );
 a13487a <=( (not A169)  and  A170 );
 a13491a <=( (not A200)  and  A166 );
 a13492a <=( (not A167)  and  a13491a );
 a13493a <=( a13492a  and  a13487a );
 a13496a <=( (not A232)  and  (not A201) );
 a13500a <=( (not A300)  and  (not A299) );
 a13501a <=( A233  and  a13500a );
 a13502a <=( a13501a  and  a13496a );
 a13505a <=( (not A169)  and  A170 );
 a13509a <=( (not A200)  and  A166 );
 a13510a <=( (not A167)  and  a13509a );
 a13511a <=( a13510a  and  a13505a );
 a13514a <=( (not A232)  and  (not A201) );
 a13518a <=( A299  and  A298 );
 a13519a <=( A233  and  a13518a );
 a13520a <=( a13519a  and  a13514a );
 a13523a <=( (not A169)  and  A170 );
 a13527a <=( (not A200)  and  A166 );
 a13528a <=( (not A167)  and  a13527a );
 a13529a <=( a13528a  and  a13523a );
 a13532a <=( (not A232)  and  (not A201) );
 a13536a <=( (not A299)  and  (not A298) );
 a13537a <=( A233  and  a13536a );
 a13538a <=( a13537a  and  a13532a );
 a13541a <=( (not A169)  and  A170 );
 a13545a <=( (not A200)  and  A166 );
 a13546a <=( (not A167)  and  a13545a );
 a13547a <=( a13546a  and  a13541a );
 a13550a <=( (not A232)  and  (not A201) );
 a13554a <=( A266  and  (not A265) );
 a13555a <=( A233  and  a13554a );
 a13556a <=( a13555a  and  a13550a );
 a13559a <=( (not A169)  and  A170 );
 a13563a <=( (not A199)  and  A166 );
 a13564a <=( (not A167)  and  a13563a );
 a13565a <=( a13564a  and  a13559a );
 a13568a <=( (not A232)  and  (not A200) );
 a13572a <=( (not A300)  and  (not A299) );
 a13573a <=( A233  and  a13572a );
 a13574a <=( a13573a  and  a13568a );
 a13577a <=( (not A169)  and  A170 );
 a13581a <=( (not A199)  and  A166 );
 a13582a <=( (not A167)  and  a13581a );
 a13583a <=( a13582a  and  a13577a );
 a13586a <=( (not A232)  and  (not A200) );
 a13590a <=( A299  and  A298 );
 a13591a <=( A233  and  a13590a );
 a13592a <=( a13591a  and  a13586a );
 a13595a <=( (not A169)  and  A170 );
 a13599a <=( (not A199)  and  A166 );
 a13600a <=( (not A167)  and  a13599a );
 a13601a <=( a13600a  and  a13595a );
 a13604a <=( (not A232)  and  (not A200) );
 a13608a <=( (not A299)  and  (not A298) );
 a13609a <=( A233  and  a13608a );
 a13610a <=( a13609a  and  a13604a );
 a13613a <=( (not A169)  and  A170 );
 a13617a <=( (not A199)  and  A166 );
 a13618a <=( (not A167)  and  a13617a );
 a13619a <=( a13618a  and  a13613a );
 a13622a <=( (not A232)  and  (not A200) );
 a13626a <=( A266  and  (not A265) );
 a13627a <=( A233  and  a13626a );
 a13628a <=( a13627a  and  a13622a );
 a13631a <=( A166  and  A168 );
 a13635a <=( A232  and  A200 );
 a13636a <=( A199  and  a13635a );
 a13637a <=( a13636a  and  a13631a );
 a13641a <=( (not A268)  and  A265 );
 a13642a <=( A233  and  a13641a );
 a13646a <=( A299  and  (not A298) );
 a13647a <=( (not A269)  and  a13646a );
 a13648a <=( a13647a  and  a13642a );
 a13651a <=( A166  and  A168 );
 a13655a <=( (not A233)  and  A200 );
 a13656a <=( A199  and  a13655a );
 a13657a <=( a13656a  and  a13651a );
 a13661a <=( A265  and  (not A236) );
 a13662a <=( (not A235)  and  a13661a );
 a13666a <=( A299  and  (not A298) );
 a13667a <=( A266  and  a13666a );
 a13668a <=( a13667a  and  a13662a );
 a13671a <=( A166  and  A168 );
 a13675a <=( (not A233)  and  A200 );
 a13676a <=( A199  and  a13675a );
 a13677a <=( a13676a  and  a13671a );
 a13681a <=( (not A266)  and  (not A236) );
 a13682a <=( (not A235)  and  a13681a );
 a13686a <=( A299  and  (not A298) );
 a13687a <=( (not A267)  and  a13686a );
 a13688a <=( a13687a  and  a13682a );
 a13691a <=( A166  and  A168 );
 a13695a <=( (not A233)  and  A200 );
 a13696a <=( A199  and  a13695a );
 a13697a <=( a13696a  and  a13691a );
 a13701a <=( (not A265)  and  (not A236) );
 a13702a <=( (not A235)  and  a13701a );
 a13706a <=( A299  and  (not A298) );
 a13707a <=( (not A266)  and  a13706a );
 a13708a <=( a13707a  and  a13702a );
 a13711a <=( A166  and  A168 );
 a13715a <=( (not A233)  and  A200 );
 a13716a <=( A199  and  a13715a );
 a13717a <=( a13716a  and  a13711a );
 a13721a <=( (not A268)  and  (not A266) );
 a13722a <=( (not A234)  and  a13721a );
 a13726a <=( A299  and  (not A298) );
 a13727a <=( (not A269)  and  a13726a );
 a13728a <=( a13727a  and  a13722a );
 a13731a <=( A166  and  A168 );
 a13735a <=( A232  and  A200 );
 a13736a <=( A199  and  a13735a );
 a13737a <=( a13736a  and  a13731a );
 a13741a <=( A235  and  A234 );
 a13742a <=( (not A233)  and  a13741a );
 a13746a <=( (not A302)  and  (not A301) );
 a13747a <=( A298  and  a13746a );
 a13748a <=( a13747a  and  a13742a );
 a13751a <=( A166  and  A168 );
 a13755a <=( A232  and  A200 );
 a13756a <=( A199  and  a13755a );
 a13757a <=( a13756a  and  a13751a );
 a13761a <=( A236  and  A234 );
 a13762a <=( (not A233)  and  a13761a );
 a13766a <=( (not A302)  and  (not A301) );
 a13767a <=( A298  and  a13766a );
 a13768a <=( a13767a  and  a13762a );
 a13771a <=( A166  and  A168 );
 a13775a <=( (not A232)  and  A200 );
 a13776a <=( A199  and  a13775a );
 a13777a <=( a13776a  and  a13771a );
 a13781a <=( (not A268)  and  (not A266) );
 a13782a <=( (not A233)  and  a13781a );
 a13786a <=( A299  and  (not A298) );
 a13787a <=( (not A269)  and  a13786a );
 a13788a <=( a13787a  and  a13782a );
 a13791a <=( A166  and  A168 );
 a13795a <=( (not A203)  and  (not A202) );
 a13796a <=( (not A200)  and  a13795a );
 a13797a <=( a13796a  and  a13791a );
 a13801a <=( A265  and  A233 );
 a13802a <=( A232  and  a13801a );
 a13806a <=( A299  and  (not A298) );
 a13807a <=( (not A267)  and  a13806a );
 a13808a <=( a13807a  and  a13802a );
 a13811a <=( A166  and  A168 );
 a13815a <=( (not A203)  and  (not A202) );
 a13816a <=( (not A200)  and  a13815a );
 a13817a <=( a13816a  and  a13811a );
 a13821a <=( A265  and  A233 );
 a13822a <=( A232  and  a13821a );
 a13826a <=( A299  and  (not A298) );
 a13827a <=( A266  and  a13826a );
 a13828a <=( a13827a  and  a13822a );
 a13831a <=( A166  and  A168 );
 a13835a <=( (not A203)  and  (not A202) );
 a13836a <=( (not A200)  and  a13835a );
 a13837a <=( a13836a  and  a13831a );
 a13841a <=( (not A265)  and  A233 );
 a13842a <=( A232  and  a13841a );
 a13846a <=( A299  and  (not A298) );
 a13847a <=( (not A266)  and  a13846a );
 a13848a <=( a13847a  and  a13842a );
 a13851a <=( A166  and  A168 );
 a13855a <=( (not A203)  and  (not A202) );
 a13856a <=( (not A200)  and  a13855a );
 a13857a <=( a13856a  and  a13851a );
 a13861a <=( A265  and  A233 );
 a13862a <=( (not A232)  and  a13861a );
 a13866a <=( A268  and  A267 );
 a13867a <=( (not A266)  and  a13866a );
 a13868a <=( a13867a  and  a13862a );
 a13871a <=( A166  and  A168 );
 a13875a <=( (not A203)  and  (not A202) );
 a13876a <=( (not A200)  and  a13875a );
 a13877a <=( a13876a  and  a13871a );
 a13881a <=( A265  and  A233 );
 a13882a <=( (not A232)  and  a13881a );
 a13886a <=( A269  and  A267 );
 a13887a <=( (not A266)  and  a13886a );
 a13888a <=( a13887a  and  a13882a );
 a13891a <=( A166  and  A168 );
 a13895a <=( (not A203)  and  (not A202) );
 a13896a <=( (not A200)  and  a13895a );
 a13897a <=( a13896a  and  a13891a );
 a13901a <=( A265  and  (not A234) );
 a13902a <=( (not A233)  and  a13901a );
 a13906a <=( A299  and  (not A298) );
 a13907a <=( A266  and  a13906a );
 a13908a <=( a13907a  and  a13902a );
 a13911a <=( A166  and  A168 );
 a13915a <=( (not A203)  and  (not A202) );
 a13916a <=( (not A200)  and  a13915a );
 a13917a <=( a13916a  and  a13911a );
 a13921a <=( (not A266)  and  (not A234) );
 a13922a <=( (not A233)  and  a13921a );
 a13926a <=( A299  and  (not A298) );
 a13927a <=( (not A267)  and  a13926a );
 a13928a <=( a13927a  and  a13922a );
 a13931a <=( A166  and  A168 );
 a13935a <=( (not A203)  and  (not A202) );
 a13936a <=( (not A200)  and  a13935a );
 a13937a <=( a13936a  and  a13931a );
 a13941a <=( (not A265)  and  (not A234) );
 a13942a <=( (not A233)  and  a13941a );
 a13946a <=( A299  and  (not A298) );
 a13947a <=( (not A266)  and  a13946a );
 a13948a <=( a13947a  and  a13942a );
 a13951a <=( A166  and  A168 );
 a13955a <=( (not A203)  and  (not A202) );
 a13956a <=( (not A200)  and  a13955a );
 a13957a <=( a13956a  and  a13951a );
 a13961a <=( A234  and  (not A233) );
 a13962a <=( A232  and  a13961a );
 a13966a <=( (not A300)  and  A298 );
 a13967a <=( A235  and  a13966a );
 a13968a <=( a13967a  and  a13962a );
 a13971a <=( A166  and  A168 );
 a13975a <=( (not A203)  and  (not A202) );
 a13976a <=( (not A200)  and  a13975a );
 a13977a <=( a13976a  and  a13971a );
 a13981a <=( A234  and  (not A233) );
 a13982a <=( A232  and  a13981a );
 a13986a <=( A299  and  A298 );
 a13987a <=( A235  and  a13986a );
 a13988a <=( a13987a  and  a13982a );
 a13991a <=( A166  and  A168 );
 a13995a <=( (not A203)  and  (not A202) );
 a13996a <=( (not A200)  and  a13995a );
 a13997a <=( a13996a  and  a13991a );
 a14001a <=( A234  and  (not A233) );
 a14002a <=( A232  and  a14001a );
 a14006a <=( (not A299)  and  (not A298) );
 a14007a <=( A235  and  a14006a );
 a14008a <=( a14007a  and  a14002a );
 a14011a <=( A166  and  A168 );
 a14015a <=( (not A203)  and  (not A202) );
 a14016a <=( (not A200)  and  a14015a );
 a14017a <=( a14016a  and  a14011a );
 a14021a <=( A234  and  (not A233) );
 a14022a <=( A232  and  a14021a );
 a14026a <=( A266  and  (not A265) );
 a14027a <=( A235  and  a14026a );
 a14028a <=( a14027a  and  a14022a );
 a14031a <=( A166  and  A168 );
 a14035a <=( (not A203)  and  (not A202) );
 a14036a <=( (not A200)  and  a14035a );
 a14037a <=( a14036a  and  a14031a );
 a14041a <=( A234  and  (not A233) );
 a14042a <=( A232  and  a14041a );
 a14046a <=( (not A300)  and  A298 );
 a14047a <=( A236  and  a14046a );
 a14048a <=( a14047a  and  a14042a );
 a14051a <=( A166  and  A168 );
 a14055a <=( (not A203)  and  (not A202) );
 a14056a <=( (not A200)  and  a14055a );
 a14057a <=( a14056a  and  a14051a );
 a14061a <=( A234  and  (not A233) );
 a14062a <=( A232  and  a14061a );
 a14066a <=( A299  and  A298 );
 a14067a <=( A236  and  a14066a );
 a14068a <=( a14067a  and  a14062a );
 a14071a <=( A166  and  A168 );
 a14075a <=( (not A203)  and  (not A202) );
 a14076a <=( (not A200)  and  a14075a );
 a14077a <=( a14076a  and  a14071a );
 a14081a <=( A234  and  (not A233) );
 a14082a <=( A232  and  a14081a );
 a14086a <=( (not A299)  and  (not A298) );
 a14087a <=( A236  and  a14086a );
 a14088a <=( a14087a  and  a14082a );
 a14091a <=( A166  and  A168 );
 a14095a <=( (not A203)  and  (not A202) );
 a14096a <=( (not A200)  and  a14095a );
 a14097a <=( a14096a  and  a14091a );
 a14101a <=( A234  and  (not A233) );
 a14102a <=( A232  and  a14101a );
 a14106a <=( A266  and  (not A265) );
 a14107a <=( A236  and  a14106a );
 a14108a <=( a14107a  and  a14102a );
 a14111a <=( A166  and  A168 );
 a14115a <=( (not A203)  and  (not A202) );
 a14116a <=( (not A200)  and  a14115a );
 a14117a <=( a14116a  and  a14111a );
 a14121a <=( A265  and  (not A233) );
 a14122a <=( (not A232)  and  a14121a );
 a14126a <=( A299  and  (not A298) );
 a14127a <=( A266  and  a14126a );
 a14128a <=( a14127a  and  a14122a );
 a14131a <=( A166  and  A168 );
 a14135a <=( (not A203)  and  (not A202) );
 a14136a <=( (not A200)  and  a14135a );
 a14137a <=( a14136a  and  a14131a );
 a14141a <=( (not A266)  and  (not A233) );
 a14142a <=( (not A232)  and  a14141a );
 a14146a <=( A299  and  (not A298) );
 a14147a <=( (not A267)  and  a14146a );
 a14148a <=( a14147a  and  a14142a );
 a14151a <=( A166  and  A168 );
 a14155a <=( (not A203)  and  (not A202) );
 a14156a <=( (not A200)  and  a14155a );
 a14157a <=( a14156a  and  a14151a );
 a14161a <=( (not A265)  and  (not A233) );
 a14162a <=( (not A232)  and  a14161a );
 a14166a <=( A299  and  (not A298) );
 a14167a <=( (not A266)  and  a14166a );
 a14168a <=( a14167a  and  a14162a );
 a14171a <=( A166  and  A168 );
 a14175a <=( A232  and  (not A201) );
 a14176a <=( (not A200)  and  a14175a );
 a14177a <=( a14176a  and  a14171a );
 a14181a <=( (not A268)  and  A265 );
 a14182a <=( A233  and  a14181a );
 a14186a <=( A299  and  (not A298) );
 a14187a <=( (not A269)  and  a14186a );
 a14188a <=( a14187a  and  a14182a );
 a14191a <=( A166  and  A168 );
 a14195a <=( (not A233)  and  (not A201) );
 a14196a <=( (not A200)  and  a14195a );
 a14197a <=( a14196a  and  a14191a );
 a14201a <=( A265  and  (not A236) );
 a14202a <=( (not A235)  and  a14201a );
 a14206a <=( A299  and  (not A298) );
 a14207a <=( A266  and  a14206a );
 a14208a <=( a14207a  and  a14202a );
 a14211a <=( A166  and  A168 );
 a14215a <=( (not A233)  and  (not A201) );
 a14216a <=( (not A200)  and  a14215a );
 a14217a <=( a14216a  and  a14211a );
 a14221a <=( (not A266)  and  (not A236) );
 a14222a <=( (not A235)  and  a14221a );
 a14226a <=( A299  and  (not A298) );
 a14227a <=( (not A267)  and  a14226a );
 a14228a <=( a14227a  and  a14222a );
 a14231a <=( A166  and  A168 );
 a14235a <=( (not A233)  and  (not A201) );
 a14236a <=( (not A200)  and  a14235a );
 a14237a <=( a14236a  and  a14231a );
 a14241a <=( (not A265)  and  (not A236) );
 a14242a <=( (not A235)  and  a14241a );
 a14246a <=( A299  and  (not A298) );
 a14247a <=( (not A266)  and  a14246a );
 a14248a <=( a14247a  and  a14242a );
 a14251a <=( A166  and  A168 );
 a14255a <=( (not A233)  and  (not A201) );
 a14256a <=( (not A200)  and  a14255a );
 a14257a <=( a14256a  and  a14251a );
 a14261a <=( (not A268)  and  (not A266) );
 a14262a <=( (not A234)  and  a14261a );
 a14266a <=( A299  and  (not A298) );
 a14267a <=( (not A269)  and  a14266a );
 a14268a <=( a14267a  and  a14262a );
 a14271a <=( A166  and  A168 );
 a14275a <=( A232  and  (not A201) );
 a14276a <=( (not A200)  and  a14275a );
 a14277a <=( a14276a  and  a14271a );
 a14281a <=( A235  and  A234 );
 a14282a <=( (not A233)  and  a14281a );
 a14286a <=( (not A302)  and  (not A301) );
 a14287a <=( A298  and  a14286a );
 a14288a <=( a14287a  and  a14282a );
 a14291a <=( A166  and  A168 );
 a14295a <=( A232  and  (not A201) );
 a14296a <=( (not A200)  and  a14295a );
 a14297a <=( a14296a  and  a14291a );
 a14301a <=( A236  and  A234 );
 a14302a <=( (not A233)  and  a14301a );
 a14306a <=( (not A302)  and  (not A301) );
 a14307a <=( A298  and  a14306a );
 a14308a <=( a14307a  and  a14302a );
 a14311a <=( A166  and  A168 );
 a14315a <=( (not A232)  and  (not A201) );
 a14316a <=( (not A200)  and  a14315a );
 a14317a <=( a14316a  and  a14311a );
 a14321a <=( (not A268)  and  (not A266) );
 a14322a <=( (not A233)  and  a14321a );
 a14326a <=( A299  and  (not A298) );
 a14327a <=( (not A269)  and  a14326a );
 a14328a <=( a14327a  and  a14322a );
 a14331a <=( A166  and  A168 );
 a14335a <=( A232  and  (not A200) );
 a14336a <=( (not A199)  and  a14335a );
 a14337a <=( a14336a  and  a14331a );
 a14341a <=( (not A268)  and  A265 );
 a14342a <=( A233  and  a14341a );
 a14346a <=( A299  and  (not A298) );
 a14347a <=( (not A269)  and  a14346a );
 a14348a <=( a14347a  and  a14342a );
 a14351a <=( A166  and  A168 );
 a14355a <=( (not A233)  and  (not A200) );
 a14356a <=( (not A199)  and  a14355a );
 a14357a <=( a14356a  and  a14351a );
 a14361a <=( A265  and  (not A236) );
 a14362a <=( (not A235)  and  a14361a );
 a14366a <=( A299  and  (not A298) );
 a14367a <=( A266  and  a14366a );
 a14368a <=( a14367a  and  a14362a );
 a14371a <=( A166  and  A168 );
 a14375a <=( (not A233)  and  (not A200) );
 a14376a <=( (not A199)  and  a14375a );
 a14377a <=( a14376a  and  a14371a );
 a14381a <=( (not A266)  and  (not A236) );
 a14382a <=( (not A235)  and  a14381a );
 a14386a <=( A299  and  (not A298) );
 a14387a <=( (not A267)  and  a14386a );
 a14388a <=( a14387a  and  a14382a );
 a14391a <=( A166  and  A168 );
 a14395a <=( (not A233)  and  (not A200) );
 a14396a <=( (not A199)  and  a14395a );
 a14397a <=( a14396a  and  a14391a );
 a14401a <=( (not A265)  and  (not A236) );
 a14402a <=( (not A235)  and  a14401a );
 a14406a <=( A299  and  (not A298) );
 a14407a <=( (not A266)  and  a14406a );
 a14408a <=( a14407a  and  a14402a );
 a14411a <=( A166  and  A168 );
 a14415a <=( (not A233)  and  (not A200) );
 a14416a <=( (not A199)  and  a14415a );
 a14417a <=( a14416a  and  a14411a );
 a14421a <=( (not A268)  and  (not A266) );
 a14422a <=( (not A234)  and  a14421a );
 a14426a <=( A299  and  (not A298) );
 a14427a <=( (not A269)  and  a14426a );
 a14428a <=( a14427a  and  a14422a );
 a14431a <=( A166  and  A168 );
 a14435a <=( A232  and  (not A200) );
 a14436a <=( (not A199)  and  a14435a );
 a14437a <=( a14436a  and  a14431a );
 a14441a <=( A235  and  A234 );
 a14442a <=( (not A233)  and  a14441a );
 a14446a <=( (not A302)  and  (not A301) );
 a14447a <=( A298  and  a14446a );
 a14448a <=( a14447a  and  a14442a );
 a14451a <=( A166  and  A168 );
 a14455a <=( A232  and  (not A200) );
 a14456a <=( (not A199)  and  a14455a );
 a14457a <=( a14456a  and  a14451a );
 a14461a <=( A236  and  A234 );
 a14462a <=( (not A233)  and  a14461a );
 a14466a <=( (not A302)  and  (not A301) );
 a14467a <=( A298  and  a14466a );
 a14468a <=( a14467a  and  a14462a );
 a14471a <=( A166  and  A168 );
 a14475a <=( (not A232)  and  (not A200) );
 a14476a <=( (not A199)  and  a14475a );
 a14477a <=( a14476a  and  a14471a );
 a14481a <=( (not A268)  and  (not A266) );
 a14482a <=( (not A233)  and  a14481a );
 a14486a <=( A299  and  (not A298) );
 a14487a <=( (not A269)  and  a14486a );
 a14488a <=( a14487a  and  a14482a );
 a14491a <=( A167  and  A168 );
 a14495a <=( A232  and  A200 );
 a14496a <=( A199  and  a14495a );
 a14497a <=( a14496a  and  a14491a );
 a14501a <=( (not A268)  and  A265 );
 a14502a <=( A233  and  a14501a );
 a14506a <=( A299  and  (not A298) );
 a14507a <=( (not A269)  and  a14506a );
 a14508a <=( a14507a  and  a14502a );
 a14511a <=( A167  and  A168 );
 a14515a <=( (not A233)  and  A200 );
 a14516a <=( A199  and  a14515a );
 a14517a <=( a14516a  and  a14511a );
 a14521a <=( A265  and  (not A236) );
 a14522a <=( (not A235)  and  a14521a );
 a14526a <=( A299  and  (not A298) );
 a14527a <=( A266  and  a14526a );
 a14528a <=( a14527a  and  a14522a );
 a14531a <=( A167  and  A168 );
 a14535a <=( (not A233)  and  A200 );
 a14536a <=( A199  and  a14535a );
 a14537a <=( a14536a  and  a14531a );
 a14541a <=( (not A266)  and  (not A236) );
 a14542a <=( (not A235)  and  a14541a );
 a14546a <=( A299  and  (not A298) );
 a14547a <=( (not A267)  and  a14546a );
 a14548a <=( a14547a  and  a14542a );
 a14551a <=( A167  and  A168 );
 a14555a <=( (not A233)  and  A200 );
 a14556a <=( A199  and  a14555a );
 a14557a <=( a14556a  and  a14551a );
 a14561a <=( (not A265)  and  (not A236) );
 a14562a <=( (not A235)  and  a14561a );
 a14566a <=( A299  and  (not A298) );
 a14567a <=( (not A266)  and  a14566a );
 a14568a <=( a14567a  and  a14562a );
 a14571a <=( A167  and  A168 );
 a14575a <=( (not A233)  and  A200 );
 a14576a <=( A199  and  a14575a );
 a14577a <=( a14576a  and  a14571a );
 a14581a <=( (not A268)  and  (not A266) );
 a14582a <=( (not A234)  and  a14581a );
 a14586a <=( A299  and  (not A298) );
 a14587a <=( (not A269)  and  a14586a );
 a14588a <=( a14587a  and  a14582a );
 a14591a <=( A167  and  A168 );
 a14595a <=( A232  and  A200 );
 a14596a <=( A199  and  a14595a );
 a14597a <=( a14596a  and  a14591a );
 a14601a <=( A235  and  A234 );
 a14602a <=( (not A233)  and  a14601a );
 a14606a <=( (not A302)  and  (not A301) );
 a14607a <=( A298  and  a14606a );
 a14608a <=( a14607a  and  a14602a );
 a14611a <=( A167  and  A168 );
 a14615a <=( A232  and  A200 );
 a14616a <=( A199  and  a14615a );
 a14617a <=( a14616a  and  a14611a );
 a14621a <=( A236  and  A234 );
 a14622a <=( (not A233)  and  a14621a );
 a14626a <=( (not A302)  and  (not A301) );
 a14627a <=( A298  and  a14626a );
 a14628a <=( a14627a  and  a14622a );
 a14631a <=( A167  and  A168 );
 a14635a <=( (not A232)  and  A200 );
 a14636a <=( A199  and  a14635a );
 a14637a <=( a14636a  and  a14631a );
 a14641a <=( (not A268)  and  (not A266) );
 a14642a <=( (not A233)  and  a14641a );
 a14646a <=( A299  and  (not A298) );
 a14647a <=( (not A269)  and  a14646a );
 a14648a <=( a14647a  and  a14642a );
 a14651a <=( A167  and  A168 );
 a14655a <=( (not A203)  and  (not A202) );
 a14656a <=( (not A200)  and  a14655a );
 a14657a <=( a14656a  and  a14651a );
 a14661a <=( A265  and  A233 );
 a14662a <=( A232  and  a14661a );
 a14666a <=( A299  and  (not A298) );
 a14667a <=( (not A267)  and  a14666a );
 a14668a <=( a14667a  and  a14662a );
 a14671a <=( A167  and  A168 );
 a14675a <=( (not A203)  and  (not A202) );
 a14676a <=( (not A200)  and  a14675a );
 a14677a <=( a14676a  and  a14671a );
 a14681a <=( A265  and  A233 );
 a14682a <=( A232  and  a14681a );
 a14686a <=( A299  and  (not A298) );
 a14687a <=( A266  and  a14686a );
 a14688a <=( a14687a  and  a14682a );
 a14691a <=( A167  and  A168 );
 a14695a <=( (not A203)  and  (not A202) );
 a14696a <=( (not A200)  and  a14695a );
 a14697a <=( a14696a  and  a14691a );
 a14701a <=( (not A265)  and  A233 );
 a14702a <=( A232  and  a14701a );
 a14706a <=( A299  and  (not A298) );
 a14707a <=( (not A266)  and  a14706a );
 a14708a <=( a14707a  and  a14702a );
 a14711a <=( A167  and  A168 );
 a14715a <=( (not A203)  and  (not A202) );
 a14716a <=( (not A200)  and  a14715a );
 a14717a <=( a14716a  and  a14711a );
 a14721a <=( A265  and  A233 );
 a14722a <=( (not A232)  and  a14721a );
 a14726a <=( A268  and  A267 );
 a14727a <=( (not A266)  and  a14726a );
 a14728a <=( a14727a  and  a14722a );
 a14731a <=( A167  and  A168 );
 a14735a <=( (not A203)  and  (not A202) );
 a14736a <=( (not A200)  and  a14735a );
 a14737a <=( a14736a  and  a14731a );
 a14741a <=( A265  and  A233 );
 a14742a <=( (not A232)  and  a14741a );
 a14746a <=( A269  and  A267 );
 a14747a <=( (not A266)  and  a14746a );
 a14748a <=( a14747a  and  a14742a );
 a14751a <=( A167  and  A168 );
 a14755a <=( (not A203)  and  (not A202) );
 a14756a <=( (not A200)  and  a14755a );
 a14757a <=( a14756a  and  a14751a );
 a14761a <=( A265  and  (not A234) );
 a14762a <=( (not A233)  and  a14761a );
 a14766a <=( A299  and  (not A298) );
 a14767a <=( A266  and  a14766a );
 a14768a <=( a14767a  and  a14762a );
 a14771a <=( A167  and  A168 );
 a14775a <=( (not A203)  and  (not A202) );
 a14776a <=( (not A200)  and  a14775a );
 a14777a <=( a14776a  and  a14771a );
 a14781a <=( (not A266)  and  (not A234) );
 a14782a <=( (not A233)  and  a14781a );
 a14786a <=( A299  and  (not A298) );
 a14787a <=( (not A267)  and  a14786a );
 a14788a <=( a14787a  and  a14782a );
 a14791a <=( A167  and  A168 );
 a14795a <=( (not A203)  and  (not A202) );
 a14796a <=( (not A200)  and  a14795a );
 a14797a <=( a14796a  and  a14791a );
 a14801a <=( (not A265)  and  (not A234) );
 a14802a <=( (not A233)  and  a14801a );
 a14806a <=( A299  and  (not A298) );
 a14807a <=( (not A266)  and  a14806a );
 a14808a <=( a14807a  and  a14802a );
 a14811a <=( A167  and  A168 );
 a14815a <=( (not A203)  and  (not A202) );
 a14816a <=( (not A200)  and  a14815a );
 a14817a <=( a14816a  and  a14811a );
 a14821a <=( A234  and  (not A233) );
 a14822a <=( A232  and  a14821a );
 a14826a <=( (not A300)  and  A298 );
 a14827a <=( A235  and  a14826a );
 a14828a <=( a14827a  and  a14822a );
 a14831a <=( A167  and  A168 );
 a14835a <=( (not A203)  and  (not A202) );
 a14836a <=( (not A200)  and  a14835a );
 a14837a <=( a14836a  and  a14831a );
 a14841a <=( A234  and  (not A233) );
 a14842a <=( A232  and  a14841a );
 a14846a <=( A299  and  A298 );
 a14847a <=( A235  and  a14846a );
 a14848a <=( a14847a  and  a14842a );
 a14851a <=( A167  and  A168 );
 a14855a <=( (not A203)  and  (not A202) );
 a14856a <=( (not A200)  and  a14855a );
 a14857a <=( a14856a  and  a14851a );
 a14861a <=( A234  and  (not A233) );
 a14862a <=( A232  and  a14861a );
 a14866a <=( (not A299)  and  (not A298) );
 a14867a <=( A235  and  a14866a );
 a14868a <=( a14867a  and  a14862a );
 a14871a <=( A167  and  A168 );
 a14875a <=( (not A203)  and  (not A202) );
 a14876a <=( (not A200)  and  a14875a );
 a14877a <=( a14876a  and  a14871a );
 a14881a <=( A234  and  (not A233) );
 a14882a <=( A232  and  a14881a );
 a14886a <=( A266  and  (not A265) );
 a14887a <=( A235  and  a14886a );
 a14888a <=( a14887a  and  a14882a );
 a14891a <=( A167  and  A168 );
 a14895a <=( (not A203)  and  (not A202) );
 a14896a <=( (not A200)  and  a14895a );
 a14897a <=( a14896a  and  a14891a );
 a14901a <=( A234  and  (not A233) );
 a14902a <=( A232  and  a14901a );
 a14906a <=( (not A300)  and  A298 );
 a14907a <=( A236  and  a14906a );
 a14908a <=( a14907a  and  a14902a );
 a14911a <=( A167  and  A168 );
 a14915a <=( (not A203)  and  (not A202) );
 a14916a <=( (not A200)  and  a14915a );
 a14917a <=( a14916a  and  a14911a );
 a14921a <=( A234  and  (not A233) );
 a14922a <=( A232  and  a14921a );
 a14926a <=( A299  and  A298 );
 a14927a <=( A236  and  a14926a );
 a14928a <=( a14927a  and  a14922a );
 a14931a <=( A167  and  A168 );
 a14935a <=( (not A203)  and  (not A202) );
 a14936a <=( (not A200)  and  a14935a );
 a14937a <=( a14936a  and  a14931a );
 a14941a <=( A234  and  (not A233) );
 a14942a <=( A232  and  a14941a );
 a14946a <=( (not A299)  and  (not A298) );
 a14947a <=( A236  and  a14946a );
 a14948a <=( a14947a  and  a14942a );
 a14951a <=( A167  and  A168 );
 a14955a <=( (not A203)  and  (not A202) );
 a14956a <=( (not A200)  and  a14955a );
 a14957a <=( a14956a  and  a14951a );
 a14961a <=( A234  and  (not A233) );
 a14962a <=( A232  and  a14961a );
 a14966a <=( A266  and  (not A265) );
 a14967a <=( A236  and  a14966a );
 a14968a <=( a14967a  and  a14962a );
 a14971a <=( A167  and  A168 );
 a14975a <=( (not A203)  and  (not A202) );
 a14976a <=( (not A200)  and  a14975a );
 a14977a <=( a14976a  and  a14971a );
 a14981a <=( A265  and  (not A233) );
 a14982a <=( (not A232)  and  a14981a );
 a14986a <=( A299  and  (not A298) );
 a14987a <=( A266  and  a14986a );
 a14988a <=( a14987a  and  a14982a );
 a14991a <=( A167  and  A168 );
 a14995a <=( (not A203)  and  (not A202) );
 a14996a <=( (not A200)  and  a14995a );
 a14997a <=( a14996a  and  a14991a );
 a15001a <=( (not A266)  and  (not A233) );
 a15002a <=( (not A232)  and  a15001a );
 a15006a <=( A299  and  (not A298) );
 a15007a <=( (not A267)  and  a15006a );
 a15008a <=( a15007a  and  a15002a );
 a15011a <=( A167  and  A168 );
 a15015a <=( (not A203)  and  (not A202) );
 a15016a <=( (not A200)  and  a15015a );
 a15017a <=( a15016a  and  a15011a );
 a15021a <=( (not A265)  and  (not A233) );
 a15022a <=( (not A232)  and  a15021a );
 a15026a <=( A299  and  (not A298) );
 a15027a <=( (not A266)  and  a15026a );
 a15028a <=( a15027a  and  a15022a );
 a15031a <=( A167  and  A168 );
 a15035a <=( A232  and  (not A201) );
 a15036a <=( (not A200)  and  a15035a );
 a15037a <=( a15036a  and  a15031a );
 a15041a <=( (not A268)  and  A265 );
 a15042a <=( A233  and  a15041a );
 a15046a <=( A299  and  (not A298) );
 a15047a <=( (not A269)  and  a15046a );
 a15048a <=( a15047a  and  a15042a );
 a15051a <=( A167  and  A168 );
 a15055a <=( (not A233)  and  (not A201) );
 a15056a <=( (not A200)  and  a15055a );
 a15057a <=( a15056a  and  a15051a );
 a15061a <=( A265  and  (not A236) );
 a15062a <=( (not A235)  and  a15061a );
 a15066a <=( A299  and  (not A298) );
 a15067a <=( A266  and  a15066a );
 a15068a <=( a15067a  and  a15062a );
 a15071a <=( A167  and  A168 );
 a15075a <=( (not A233)  and  (not A201) );
 a15076a <=( (not A200)  and  a15075a );
 a15077a <=( a15076a  and  a15071a );
 a15081a <=( (not A266)  and  (not A236) );
 a15082a <=( (not A235)  and  a15081a );
 a15086a <=( A299  and  (not A298) );
 a15087a <=( (not A267)  and  a15086a );
 a15088a <=( a15087a  and  a15082a );
 a15091a <=( A167  and  A168 );
 a15095a <=( (not A233)  and  (not A201) );
 a15096a <=( (not A200)  and  a15095a );
 a15097a <=( a15096a  and  a15091a );
 a15101a <=( (not A265)  and  (not A236) );
 a15102a <=( (not A235)  and  a15101a );
 a15106a <=( A299  and  (not A298) );
 a15107a <=( (not A266)  and  a15106a );
 a15108a <=( a15107a  and  a15102a );
 a15111a <=( A167  and  A168 );
 a15115a <=( (not A233)  and  (not A201) );
 a15116a <=( (not A200)  and  a15115a );
 a15117a <=( a15116a  and  a15111a );
 a15121a <=( (not A268)  and  (not A266) );
 a15122a <=( (not A234)  and  a15121a );
 a15126a <=( A299  and  (not A298) );
 a15127a <=( (not A269)  and  a15126a );
 a15128a <=( a15127a  and  a15122a );
 a15131a <=( A167  and  A168 );
 a15135a <=( A232  and  (not A201) );
 a15136a <=( (not A200)  and  a15135a );
 a15137a <=( a15136a  and  a15131a );
 a15141a <=( A235  and  A234 );
 a15142a <=( (not A233)  and  a15141a );
 a15146a <=( (not A302)  and  (not A301) );
 a15147a <=( A298  and  a15146a );
 a15148a <=( a15147a  and  a15142a );
 a15151a <=( A167  and  A168 );
 a15155a <=( A232  and  (not A201) );
 a15156a <=( (not A200)  and  a15155a );
 a15157a <=( a15156a  and  a15151a );
 a15161a <=( A236  and  A234 );
 a15162a <=( (not A233)  and  a15161a );
 a15166a <=( (not A302)  and  (not A301) );
 a15167a <=( A298  and  a15166a );
 a15168a <=( a15167a  and  a15162a );
 a15171a <=( A167  and  A168 );
 a15175a <=( (not A232)  and  (not A201) );
 a15176a <=( (not A200)  and  a15175a );
 a15177a <=( a15176a  and  a15171a );
 a15181a <=( (not A268)  and  (not A266) );
 a15182a <=( (not A233)  and  a15181a );
 a15186a <=( A299  and  (not A298) );
 a15187a <=( (not A269)  and  a15186a );
 a15188a <=( a15187a  and  a15182a );
 a15191a <=( A167  and  A168 );
 a15195a <=( A232  and  (not A200) );
 a15196a <=( (not A199)  and  a15195a );
 a15197a <=( a15196a  and  a15191a );
 a15201a <=( (not A268)  and  A265 );
 a15202a <=( A233  and  a15201a );
 a15206a <=( A299  and  (not A298) );
 a15207a <=( (not A269)  and  a15206a );
 a15208a <=( a15207a  and  a15202a );
 a15211a <=( A167  and  A168 );
 a15215a <=( (not A233)  and  (not A200) );
 a15216a <=( (not A199)  and  a15215a );
 a15217a <=( a15216a  and  a15211a );
 a15221a <=( A265  and  (not A236) );
 a15222a <=( (not A235)  and  a15221a );
 a15226a <=( A299  and  (not A298) );
 a15227a <=( A266  and  a15226a );
 a15228a <=( a15227a  and  a15222a );
 a15231a <=( A167  and  A168 );
 a15235a <=( (not A233)  and  (not A200) );
 a15236a <=( (not A199)  and  a15235a );
 a15237a <=( a15236a  and  a15231a );
 a15241a <=( (not A266)  and  (not A236) );
 a15242a <=( (not A235)  and  a15241a );
 a15246a <=( A299  and  (not A298) );
 a15247a <=( (not A267)  and  a15246a );
 a15248a <=( a15247a  and  a15242a );
 a15251a <=( A167  and  A168 );
 a15255a <=( (not A233)  and  (not A200) );
 a15256a <=( (not A199)  and  a15255a );
 a15257a <=( a15256a  and  a15251a );
 a15261a <=( (not A265)  and  (not A236) );
 a15262a <=( (not A235)  and  a15261a );
 a15266a <=( A299  and  (not A298) );
 a15267a <=( (not A266)  and  a15266a );
 a15268a <=( a15267a  and  a15262a );
 a15271a <=( A167  and  A168 );
 a15275a <=( (not A233)  and  (not A200) );
 a15276a <=( (not A199)  and  a15275a );
 a15277a <=( a15276a  and  a15271a );
 a15281a <=( (not A268)  and  (not A266) );
 a15282a <=( (not A234)  and  a15281a );
 a15286a <=( A299  and  (not A298) );
 a15287a <=( (not A269)  and  a15286a );
 a15288a <=( a15287a  and  a15282a );
 a15291a <=( A167  and  A168 );
 a15295a <=( A232  and  (not A200) );
 a15296a <=( (not A199)  and  a15295a );
 a15297a <=( a15296a  and  a15291a );
 a15301a <=( A235  and  A234 );
 a15302a <=( (not A233)  and  a15301a );
 a15306a <=( (not A302)  and  (not A301) );
 a15307a <=( A298  and  a15306a );
 a15308a <=( a15307a  and  a15302a );
 a15311a <=( A167  and  A168 );
 a15315a <=( A232  and  (not A200) );
 a15316a <=( (not A199)  and  a15315a );
 a15317a <=( a15316a  and  a15311a );
 a15321a <=( A236  and  A234 );
 a15322a <=( (not A233)  and  a15321a );
 a15326a <=( (not A302)  and  (not A301) );
 a15327a <=( A298  and  a15326a );
 a15328a <=( a15327a  and  a15322a );
 a15331a <=( A167  and  A168 );
 a15335a <=( (not A232)  and  (not A200) );
 a15336a <=( (not A199)  and  a15335a );
 a15337a <=( a15336a  and  a15331a );
 a15341a <=( (not A268)  and  (not A266) );
 a15342a <=( (not A233)  and  a15341a );
 a15346a <=( A299  and  (not A298) );
 a15347a <=( (not A269)  and  a15346a );
 a15348a <=( a15347a  and  a15342a );
 a15351a <=( (not A167)  and  A170 );
 a15355a <=( A200  and  (not A199) );
 a15356a <=( (not A166)  and  a15355a );
 a15357a <=( a15356a  and  a15351a );
 a15361a <=( A265  and  A233 );
 a15362a <=( A232  and  a15361a );
 a15366a <=( A299  and  (not A298) );
 a15367a <=( (not A267)  and  a15366a );
 a15368a <=( a15367a  and  a15362a );
 a15371a <=( (not A167)  and  A170 );
 a15375a <=( A200  and  (not A199) );
 a15376a <=( (not A166)  and  a15375a );
 a15377a <=( a15376a  and  a15371a );
 a15381a <=( A265  and  A233 );
 a15382a <=( A232  and  a15381a );
 a15386a <=( A299  and  (not A298) );
 a15387a <=( A266  and  a15386a );
 a15388a <=( a15387a  and  a15382a );
 a15391a <=( (not A167)  and  A170 );
 a15395a <=( A200  and  (not A199) );
 a15396a <=( (not A166)  and  a15395a );
 a15397a <=( a15396a  and  a15391a );
 a15401a <=( (not A265)  and  A233 );
 a15402a <=( A232  and  a15401a );
 a15406a <=( A299  and  (not A298) );
 a15407a <=( (not A266)  and  a15406a );
 a15408a <=( a15407a  and  a15402a );
 a15411a <=( (not A167)  and  A170 );
 a15415a <=( A200  and  (not A199) );
 a15416a <=( (not A166)  and  a15415a );
 a15417a <=( a15416a  and  a15411a );
 a15421a <=( A265  and  A233 );
 a15422a <=( (not A232)  and  a15421a );
 a15426a <=( A268  and  A267 );
 a15427a <=( (not A266)  and  a15426a );
 a15428a <=( a15427a  and  a15422a );
 a15431a <=( (not A167)  and  A170 );
 a15435a <=( A200  and  (not A199) );
 a15436a <=( (not A166)  and  a15435a );
 a15437a <=( a15436a  and  a15431a );
 a15441a <=( A265  and  A233 );
 a15442a <=( (not A232)  and  a15441a );
 a15446a <=( A269  and  A267 );
 a15447a <=( (not A266)  and  a15446a );
 a15448a <=( a15447a  and  a15442a );
 a15451a <=( (not A167)  and  A170 );
 a15455a <=( A200  and  (not A199) );
 a15456a <=( (not A166)  and  a15455a );
 a15457a <=( a15456a  and  a15451a );
 a15461a <=( A265  and  (not A234) );
 a15462a <=( (not A233)  and  a15461a );
 a15466a <=( A299  and  (not A298) );
 a15467a <=( A266  and  a15466a );
 a15468a <=( a15467a  and  a15462a );
 a15471a <=( (not A167)  and  A170 );
 a15475a <=( A200  and  (not A199) );
 a15476a <=( (not A166)  and  a15475a );
 a15477a <=( a15476a  and  a15471a );
 a15481a <=( (not A266)  and  (not A234) );
 a15482a <=( (not A233)  and  a15481a );
 a15486a <=( A299  and  (not A298) );
 a15487a <=( (not A267)  and  a15486a );
 a15488a <=( a15487a  and  a15482a );
 a15491a <=( (not A167)  and  A170 );
 a15495a <=( A200  and  (not A199) );
 a15496a <=( (not A166)  and  a15495a );
 a15497a <=( a15496a  and  a15491a );
 a15501a <=( (not A265)  and  (not A234) );
 a15502a <=( (not A233)  and  a15501a );
 a15506a <=( A299  and  (not A298) );
 a15507a <=( (not A266)  and  a15506a );
 a15508a <=( a15507a  and  a15502a );
 a15511a <=( (not A167)  and  A170 );
 a15515a <=( A200  and  (not A199) );
 a15516a <=( (not A166)  and  a15515a );
 a15517a <=( a15516a  and  a15511a );
 a15521a <=( A234  and  (not A233) );
 a15522a <=( A232  and  a15521a );
 a15526a <=( (not A300)  and  A298 );
 a15527a <=( A235  and  a15526a );
 a15528a <=( a15527a  and  a15522a );
 a15531a <=( (not A167)  and  A170 );
 a15535a <=( A200  and  (not A199) );
 a15536a <=( (not A166)  and  a15535a );
 a15537a <=( a15536a  and  a15531a );
 a15541a <=( A234  and  (not A233) );
 a15542a <=( A232  and  a15541a );
 a15546a <=( A299  and  A298 );
 a15547a <=( A235  and  a15546a );
 a15548a <=( a15547a  and  a15542a );
 a15551a <=( (not A167)  and  A170 );
 a15555a <=( A200  and  (not A199) );
 a15556a <=( (not A166)  and  a15555a );
 a15557a <=( a15556a  and  a15551a );
 a15561a <=( A234  and  (not A233) );
 a15562a <=( A232  and  a15561a );
 a15566a <=( (not A299)  and  (not A298) );
 a15567a <=( A235  and  a15566a );
 a15568a <=( a15567a  and  a15562a );
 a15571a <=( (not A167)  and  A170 );
 a15575a <=( A200  and  (not A199) );
 a15576a <=( (not A166)  and  a15575a );
 a15577a <=( a15576a  and  a15571a );
 a15581a <=( A234  and  (not A233) );
 a15582a <=( A232  and  a15581a );
 a15586a <=( A266  and  (not A265) );
 a15587a <=( A235  and  a15586a );
 a15588a <=( a15587a  and  a15582a );
 a15591a <=( (not A167)  and  A170 );
 a15595a <=( A200  and  (not A199) );
 a15596a <=( (not A166)  and  a15595a );
 a15597a <=( a15596a  and  a15591a );
 a15601a <=( A234  and  (not A233) );
 a15602a <=( A232  and  a15601a );
 a15606a <=( (not A300)  and  A298 );
 a15607a <=( A236  and  a15606a );
 a15608a <=( a15607a  and  a15602a );
 a15611a <=( (not A167)  and  A170 );
 a15615a <=( A200  and  (not A199) );
 a15616a <=( (not A166)  and  a15615a );
 a15617a <=( a15616a  and  a15611a );
 a15621a <=( A234  and  (not A233) );
 a15622a <=( A232  and  a15621a );
 a15626a <=( A299  and  A298 );
 a15627a <=( A236  and  a15626a );
 a15628a <=( a15627a  and  a15622a );
 a15631a <=( (not A167)  and  A170 );
 a15635a <=( A200  and  (not A199) );
 a15636a <=( (not A166)  and  a15635a );
 a15637a <=( a15636a  and  a15631a );
 a15641a <=( A234  and  (not A233) );
 a15642a <=( A232  and  a15641a );
 a15646a <=( (not A299)  and  (not A298) );
 a15647a <=( A236  and  a15646a );
 a15648a <=( a15647a  and  a15642a );
 a15651a <=( (not A167)  and  A170 );
 a15655a <=( A200  and  (not A199) );
 a15656a <=( (not A166)  and  a15655a );
 a15657a <=( a15656a  and  a15651a );
 a15661a <=( A234  and  (not A233) );
 a15662a <=( A232  and  a15661a );
 a15666a <=( A266  and  (not A265) );
 a15667a <=( A236  and  a15666a );
 a15668a <=( a15667a  and  a15662a );
 a15671a <=( (not A167)  and  A170 );
 a15675a <=( A200  and  (not A199) );
 a15676a <=( (not A166)  and  a15675a );
 a15677a <=( a15676a  and  a15671a );
 a15681a <=( A265  and  (not A233) );
 a15682a <=( (not A232)  and  a15681a );
 a15686a <=( A299  and  (not A298) );
 a15687a <=( A266  and  a15686a );
 a15688a <=( a15687a  and  a15682a );
 a15691a <=( (not A167)  and  A170 );
 a15695a <=( A200  and  (not A199) );
 a15696a <=( (not A166)  and  a15695a );
 a15697a <=( a15696a  and  a15691a );
 a15701a <=( (not A266)  and  (not A233) );
 a15702a <=( (not A232)  and  a15701a );
 a15706a <=( A299  and  (not A298) );
 a15707a <=( (not A267)  and  a15706a );
 a15708a <=( a15707a  and  a15702a );
 a15711a <=( (not A167)  and  A170 );
 a15715a <=( A200  and  (not A199) );
 a15716a <=( (not A166)  and  a15715a );
 a15717a <=( a15716a  and  a15711a );
 a15721a <=( (not A265)  and  (not A233) );
 a15722a <=( (not A232)  and  a15721a );
 a15726a <=( A299  and  (not A298) );
 a15727a <=( (not A266)  and  a15726a );
 a15728a <=( a15727a  and  a15722a );
 a15731a <=( (not A167)  and  A170 );
 a15735a <=( (not A200)  and  A199 );
 a15736a <=( (not A166)  and  a15735a );
 a15737a <=( a15736a  and  a15731a );
 a15741a <=( (not A232)  and  A202 );
 a15742a <=( A201  and  a15741a );
 a15746a <=( (not A300)  and  (not A299) );
 a15747a <=( A233  and  a15746a );
 a15748a <=( a15747a  and  a15742a );
 a15751a <=( (not A167)  and  A170 );
 a15755a <=( (not A200)  and  A199 );
 a15756a <=( (not A166)  and  a15755a );
 a15757a <=( a15756a  and  a15751a );
 a15761a <=( (not A232)  and  A202 );
 a15762a <=( A201  and  a15761a );
 a15766a <=( A299  and  A298 );
 a15767a <=( A233  and  a15766a );
 a15768a <=( a15767a  and  a15762a );
 a15771a <=( (not A167)  and  A170 );
 a15775a <=( (not A200)  and  A199 );
 a15776a <=( (not A166)  and  a15775a );
 a15777a <=( a15776a  and  a15771a );
 a15781a <=( (not A232)  and  A202 );
 a15782a <=( A201  and  a15781a );
 a15786a <=( (not A299)  and  (not A298) );
 a15787a <=( A233  and  a15786a );
 a15788a <=( a15787a  and  a15782a );
 a15791a <=( (not A167)  and  A170 );
 a15795a <=( (not A200)  and  A199 );
 a15796a <=( (not A166)  and  a15795a );
 a15797a <=( a15796a  and  a15791a );
 a15801a <=( (not A232)  and  A202 );
 a15802a <=( A201  and  a15801a );
 a15806a <=( A266  and  (not A265) );
 a15807a <=( A233  and  a15806a );
 a15808a <=( a15807a  and  a15802a );
 a15811a <=( (not A167)  and  A170 );
 a15815a <=( (not A200)  and  A199 );
 a15816a <=( (not A166)  and  a15815a );
 a15817a <=( a15816a  and  a15811a );
 a15821a <=( (not A232)  and  A203 );
 a15822a <=( A201  and  a15821a );
 a15826a <=( (not A300)  and  (not A299) );
 a15827a <=( A233  and  a15826a );
 a15828a <=( a15827a  and  a15822a );
 a15831a <=( (not A167)  and  A170 );
 a15835a <=( (not A200)  and  A199 );
 a15836a <=( (not A166)  and  a15835a );
 a15837a <=( a15836a  and  a15831a );
 a15841a <=( (not A232)  and  A203 );
 a15842a <=( A201  and  a15841a );
 a15846a <=( A299  and  A298 );
 a15847a <=( A233  and  a15846a );
 a15848a <=( a15847a  and  a15842a );
 a15851a <=( (not A167)  and  A170 );
 a15855a <=( (not A200)  and  A199 );
 a15856a <=( (not A166)  and  a15855a );
 a15857a <=( a15856a  and  a15851a );
 a15861a <=( (not A232)  and  A203 );
 a15862a <=( A201  and  a15861a );
 a15866a <=( (not A299)  and  (not A298) );
 a15867a <=( A233  and  a15866a );
 a15868a <=( a15867a  and  a15862a );
 a15871a <=( (not A167)  and  A170 );
 a15875a <=( (not A200)  and  A199 );
 a15876a <=( (not A166)  and  a15875a );
 a15877a <=( a15876a  and  a15871a );
 a15881a <=( (not A232)  and  A203 );
 a15882a <=( A201  and  a15881a );
 a15886a <=( A266  and  (not A265) );
 a15887a <=( A233  and  a15886a );
 a15888a <=( a15887a  and  a15882a );
 a15891a <=( (not A168)  and  A170 );
 a15895a <=( (not A199)  and  A166 );
 a15896a <=( A167  and  a15895a );
 a15897a <=( a15896a  and  a15891a );
 a15901a <=( A233  and  (not A232) );
 a15902a <=( A200  and  a15901a );
 a15906a <=( (not A302)  and  (not A301) );
 a15907a <=( (not A299)  and  a15906a );
 a15908a <=( a15907a  and  a15902a );
 a15911a <=( (not A168)  and  (not A170) );
 a15915a <=( (not A199)  and  (not A166) );
 a15916a <=( A167  and  a15915a );
 a15917a <=( a15916a  and  a15911a );
 a15921a <=( A233  and  (not A232) );
 a15922a <=( A200  and  a15921a );
 a15926a <=( (not A302)  and  (not A301) );
 a15927a <=( (not A299)  and  a15926a );
 a15928a <=( a15927a  and  a15922a );
 a15931a <=( (not A168)  and  (not A170) );
 a15935a <=( (not A199)  and  A166 );
 a15936a <=( (not A167)  and  a15935a );
 a15937a <=( a15936a  and  a15931a );
 a15941a <=( A233  and  (not A232) );
 a15942a <=( A200  and  a15941a );
 a15946a <=( (not A302)  and  (not A301) );
 a15947a <=( (not A299)  and  a15946a );
 a15948a <=( a15947a  and  a15942a );
 a15951a <=( (not A168)  and  A169 );
 a15955a <=( (not A199)  and  (not A166) );
 a15956a <=( A167  and  a15955a );
 a15957a <=( a15956a  and  a15951a );
 a15961a <=( A233  and  (not A232) );
 a15962a <=( A200  and  a15961a );
 a15966a <=( (not A302)  and  (not A301) );
 a15967a <=( (not A299)  and  a15966a );
 a15968a <=( a15967a  and  a15962a );
 a15971a <=( (not A168)  and  A169 );
 a15975a <=( (not A199)  and  A166 );
 a15976a <=( (not A167)  and  a15975a );
 a15977a <=( a15976a  and  a15971a );
 a15981a <=( A233  and  (not A232) );
 a15982a <=( A200  and  a15981a );
 a15986a <=( (not A302)  and  (not A301) );
 a15987a <=( (not A299)  and  a15986a );
 a15988a <=( a15987a  and  a15982a );
 a15991a <=( A169  and  A170 );
 a15995a <=( (not A200)  and  A199 );
 a15996a <=( (not A168)  and  a15995a );
 a15997a <=( a15996a  and  a15991a );
 a16001a <=( (not A232)  and  A202 );
 a16002a <=( A201  and  a16001a );
 a16006a <=( (not A300)  and  (not A299) );
 a16007a <=( A233  and  a16006a );
 a16008a <=( a16007a  and  a16002a );
 a16011a <=( A169  and  A170 );
 a16015a <=( (not A200)  and  A199 );
 a16016a <=( (not A168)  and  a16015a );
 a16017a <=( a16016a  and  a16011a );
 a16021a <=( (not A232)  and  A202 );
 a16022a <=( A201  and  a16021a );
 a16026a <=( A299  and  A298 );
 a16027a <=( A233  and  a16026a );
 a16028a <=( a16027a  and  a16022a );
 a16031a <=( A169  and  A170 );
 a16035a <=( (not A200)  and  A199 );
 a16036a <=( (not A168)  and  a16035a );
 a16037a <=( a16036a  and  a16031a );
 a16041a <=( (not A232)  and  A202 );
 a16042a <=( A201  and  a16041a );
 a16046a <=( (not A299)  and  (not A298) );
 a16047a <=( A233  and  a16046a );
 a16048a <=( a16047a  and  a16042a );
 a16051a <=( A169  and  A170 );
 a16055a <=( (not A200)  and  A199 );
 a16056a <=( (not A168)  and  a16055a );
 a16057a <=( a16056a  and  a16051a );
 a16061a <=( (not A232)  and  A202 );
 a16062a <=( A201  and  a16061a );
 a16066a <=( A266  and  (not A265) );
 a16067a <=( A233  and  a16066a );
 a16068a <=( a16067a  and  a16062a );
 a16071a <=( A169  and  A170 );
 a16075a <=( (not A200)  and  A199 );
 a16076a <=( (not A168)  and  a16075a );
 a16077a <=( a16076a  and  a16071a );
 a16081a <=( (not A232)  and  A203 );
 a16082a <=( A201  and  a16081a );
 a16086a <=( (not A300)  and  (not A299) );
 a16087a <=( A233  and  a16086a );
 a16088a <=( a16087a  and  a16082a );
 a16091a <=( A169  and  A170 );
 a16095a <=( (not A200)  and  A199 );
 a16096a <=( (not A168)  and  a16095a );
 a16097a <=( a16096a  and  a16091a );
 a16101a <=( (not A232)  and  A203 );
 a16102a <=( A201  and  a16101a );
 a16106a <=( A299  and  A298 );
 a16107a <=( A233  and  a16106a );
 a16108a <=( a16107a  and  a16102a );
 a16111a <=( A169  and  A170 );
 a16115a <=( (not A200)  and  A199 );
 a16116a <=( (not A168)  and  a16115a );
 a16117a <=( a16116a  and  a16111a );
 a16121a <=( (not A232)  and  A203 );
 a16122a <=( A201  and  a16121a );
 a16126a <=( (not A299)  and  (not A298) );
 a16127a <=( A233  and  a16126a );
 a16128a <=( a16127a  and  a16122a );
 a16131a <=( A169  and  A170 );
 a16135a <=( (not A200)  and  A199 );
 a16136a <=( (not A168)  and  a16135a );
 a16137a <=( a16136a  and  a16131a );
 a16141a <=( (not A232)  and  A203 );
 a16142a <=( A201  and  a16141a );
 a16146a <=( A266  and  (not A265) );
 a16147a <=( A233  and  a16146a );
 a16148a <=( a16147a  and  a16142a );
 a16151a <=( A169  and  (not A170) );
 a16155a <=( A199  and  A166 );
 a16156a <=( A167  and  a16155a );
 a16157a <=( a16156a  and  a16151a );
 a16161a <=( A233  and  (not A232) );
 a16162a <=( A200  and  a16161a );
 a16166a <=( (not A302)  and  (not A301) );
 a16167a <=( (not A299)  and  a16166a );
 a16168a <=( a16167a  and  a16162a );
 a16171a <=( A169  and  (not A170) );
 a16175a <=( (not A200)  and  A166 );
 a16176a <=( A167  and  a16175a );
 a16177a <=( a16176a  and  a16171a );
 a16181a <=( (not A232)  and  (not A203) );
 a16182a <=( (not A202)  and  a16181a );
 a16186a <=( (not A300)  and  (not A299) );
 a16187a <=( A233  and  a16186a );
 a16188a <=( a16187a  and  a16182a );
 a16191a <=( A169  and  (not A170) );
 a16195a <=( (not A200)  and  A166 );
 a16196a <=( A167  and  a16195a );
 a16197a <=( a16196a  and  a16191a );
 a16201a <=( (not A232)  and  (not A203) );
 a16202a <=( (not A202)  and  a16201a );
 a16206a <=( A299  and  A298 );
 a16207a <=( A233  and  a16206a );
 a16208a <=( a16207a  and  a16202a );
 a16211a <=( A169  and  (not A170) );
 a16215a <=( (not A200)  and  A166 );
 a16216a <=( A167  and  a16215a );
 a16217a <=( a16216a  and  a16211a );
 a16221a <=( (not A232)  and  (not A203) );
 a16222a <=( (not A202)  and  a16221a );
 a16226a <=( (not A299)  and  (not A298) );
 a16227a <=( A233  and  a16226a );
 a16228a <=( a16227a  and  a16222a );
 a16231a <=( A169  and  (not A170) );
 a16235a <=( (not A200)  and  A166 );
 a16236a <=( A167  and  a16235a );
 a16237a <=( a16236a  and  a16231a );
 a16241a <=( (not A232)  and  (not A203) );
 a16242a <=( (not A202)  and  a16241a );
 a16246a <=( A266  and  (not A265) );
 a16247a <=( A233  and  a16246a );
 a16248a <=( a16247a  and  a16242a );
 a16251a <=( A169  and  (not A170) );
 a16255a <=( (not A200)  and  A166 );
 a16256a <=( A167  and  a16255a );
 a16257a <=( a16256a  and  a16251a );
 a16261a <=( A233  and  (not A232) );
 a16262a <=( (not A201)  and  a16261a );
 a16266a <=( (not A302)  and  (not A301) );
 a16267a <=( (not A299)  and  a16266a );
 a16268a <=( a16267a  and  a16262a );
 a16271a <=( A169  and  (not A170) );
 a16275a <=( (not A199)  and  A166 );
 a16276a <=( A167  and  a16275a );
 a16277a <=( a16276a  and  a16271a );
 a16281a <=( A233  and  (not A232) );
 a16282a <=( (not A200)  and  a16281a );
 a16286a <=( (not A302)  and  (not A301) );
 a16287a <=( (not A299)  and  a16286a );
 a16288a <=( a16287a  and  a16282a );
 a16291a <=( A169  and  (not A170) );
 a16295a <=( A199  and  (not A166) );
 a16296a <=( (not A167)  and  a16295a );
 a16297a <=( a16296a  and  a16291a );
 a16301a <=( A233  and  (not A232) );
 a16302a <=( A200  and  a16301a );
 a16306a <=( (not A302)  and  (not A301) );
 a16307a <=( (not A299)  and  a16306a );
 a16308a <=( a16307a  and  a16302a );
 a16311a <=( A169  and  (not A170) );
 a16315a <=( (not A200)  and  (not A166) );
 a16316a <=( (not A167)  and  a16315a );
 a16317a <=( a16316a  and  a16311a );
 a16321a <=( (not A232)  and  (not A203) );
 a16322a <=( (not A202)  and  a16321a );
 a16326a <=( (not A300)  and  (not A299) );
 a16327a <=( A233  and  a16326a );
 a16328a <=( a16327a  and  a16322a );
 a16331a <=( A169  and  (not A170) );
 a16335a <=( (not A200)  and  (not A166) );
 a16336a <=( (not A167)  and  a16335a );
 a16337a <=( a16336a  and  a16331a );
 a16341a <=( (not A232)  and  (not A203) );
 a16342a <=( (not A202)  and  a16341a );
 a16346a <=( A299  and  A298 );
 a16347a <=( A233  and  a16346a );
 a16348a <=( a16347a  and  a16342a );
 a16351a <=( A169  and  (not A170) );
 a16355a <=( (not A200)  and  (not A166) );
 a16356a <=( (not A167)  and  a16355a );
 a16357a <=( a16356a  and  a16351a );
 a16361a <=( (not A232)  and  (not A203) );
 a16362a <=( (not A202)  and  a16361a );
 a16366a <=( (not A299)  and  (not A298) );
 a16367a <=( A233  and  a16366a );
 a16368a <=( a16367a  and  a16362a );
 a16371a <=( A169  and  (not A170) );
 a16375a <=( (not A200)  and  (not A166) );
 a16376a <=( (not A167)  and  a16375a );
 a16377a <=( a16376a  and  a16371a );
 a16381a <=( (not A232)  and  (not A203) );
 a16382a <=( (not A202)  and  a16381a );
 a16386a <=( A266  and  (not A265) );
 a16387a <=( A233  and  a16386a );
 a16388a <=( a16387a  and  a16382a );
 a16391a <=( A169  and  (not A170) );
 a16395a <=( (not A200)  and  (not A166) );
 a16396a <=( (not A167)  and  a16395a );
 a16397a <=( a16396a  and  a16391a );
 a16401a <=( A233  and  (not A232) );
 a16402a <=( (not A201)  and  a16401a );
 a16406a <=( (not A302)  and  (not A301) );
 a16407a <=( (not A299)  and  a16406a );
 a16408a <=( a16407a  and  a16402a );
 a16411a <=( A169  and  (not A170) );
 a16415a <=( (not A199)  and  (not A166) );
 a16416a <=( (not A167)  and  a16415a );
 a16417a <=( a16416a  and  a16411a );
 a16421a <=( A233  and  (not A232) );
 a16422a <=( (not A200)  and  a16421a );
 a16426a <=( (not A302)  and  (not A301) );
 a16427a <=( (not A299)  and  a16426a );
 a16428a <=( a16427a  and  a16422a );
 a16431a <=( (not A167)  and  (not A169) );
 a16435a <=( A200  and  (not A199) );
 a16436a <=( (not A166)  and  a16435a );
 a16437a <=( a16436a  and  a16431a );
 a16441a <=( A265  and  A233 );
 a16442a <=( A232  and  a16441a );
 a16446a <=( A299  and  (not A298) );
 a16447a <=( (not A267)  and  a16446a );
 a16448a <=( a16447a  and  a16442a );
 a16451a <=( (not A167)  and  (not A169) );
 a16455a <=( A200  and  (not A199) );
 a16456a <=( (not A166)  and  a16455a );
 a16457a <=( a16456a  and  a16451a );
 a16461a <=( A265  and  A233 );
 a16462a <=( A232  and  a16461a );
 a16466a <=( A299  and  (not A298) );
 a16467a <=( A266  and  a16466a );
 a16468a <=( a16467a  and  a16462a );
 a16471a <=( (not A167)  and  (not A169) );
 a16475a <=( A200  and  (not A199) );
 a16476a <=( (not A166)  and  a16475a );
 a16477a <=( a16476a  and  a16471a );
 a16481a <=( (not A265)  and  A233 );
 a16482a <=( A232  and  a16481a );
 a16486a <=( A299  and  (not A298) );
 a16487a <=( (not A266)  and  a16486a );
 a16488a <=( a16487a  and  a16482a );
 a16491a <=( (not A167)  and  (not A169) );
 a16495a <=( A200  and  (not A199) );
 a16496a <=( (not A166)  and  a16495a );
 a16497a <=( a16496a  and  a16491a );
 a16501a <=( A265  and  A233 );
 a16502a <=( (not A232)  and  a16501a );
 a16506a <=( A268  and  A267 );
 a16507a <=( (not A266)  and  a16506a );
 a16508a <=( a16507a  and  a16502a );
 a16511a <=( (not A167)  and  (not A169) );
 a16515a <=( A200  and  (not A199) );
 a16516a <=( (not A166)  and  a16515a );
 a16517a <=( a16516a  and  a16511a );
 a16521a <=( A265  and  A233 );
 a16522a <=( (not A232)  and  a16521a );
 a16526a <=( A269  and  A267 );
 a16527a <=( (not A266)  and  a16526a );
 a16528a <=( a16527a  and  a16522a );
 a16531a <=( (not A167)  and  (not A169) );
 a16535a <=( A200  and  (not A199) );
 a16536a <=( (not A166)  and  a16535a );
 a16537a <=( a16536a  and  a16531a );
 a16541a <=( A265  and  (not A234) );
 a16542a <=( (not A233)  and  a16541a );
 a16546a <=( A299  and  (not A298) );
 a16547a <=( A266  and  a16546a );
 a16548a <=( a16547a  and  a16542a );
 a16551a <=( (not A167)  and  (not A169) );
 a16555a <=( A200  and  (not A199) );
 a16556a <=( (not A166)  and  a16555a );
 a16557a <=( a16556a  and  a16551a );
 a16561a <=( (not A266)  and  (not A234) );
 a16562a <=( (not A233)  and  a16561a );
 a16566a <=( A299  and  (not A298) );
 a16567a <=( (not A267)  and  a16566a );
 a16568a <=( a16567a  and  a16562a );
 a16571a <=( (not A167)  and  (not A169) );
 a16575a <=( A200  and  (not A199) );
 a16576a <=( (not A166)  and  a16575a );
 a16577a <=( a16576a  and  a16571a );
 a16581a <=( (not A265)  and  (not A234) );
 a16582a <=( (not A233)  and  a16581a );
 a16586a <=( A299  and  (not A298) );
 a16587a <=( (not A266)  and  a16586a );
 a16588a <=( a16587a  and  a16582a );
 a16591a <=( (not A167)  and  (not A169) );
 a16595a <=( A200  and  (not A199) );
 a16596a <=( (not A166)  and  a16595a );
 a16597a <=( a16596a  and  a16591a );
 a16601a <=( A234  and  (not A233) );
 a16602a <=( A232  and  a16601a );
 a16606a <=( (not A300)  and  A298 );
 a16607a <=( A235  and  a16606a );
 a16608a <=( a16607a  and  a16602a );
 a16611a <=( (not A167)  and  (not A169) );
 a16615a <=( A200  and  (not A199) );
 a16616a <=( (not A166)  and  a16615a );
 a16617a <=( a16616a  and  a16611a );
 a16621a <=( A234  and  (not A233) );
 a16622a <=( A232  and  a16621a );
 a16626a <=( A299  and  A298 );
 a16627a <=( A235  and  a16626a );
 a16628a <=( a16627a  and  a16622a );
 a16631a <=( (not A167)  and  (not A169) );
 a16635a <=( A200  and  (not A199) );
 a16636a <=( (not A166)  and  a16635a );
 a16637a <=( a16636a  and  a16631a );
 a16641a <=( A234  and  (not A233) );
 a16642a <=( A232  and  a16641a );
 a16646a <=( (not A299)  and  (not A298) );
 a16647a <=( A235  and  a16646a );
 a16648a <=( a16647a  and  a16642a );
 a16651a <=( (not A167)  and  (not A169) );
 a16655a <=( A200  and  (not A199) );
 a16656a <=( (not A166)  and  a16655a );
 a16657a <=( a16656a  and  a16651a );
 a16661a <=( A234  and  (not A233) );
 a16662a <=( A232  and  a16661a );
 a16666a <=( A266  and  (not A265) );
 a16667a <=( A235  and  a16666a );
 a16668a <=( a16667a  and  a16662a );
 a16671a <=( (not A167)  and  (not A169) );
 a16675a <=( A200  and  (not A199) );
 a16676a <=( (not A166)  and  a16675a );
 a16677a <=( a16676a  and  a16671a );
 a16681a <=( A234  and  (not A233) );
 a16682a <=( A232  and  a16681a );
 a16686a <=( (not A300)  and  A298 );
 a16687a <=( A236  and  a16686a );
 a16688a <=( a16687a  and  a16682a );
 a16691a <=( (not A167)  and  (not A169) );
 a16695a <=( A200  and  (not A199) );
 a16696a <=( (not A166)  and  a16695a );
 a16697a <=( a16696a  and  a16691a );
 a16701a <=( A234  and  (not A233) );
 a16702a <=( A232  and  a16701a );
 a16706a <=( A299  and  A298 );
 a16707a <=( A236  and  a16706a );
 a16708a <=( a16707a  and  a16702a );
 a16711a <=( (not A167)  and  (not A169) );
 a16715a <=( A200  and  (not A199) );
 a16716a <=( (not A166)  and  a16715a );
 a16717a <=( a16716a  and  a16711a );
 a16721a <=( A234  and  (not A233) );
 a16722a <=( A232  and  a16721a );
 a16726a <=( (not A299)  and  (not A298) );
 a16727a <=( A236  and  a16726a );
 a16728a <=( a16727a  and  a16722a );
 a16731a <=( (not A167)  and  (not A169) );
 a16735a <=( A200  and  (not A199) );
 a16736a <=( (not A166)  and  a16735a );
 a16737a <=( a16736a  and  a16731a );
 a16741a <=( A234  and  (not A233) );
 a16742a <=( A232  and  a16741a );
 a16746a <=( A266  and  (not A265) );
 a16747a <=( A236  and  a16746a );
 a16748a <=( a16747a  and  a16742a );
 a16751a <=( (not A167)  and  (not A169) );
 a16755a <=( A200  and  (not A199) );
 a16756a <=( (not A166)  and  a16755a );
 a16757a <=( a16756a  and  a16751a );
 a16761a <=( A265  and  (not A233) );
 a16762a <=( (not A232)  and  a16761a );
 a16766a <=( A299  and  (not A298) );
 a16767a <=( A266  and  a16766a );
 a16768a <=( a16767a  and  a16762a );
 a16771a <=( (not A167)  and  (not A169) );
 a16775a <=( A200  and  (not A199) );
 a16776a <=( (not A166)  and  a16775a );
 a16777a <=( a16776a  and  a16771a );
 a16781a <=( (not A266)  and  (not A233) );
 a16782a <=( (not A232)  and  a16781a );
 a16786a <=( A299  and  (not A298) );
 a16787a <=( (not A267)  and  a16786a );
 a16788a <=( a16787a  and  a16782a );
 a16791a <=( (not A167)  and  (not A169) );
 a16795a <=( A200  and  (not A199) );
 a16796a <=( (not A166)  and  a16795a );
 a16797a <=( a16796a  and  a16791a );
 a16801a <=( (not A265)  and  (not A233) );
 a16802a <=( (not A232)  and  a16801a );
 a16806a <=( A299  and  (not A298) );
 a16807a <=( (not A266)  and  a16806a );
 a16808a <=( a16807a  and  a16802a );
 a16811a <=( (not A167)  and  (not A169) );
 a16815a <=( (not A200)  and  A199 );
 a16816a <=( (not A166)  and  a16815a );
 a16817a <=( a16816a  and  a16811a );
 a16821a <=( (not A232)  and  A202 );
 a16822a <=( A201  and  a16821a );
 a16826a <=( (not A300)  and  (not A299) );
 a16827a <=( A233  and  a16826a );
 a16828a <=( a16827a  and  a16822a );
 a16831a <=( (not A167)  and  (not A169) );
 a16835a <=( (not A200)  and  A199 );
 a16836a <=( (not A166)  and  a16835a );
 a16837a <=( a16836a  and  a16831a );
 a16841a <=( (not A232)  and  A202 );
 a16842a <=( A201  and  a16841a );
 a16846a <=( A299  and  A298 );
 a16847a <=( A233  and  a16846a );
 a16848a <=( a16847a  and  a16842a );
 a16851a <=( (not A167)  and  (not A169) );
 a16855a <=( (not A200)  and  A199 );
 a16856a <=( (not A166)  and  a16855a );
 a16857a <=( a16856a  and  a16851a );
 a16861a <=( (not A232)  and  A202 );
 a16862a <=( A201  and  a16861a );
 a16866a <=( (not A299)  and  (not A298) );
 a16867a <=( A233  and  a16866a );
 a16868a <=( a16867a  and  a16862a );
 a16871a <=( (not A167)  and  (not A169) );
 a16875a <=( (not A200)  and  A199 );
 a16876a <=( (not A166)  and  a16875a );
 a16877a <=( a16876a  and  a16871a );
 a16881a <=( (not A232)  and  A202 );
 a16882a <=( A201  and  a16881a );
 a16886a <=( A266  and  (not A265) );
 a16887a <=( A233  and  a16886a );
 a16888a <=( a16887a  and  a16882a );
 a16891a <=( (not A167)  and  (not A169) );
 a16895a <=( (not A200)  and  A199 );
 a16896a <=( (not A166)  and  a16895a );
 a16897a <=( a16896a  and  a16891a );
 a16901a <=( (not A232)  and  A203 );
 a16902a <=( A201  and  a16901a );
 a16906a <=( (not A300)  and  (not A299) );
 a16907a <=( A233  and  a16906a );
 a16908a <=( a16907a  and  a16902a );
 a16911a <=( (not A167)  and  (not A169) );
 a16915a <=( (not A200)  and  A199 );
 a16916a <=( (not A166)  and  a16915a );
 a16917a <=( a16916a  and  a16911a );
 a16921a <=( (not A232)  and  A203 );
 a16922a <=( A201  and  a16921a );
 a16926a <=( A299  and  A298 );
 a16927a <=( A233  and  a16926a );
 a16928a <=( a16927a  and  a16922a );
 a16931a <=( (not A167)  and  (not A169) );
 a16935a <=( (not A200)  and  A199 );
 a16936a <=( (not A166)  and  a16935a );
 a16937a <=( a16936a  and  a16931a );
 a16941a <=( (not A232)  and  A203 );
 a16942a <=( A201  and  a16941a );
 a16946a <=( (not A299)  and  (not A298) );
 a16947a <=( A233  and  a16946a );
 a16948a <=( a16947a  and  a16942a );
 a16951a <=( (not A167)  and  (not A169) );
 a16955a <=( (not A200)  and  A199 );
 a16956a <=( (not A166)  and  a16955a );
 a16957a <=( a16956a  and  a16951a );
 a16961a <=( (not A232)  and  A203 );
 a16962a <=( A201  and  a16961a );
 a16966a <=( A266  and  (not A265) );
 a16967a <=( A233  and  a16966a );
 a16968a <=( a16967a  and  a16962a );
 a16971a <=( (not A168)  and  (not A169) );
 a16975a <=( (not A199)  and  A166 );
 a16976a <=( A167  and  a16975a );
 a16977a <=( a16976a  and  a16971a );
 a16981a <=( A233  and  (not A232) );
 a16982a <=( A200  and  a16981a );
 a16986a <=( (not A302)  and  (not A301) );
 a16987a <=( (not A299)  and  a16986a );
 a16988a <=( a16987a  and  a16982a );
 a16991a <=( (not A169)  and  A170 );
 a16995a <=( A199  and  (not A166) );
 a16996a <=( A167  and  a16995a );
 a16997a <=( a16996a  and  a16991a );
 a17001a <=( A233  and  (not A232) );
 a17002a <=( A200  and  a17001a );
 a17006a <=( (not A302)  and  (not A301) );
 a17007a <=( (not A299)  and  a17006a );
 a17008a <=( a17007a  and  a17002a );
 a17011a <=( (not A169)  and  A170 );
 a17015a <=( (not A200)  and  (not A166) );
 a17016a <=( A167  and  a17015a );
 a17017a <=( a17016a  and  a17011a );
 a17021a <=( (not A232)  and  (not A203) );
 a17022a <=( (not A202)  and  a17021a );
 a17026a <=( (not A300)  and  (not A299) );
 a17027a <=( A233  and  a17026a );
 a17028a <=( a17027a  and  a17022a );
 a17031a <=( (not A169)  and  A170 );
 a17035a <=( (not A200)  and  (not A166) );
 a17036a <=( A167  and  a17035a );
 a17037a <=( a17036a  and  a17031a );
 a17041a <=( (not A232)  and  (not A203) );
 a17042a <=( (not A202)  and  a17041a );
 a17046a <=( A299  and  A298 );
 a17047a <=( A233  and  a17046a );
 a17048a <=( a17047a  and  a17042a );
 a17051a <=( (not A169)  and  A170 );
 a17055a <=( (not A200)  and  (not A166) );
 a17056a <=( A167  and  a17055a );
 a17057a <=( a17056a  and  a17051a );
 a17061a <=( (not A232)  and  (not A203) );
 a17062a <=( (not A202)  and  a17061a );
 a17066a <=( (not A299)  and  (not A298) );
 a17067a <=( A233  and  a17066a );
 a17068a <=( a17067a  and  a17062a );
 a17071a <=( (not A169)  and  A170 );
 a17075a <=( (not A200)  and  (not A166) );
 a17076a <=( A167  and  a17075a );
 a17077a <=( a17076a  and  a17071a );
 a17081a <=( (not A232)  and  (not A203) );
 a17082a <=( (not A202)  and  a17081a );
 a17086a <=( A266  and  (not A265) );
 a17087a <=( A233  and  a17086a );
 a17088a <=( a17087a  and  a17082a );
 a17091a <=( (not A169)  and  A170 );
 a17095a <=( (not A200)  and  (not A166) );
 a17096a <=( A167  and  a17095a );
 a17097a <=( a17096a  and  a17091a );
 a17101a <=( A233  and  (not A232) );
 a17102a <=( (not A201)  and  a17101a );
 a17106a <=( (not A302)  and  (not A301) );
 a17107a <=( (not A299)  and  a17106a );
 a17108a <=( a17107a  and  a17102a );
 a17111a <=( (not A169)  and  A170 );
 a17115a <=( (not A199)  and  (not A166) );
 a17116a <=( A167  and  a17115a );
 a17117a <=( a17116a  and  a17111a );
 a17121a <=( A233  and  (not A232) );
 a17122a <=( (not A200)  and  a17121a );
 a17126a <=( (not A302)  and  (not A301) );
 a17127a <=( (not A299)  and  a17126a );
 a17128a <=( a17127a  and  a17122a );
 a17131a <=( (not A169)  and  A170 );
 a17135a <=( A199  and  A166 );
 a17136a <=( (not A167)  and  a17135a );
 a17137a <=( a17136a  and  a17131a );
 a17141a <=( A233  and  (not A232) );
 a17142a <=( A200  and  a17141a );
 a17146a <=( (not A302)  and  (not A301) );
 a17147a <=( (not A299)  and  a17146a );
 a17148a <=( a17147a  and  a17142a );
 a17151a <=( (not A169)  and  A170 );
 a17155a <=( (not A200)  and  A166 );
 a17156a <=( (not A167)  and  a17155a );
 a17157a <=( a17156a  and  a17151a );
 a17161a <=( (not A232)  and  (not A203) );
 a17162a <=( (not A202)  and  a17161a );
 a17166a <=( (not A300)  and  (not A299) );
 a17167a <=( A233  and  a17166a );
 a17168a <=( a17167a  and  a17162a );
 a17171a <=( (not A169)  and  A170 );
 a17175a <=( (not A200)  and  A166 );
 a17176a <=( (not A167)  and  a17175a );
 a17177a <=( a17176a  and  a17171a );
 a17181a <=( (not A232)  and  (not A203) );
 a17182a <=( (not A202)  and  a17181a );
 a17186a <=( A299  and  A298 );
 a17187a <=( A233  and  a17186a );
 a17188a <=( a17187a  and  a17182a );
 a17191a <=( (not A169)  and  A170 );
 a17195a <=( (not A200)  and  A166 );
 a17196a <=( (not A167)  and  a17195a );
 a17197a <=( a17196a  and  a17191a );
 a17201a <=( (not A232)  and  (not A203) );
 a17202a <=( (not A202)  and  a17201a );
 a17206a <=( (not A299)  and  (not A298) );
 a17207a <=( A233  and  a17206a );
 a17208a <=( a17207a  and  a17202a );
 a17211a <=( (not A169)  and  A170 );
 a17215a <=( (not A200)  and  A166 );
 a17216a <=( (not A167)  and  a17215a );
 a17217a <=( a17216a  and  a17211a );
 a17221a <=( (not A232)  and  (not A203) );
 a17222a <=( (not A202)  and  a17221a );
 a17226a <=( A266  and  (not A265) );
 a17227a <=( A233  and  a17226a );
 a17228a <=( a17227a  and  a17222a );
 a17231a <=( (not A169)  and  A170 );
 a17235a <=( (not A200)  and  A166 );
 a17236a <=( (not A167)  and  a17235a );
 a17237a <=( a17236a  and  a17231a );
 a17241a <=( A233  and  (not A232) );
 a17242a <=( (not A201)  and  a17241a );
 a17246a <=( (not A302)  and  (not A301) );
 a17247a <=( (not A299)  and  a17246a );
 a17248a <=( a17247a  and  a17242a );
 a17251a <=( (not A169)  and  A170 );
 a17255a <=( (not A199)  and  A166 );
 a17256a <=( (not A167)  and  a17255a );
 a17257a <=( a17256a  and  a17251a );
 a17261a <=( A233  and  (not A232) );
 a17262a <=( (not A200)  and  a17261a );
 a17266a <=( (not A302)  and  (not A301) );
 a17267a <=( (not A299)  and  a17266a );
 a17268a <=( a17267a  and  a17262a );
 a17271a <=( (not A169)  and  (not A170) );
 a17275a <=( (not A200)  and  A199 );
 a17276a <=( (not A168)  and  a17275a );
 a17277a <=( a17276a  and  a17271a );
 a17281a <=( (not A232)  and  A202 );
 a17282a <=( A201  and  a17281a );
 a17286a <=( (not A300)  and  (not A299) );
 a17287a <=( A233  and  a17286a );
 a17288a <=( a17287a  and  a17282a );
 a17291a <=( (not A169)  and  (not A170) );
 a17295a <=( (not A200)  and  A199 );
 a17296a <=( (not A168)  and  a17295a );
 a17297a <=( a17296a  and  a17291a );
 a17301a <=( (not A232)  and  A202 );
 a17302a <=( A201  and  a17301a );
 a17306a <=( A299  and  A298 );
 a17307a <=( A233  and  a17306a );
 a17308a <=( a17307a  and  a17302a );
 a17311a <=( (not A169)  and  (not A170) );
 a17315a <=( (not A200)  and  A199 );
 a17316a <=( (not A168)  and  a17315a );
 a17317a <=( a17316a  and  a17311a );
 a17321a <=( (not A232)  and  A202 );
 a17322a <=( A201  and  a17321a );
 a17326a <=( (not A299)  and  (not A298) );
 a17327a <=( A233  and  a17326a );
 a17328a <=( a17327a  and  a17322a );
 a17331a <=( (not A169)  and  (not A170) );
 a17335a <=( (not A200)  and  A199 );
 a17336a <=( (not A168)  and  a17335a );
 a17337a <=( a17336a  and  a17331a );
 a17341a <=( (not A232)  and  A202 );
 a17342a <=( A201  and  a17341a );
 a17346a <=( A266  and  (not A265) );
 a17347a <=( A233  and  a17346a );
 a17348a <=( a17347a  and  a17342a );
 a17351a <=( (not A169)  and  (not A170) );
 a17355a <=( (not A200)  and  A199 );
 a17356a <=( (not A168)  and  a17355a );
 a17357a <=( a17356a  and  a17351a );
 a17361a <=( (not A232)  and  A203 );
 a17362a <=( A201  and  a17361a );
 a17366a <=( (not A300)  and  (not A299) );
 a17367a <=( A233  and  a17366a );
 a17368a <=( a17367a  and  a17362a );
 a17371a <=( (not A169)  and  (not A170) );
 a17375a <=( (not A200)  and  A199 );
 a17376a <=( (not A168)  and  a17375a );
 a17377a <=( a17376a  and  a17371a );
 a17381a <=( (not A232)  and  A203 );
 a17382a <=( A201  and  a17381a );
 a17386a <=( A299  and  A298 );
 a17387a <=( A233  and  a17386a );
 a17388a <=( a17387a  and  a17382a );
 a17391a <=( (not A169)  and  (not A170) );
 a17395a <=( (not A200)  and  A199 );
 a17396a <=( (not A168)  and  a17395a );
 a17397a <=( a17396a  and  a17391a );
 a17401a <=( (not A232)  and  A203 );
 a17402a <=( A201  and  a17401a );
 a17406a <=( (not A299)  and  (not A298) );
 a17407a <=( A233  and  a17406a );
 a17408a <=( a17407a  and  a17402a );
 a17411a <=( (not A169)  and  (not A170) );
 a17415a <=( (not A200)  and  A199 );
 a17416a <=( (not A168)  and  a17415a );
 a17417a <=( a17416a  and  a17411a );
 a17421a <=( (not A232)  and  A203 );
 a17422a <=( A201  and  a17421a );
 a17426a <=( A266  and  (not A265) );
 a17427a <=( A233  and  a17426a );
 a17428a <=( a17427a  and  a17422a );
 a17432a <=( A199  and  A166 );
 a17433a <=( A168  and  a17432a );
 a17437a <=( A233  and  A232 );
 a17438a <=( A200  and  a17437a );
 a17439a <=( a17438a  and  a17433a );
 a17443a <=( A298  and  (not A267) );
 a17444a <=( A265  and  a17443a );
 a17448a <=( A301  and  A300 );
 a17449a <=( (not A299)  and  a17448a );
 a17450a <=( a17449a  and  a17444a );
 a17454a <=( A199  and  A166 );
 a17455a <=( A168  and  a17454a );
 a17459a <=( A233  and  A232 );
 a17460a <=( A200  and  a17459a );
 a17461a <=( a17460a  and  a17455a );
 a17465a <=( A298  and  (not A267) );
 a17466a <=( A265  and  a17465a );
 a17470a <=( A302  and  A300 );
 a17471a <=( (not A299)  and  a17470a );
 a17472a <=( a17471a  and  a17466a );
 a17476a <=( A199  and  A166 );
 a17477a <=( A168  and  a17476a );
 a17481a <=( A233  and  A232 );
 a17482a <=( A200  and  a17481a );
 a17483a <=( a17482a  and  a17477a );
 a17487a <=( A298  and  A266 );
 a17488a <=( A265  and  a17487a );
 a17492a <=( A301  and  A300 );
 a17493a <=( (not A299)  and  a17492a );
 a17494a <=( a17493a  and  a17488a );
 a17498a <=( A199  and  A166 );
 a17499a <=( A168  and  a17498a );
 a17503a <=( A233  and  A232 );
 a17504a <=( A200  and  a17503a );
 a17505a <=( a17504a  and  a17499a );
 a17509a <=( A298  and  A266 );
 a17510a <=( A265  and  a17509a );
 a17514a <=( A302  and  A300 );
 a17515a <=( (not A299)  and  a17514a );
 a17516a <=( a17515a  and  a17510a );
 a17520a <=( A199  and  A166 );
 a17521a <=( A168  and  a17520a );
 a17525a <=( A233  and  A232 );
 a17526a <=( A200  and  a17525a );
 a17527a <=( a17526a  and  a17521a );
 a17531a <=( A298  and  (not A266) );
 a17532a <=( (not A265)  and  a17531a );
 a17536a <=( A301  and  A300 );
 a17537a <=( (not A299)  and  a17536a );
 a17538a <=( a17537a  and  a17532a );
 a17542a <=( A199  and  A166 );
 a17543a <=( A168  and  a17542a );
 a17547a <=( A233  and  A232 );
 a17548a <=( A200  and  a17547a );
 a17549a <=( a17548a  and  a17543a );
 a17553a <=( A298  and  (not A266) );
 a17554a <=( (not A265)  and  a17553a );
 a17558a <=( A302  and  A300 );
 a17559a <=( (not A299)  and  a17558a );
 a17560a <=( a17559a  and  a17554a );
 a17564a <=( A199  and  A166 );
 a17565a <=( A168  and  a17564a );
 a17569a <=( (not A235)  and  (not A233) );
 a17570a <=( A200  and  a17569a );
 a17571a <=( a17570a  and  a17565a );
 a17575a <=( (not A268)  and  (not A266) );
 a17576a <=( (not A236)  and  a17575a );
 a17580a <=( A299  and  (not A298) );
 a17581a <=( (not A269)  and  a17580a );
 a17582a <=( a17581a  and  a17576a );
 a17586a <=( A199  and  A166 );
 a17587a <=( A168  and  a17586a );
 a17591a <=( (not A234)  and  (not A233) );
 a17592a <=( A200  and  a17591a );
 a17593a <=( a17592a  and  a17587a );
 a17597a <=( A298  and  A266 );
 a17598a <=( A265  and  a17597a );
 a17602a <=( A301  and  A300 );
 a17603a <=( (not A299)  and  a17602a );
 a17604a <=( a17603a  and  a17598a );
 a17608a <=( A199  and  A166 );
 a17609a <=( A168  and  a17608a );
 a17613a <=( (not A234)  and  (not A233) );
 a17614a <=( A200  and  a17613a );
 a17615a <=( a17614a  and  a17609a );
 a17619a <=( A298  and  A266 );
 a17620a <=( A265  and  a17619a );
 a17624a <=( A302  and  A300 );
 a17625a <=( (not A299)  and  a17624a );
 a17626a <=( a17625a  and  a17620a );
 a17630a <=( A199  and  A166 );
 a17631a <=( A168  and  a17630a );
 a17635a <=( (not A234)  and  (not A233) );
 a17636a <=( A200  and  a17635a );
 a17637a <=( a17636a  and  a17631a );
 a17641a <=( A298  and  (not A267) );
 a17642a <=( (not A266)  and  a17641a );
 a17646a <=( A301  and  A300 );
 a17647a <=( (not A299)  and  a17646a );
 a17648a <=( a17647a  and  a17642a );
 a17652a <=( A199  and  A166 );
 a17653a <=( A168  and  a17652a );
 a17657a <=( (not A234)  and  (not A233) );
 a17658a <=( A200  and  a17657a );
 a17659a <=( a17658a  and  a17653a );
 a17663a <=( A298  and  (not A267) );
 a17664a <=( (not A266)  and  a17663a );
 a17668a <=( A302  and  A300 );
 a17669a <=( (not A299)  and  a17668a );
 a17670a <=( a17669a  and  a17664a );
 a17674a <=( A199  and  A166 );
 a17675a <=( A168  and  a17674a );
 a17679a <=( (not A234)  and  (not A233) );
 a17680a <=( A200  and  a17679a );
 a17681a <=( a17680a  and  a17675a );
 a17685a <=( A298  and  (not A266) );
 a17686a <=( (not A265)  and  a17685a );
 a17690a <=( A301  and  A300 );
 a17691a <=( (not A299)  and  a17690a );
 a17692a <=( a17691a  and  a17686a );
 a17696a <=( A199  and  A166 );
 a17697a <=( A168  and  a17696a );
 a17701a <=( (not A234)  and  (not A233) );
 a17702a <=( A200  and  a17701a );
 a17703a <=( a17702a  and  a17697a );
 a17707a <=( A298  and  (not A266) );
 a17708a <=( (not A265)  and  a17707a );
 a17712a <=( A302  and  A300 );
 a17713a <=( (not A299)  and  a17712a );
 a17714a <=( a17713a  and  a17708a );
 a17718a <=( A199  and  A166 );
 a17719a <=( A168  and  a17718a );
 a17723a <=( (not A233)  and  A232 );
 a17724a <=( A200  and  a17723a );
 a17725a <=( a17724a  and  a17719a );
 a17729a <=( A265  and  A235 );
 a17730a <=( A234  and  a17729a );
 a17734a <=( A268  and  A267 );
 a17735a <=( (not A266)  and  a17734a );
 a17736a <=( a17735a  and  a17730a );
 a17740a <=( A199  and  A166 );
 a17741a <=( A168  and  a17740a );
 a17745a <=( (not A233)  and  A232 );
 a17746a <=( A200  and  a17745a );
 a17747a <=( a17746a  and  a17741a );
 a17751a <=( A265  and  A235 );
 a17752a <=( A234  and  a17751a );
 a17756a <=( A269  and  A267 );
 a17757a <=( (not A266)  and  a17756a );
 a17758a <=( a17757a  and  a17752a );
 a17762a <=( A199  and  A166 );
 a17763a <=( A168  and  a17762a );
 a17767a <=( (not A233)  and  A232 );
 a17768a <=( A200  and  a17767a );
 a17769a <=( a17768a  and  a17763a );
 a17773a <=( A265  and  A236 );
 a17774a <=( A234  and  a17773a );
 a17778a <=( A268  and  A267 );
 a17779a <=( (not A266)  and  a17778a );
 a17780a <=( a17779a  and  a17774a );
 a17784a <=( A199  and  A166 );
 a17785a <=( A168  and  a17784a );
 a17789a <=( (not A233)  and  A232 );
 a17790a <=( A200  and  a17789a );
 a17791a <=( a17790a  and  a17785a );
 a17795a <=( A265  and  A236 );
 a17796a <=( A234  and  a17795a );
 a17800a <=( A269  and  A267 );
 a17801a <=( (not A266)  and  a17800a );
 a17802a <=( a17801a  and  a17796a );
 a17806a <=( A199  and  A166 );
 a17807a <=( A168  and  a17806a );
 a17811a <=( (not A233)  and  (not A232) );
 a17812a <=( A200  and  a17811a );
 a17813a <=( a17812a  and  a17807a );
 a17817a <=( A298  and  A266 );
 a17818a <=( A265  and  a17817a );
 a17822a <=( A301  and  A300 );
 a17823a <=( (not A299)  and  a17822a );
 a17824a <=( a17823a  and  a17818a );
 a17828a <=( A199  and  A166 );
 a17829a <=( A168  and  a17828a );
 a17833a <=( (not A233)  and  (not A232) );
 a17834a <=( A200  and  a17833a );
 a17835a <=( a17834a  and  a17829a );
 a17839a <=( A298  and  A266 );
 a17840a <=( A265  and  a17839a );
 a17844a <=( A302  and  A300 );
 a17845a <=( (not A299)  and  a17844a );
 a17846a <=( a17845a  and  a17840a );
 a17850a <=( A199  and  A166 );
 a17851a <=( A168  and  a17850a );
 a17855a <=( (not A233)  and  (not A232) );
 a17856a <=( A200  and  a17855a );
 a17857a <=( a17856a  and  a17851a );
 a17861a <=( A298  and  (not A267) );
 a17862a <=( (not A266)  and  a17861a );
 a17866a <=( A301  and  A300 );
 a17867a <=( (not A299)  and  a17866a );
 a17868a <=( a17867a  and  a17862a );
 a17872a <=( A199  and  A166 );
 a17873a <=( A168  and  a17872a );
 a17877a <=( (not A233)  and  (not A232) );
 a17878a <=( A200  and  a17877a );
 a17879a <=( a17878a  and  a17873a );
 a17883a <=( A298  and  (not A267) );
 a17884a <=( (not A266)  and  a17883a );
 a17888a <=( A302  and  A300 );
 a17889a <=( (not A299)  and  a17888a );
 a17890a <=( a17889a  and  a17884a );
 a17894a <=( A199  and  A166 );
 a17895a <=( A168  and  a17894a );
 a17899a <=( (not A233)  and  (not A232) );
 a17900a <=( A200  and  a17899a );
 a17901a <=( a17900a  and  a17895a );
 a17905a <=( A298  and  (not A266) );
 a17906a <=( (not A265)  and  a17905a );
 a17910a <=( A301  and  A300 );
 a17911a <=( (not A299)  and  a17910a );
 a17912a <=( a17911a  and  a17906a );
 a17916a <=( A199  and  A166 );
 a17917a <=( A168  and  a17916a );
 a17921a <=( (not A233)  and  (not A232) );
 a17922a <=( A200  and  a17921a );
 a17923a <=( a17922a  and  a17917a );
 a17927a <=( A298  and  (not A266) );
 a17928a <=( (not A265)  and  a17927a );
 a17932a <=( A302  and  A300 );
 a17933a <=( (not A299)  and  a17932a );
 a17934a <=( a17933a  and  a17928a );
 a17938a <=( (not A200)  and  A166 );
 a17939a <=( A168  and  a17938a );
 a17943a <=( A232  and  (not A203) );
 a17944a <=( (not A202)  and  a17943a );
 a17945a <=( a17944a  and  a17939a );
 a17949a <=( (not A268)  and  A265 );
 a17950a <=( A233  and  a17949a );
 a17954a <=( A299  and  (not A298) );
 a17955a <=( (not A269)  and  a17954a );
 a17956a <=( a17955a  and  a17950a );
 a17960a <=( (not A200)  and  A166 );
 a17961a <=( A168  and  a17960a );
 a17965a <=( (not A233)  and  (not A203) );
 a17966a <=( (not A202)  and  a17965a );
 a17967a <=( a17966a  and  a17961a );
 a17971a <=( A265  and  (not A236) );
 a17972a <=( (not A235)  and  a17971a );
 a17976a <=( A299  and  (not A298) );
 a17977a <=( A266  and  a17976a );
 a17978a <=( a17977a  and  a17972a );
 a17982a <=( (not A200)  and  A166 );
 a17983a <=( A168  and  a17982a );
 a17987a <=( (not A233)  and  (not A203) );
 a17988a <=( (not A202)  and  a17987a );
 a17989a <=( a17988a  and  a17983a );
 a17993a <=( (not A266)  and  (not A236) );
 a17994a <=( (not A235)  and  a17993a );
 a17998a <=( A299  and  (not A298) );
 a17999a <=( (not A267)  and  a17998a );
 a18000a <=( a17999a  and  a17994a );
 a18004a <=( (not A200)  and  A166 );
 a18005a <=( A168  and  a18004a );
 a18009a <=( (not A233)  and  (not A203) );
 a18010a <=( (not A202)  and  a18009a );
 a18011a <=( a18010a  and  a18005a );
 a18015a <=( (not A265)  and  (not A236) );
 a18016a <=( (not A235)  and  a18015a );
 a18020a <=( A299  and  (not A298) );
 a18021a <=( (not A266)  and  a18020a );
 a18022a <=( a18021a  and  a18016a );
 a18026a <=( (not A200)  and  A166 );
 a18027a <=( A168  and  a18026a );
 a18031a <=( (not A233)  and  (not A203) );
 a18032a <=( (not A202)  and  a18031a );
 a18033a <=( a18032a  and  a18027a );
 a18037a <=( (not A268)  and  (not A266) );
 a18038a <=( (not A234)  and  a18037a );
 a18042a <=( A299  and  (not A298) );
 a18043a <=( (not A269)  and  a18042a );
 a18044a <=( a18043a  and  a18038a );
 a18048a <=( (not A200)  and  A166 );
 a18049a <=( A168  and  a18048a );
 a18053a <=( A232  and  (not A203) );
 a18054a <=( (not A202)  and  a18053a );
 a18055a <=( a18054a  and  a18049a );
 a18059a <=( A235  and  A234 );
 a18060a <=( (not A233)  and  a18059a );
 a18064a <=( (not A302)  and  (not A301) );
 a18065a <=( A298  and  a18064a );
 a18066a <=( a18065a  and  a18060a );
 a18070a <=( (not A200)  and  A166 );
 a18071a <=( A168  and  a18070a );
 a18075a <=( A232  and  (not A203) );
 a18076a <=( (not A202)  and  a18075a );
 a18077a <=( a18076a  and  a18071a );
 a18081a <=( A236  and  A234 );
 a18082a <=( (not A233)  and  a18081a );
 a18086a <=( (not A302)  and  (not A301) );
 a18087a <=( A298  and  a18086a );
 a18088a <=( a18087a  and  a18082a );
 a18092a <=( (not A200)  and  A166 );
 a18093a <=( A168  and  a18092a );
 a18097a <=( (not A232)  and  (not A203) );
 a18098a <=( (not A202)  and  a18097a );
 a18099a <=( a18098a  and  a18093a );
 a18103a <=( (not A268)  and  (not A266) );
 a18104a <=( (not A233)  and  a18103a );
 a18108a <=( A299  and  (not A298) );
 a18109a <=( (not A269)  and  a18108a );
 a18110a <=( a18109a  and  a18104a );
 a18114a <=( (not A200)  and  A166 );
 a18115a <=( A168  and  a18114a );
 a18119a <=( A233  and  A232 );
 a18120a <=( (not A201)  and  a18119a );
 a18121a <=( a18120a  and  a18115a );
 a18125a <=( A298  and  (not A267) );
 a18126a <=( A265  and  a18125a );
 a18130a <=( A301  and  A300 );
 a18131a <=( (not A299)  and  a18130a );
 a18132a <=( a18131a  and  a18126a );
 a18136a <=( (not A200)  and  A166 );
 a18137a <=( A168  and  a18136a );
 a18141a <=( A233  and  A232 );
 a18142a <=( (not A201)  and  a18141a );
 a18143a <=( a18142a  and  a18137a );
 a18147a <=( A298  and  (not A267) );
 a18148a <=( A265  and  a18147a );
 a18152a <=( A302  and  A300 );
 a18153a <=( (not A299)  and  a18152a );
 a18154a <=( a18153a  and  a18148a );
 a18158a <=( (not A200)  and  A166 );
 a18159a <=( A168  and  a18158a );
 a18163a <=( A233  and  A232 );
 a18164a <=( (not A201)  and  a18163a );
 a18165a <=( a18164a  and  a18159a );
 a18169a <=( A298  and  A266 );
 a18170a <=( A265  and  a18169a );
 a18174a <=( A301  and  A300 );
 a18175a <=( (not A299)  and  a18174a );
 a18176a <=( a18175a  and  a18170a );
 a18180a <=( (not A200)  and  A166 );
 a18181a <=( A168  and  a18180a );
 a18185a <=( A233  and  A232 );
 a18186a <=( (not A201)  and  a18185a );
 a18187a <=( a18186a  and  a18181a );
 a18191a <=( A298  and  A266 );
 a18192a <=( A265  and  a18191a );
 a18196a <=( A302  and  A300 );
 a18197a <=( (not A299)  and  a18196a );
 a18198a <=( a18197a  and  a18192a );
 a18202a <=( (not A200)  and  A166 );
 a18203a <=( A168  and  a18202a );
 a18207a <=( A233  and  A232 );
 a18208a <=( (not A201)  and  a18207a );
 a18209a <=( a18208a  and  a18203a );
 a18213a <=( A298  and  (not A266) );
 a18214a <=( (not A265)  and  a18213a );
 a18218a <=( A301  and  A300 );
 a18219a <=( (not A299)  and  a18218a );
 a18220a <=( a18219a  and  a18214a );
 a18224a <=( (not A200)  and  A166 );
 a18225a <=( A168  and  a18224a );
 a18229a <=( A233  and  A232 );
 a18230a <=( (not A201)  and  a18229a );
 a18231a <=( a18230a  and  a18225a );
 a18235a <=( A298  and  (not A266) );
 a18236a <=( (not A265)  and  a18235a );
 a18240a <=( A302  and  A300 );
 a18241a <=( (not A299)  and  a18240a );
 a18242a <=( a18241a  and  a18236a );
 a18246a <=( (not A200)  and  A166 );
 a18247a <=( A168  and  a18246a );
 a18251a <=( (not A235)  and  (not A233) );
 a18252a <=( (not A201)  and  a18251a );
 a18253a <=( a18252a  and  a18247a );
 a18257a <=( (not A268)  and  (not A266) );
 a18258a <=( (not A236)  and  a18257a );
 a18262a <=( A299  and  (not A298) );
 a18263a <=( (not A269)  and  a18262a );
 a18264a <=( a18263a  and  a18258a );
 a18268a <=( (not A200)  and  A166 );
 a18269a <=( A168  and  a18268a );
 a18273a <=( (not A234)  and  (not A233) );
 a18274a <=( (not A201)  and  a18273a );
 a18275a <=( a18274a  and  a18269a );
 a18279a <=( A298  and  A266 );
 a18280a <=( A265  and  a18279a );
 a18284a <=( A301  and  A300 );
 a18285a <=( (not A299)  and  a18284a );
 a18286a <=( a18285a  and  a18280a );
 a18290a <=( (not A200)  and  A166 );
 a18291a <=( A168  and  a18290a );
 a18295a <=( (not A234)  and  (not A233) );
 a18296a <=( (not A201)  and  a18295a );
 a18297a <=( a18296a  and  a18291a );
 a18301a <=( A298  and  A266 );
 a18302a <=( A265  and  a18301a );
 a18306a <=( A302  and  A300 );
 a18307a <=( (not A299)  and  a18306a );
 a18308a <=( a18307a  and  a18302a );
 a18312a <=( (not A200)  and  A166 );
 a18313a <=( A168  and  a18312a );
 a18317a <=( (not A234)  and  (not A233) );
 a18318a <=( (not A201)  and  a18317a );
 a18319a <=( a18318a  and  a18313a );
 a18323a <=( A298  and  (not A267) );
 a18324a <=( (not A266)  and  a18323a );
 a18328a <=( A301  and  A300 );
 a18329a <=( (not A299)  and  a18328a );
 a18330a <=( a18329a  and  a18324a );
 a18334a <=( (not A200)  and  A166 );
 a18335a <=( A168  and  a18334a );
 a18339a <=( (not A234)  and  (not A233) );
 a18340a <=( (not A201)  and  a18339a );
 a18341a <=( a18340a  and  a18335a );
 a18345a <=( A298  and  (not A267) );
 a18346a <=( (not A266)  and  a18345a );
 a18350a <=( A302  and  A300 );
 a18351a <=( (not A299)  and  a18350a );
 a18352a <=( a18351a  and  a18346a );
 a18356a <=( (not A200)  and  A166 );
 a18357a <=( A168  and  a18356a );
 a18361a <=( (not A234)  and  (not A233) );
 a18362a <=( (not A201)  and  a18361a );
 a18363a <=( a18362a  and  a18357a );
 a18367a <=( A298  and  (not A266) );
 a18368a <=( (not A265)  and  a18367a );
 a18372a <=( A301  and  A300 );
 a18373a <=( (not A299)  and  a18372a );
 a18374a <=( a18373a  and  a18368a );
 a18378a <=( (not A200)  and  A166 );
 a18379a <=( A168  and  a18378a );
 a18383a <=( (not A234)  and  (not A233) );
 a18384a <=( (not A201)  and  a18383a );
 a18385a <=( a18384a  and  a18379a );
 a18389a <=( A298  and  (not A266) );
 a18390a <=( (not A265)  and  a18389a );
 a18394a <=( A302  and  A300 );
 a18395a <=( (not A299)  and  a18394a );
 a18396a <=( a18395a  and  a18390a );
 a18400a <=( (not A200)  and  A166 );
 a18401a <=( A168  and  a18400a );
 a18405a <=( (not A233)  and  A232 );
 a18406a <=( (not A201)  and  a18405a );
 a18407a <=( a18406a  and  a18401a );
 a18411a <=( A265  and  A235 );
 a18412a <=( A234  and  a18411a );
 a18416a <=( A268  and  A267 );
 a18417a <=( (not A266)  and  a18416a );
 a18418a <=( a18417a  and  a18412a );
 a18422a <=( (not A200)  and  A166 );
 a18423a <=( A168  and  a18422a );
 a18427a <=( (not A233)  and  A232 );
 a18428a <=( (not A201)  and  a18427a );
 a18429a <=( a18428a  and  a18423a );
 a18433a <=( A265  and  A235 );
 a18434a <=( A234  and  a18433a );
 a18438a <=( A269  and  A267 );
 a18439a <=( (not A266)  and  a18438a );
 a18440a <=( a18439a  and  a18434a );
 a18444a <=( (not A200)  and  A166 );
 a18445a <=( A168  and  a18444a );
 a18449a <=( (not A233)  and  A232 );
 a18450a <=( (not A201)  and  a18449a );
 a18451a <=( a18450a  and  a18445a );
 a18455a <=( A265  and  A236 );
 a18456a <=( A234  and  a18455a );
 a18460a <=( A268  and  A267 );
 a18461a <=( (not A266)  and  a18460a );
 a18462a <=( a18461a  and  a18456a );
 a18466a <=( (not A200)  and  A166 );
 a18467a <=( A168  and  a18466a );
 a18471a <=( (not A233)  and  A232 );
 a18472a <=( (not A201)  and  a18471a );
 a18473a <=( a18472a  and  a18467a );
 a18477a <=( A265  and  A236 );
 a18478a <=( A234  and  a18477a );
 a18482a <=( A269  and  A267 );
 a18483a <=( (not A266)  and  a18482a );
 a18484a <=( a18483a  and  a18478a );
 a18488a <=( (not A200)  and  A166 );
 a18489a <=( A168  and  a18488a );
 a18493a <=( (not A233)  and  (not A232) );
 a18494a <=( (not A201)  and  a18493a );
 a18495a <=( a18494a  and  a18489a );
 a18499a <=( A298  and  A266 );
 a18500a <=( A265  and  a18499a );
 a18504a <=( A301  and  A300 );
 a18505a <=( (not A299)  and  a18504a );
 a18506a <=( a18505a  and  a18500a );
 a18510a <=( (not A200)  and  A166 );
 a18511a <=( A168  and  a18510a );
 a18515a <=( (not A233)  and  (not A232) );
 a18516a <=( (not A201)  and  a18515a );
 a18517a <=( a18516a  and  a18511a );
 a18521a <=( A298  and  A266 );
 a18522a <=( A265  and  a18521a );
 a18526a <=( A302  and  A300 );
 a18527a <=( (not A299)  and  a18526a );
 a18528a <=( a18527a  and  a18522a );
 a18532a <=( (not A200)  and  A166 );
 a18533a <=( A168  and  a18532a );
 a18537a <=( (not A233)  and  (not A232) );
 a18538a <=( (not A201)  and  a18537a );
 a18539a <=( a18538a  and  a18533a );
 a18543a <=( A298  and  (not A267) );
 a18544a <=( (not A266)  and  a18543a );
 a18548a <=( A301  and  A300 );
 a18549a <=( (not A299)  and  a18548a );
 a18550a <=( a18549a  and  a18544a );
 a18554a <=( (not A200)  and  A166 );
 a18555a <=( A168  and  a18554a );
 a18559a <=( (not A233)  and  (not A232) );
 a18560a <=( (not A201)  and  a18559a );
 a18561a <=( a18560a  and  a18555a );
 a18565a <=( A298  and  (not A267) );
 a18566a <=( (not A266)  and  a18565a );
 a18570a <=( A302  and  A300 );
 a18571a <=( (not A299)  and  a18570a );
 a18572a <=( a18571a  and  a18566a );
 a18576a <=( (not A200)  and  A166 );
 a18577a <=( A168  and  a18576a );
 a18581a <=( (not A233)  and  (not A232) );
 a18582a <=( (not A201)  and  a18581a );
 a18583a <=( a18582a  and  a18577a );
 a18587a <=( A298  and  (not A266) );
 a18588a <=( (not A265)  and  a18587a );
 a18592a <=( A301  and  A300 );
 a18593a <=( (not A299)  and  a18592a );
 a18594a <=( a18593a  and  a18588a );
 a18598a <=( (not A200)  and  A166 );
 a18599a <=( A168  and  a18598a );
 a18603a <=( (not A233)  and  (not A232) );
 a18604a <=( (not A201)  and  a18603a );
 a18605a <=( a18604a  and  a18599a );
 a18609a <=( A298  and  (not A266) );
 a18610a <=( (not A265)  and  a18609a );
 a18614a <=( A302  and  A300 );
 a18615a <=( (not A299)  and  a18614a );
 a18616a <=( a18615a  and  a18610a );
 a18620a <=( (not A199)  and  A166 );
 a18621a <=( A168  and  a18620a );
 a18625a <=( A233  and  A232 );
 a18626a <=( (not A200)  and  a18625a );
 a18627a <=( a18626a  and  a18621a );
 a18631a <=( A298  and  (not A267) );
 a18632a <=( A265  and  a18631a );
 a18636a <=( A301  and  A300 );
 a18637a <=( (not A299)  and  a18636a );
 a18638a <=( a18637a  and  a18632a );
 a18642a <=( (not A199)  and  A166 );
 a18643a <=( A168  and  a18642a );
 a18647a <=( A233  and  A232 );
 a18648a <=( (not A200)  and  a18647a );
 a18649a <=( a18648a  and  a18643a );
 a18653a <=( A298  and  (not A267) );
 a18654a <=( A265  and  a18653a );
 a18658a <=( A302  and  A300 );
 a18659a <=( (not A299)  and  a18658a );
 a18660a <=( a18659a  and  a18654a );
 a18664a <=( (not A199)  and  A166 );
 a18665a <=( A168  and  a18664a );
 a18669a <=( A233  and  A232 );
 a18670a <=( (not A200)  and  a18669a );
 a18671a <=( a18670a  and  a18665a );
 a18675a <=( A298  and  A266 );
 a18676a <=( A265  and  a18675a );
 a18680a <=( A301  and  A300 );
 a18681a <=( (not A299)  and  a18680a );
 a18682a <=( a18681a  and  a18676a );
 a18686a <=( (not A199)  and  A166 );
 a18687a <=( A168  and  a18686a );
 a18691a <=( A233  and  A232 );
 a18692a <=( (not A200)  and  a18691a );
 a18693a <=( a18692a  and  a18687a );
 a18697a <=( A298  and  A266 );
 a18698a <=( A265  and  a18697a );
 a18702a <=( A302  and  A300 );
 a18703a <=( (not A299)  and  a18702a );
 a18704a <=( a18703a  and  a18698a );
 a18708a <=( (not A199)  and  A166 );
 a18709a <=( A168  and  a18708a );
 a18713a <=( A233  and  A232 );
 a18714a <=( (not A200)  and  a18713a );
 a18715a <=( a18714a  and  a18709a );
 a18719a <=( A298  and  (not A266) );
 a18720a <=( (not A265)  and  a18719a );
 a18724a <=( A301  and  A300 );
 a18725a <=( (not A299)  and  a18724a );
 a18726a <=( a18725a  and  a18720a );
 a18730a <=( (not A199)  and  A166 );
 a18731a <=( A168  and  a18730a );
 a18735a <=( A233  and  A232 );
 a18736a <=( (not A200)  and  a18735a );
 a18737a <=( a18736a  and  a18731a );
 a18741a <=( A298  and  (not A266) );
 a18742a <=( (not A265)  and  a18741a );
 a18746a <=( A302  and  A300 );
 a18747a <=( (not A299)  and  a18746a );
 a18748a <=( a18747a  and  a18742a );
 a18752a <=( (not A199)  and  A166 );
 a18753a <=( A168  and  a18752a );
 a18757a <=( (not A235)  and  (not A233) );
 a18758a <=( (not A200)  and  a18757a );
 a18759a <=( a18758a  and  a18753a );
 a18763a <=( (not A268)  and  (not A266) );
 a18764a <=( (not A236)  and  a18763a );
 a18768a <=( A299  and  (not A298) );
 a18769a <=( (not A269)  and  a18768a );
 a18770a <=( a18769a  and  a18764a );
 a18774a <=( (not A199)  and  A166 );
 a18775a <=( A168  and  a18774a );
 a18779a <=( (not A234)  and  (not A233) );
 a18780a <=( (not A200)  and  a18779a );
 a18781a <=( a18780a  and  a18775a );
 a18785a <=( A298  and  A266 );
 a18786a <=( A265  and  a18785a );
 a18790a <=( A301  and  A300 );
 a18791a <=( (not A299)  and  a18790a );
 a18792a <=( a18791a  and  a18786a );
 a18796a <=( (not A199)  and  A166 );
 a18797a <=( A168  and  a18796a );
 a18801a <=( (not A234)  and  (not A233) );
 a18802a <=( (not A200)  and  a18801a );
 a18803a <=( a18802a  and  a18797a );
 a18807a <=( A298  and  A266 );
 a18808a <=( A265  and  a18807a );
 a18812a <=( A302  and  A300 );
 a18813a <=( (not A299)  and  a18812a );
 a18814a <=( a18813a  and  a18808a );
 a18818a <=( (not A199)  and  A166 );
 a18819a <=( A168  and  a18818a );
 a18823a <=( (not A234)  and  (not A233) );
 a18824a <=( (not A200)  and  a18823a );
 a18825a <=( a18824a  and  a18819a );
 a18829a <=( A298  and  (not A267) );
 a18830a <=( (not A266)  and  a18829a );
 a18834a <=( A301  and  A300 );
 a18835a <=( (not A299)  and  a18834a );
 a18836a <=( a18835a  and  a18830a );
 a18840a <=( (not A199)  and  A166 );
 a18841a <=( A168  and  a18840a );
 a18845a <=( (not A234)  and  (not A233) );
 a18846a <=( (not A200)  and  a18845a );
 a18847a <=( a18846a  and  a18841a );
 a18851a <=( A298  and  (not A267) );
 a18852a <=( (not A266)  and  a18851a );
 a18856a <=( A302  and  A300 );
 a18857a <=( (not A299)  and  a18856a );
 a18858a <=( a18857a  and  a18852a );
 a18862a <=( (not A199)  and  A166 );
 a18863a <=( A168  and  a18862a );
 a18867a <=( (not A234)  and  (not A233) );
 a18868a <=( (not A200)  and  a18867a );
 a18869a <=( a18868a  and  a18863a );
 a18873a <=( A298  and  (not A266) );
 a18874a <=( (not A265)  and  a18873a );
 a18878a <=( A301  and  A300 );
 a18879a <=( (not A299)  and  a18878a );
 a18880a <=( a18879a  and  a18874a );
 a18884a <=( (not A199)  and  A166 );
 a18885a <=( A168  and  a18884a );
 a18889a <=( (not A234)  and  (not A233) );
 a18890a <=( (not A200)  and  a18889a );
 a18891a <=( a18890a  and  a18885a );
 a18895a <=( A298  and  (not A266) );
 a18896a <=( (not A265)  and  a18895a );
 a18900a <=( A302  and  A300 );
 a18901a <=( (not A299)  and  a18900a );
 a18902a <=( a18901a  and  a18896a );
 a18906a <=( (not A199)  and  A166 );
 a18907a <=( A168  and  a18906a );
 a18911a <=( (not A233)  and  A232 );
 a18912a <=( (not A200)  and  a18911a );
 a18913a <=( a18912a  and  a18907a );
 a18917a <=( A265  and  A235 );
 a18918a <=( A234  and  a18917a );
 a18922a <=( A268  and  A267 );
 a18923a <=( (not A266)  and  a18922a );
 a18924a <=( a18923a  and  a18918a );
 a18928a <=( (not A199)  and  A166 );
 a18929a <=( A168  and  a18928a );
 a18933a <=( (not A233)  and  A232 );
 a18934a <=( (not A200)  and  a18933a );
 a18935a <=( a18934a  and  a18929a );
 a18939a <=( A265  and  A235 );
 a18940a <=( A234  and  a18939a );
 a18944a <=( A269  and  A267 );
 a18945a <=( (not A266)  and  a18944a );
 a18946a <=( a18945a  and  a18940a );
 a18950a <=( (not A199)  and  A166 );
 a18951a <=( A168  and  a18950a );
 a18955a <=( (not A233)  and  A232 );
 a18956a <=( (not A200)  and  a18955a );
 a18957a <=( a18956a  and  a18951a );
 a18961a <=( A265  and  A236 );
 a18962a <=( A234  and  a18961a );
 a18966a <=( A268  and  A267 );
 a18967a <=( (not A266)  and  a18966a );
 a18968a <=( a18967a  and  a18962a );
 a18972a <=( (not A199)  and  A166 );
 a18973a <=( A168  and  a18972a );
 a18977a <=( (not A233)  and  A232 );
 a18978a <=( (not A200)  and  a18977a );
 a18979a <=( a18978a  and  a18973a );
 a18983a <=( A265  and  A236 );
 a18984a <=( A234  and  a18983a );
 a18988a <=( A269  and  A267 );
 a18989a <=( (not A266)  and  a18988a );
 a18990a <=( a18989a  and  a18984a );
 a18994a <=( (not A199)  and  A166 );
 a18995a <=( A168  and  a18994a );
 a18999a <=( (not A233)  and  (not A232) );
 a19000a <=( (not A200)  and  a18999a );
 a19001a <=( a19000a  and  a18995a );
 a19005a <=( A298  and  A266 );
 a19006a <=( A265  and  a19005a );
 a19010a <=( A301  and  A300 );
 a19011a <=( (not A299)  and  a19010a );
 a19012a <=( a19011a  and  a19006a );
 a19016a <=( (not A199)  and  A166 );
 a19017a <=( A168  and  a19016a );
 a19021a <=( (not A233)  and  (not A232) );
 a19022a <=( (not A200)  and  a19021a );
 a19023a <=( a19022a  and  a19017a );
 a19027a <=( A298  and  A266 );
 a19028a <=( A265  and  a19027a );
 a19032a <=( A302  and  A300 );
 a19033a <=( (not A299)  and  a19032a );
 a19034a <=( a19033a  and  a19028a );
 a19038a <=( (not A199)  and  A166 );
 a19039a <=( A168  and  a19038a );
 a19043a <=( (not A233)  and  (not A232) );
 a19044a <=( (not A200)  and  a19043a );
 a19045a <=( a19044a  and  a19039a );
 a19049a <=( A298  and  (not A267) );
 a19050a <=( (not A266)  and  a19049a );
 a19054a <=( A301  and  A300 );
 a19055a <=( (not A299)  and  a19054a );
 a19056a <=( a19055a  and  a19050a );
 a19060a <=( (not A199)  and  A166 );
 a19061a <=( A168  and  a19060a );
 a19065a <=( (not A233)  and  (not A232) );
 a19066a <=( (not A200)  and  a19065a );
 a19067a <=( a19066a  and  a19061a );
 a19071a <=( A298  and  (not A267) );
 a19072a <=( (not A266)  and  a19071a );
 a19076a <=( A302  and  A300 );
 a19077a <=( (not A299)  and  a19076a );
 a19078a <=( a19077a  and  a19072a );
 a19082a <=( (not A199)  and  A166 );
 a19083a <=( A168  and  a19082a );
 a19087a <=( (not A233)  and  (not A232) );
 a19088a <=( (not A200)  and  a19087a );
 a19089a <=( a19088a  and  a19083a );
 a19093a <=( A298  and  (not A266) );
 a19094a <=( (not A265)  and  a19093a );
 a19098a <=( A301  and  A300 );
 a19099a <=( (not A299)  and  a19098a );
 a19100a <=( a19099a  and  a19094a );
 a19104a <=( (not A199)  and  A166 );
 a19105a <=( A168  and  a19104a );
 a19109a <=( (not A233)  and  (not A232) );
 a19110a <=( (not A200)  and  a19109a );
 a19111a <=( a19110a  and  a19105a );
 a19115a <=( A298  and  (not A266) );
 a19116a <=( (not A265)  and  a19115a );
 a19120a <=( A302  and  A300 );
 a19121a <=( (not A299)  and  a19120a );
 a19122a <=( a19121a  and  a19116a );
 a19126a <=( A199  and  A167 );
 a19127a <=( A168  and  a19126a );
 a19131a <=( A233  and  A232 );
 a19132a <=( A200  and  a19131a );
 a19133a <=( a19132a  and  a19127a );
 a19137a <=( A298  and  (not A267) );
 a19138a <=( A265  and  a19137a );
 a19142a <=( A301  and  A300 );
 a19143a <=( (not A299)  and  a19142a );
 a19144a <=( a19143a  and  a19138a );
 a19148a <=( A199  and  A167 );
 a19149a <=( A168  and  a19148a );
 a19153a <=( A233  and  A232 );
 a19154a <=( A200  and  a19153a );
 a19155a <=( a19154a  and  a19149a );
 a19159a <=( A298  and  (not A267) );
 a19160a <=( A265  and  a19159a );
 a19164a <=( A302  and  A300 );
 a19165a <=( (not A299)  and  a19164a );
 a19166a <=( a19165a  and  a19160a );
 a19170a <=( A199  and  A167 );
 a19171a <=( A168  and  a19170a );
 a19175a <=( A233  and  A232 );
 a19176a <=( A200  and  a19175a );
 a19177a <=( a19176a  and  a19171a );
 a19181a <=( A298  and  A266 );
 a19182a <=( A265  and  a19181a );
 a19186a <=( A301  and  A300 );
 a19187a <=( (not A299)  and  a19186a );
 a19188a <=( a19187a  and  a19182a );
 a19192a <=( A199  and  A167 );
 a19193a <=( A168  and  a19192a );
 a19197a <=( A233  and  A232 );
 a19198a <=( A200  and  a19197a );
 a19199a <=( a19198a  and  a19193a );
 a19203a <=( A298  and  A266 );
 a19204a <=( A265  and  a19203a );
 a19208a <=( A302  and  A300 );
 a19209a <=( (not A299)  and  a19208a );
 a19210a <=( a19209a  and  a19204a );
 a19214a <=( A199  and  A167 );
 a19215a <=( A168  and  a19214a );
 a19219a <=( A233  and  A232 );
 a19220a <=( A200  and  a19219a );
 a19221a <=( a19220a  and  a19215a );
 a19225a <=( A298  and  (not A266) );
 a19226a <=( (not A265)  and  a19225a );
 a19230a <=( A301  and  A300 );
 a19231a <=( (not A299)  and  a19230a );
 a19232a <=( a19231a  and  a19226a );
 a19236a <=( A199  and  A167 );
 a19237a <=( A168  and  a19236a );
 a19241a <=( A233  and  A232 );
 a19242a <=( A200  and  a19241a );
 a19243a <=( a19242a  and  a19237a );
 a19247a <=( A298  and  (not A266) );
 a19248a <=( (not A265)  and  a19247a );
 a19252a <=( A302  and  A300 );
 a19253a <=( (not A299)  and  a19252a );
 a19254a <=( a19253a  and  a19248a );
 a19258a <=( A199  and  A167 );
 a19259a <=( A168  and  a19258a );
 a19263a <=( (not A235)  and  (not A233) );
 a19264a <=( A200  and  a19263a );
 a19265a <=( a19264a  and  a19259a );
 a19269a <=( (not A268)  and  (not A266) );
 a19270a <=( (not A236)  and  a19269a );
 a19274a <=( A299  and  (not A298) );
 a19275a <=( (not A269)  and  a19274a );
 a19276a <=( a19275a  and  a19270a );
 a19280a <=( A199  and  A167 );
 a19281a <=( A168  and  a19280a );
 a19285a <=( (not A234)  and  (not A233) );
 a19286a <=( A200  and  a19285a );
 a19287a <=( a19286a  and  a19281a );
 a19291a <=( A298  and  A266 );
 a19292a <=( A265  and  a19291a );
 a19296a <=( A301  and  A300 );
 a19297a <=( (not A299)  and  a19296a );
 a19298a <=( a19297a  and  a19292a );
 a19302a <=( A199  and  A167 );
 a19303a <=( A168  and  a19302a );
 a19307a <=( (not A234)  and  (not A233) );
 a19308a <=( A200  and  a19307a );
 a19309a <=( a19308a  and  a19303a );
 a19313a <=( A298  and  A266 );
 a19314a <=( A265  and  a19313a );
 a19318a <=( A302  and  A300 );
 a19319a <=( (not A299)  and  a19318a );
 a19320a <=( a19319a  and  a19314a );
 a19324a <=( A199  and  A167 );
 a19325a <=( A168  and  a19324a );
 a19329a <=( (not A234)  and  (not A233) );
 a19330a <=( A200  and  a19329a );
 a19331a <=( a19330a  and  a19325a );
 a19335a <=( A298  and  (not A267) );
 a19336a <=( (not A266)  and  a19335a );
 a19340a <=( A301  and  A300 );
 a19341a <=( (not A299)  and  a19340a );
 a19342a <=( a19341a  and  a19336a );
 a19346a <=( A199  and  A167 );
 a19347a <=( A168  and  a19346a );
 a19351a <=( (not A234)  and  (not A233) );
 a19352a <=( A200  and  a19351a );
 a19353a <=( a19352a  and  a19347a );
 a19357a <=( A298  and  (not A267) );
 a19358a <=( (not A266)  and  a19357a );
 a19362a <=( A302  and  A300 );
 a19363a <=( (not A299)  and  a19362a );
 a19364a <=( a19363a  and  a19358a );
 a19368a <=( A199  and  A167 );
 a19369a <=( A168  and  a19368a );
 a19373a <=( (not A234)  and  (not A233) );
 a19374a <=( A200  and  a19373a );
 a19375a <=( a19374a  and  a19369a );
 a19379a <=( A298  and  (not A266) );
 a19380a <=( (not A265)  and  a19379a );
 a19384a <=( A301  and  A300 );
 a19385a <=( (not A299)  and  a19384a );
 a19386a <=( a19385a  and  a19380a );
 a19390a <=( A199  and  A167 );
 a19391a <=( A168  and  a19390a );
 a19395a <=( (not A234)  and  (not A233) );
 a19396a <=( A200  and  a19395a );
 a19397a <=( a19396a  and  a19391a );
 a19401a <=( A298  and  (not A266) );
 a19402a <=( (not A265)  and  a19401a );
 a19406a <=( A302  and  A300 );
 a19407a <=( (not A299)  and  a19406a );
 a19408a <=( a19407a  and  a19402a );
 a19412a <=( A199  and  A167 );
 a19413a <=( A168  and  a19412a );
 a19417a <=( (not A233)  and  A232 );
 a19418a <=( A200  and  a19417a );
 a19419a <=( a19418a  and  a19413a );
 a19423a <=( A265  and  A235 );
 a19424a <=( A234  and  a19423a );
 a19428a <=( A268  and  A267 );
 a19429a <=( (not A266)  and  a19428a );
 a19430a <=( a19429a  and  a19424a );
 a19434a <=( A199  and  A167 );
 a19435a <=( A168  and  a19434a );
 a19439a <=( (not A233)  and  A232 );
 a19440a <=( A200  and  a19439a );
 a19441a <=( a19440a  and  a19435a );
 a19445a <=( A265  and  A235 );
 a19446a <=( A234  and  a19445a );
 a19450a <=( A269  and  A267 );
 a19451a <=( (not A266)  and  a19450a );
 a19452a <=( a19451a  and  a19446a );
 a19456a <=( A199  and  A167 );
 a19457a <=( A168  and  a19456a );
 a19461a <=( (not A233)  and  A232 );
 a19462a <=( A200  and  a19461a );
 a19463a <=( a19462a  and  a19457a );
 a19467a <=( A265  and  A236 );
 a19468a <=( A234  and  a19467a );
 a19472a <=( A268  and  A267 );
 a19473a <=( (not A266)  and  a19472a );
 a19474a <=( a19473a  and  a19468a );
 a19478a <=( A199  and  A167 );
 a19479a <=( A168  and  a19478a );
 a19483a <=( (not A233)  and  A232 );
 a19484a <=( A200  and  a19483a );
 a19485a <=( a19484a  and  a19479a );
 a19489a <=( A265  and  A236 );
 a19490a <=( A234  and  a19489a );
 a19494a <=( A269  and  A267 );
 a19495a <=( (not A266)  and  a19494a );
 a19496a <=( a19495a  and  a19490a );
 a19500a <=( A199  and  A167 );
 a19501a <=( A168  and  a19500a );
 a19505a <=( (not A233)  and  (not A232) );
 a19506a <=( A200  and  a19505a );
 a19507a <=( a19506a  and  a19501a );
 a19511a <=( A298  and  A266 );
 a19512a <=( A265  and  a19511a );
 a19516a <=( A301  and  A300 );
 a19517a <=( (not A299)  and  a19516a );
 a19518a <=( a19517a  and  a19512a );
 a19522a <=( A199  and  A167 );
 a19523a <=( A168  and  a19522a );
 a19527a <=( (not A233)  and  (not A232) );
 a19528a <=( A200  and  a19527a );
 a19529a <=( a19528a  and  a19523a );
 a19533a <=( A298  and  A266 );
 a19534a <=( A265  and  a19533a );
 a19538a <=( A302  and  A300 );
 a19539a <=( (not A299)  and  a19538a );
 a19540a <=( a19539a  and  a19534a );
 a19544a <=( A199  and  A167 );
 a19545a <=( A168  and  a19544a );
 a19549a <=( (not A233)  and  (not A232) );
 a19550a <=( A200  and  a19549a );
 a19551a <=( a19550a  and  a19545a );
 a19555a <=( A298  and  (not A267) );
 a19556a <=( (not A266)  and  a19555a );
 a19560a <=( A301  and  A300 );
 a19561a <=( (not A299)  and  a19560a );
 a19562a <=( a19561a  and  a19556a );
 a19566a <=( A199  and  A167 );
 a19567a <=( A168  and  a19566a );
 a19571a <=( (not A233)  and  (not A232) );
 a19572a <=( A200  and  a19571a );
 a19573a <=( a19572a  and  a19567a );
 a19577a <=( A298  and  (not A267) );
 a19578a <=( (not A266)  and  a19577a );
 a19582a <=( A302  and  A300 );
 a19583a <=( (not A299)  and  a19582a );
 a19584a <=( a19583a  and  a19578a );
 a19588a <=( A199  and  A167 );
 a19589a <=( A168  and  a19588a );
 a19593a <=( (not A233)  and  (not A232) );
 a19594a <=( A200  and  a19593a );
 a19595a <=( a19594a  and  a19589a );
 a19599a <=( A298  and  (not A266) );
 a19600a <=( (not A265)  and  a19599a );
 a19604a <=( A301  and  A300 );
 a19605a <=( (not A299)  and  a19604a );
 a19606a <=( a19605a  and  a19600a );
 a19610a <=( A199  and  A167 );
 a19611a <=( A168  and  a19610a );
 a19615a <=( (not A233)  and  (not A232) );
 a19616a <=( A200  and  a19615a );
 a19617a <=( a19616a  and  a19611a );
 a19621a <=( A298  and  (not A266) );
 a19622a <=( (not A265)  and  a19621a );
 a19626a <=( A302  and  A300 );
 a19627a <=( (not A299)  and  a19626a );
 a19628a <=( a19627a  and  a19622a );
 a19632a <=( (not A200)  and  A167 );
 a19633a <=( A168  and  a19632a );
 a19637a <=( A232  and  (not A203) );
 a19638a <=( (not A202)  and  a19637a );
 a19639a <=( a19638a  and  a19633a );
 a19643a <=( (not A268)  and  A265 );
 a19644a <=( A233  and  a19643a );
 a19648a <=( A299  and  (not A298) );
 a19649a <=( (not A269)  and  a19648a );
 a19650a <=( a19649a  and  a19644a );
 a19654a <=( (not A200)  and  A167 );
 a19655a <=( A168  and  a19654a );
 a19659a <=( (not A233)  and  (not A203) );
 a19660a <=( (not A202)  and  a19659a );
 a19661a <=( a19660a  and  a19655a );
 a19665a <=( A265  and  (not A236) );
 a19666a <=( (not A235)  and  a19665a );
 a19670a <=( A299  and  (not A298) );
 a19671a <=( A266  and  a19670a );
 a19672a <=( a19671a  and  a19666a );
 a19676a <=( (not A200)  and  A167 );
 a19677a <=( A168  and  a19676a );
 a19681a <=( (not A233)  and  (not A203) );
 a19682a <=( (not A202)  and  a19681a );
 a19683a <=( a19682a  and  a19677a );
 a19687a <=( (not A266)  and  (not A236) );
 a19688a <=( (not A235)  and  a19687a );
 a19692a <=( A299  and  (not A298) );
 a19693a <=( (not A267)  and  a19692a );
 a19694a <=( a19693a  and  a19688a );
 a19698a <=( (not A200)  and  A167 );
 a19699a <=( A168  and  a19698a );
 a19703a <=( (not A233)  and  (not A203) );
 a19704a <=( (not A202)  and  a19703a );
 a19705a <=( a19704a  and  a19699a );
 a19709a <=( (not A265)  and  (not A236) );
 a19710a <=( (not A235)  and  a19709a );
 a19714a <=( A299  and  (not A298) );
 a19715a <=( (not A266)  and  a19714a );
 a19716a <=( a19715a  and  a19710a );
 a19720a <=( (not A200)  and  A167 );
 a19721a <=( A168  and  a19720a );
 a19725a <=( (not A233)  and  (not A203) );
 a19726a <=( (not A202)  and  a19725a );
 a19727a <=( a19726a  and  a19721a );
 a19731a <=( (not A268)  and  (not A266) );
 a19732a <=( (not A234)  and  a19731a );
 a19736a <=( A299  and  (not A298) );
 a19737a <=( (not A269)  and  a19736a );
 a19738a <=( a19737a  and  a19732a );
 a19742a <=( (not A200)  and  A167 );
 a19743a <=( A168  and  a19742a );
 a19747a <=( A232  and  (not A203) );
 a19748a <=( (not A202)  and  a19747a );
 a19749a <=( a19748a  and  a19743a );
 a19753a <=( A235  and  A234 );
 a19754a <=( (not A233)  and  a19753a );
 a19758a <=( (not A302)  and  (not A301) );
 a19759a <=( A298  and  a19758a );
 a19760a <=( a19759a  and  a19754a );
 a19764a <=( (not A200)  and  A167 );
 a19765a <=( A168  and  a19764a );
 a19769a <=( A232  and  (not A203) );
 a19770a <=( (not A202)  and  a19769a );
 a19771a <=( a19770a  and  a19765a );
 a19775a <=( A236  and  A234 );
 a19776a <=( (not A233)  and  a19775a );
 a19780a <=( (not A302)  and  (not A301) );
 a19781a <=( A298  and  a19780a );
 a19782a <=( a19781a  and  a19776a );
 a19786a <=( (not A200)  and  A167 );
 a19787a <=( A168  and  a19786a );
 a19791a <=( (not A232)  and  (not A203) );
 a19792a <=( (not A202)  and  a19791a );
 a19793a <=( a19792a  and  a19787a );
 a19797a <=( (not A268)  and  (not A266) );
 a19798a <=( (not A233)  and  a19797a );
 a19802a <=( A299  and  (not A298) );
 a19803a <=( (not A269)  and  a19802a );
 a19804a <=( a19803a  and  a19798a );
 a19808a <=( (not A200)  and  A167 );
 a19809a <=( A168  and  a19808a );
 a19813a <=( A233  and  A232 );
 a19814a <=( (not A201)  and  a19813a );
 a19815a <=( a19814a  and  a19809a );
 a19819a <=( A298  and  (not A267) );
 a19820a <=( A265  and  a19819a );
 a19824a <=( A301  and  A300 );
 a19825a <=( (not A299)  and  a19824a );
 a19826a <=( a19825a  and  a19820a );
 a19830a <=( (not A200)  and  A167 );
 a19831a <=( A168  and  a19830a );
 a19835a <=( A233  and  A232 );
 a19836a <=( (not A201)  and  a19835a );
 a19837a <=( a19836a  and  a19831a );
 a19841a <=( A298  and  (not A267) );
 a19842a <=( A265  and  a19841a );
 a19846a <=( A302  and  A300 );
 a19847a <=( (not A299)  and  a19846a );
 a19848a <=( a19847a  and  a19842a );
 a19852a <=( (not A200)  and  A167 );
 a19853a <=( A168  and  a19852a );
 a19857a <=( A233  and  A232 );
 a19858a <=( (not A201)  and  a19857a );
 a19859a <=( a19858a  and  a19853a );
 a19863a <=( A298  and  A266 );
 a19864a <=( A265  and  a19863a );
 a19868a <=( A301  and  A300 );
 a19869a <=( (not A299)  and  a19868a );
 a19870a <=( a19869a  and  a19864a );
 a19874a <=( (not A200)  and  A167 );
 a19875a <=( A168  and  a19874a );
 a19879a <=( A233  and  A232 );
 a19880a <=( (not A201)  and  a19879a );
 a19881a <=( a19880a  and  a19875a );
 a19885a <=( A298  and  A266 );
 a19886a <=( A265  and  a19885a );
 a19890a <=( A302  and  A300 );
 a19891a <=( (not A299)  and  a19890a );
 a19892a <=( a19891a  and  a19886a );
 a19896a <=( (not A200)  and  A167 );
 a19897a <=( A168  and  a19896a );
 a19901a <=( A233  and  A232 );
 a19902a <=( (not A201)  and  a19901a );
 a19903a <=( a19902a  and  a19897a );
 a19907a <=( A298  and  (not A266) );
 a19908a <=( (not A265)  and  a19907a );
 a19912a <=( A301  and  A300 );
 a19913a <=( (not A299)  and  a19912a );
 a19914a <=( a19913a  and  a19908a );
 a19918a <=( (not A200)  and  A167 );
 a19919a <=( A168  and  a19918a );
 a19923a <=( A233  and  A232 );
 a19924a <=( (not A201)  and  a19923a );
 a19925a <=( a19924a  and  a19919a );
 a19929a <=( A298  and  (not A266) );
 a19930a <=( (not A265)  and  a19929a );
 a19934a <=( A302  and  A300 );
 a19935a <=( (not A299)  and  a19934a );
 a19936a <=( a19935a  and  a19930a );
 a19940a <=( (not A200)  and  A167 );
 a19941a <=( A168  and  a19940a );
 a19945a <=( (not A235)  and  (not A233) );
 a19946a <=( (not A201)  and  a19945a );
 a19947a <=( a19946a  and  a19941a );
 a19951a <=( (not A268)  and  (not A266) );
 a19952a <=( (not A236)  and  a19951a );
 a19956a <=( A299  and  (not A298) );
 a19957a <=( (not A269)  and  a19956a );
 a19958a <=( a19957a  and  a19952a );
 a19962a <=( (not A200)  and  A167 );
 a19963a <=( A168  and  a19962a );
 a19967a <=( (not A234)  and  (not A233) );
 a19968a <=( (not A201)  and  a19967a );
 a19969a <=( a19968a  and  a19963a );
 a19973a <=( A298  and  A266 );
 a19974a <=( A265  and  a19973a );
 a19978a <=( A301  and  A300 );
 a19979a <=( (not A299)  and  a19978a );
 a19980a <=( a19979a  and  a19974a );
 a19984a <=( (not A200)  and  A167 );
 a19985a <=( A168  and  a19984a );
 a19989a <=( (not A234)  and  (not A233) );
 a19990a <=( (not A201)  and  a19989a );
 a19991a <=( a19990a  and  a19985a );
 a19995a <=( A298  and  A266 );
 a19996a <=( A265  and  a19995a );
 a20000a <=( A302  and  A300 );
 a20001a <=( (not A299)  and  a20000a );
 a20002a <=( a20001a  and  a19996a );
 a20006a <=( (not A200)  and  A167 );
 a20007a <=( A168  and  a20006a );
 a20011a <=( (not A234)  and  (not A233) );
 a20012a <=( (not A201)  and  a20011a );
 a20013a <=( a20012a  and  a20007a );
 a20017a <=( A298  and  (not A267) );
 a20018a <=( (not A266)  and  a20017a );
 a20022a <=( A301  and  A300 );
 a20023a <=( (not A299)  and  a20022a );
 a20024a <=( a20023a  and  a20018a );
 a20028a <=( (not A200)  and  A167 );
 a20029a <=( A168  and  a20028a );
 a20033a <=( (not A234)  and  (not A233) );
 a20034a <=( (not A201)  and  a20033a );
 a20035a <=( a20034a  and  a20029a );
 a20039a <=( A298  and  (not A267) );
 a20040a <=( (not A266)  and  a20039a );
 a20044a <=( A302  and  A300 );
 a20045a <=( (not A299)  and  a20044a );
 a20046a <=( a20045a  and  a20040a );
 a20050a <=( (not A200)  and  A167 );
 a20051a <=( A168  and  a20050a );
 a20055a <=( (not A234)  and  (not A233) );
 a20056a <=( (not A201)  and  a20055a );
 a20057a <=( a20056a  and  a20051a );
 a20061a <=( A298  and  (not A266) );
 a20062a <=( (not A265)  and  a20061a );
 a20066a <=( A301  and  A300 );
 a20067a <=( (not A299)  and  a20066a );
 a20068a <=( a20067a  and  a20062a );
 a20072a <=( (not A200)  and  A167 );
 a20073a <=( A168  and  a20072a );
 a20077a <=( (not A234)  and  (not A233) );
 a20078a <=( (not A201)  and  a20077a );
 a20079a <=( a20078a  and  a20073a );
 a20083a <=( A298  and  (not A266) );
 a20084a <=( (not A265)  and  a20083a );
 a20088a <=( A302  and  A300 );
 a20089a <=( (not A299)  and  a20088a );
 a20090a <=( a20089a  and  a20084a );
 a20094a <=( (not A200)  and  A167 );
 a20095a <=( A168  and  a20094a );
 a20099a <=( (not A233)  and  A232 );
 a20100a <=( (not A201)  and  a20099a );
 a20101a <=( a20100a  and  a20095a );
 a20105a <=( A265  and  A235 );
 a20106a <=( A234  and  a20105a );
 a20110a <=( A268  and  A267 );
 a20111a <=( (not A266)  and  a20110a );
 a20112a <=( a20111a  and  a20106a );
 a20116a <=( (not A200)  and  A167 );
 a20117a <=( A168  and  a20116a );
 a20121a <=( (not A233)  and  A232 );
 a20122a <=( (not A201)  and  a20121a );
 a20123a <=( a20122a  and  a20117a );
 a20127a <=( A265  and  A235 );
 a20128a <=( A234  and  a20127a );
 a20132a <=( A269  and  A267 );
 a20133a <=( (not A266)  and  a20132a );
 a20134a <=( a20133a  and  a20128a );
 a20138a <=( (not A200)  and  A167 );
 a20139a <=( A168  and  a20138a );
 a20143a <=( (not A233)  and  A232 );
 a20144a <=( (not A201)  and  a20143a );
 a20145a <=( a20144a  and  a20139a );
 a20149a <=( A265  and  A236 );
 a20150a <=( A234  and  a20149a );
 a20154a <=( A268  and  A267 );
 a20155a <=( (not A266)  and  a20154a );
 a20156a <=( a20155a  and  a20150a );
 a20160a <=( (not A200)  and  A167 );
 a20161a <=( A168  and  a20160a );
 a20165a <=( (not A233)  and  A232 );
 a20166a <=( (not A201)  and  a20165a );
 a20167a <=( a20166a  and  a20161a );
 a20171a <=( A265  and  A236 );
 a20172a <=( A234  and  a20171a );
 a20176a <=( A269  and  A267 );
 a20177a <=( (not A266)  and  a20176a );
 a20178a <=( a20177a  and  a20172a );
 a20182a <=( (not A200)  and  A167 );
 a20183a <=( A168  and  a20182a );
 a20187a <=( (not A233)  and  (not A232) );
 a20188a <=( (not A201)  and  a20187a );
 a20189a <=( a20188a  and  a20183a );
 a20193a <=( A298  and  A266 );
 a20194a <=( A265  and  a20193a );
 a20198a <=( A301  and  A300 );
 a20199a <=( (not A299)  and  a20198a );
 a20200a <=( a20199a  and  a20194a );
 a20204a <=( (not A200)  and  A167 );
 a20205a <=( A168  and  a20204a );
 a20209a <=( (not A233)  and  (not A232) );
 a20210a <=( (not A201)  and  a20209a );
 a20211a <=( a20210a  and  a20205a );
 a20215a <=( A298  and  A266 );
 a20216a <=( A265  and  a20215a );
 a20220a <=( A302  and  A300 );
 a20221a <=( (not A299)  and  a20220a );
 a20222a <=( a20221a  and  a20216a );
 a20226a <=( (not A200)  and  A167 );
 a20227a <=( A168  and  a20226a );
 a20231a <=( (not A233)  and  (not A232) );
 a20232a <=( (not A201)  and  a20231a );
 a20233a <=( a20232a  and  a20227a );
 a20237a <=( A298  and  (not A267) );
 a20238a <=( (not A266)  and  a20237a );
 a20242a <=( A301  and  A300 );
 a20243a <=( (not A299)  and  a20242a );
 a20244a <=( a20243a  and  a20238a );
 a20248a <=( (not A200)  and  A167 );
 a20249a <=( A168  and  a20248a );
 a20253a <=( (not A233)  and  (not A232) );
 a20254a <=( (not A201)  and  a20253a );
 a20255a <=( a20254a  and  a20249a );
 a20259a <=( A298  and  (not A267) );
 a20260a <=( (not A266)  and  a20259a );
 a20264a <=( A302  and  A300 );
 a20265a <=( (not A299)  and  a20264a );
 a20266a <=( a20265a  and  a20260a );
 a20270a <=( (not A200)  and  A167 );
 a20271a <=( A168  and  a20270a );
 a20275a <=( (not A233)  and  (not A232) );
 a20276a <=( (not A201)  and  a20275a );
 a20277a <=( a20276a  and  a20271a );
 a20281a <=( A298  and  (not A266) );
 a20282a <=( (not A265)  and  a20281a );
 a20286a <=( A301  and  A300 );
 a20287a <=( (not A299)  and  a20286a );
 a20288a <=( a20287a  and  a20282a );
 a20292a <=( (not A200)  and  A167 );
 a20293a <=( A168  and  a20292a );
 a20297a <=( (not A233)  and  (not A232) );
 a20298a <=( (not A201)  and  a20297a );
 a20299a <=( a20298a  and  a20293a );
 a20303a <=( A298  and  (not A266) );
 a20304a <=( (not A265)  and  a20303a );
 a20308a <=( A302  and  A300 );
 a20309a <=( (not A299)  and  a20308a );
 a20310a <=( a20309a  and  a20304a );
 a20314a <=( (not A199)  and  A167 );
 a20315a <=( A168  and  a20314a );
 a20319a <=( A233  and  A232 );
 a20320a <=( (not A200)  and  a20319a );
 a20321a <=( a20320a  and  a20315a );
 a20325a <=( A298  and  (not A267) );
 a20326a <=( A265  and  a20325a );
 a20330a <=( A301  and  A300 );
 a20331a <=( (not A299)  and  a20330a );
 a20332a <=( a20331a  and  a20326a );
 a20336a <=( (not A199)  and  A167 );
 a20337a <=( A168  and  a20336a );
 a20341a <=( A233  and  A232 );
 a20342a <=( (not A200)  and  a20341a );
 a20343a <=( a20342a  and  a20337a );
 a20347a <=( A298  and  (not A267) );
 a20348a <=( A265  and  a20347a );
 a20352a <=( A302  and  A300 );
 a20353a <=( (not A299)  and  a20352a );
 a20354a <=( a20353a  and  a20348a );
 a20358a <=( (not A199)  and  A167 );
 a20359a <=( A168  and  a20358a );
 a20363a <=( A233  and  A232 );
 a20364a <=( (not A200)  and  a20363a );
 a20365a <=( a20364a  and  a20359a );
 a20369a <=( A298  and  A266 );
 a20370a <=( A265  and  a20369a );
 a20374a <=( A301  and  A300 );
 a20375a <=( (not A299)  and  a20374a );
 a20376a <=( a20375a  and  a20370a );
 a20380a <=( (not A199)  and  A167 );
 a20381a <=( A168  and  a20380a );
 a20385a <=( A233  and  A232 );
 a20386a <=( (not A200)  and  a20385a );
 a20387a <=( a20386a  and  a20381a );
 a20391a <=( A298  and  A266 );
 a20392a <=( A265  and  a20391a );
 a20396a <=( A302  and  A300 );
 a20397a <=( (not A299)  and  a20396a );
 a20398a <=( a20397a  and  a20392a );
 a20402a <=( (not A199)  and  A167 );
 a20403a <=( A168  and  a20402a );
 a20407a <=( A233  and  A232 );
 a20408a <=( (not A200)  and  a20407a );
 a20409a <=( a20408a  and  a20403a );
 a20413a <=( A298  and  (not A266) );
 a20414a <=( (not A265)  and  a20413a );
 a20418a <=( A301  and  A300 );
 a20419a <=( (not A299)  and  a20418a );
 a20420a <=( a20419a  and  a20414a );
 a20424a <=( (not A199)  and  A167 );
 a20425a <=( A168  and  a20424a );
 a20429a <=( A233  and  A232 );
 a20430a <=( (not A200)  and  a20429a );
 a20431a <=( a20430a  and  a20425a );
 a20435a <=( A298  and  (not A266) );
 a20436a <=( (not A265)  and  a20435a );
 a20440a <=( A302  and  A300 );
 a20441a <=( (not A299)  and  a20440a );
 a20442a <=( a20441a  and  a20436a );
 a20446a <=( (not A199)  and  A167 );
 a20447a <=( A168  and  a20446a );
 a20451a <=( (not A235)  and  (not A233) );
 a20452a <=( (not A200)  and  a20451a );
 a20453a <=( a20452a  and  a20447a );
 a20457a <=( (not A268)  and  (not A266) );
 a20458a <=( (not A236)  and  a20457a );
 a20462a <=( A299  and  (not A298) );
 a20463a <=( (not A269)  and  a20462a );
 a20464a <=( a20463a  and  a20458a );
 a20468a <=( (not A199)  and  A167 );
 a20469a <=( A168  and  a20468a );
 a20473a <=( (not A234)  and  (not A233) );
 a20474a <=( (not A200)  and  a20473a );
 a20475a <=( a20474a  and  a20469a );
 a20479a <=( A298  and  A266 );
 a20480a <=( A265  and  a20479a );
 a20484a <=( A301  and  A300 );
 a20485a <=( (not A299)  and  a20484a );
 a20486a <=( a20485a  and  a20480a );
 a20490a <=( (not A199)  and  A167 );
 a20491a <=( A168  and  a20490a );
 a20495a <=( (not A234)  and  (not A233) );
 a20496a <=( (not A200)  and  a20495a );
 a20497a <=( a20496a  and  a20491a );
 a20501a <=( A298  and  A266 );
 a20502a <=( A265  and  a20501a );
 a20506a <=( A302  and  A300 );
 a20507a <=( (not A299)  and  a20506a );
 a20508a <=( a20507a  and  a20502a );
 a20512a <=( (not A199)  and  A167 );
 a20513a <=( A168  and  a20512a );
 a20517a <=( (not A234)  and  (not A233) );
 a20518a <=( (not A200)  and  a20517a );
 a20519a <=( a20518a  and  a20513a );
 a20523a <=( A298  and  (not A267) );
 a20524a <=( (not A266)  and  a20523a );
 a20528a <=( A301  and  A300 );
 a20529a <=( (not A299)  and  a20528a );
 a20530a <=( a20529a  and  a20524a );
 a20534a <=( (not A199)  and  A167 );
 a20535a <=( A168  and  a20534a );
 a20539a <=( (not A234)  and  (not A233) );
 a20540a <=( (not A200)  and  a20539a );
 a20541a <=( a20540a  and  a20535a );
 a20545a <=( A298  and  (not A267) );
 a20546a <=( (not A266)  and  a20545a );
 a20550a <=( A302  and  A300 );
 a20551a <=( (not A299)  and  a20550a );
 a20552a <=( a20551a  and  a20546a );
 a20556a <=( (not A199)  and  A167 );
 a20557a <=( A168  and  a20556a );
 a20561a <=( (not A234)  and  (not A233) );
 a20562a <=( (not A200)  and  a20561a );
 a20563a <=( a20562a  and  a20557a );
 a20567a <=( A298  and  (not A266) );
 a20568a <=( (not A265)  and  a20567a );
 a20572a <=( A301  and  A300 );
 a20573a <=( (not A299)  and  a20572a );
 a20574a <=( a20573a  and  a20568a );
 a20578a <=( (not A199)  and  A167 );
 a20579a <=( A168  and  a20578a );
 a20583a <=( (not A234)  and  (not A233) );
 a20584a <=( (not A200)  and  a20583a );
 a20585a <=( a20584a  and  a20579a );
 a20589a <=( A298  and  (not A266) );
 a20590a <=( (not A265)  and  a20589a );
 a20594a <=( A302  and  A300 );
 a20595a <=( (not A299)  and  a20594a );
 a20596a <=( a20595a  and  a20590a );
 a20600a <=( (not A199)  and  A167 );
 a20601a <=( A168  and  a20600a );
 a20605a <=( (not A233)  and  A232 );
 a20606a <=( (not A200)  and  a20605a );
 a20607a <=( a20606a  and  a20601a );
 a20611a <=( A265  and  A235 );
 a20612a <=( A234  and  a20611a );
 a20616a <=( A268  and  A267 );
 a20617a <=( (not A266)  and  a20616a );
 a20618a <=( a20617a  and  a20612a );
 a20622a <=( (not A199)  and  A167 );
 a20623a <=( A168  and  a20622a );
 a20627a <=( (not A233)  and  A232 );
 a20628a <=( (not A200)  and  a20627a );
 a20629a <=( a20628a  and  a20623a );
 a20633a <=( A265  and  A235 );
 a20634a <=( A234  and  a20633a );
 a20638a <=( A269  and  A267 );
 a20639a <=( (not A266)  and  a20638a );
 a20640a <=( a20639a  and  a20634a );
 a20644a <=( (not A199)  and  A167 );
 a20645a <=( A168  and  a20644a );
 a20649a <=( (not A233)  and  A232 );
 a20650a <=( (not A200)  and  a20649a );
 a20651a <=( a20650a  and  a20645a );
 a20655a <=( A265  and  A236 );
 a20656a <=( A234  and  a20655a );
 a20660a <=( A268  and  A267 );
 a20661a <=( (not A266)  and  a20660a );
 a20662a <=( a20661a  and  a20656a );
 a20666a <=( (not A199)  and  A167 );
 a20667a <=( A168  and  a20666a );
 a20671a <=( (not A233)  and  A232 );
 a20672a <=( (not A200)  and  a20671a );
 a20673a <=( a20672a  and  a20667a );
 a20677a <=( A265  and  A236 );
 a20678a <=( A234  and  a20677a );
 a20682a <=( A269  and  A267 );
 a20683a <=( (not A266)  and  a20682a );
 a20684a <=( a20683a  and  a20678a );
 a20688a <=( (not A199)  and  A167 );
 a20689a <=( A168  and  a20688a );
 a20693a <=( (not A233)  and  (not A232) );
 a20694a <=( (not A200)  and  a20693a );
 a20695a <=( a20694a  and  a20689a );
 a20699a <=( A298  and  A266 );
 a20700a <=( A265  and  a20699a );
 a20704a <=( A301  and  A300 );
 a20705a <=( (not A299)  and  a20704a );
 a20706a <=( a20705a  and  a20700a );
 a20710a <=( (not A199)  and  A167 );
 a20711a <=( A168  and  a20710a );
 a20715a <=( (not A233)  and  (not A232) );
 a20716a <=( (not A200)  and  a20715a );
 a20717a <=( a20716a  and  a20711a );
 a20721a <=( A298  and  A266 );
 a20722a <=( A265  and  a20721a );
 a20726a <=( A302  and  A300 );
 a20727a <=( (not A299)  and  a20726a );
 a20728a <=( a20727a  and  a20722a );
 a20732a <=( (not A199)  and  A167 );
 a20733a <=( A168  and  a20732a );
 a20737a <=( (not A233)  and  (not A232) );
 a20738a <=( (not A200)  and  a20737a );
 a20739a <=( a20738a  and  a20733a );
 a20743a <=( A298  and  (not A267) );
 a20744a <=( (not A266)  and  a20743a );
 a20748a <=( A301  and  A300 );
 a20749a <=( (not A299)  and  a20748a );
 a20750a <=( a20749a  and  a20744a );
 a20754a <=( (not A199)  and  A167 );
 a20755a <=( A168  and  a20754a );
 a20759a <=( (not A233)  and  (not A232) );
 a20760a <=( (not A200)  and  a20759a );
 a20761a <=( a20760a  and  a20755a );
 a20765a <=( A298  and  (not A267) );
 a20766a <=( (not A266)  and  a20765a );
 a20770a <=( A302  and  A300 );
 a20771a <=( (not A299)  and  a20770a );
 a20772a <=( a20771a  and  a20766a );
 a20776a <=( (not A199)  and  A167 );
 a20777a <=( A168  and  a20776a );
 a20781a <=( (not A233)  and  (not A232) );
 a20782a <=( (not A200)  and  a20781a );
 a20783a <=( a20782a  and  a20777a );
 a20787a <=( A298  and  (not A266) );
 a20788a <=( (not A265)  and  a20787a );
 a20792a <=( A301  and  A300 );
 a20793a <=( (not A299)  and  a20792a );
 a20794a <=( a20793a  and  a20788a );
 a20798a <=( (not A199)  and  A167 );
 a20799a <=( A168  and  a20798a );
 a20803a <=( (not A233)  and  (not A232) );
 a20804a <=( (not A200)  and  a20803a );
 a20805a <=( a20804a  and  a20799a );
 a20809a <=( A298  and  (not A266) );
 a20810a <=( (not A265)  and  a20809a );
 a20814a <=( A302  and  A300 );
 a20815a <=( (not A299)  and  a20814a );
 a20816a <=( a20815a  and  a20810a );
 a20820a <=( (not A166)  and  (not A167) );
 a20821a <=( A170  and  a20820a );
 a20825a <=( A232  and  A200 );
 a20826a <=( (not A199)  and  a20825a );
 a20827a <=( a20826a  and  a20821a );
 a20831a <=( (not A268)  and  A265 );
 a20832a <=( A233  and  a20831a );
 a20836a <=( A299  and  (not A298) );
 a20837a <=( (not A269)  and  a20836a );
 a20838a <=( a20837a  and  a20832a );
 a20842a <=( (not A166)  and  (not A167) );
 a20843a <=( A170  and  a20842a );
 a20847a <=( (not A233)  and  A200 );
 a20848a <=( (not A199)  and  a20847a );
 a20849a <=( a20848a  and  a20843a );
 a20853a <=( A265  and  (not A236) );
 a20854a <=( (not A235)  and  a20853a );
 a20858a <=( A299  and  (not A298) );
 a20859a <=( A266  and  a20858a );
 a20860a <=( a20859a  and  a20854a );
 a20864a <=( (not A166)  and  (not A167) );
 a20865a <=( A170  and  a20864a );
 a20869a <=( (not A233)  and  A200 );
 a20870a <=( (not A199)  and  a20869a );
 a20871a <=( a20870a  and  a20865a );
 a20875a <=( (not A266)  and  (not A236) );
 a20876a <=( (not A235)  and  a20875a );
 a20880a <=( A299  and  (not A298) );
 a20881a <=( (not A267)  and  a20880a );
 a20882a <=( a20881a  and  a20876a );
 a20886a <=( (not A166)  and  (not A167) );
 a20887a <=( A170  and  a20886a );
 a20891a <=( (not A233)  and  A200 );
 a20892a <=( (not A199)  and  a20891a );
 a20893a <=( a20892a  and  a20887a );
 a20897a <=( (not A265)  and  (not A236) );
 a20898a <=( (not A235)  and  a20897a );
 a20902a <=( A299  and  (not A298) );
 a20903a <=( (not A266)  and  a20902a );
 a20904a <=( a20903a  and  a20898a );
 a20908a <=( (not A166)  and  (not A167) );
 a20909a <=( A170  and  a20908a );
 a20913a <=( (not A233)  and  A200 );
 a20914a <=( (not A199)  and  a20913a );
 a20915a <=( a20914a  and  a20909a );
 a20919a <=( (not A268)  and  (not A266) );
 a20920a <=( (not A234)  and  a20919a );
 a20924a <=( A299  and  (not A298) );
 a20925a <=( (not A269)  and  a20924a );
 a20926a <=( a20925a  and  a20920a );
 a20930a <=( (not A166)  and  (not A167) );
 a20931a <=( A170  and  a20930a );
 a20935a <=( A232  and  A200 );
 a20936a <=( (not A199)  and  a20935a );
 a20937a <=( a20936a  and  a20931a );
 a20941a <=( A235  and  A234 );
 a20942a <=( (not A233)  and  a20941a );
 a20946a <=( (not A302)  and  (not A301) );
 a20947a <=( A298  and  a20946a );
 a20948a <=( a20947a  and  a20942a );
 a20952a <=( (not A166)  and  (not A167) );
 a20953a <=( A170  and  a20952a );
 a20957a <=( A232  and  A200 );
 a20958a <=( (not A199)  and  a20957a );
 a20959a <=( a20958a  and  a20953a );
 a20963a <=( A236  and  A234 );
 a20964a <=( (not A233)  and  a20963a );
 a20968a <=( (not A302)  and  (not A301) );
 a20969a <=( A298  and  a20968a );
 a20970a <=( a20969a  and  a20964a );
 a20974a <=( (not A166)  and  (not A167) );
 a20975a <=( A170  and  a20974a );
 a20979a <=( (not A232)  and  A200 );
 a20980a <=( (not A199)  and  a20979a );
 a20981a <=( a20980a  and  a20975a );
 a20985a <=( (not A268)  and  (not A266) );
 a20986a <=( (not A233)  and  a20985a );
 a20990a <=( A299  and  (not A298) );
 a20991a <=( (not A269)  and  a20990a );
 a20992a <=( a20991a  and  a20986a );
 a20996a <=( (not A166)  and  (not A167) );
 a20997a <=( A170  and  a20996a );
 a21001a <=( A201  and  (not A200) );
 a21002a <=( A199  and  a21001a );
 a21003a <=( a21002a  and  a20997a );
 a21007a <=( A233  and  (not A232) );
 a21008a <=( A202  and  a21007a );
 a21012a <=( (not A302)  and  (not A301) );
 a21013a <=( (not A299)  and  a21012a );
 a21014a <=( a21013a  and  a21008a );
 a21018a <=( (not A166)  and  (not A167) );
 a21019a <=( A170  and  a21018a );
 a21023a <=( A201  and  (not A200) );
 a21024a <=( A199  and  a21023a );
 a21025a <=( a21024a  and  a21019a );
 a21029a <=( A233  and  (not A232) );
 a21030a <=( A203  and  a21029a );
 a21034a <=( (not A302)  and  (not A301) );
 a21035a <=( (not A299)  and  a21034a );
 a21036a <=( a21035a  and  a21030a );
 a21040a <=( A167  and  (not A168) );
 a21041a <=( A170  and  a21040a );
 a21045a <=( A200  and  (not A199) );
 a21046a <=( A166  and  a21045a );
 a21047a <=( a21046a  and  a21041a );
 a21051a <=( A265  and  A233 );
 a21052a <=( A232  and  a21051a );
 a21056a <=( A299  and  (not A298) );
 a21057a <=( (not A267)  and  a21056a );
 a21058a <=( a21057a  and  a21052a );
 a21062a <=( A167  and  (not A168) );
 a21063a <=( A170  and  a21062a );
 a21067a <=( A200  and  (not A199) );
 a21068a <=( A166  and  a21067a );
 a21069a <=( a21068a  and  a21063a );
 a21073a <=( A265  and  A233 );
 a21074a <=( A232  and  a21073a );
 a21078a <=( A299  and  (not A298) );
 a21079a <=( A266  and  a21078a );
 a21080a <=( a21079a  and  a21074a );
 a21084a <=( A167  and  (not A168) );
 a21085a <=( A170  and  a21084a );
 a21089a <=( A200  and  (not A199) );
 a21090a <=( A166  and  a21089a );
 a21091a <=( a21090a  and  a21085a );
 a21095a <=( (not A265)  and  A233 );
 a21096a <=( A232  and  a21095a );
 a21100a <=( A299  and  (not A298) );
 a21101a <=( (not A266)  and  a21100a );
 a21102a <=( a21101a  and  a21096a );
 a21106a <=( A167  and  (not A168) );
 a21107a <=( A170  and  a21106a );
 a21111a <=( A200  and  (not A199) );
 a21112a <=( A166  and  a21111a );
 a21113a <=( a21112a  and  a21107a );
 a21117a <=( A265  and  A233 );
 a21118a <=( (not A232)  and  a21117a );
 a21122a <=( A268  and  A267 );
 a21123a <=( (not A266)  and  a21122a );
 a21124a <=( a21123a  and  a21118a );
 a21128a <=( A167  and  (not A168) );
 a21129a <=( A170  and  a21128a );
 a21133a <=( A200  and  (not A199) );
 a21134a <=( A166  and  a21133a );
 a21135a <=( a21134a  and  a21129a );
 a21139a <=( A265  and  A233 );
 a21140a <=( (not A232)  and  a21139a );
 a21144a <=( A269  and  A267 );
 a21145a <=( (not A266)  and  a21144a );
 a21146a <=( a21145a  and  a21140a );
 a21150a <=( A167  and  (not A168) );
 a21151a <=( A170  and  a21150a );
 a21155a <=( A200  and  (not A199) );
 a21156a <=( A166  and  a21155a );
 a21157a <=( a21156a  and  a21151a );
 a21161a <=( A265  and  (not A234) );
 a21162a <=( (not A233)  and  a21161a );
 a21166a <=( A299  and  (not A298) );
 a21167a <=( A266  and  a21166a );
 a21168a <=( a21167a  and  a21162a );
 a21172a <=( A167  and  (not A168) );
 a21173a <=( A170  and  a21172a );
 a21177a <=( A200  and  (not A199) );
 a21178a <=( A166  and  a21177a );
 a21179a <=( a21178a  and  a21173a );
 a21183a <=( (not A266)  and  (not A234) );
 a21184a <=( (not A233)  and  a21183a );
 a21188a <=( A299  and  (not A298) );
 a21189a <=( (not A267)  and  a21188a );
 a21190a <=( a21189a  and  a21184a );
 a21194a <=( A167  and  (not A168) );
 a21195a <=( A170  and  a21194a );
 a21199a <=( A200  and  (not A199) );
 a21200a <=( A166  and  a21199a );
 a21201a <=( a21200a  and  a21195a );
 a21205a <=( (not A265)  and  (not A234) );
 a21206a <=( (not A233)  and  a21205a );
 a21210a <=( A299  and  (not A298) );
 a21211a <=( (not A266)  and  a21210a );
 a21212a <=( a21211a  and  a21206a );
 a21216a <=( A167  and  (not A168) );
 a21217a <=( A170  and  a21216a );
 a21221a <=( A200  and  (not A199) );
 a21222a <=( A166  and  a21221a );
 a21223a <=( a21222a  and  a21217a );
 a21227a <=( A234  and  (not A233) );
 a21228a <=( A232  and  a21227a );
 a21232a <=( (not A300)  and  A298 );
 a21233a <=( A235  and  a21232a );
 a21234a <=( a21233a  and  a21228a );
 a21238a <=( A167  and  (not A168) );
 a21239a <=( A170  and  a21238a );
 a21243a <=( A200  and  (not A199) );
 a21244a <=( A166  and  a21243a );
 a21245a <=( a21244a  and  a21239a );
 a21249a <=( A234  and  (not A233) );
 a21250a <=( A232  and  a21249a );
 a21254a <=( A299  and  A298 );
 a21255a <=( A235  and  a21254a );
 a21256a <=( a21255a  and  a21250a );
 a21260a <=( A167  and  (not A168) );
 a21261a <=( A170  and  a21260a );
 a21265a <=( A200  and  (not A199) );
 a21266a <=( A166  and  a21265a );
 a21267a <=( a21266a  and  a21261a );
 a21271a <=( A234  and  (not A233) );
 a21272a <=( A232  and  a21271a );
 a21276a <=( (not A299)  and  (not A298) );
 a21277a <=( A235  and  a21276a );
 a21278a <=( a21277a  and  a21272a );
 a21282a <=( A167  and  (not A168) );
 a21283a <=( A170  and  a21282a );
 a21287a <=( A200  and  (not A199) );
 a21288a <=( A166  and  a21287a );
 a21289a <=( a21288a  and  a21283a );
 a21293a <=( A234  and  (not A233) );
 a21294a <=( A232  and  a21293a );
 a21298a <=( A266  and  (not A265) );
 a21299a <=( A235  and  a21298a );
 a21300a <=( a21299a  and  a21294a );
 a21304a <=( A167  and  (not A168) );
 a21305a <=( A170  and  a21304a );
 a21309a <=( A200  and  (not A199) );
 a21310a <=( A166  and  a21309a );
 a21311a <=( a21310a  and  a21305a );
 a21315a <=( A234  and  (not A233) );
 a21316a <=( A232  and  a21315a );
 a21320a <=( (not A300)  and  A298 );
 a21321a <=( A236  and  a21320a );
 a21322a <=( a21321a  and  a21316a );
 a21326a <=( A167  and  (not A168) );
 a21327a <=( A170  and  a21326a );
 a21331a <=( A200  and  (not A199) );
 a21332a <=( A166  and  a21331a );
 a21333a <=( a21332a  and  a21327a );
 a21337a <=( A234  and  (not A233) );
 a21338a <=( A232  and  a21337a );
 a21342a <=( A299  and  A298 );
 a21343a <=( A236  and  a21342a );
 a21344a <=( a21343a  and  a21338a );
 a21348a <=( A167  and  (not A168) );
 a21349a <=( A170  and  a21348a );
 a21353a <=( A200  and  (not A199) );
 a21354a <=( A166  and  a21353a );
 a21355a <=( a21354a  and  a21349a );
 a21359a <=( A234  and  (not A233) );
 a21360a <=( A232  and  a21359a );
 a21364a <=( (not A299)  and  (not A298) );
 a21365a <=( A236  and  a21364a );
 a21366a <=( a21365a  and  a21360a );
 a21370a <=( A167  and  (not A168) );
 a21371a <=( A170  and  a21370a );
 a21375a <=( A200  and  (not A199) );
 a21376a <=( A166  and  a21375a );
 a21377a <=( a21376a  and  a21371a );
 a21381a <=( A234  and  (not A233) );
 a21382a <=( A232  and  a21381a );
 a21386a <=( A266  and  (not A265) );
 a21387a <=( A236  and  a21386a );
 a21388a <=( a21387a  and  a21382a );
 a21392a <=( A167  and  (not A168) );
 a21393a <=( A170  and  a21392a );
 a21397a <=( A200  and  (not A199) );
 a21398a <=( A166  and  a21397a );
 a21399a <=( a21398a  and  a21393a );
 a21403a <=( A265  and  (not A233) );
 a21404a <=( (not A232)  and  a21403a );
 a21408a <=( A299  and  (not A298) );
 a21409a <=( A266  and  a21408a );
 a21410a <=( a21409a  and  a21404a );
 a21414a <=( A167  and  (not A168) );
 a21415a <=( A170  and  a21414a );
 a21419a <=( A200  and  (not A199) );
 a21420a <=( A166  and  a21419a );
 a21421a <=( a21420a  and  a21415a );
 a21425a <=( (not A266)  and  (not A233) );
 a21426a <=( (not A232)  and  a21425a );
 a21430a <=( A299  and  (not A298) );
 a21431a <=( (not A267)  and  a21430a );
 a21432a <=( a21431a  and  a21426a );
 a21436a <=( A167  and  (not A168) );
 a21437a <=( A170  and  a21436a );
 a21441a <=( A200  and  (not A199) );
 a21442a <=( A166  and  a21441a );
 a21443a <=( a21442a  and  a21437a );
 a21447a <=( (not A265)  and  (not A233) );
 a21448a <=( (not A232)  and  a21447a );
 a21452a <=( A299  and  (not A298) );
 a21453a <=( (not A266)  and  a21452a );
 a21454a <=( a21453a  and  a21448a );
 a21458a <=( A167  and  (not A168) );
 a21459a <=( (not A170)  and  a21458a );
 a21463a <=( A200  and  (not A199) );
 a21464a <=( (not A166)  and  a21463a );
 a21465a <=( a21464a  and  a21459a );
 a21469a <=( A265  and  A233 );
 a21470a <=( A232  and  a21469a );
 a21474a <=( A299  and  (not A298) );
 a21475a <=( (not A267)  and  a21474a );
 a21476a <=( a21475a  and  a21470a );
 a21480a <=( A167  and  (not A168) );
 a21481a <=( (not A170)  and  a21480a );
 a21485a <=( A200  and  (not A199) );
 a21486a <=( (not A166)  and  a21485a );
 a21487a <=( a21486a  and  a21481a );
 a21491a <=( A265  and  A233 );
 a21492a <=( A232  and  a21491a );
 a21496a <=( A299  and  (not A298) );
 a21497a <=( A266  and  a21496a );
 a21498a <=( a21497a  and  a21492a );
 a21502a <=( A167  and  (not A168) );
 a21503a <=( (not A170)  and  a21502a );
 a21507a <=( A200  and  (not A199) );
 a21508a <=( (not A166)  and  a21507a );
 a21509a <=( a21508a  and  a21503a );
 a21513a <=( (not A265)  and  A233 );
 a21514a <=( A232  and  a21513a );
 a21518a <=( A299  and  (not A298) );
 a21519a <=( (not A266)  and  a21518a );
 a21520a <=( a21519a  and  a21514a );
 a21524a <=( A167  and  (not A168) );
 a21525a <=( (not A170)  and  a21524a );
 a21529a <=( A200  and  (not A199) );
 a21530a <=( (not A166)  and  a21529a );
 a21531a <=( a21530a  and  a21525a );
 a21535a <=( A265  and  A233 );
 a21536a <=( (not A232)  and  a21535a );
 a21540a <=( A268  and  A267 );
 a21541a <=( (not A266)  and  a21540a );
 a21542a <=( a21541a  and  a21536a );
 a21546a <=( A167  and  (not A168) );
 a21547a <=( (not A170)  and  a21546a );
 a21551a <=( A200  and  (not A199) );
 a21552a <=( (not A166)  and  a21551a );
 a21553a <=( a21552a  and  a21547a );
 a21557a <=( A265  and  A233 );
 a21558a <=( (not A232)  and  a21557a );
 a21562a <=( A269  and  A267 );
 a21563a <=( (not A266)  and  a21562a );
 a21564a <=( a21563a  and  a21558a );
 a21568a <=( A167  and  (not A168) );
 a21569a <=( (not A170)  and  a21568a );
 a21573a <=( A200  and  (not A199) );
 a21574a <=( (not A166)  and  a21573a );
 a21575a <=( a21574a  and  a21569a );
 a21579a <=( A265  and  (not A234) );
 a21580a <=( (not A233)  and  a21579a );
 a21584a <=( A299  and  (not A298) );
 a21585a <=( A266  and  a21584a );
 a21586a <=( a21585a  and  a21580a );
 a21590a <=( A167  and  (not A168) );
 a21591a <=( (not A170)  and  a21590a );
 a21595a <=( A200  and  (not A199) );
 a21596a <=( (not A166)  and  a21595a );
 a21597a <=( a21596a  and  a21591a );
 a21601a <=( (not A266)  and  (not A234) );
 a21602a <=( (not A233)  and  a21601a );
 a21606a <=( A299  and  (not A298) );
 a21607a <=( (not A267)  and  a21606a );
 a21608a <=( a21607a  and  a21602a );
 a21612a <=( A167  and  (not A168) );
 a21613a <=( (not A170)  and  a21612a );
 a21617a <=( A200  and  (not A199) );
 a21618a <=( (not A166)  and  a21617a );
 a21619a <=( a21618a  and  a21613a );
 a21623a <=( (not A265)  and  (not A234) );
 a21624a <=( (not A233)  and  a21623a );
 a21628a <=( A299  and  (not A298) );
 a21629a <=( (not A266)  and  a21628a );
 a21630a <=( a21629a  and  a21624a );
 a21634a <=( A167  and  (not A168) );
 a21635a <=( (not A170)  and  a21634a );
 a21639a <=( A200  and  (not A199) );
 a21640a <=( (not A166)  and  a21639a );
 a21641a <=( a21640a  and  a21635a );
 a21645a <=( A234  and  (not A233) );
 a21646a <=( A232  and  a21645a );
 a21650a <=( (not A300)  and  A298 );
 a21651a <=( A235  and  a21650a );
 a21652a <=( a21651a  and  a21646a );
 a21656a <=( A167  and  (not A168) );
 a21657a <=( (not A170)  and  a21656a );
 a21661a <=( A200  and  (not A199) );
 a21662a <=( (not A166)  and  a21661a );
 a21663a <=( a21662a  and  a21657a );
 a21667a <=( A234  and  (not A233) );
 a21668a <=( A232  and  a21667a );
 a21672a <=( A299  and  A298 );
 a21673a <=( A235  and  a21672a );
 a21674a <=( a21673a  and  a21668a );
 a21678a <=( A167  and  (not A168) );
 a21679a <=( (not A170)  and  a21678a );
 a21683a <=( A200  and  (not A199) );
 a21684a <=( (not A166)  and  a21683a );
 a21685a <=( a21684a  and  a21679a );
 a21689a <=( A234  and  (not A233) );
 a21690a <=( A232  and  a21689a );
 a21694a <=( (not A299)  and  (not A298) );
 a21695a <=( A235  and  a21694a );
 a21696a <=( a21695a  and  a21690a );
 a21700a <=( A167  and  (not A168) );
 a21701a <=( (not A170)  and  a21700a );
 a21705a <=( A200  and  (not A199) );
 a21706a <=( (not A166)  and  a21705a );
 a21707a <=( a21706a  and  a21701a );
 a21711a <=( A234  and  (not A233) );
 a21712a <=( A232  and  a21711a );
 a21716a <=( A266  and  (not A265) );
 a21717a <=( A235  and  a21716a );
 a21718a <=( a21717a  and  a21712a );
 a21722a <=( A167  and  (not A168) );
 a21723a <=( (not A170)  and  a21722a );
 a21727a <=( A200  and  (not A199) );
 a21728a <=( (not A166)  and  a21727a );
 a21729a <=( a21728a  and  a21723a );
 a21733a <=( A234  and  (not A233) );
 a21734a <=( A232  and  a21733a );
 a21738a <=( (not A300)  and  A298 );
 a21739a <=( A236  and  a21738a );
 a21740a <=( a21739a  and  a21734a );
 a21744a <=( A167  and  (not A168) );
 a21745a <=( (not A170)  and  a21744a );
 a21749a <=( A200  and  (not A199) );
 a21750a <=( (not A166)  and  a21749a );
 a21751a <=( a21750a  and  a21745a );
 a21755a <=( A234  and  (not A233) );
 a21756a <=( A232  and  a21755a );
 a21760a <=( A299  and  A298 );
 a21761a <=( A236  and  a21760a );
 a21762a <=( a21761a  and  a21756a );
 a21766a <=( A167  and  (not A168) );
 a21767a <=( (not A170)  and  a21766a );
 a21771a <=( A200  and  (not A199) );
 a21772a <=( (not A166)  and  a21771a );
 a21773a <=( a21772a  and  a21767a );
 a21777a <=( A234  and  (not A233) );
 a21778a <=( A232  and  a21777a );
 a21782a <=( (not A299)  and  (not A298) );
 a21783a <=( A236  and  a21782a );
 a21784a <=( a21783a  and  a21778a );
 a21788a <=( A167  and  (not A168) );
 a21789a <=( (not A170)  and  a21788a );
 a21793a <=( A200  and  (not A199) );
 a21794a <=( (not A166)  and  a21793a );
 a21795a <=( a21794a  and  a21789a );
 a21799a <=( A234  and  (not A233) );
 a21800a <=( A232  and  a21799a );
 a21804a <=( A266  and  (not A265) );
 a21805a <=( A236  and  a21804a );
 a21806a <=( a21805a  and  a21800a );
 a21810a <=( A167  and  (not A168) );
 a21811a <=( (not A170)  and  a21810a );
 a21815a <=( A200  and  (not A199) );
 a21816a <=( (not A166)  and  a21815a );
 a21817a <=( a21816a  and  a21811a );
 a21821a <=( A265  and  (not A233) );
 a21822a <=( (not A232)  and  a21821a );
 a21826a <=( A299  and  (not A298) );
 a21827a <=( A266  and  a21826a );
 a21828a <=( a21827a  and  a21822a );
 a21832a <=( A167  and  (not A168) );
 a21833a <=( (not A170)  and  a21832a );
 a21837a <=( A200  and  (not A199) );
 a21838a <=( (not A166)  and  a21837a );
 a21839a <=( a21838a  and  a21833a );
 a21843a <=( (not A266)  and  (not A233) );
 a21844a <=( (not A232)  and  a21843a );
 a21848a <=( A299  and  (not A298) );
 a21849a <=( (not A267)  and  a21848a );
 a21850a <=( a21849a  and  a21844a );
 a21854a <=( A167  and  (not A168) );
 a21855a <=( (not A170)  and  a21854a );
 a21859a <=( A200  and  (not A199) );
 a21860a <=( (not A166)  and  a21859a );
 a21861a <=( a21860a  and  a21855a );
 a21865a <=( (not A265)  and  (not A233) );
 a21866a <=( (not A232)  and  a21865a );
 a21870a <=( A299  and  (not A298) );
 a21871a <=( (not A266)  and  a21870a );
 a21872a <=( a21871a  and  a21866a );
 a21876a <=( (not A167)  and  (not A168) );
 a21877a <=( (not A170)  and  a21876a );
 a21881a <=( A200  and  (not A199) );
 a21882a <=( A166  and  a21881a );
 a21883a <=( a21882a  and  a21877a );
 a21887a <=( A265  and  A233 );
 a21888a <=( A232  and  a21887a );
 a21892a <=( A299  and  (not A298) );
 a21893a <=( (not A267)  and  a21892a );
 a21894a <=( a21893a  and  a21888a );
 a21898a <=( (not A167)  and  (not A168) );
 a21899a <=( (not A170)  and  a21898a );
 a21903a <=( A200  and  (not A199) );
 a21904a <=( A166  and  a21903a );
 a21905a <=( a21904a  and  a21899a );
 a21909a <=( A265  and  A233 );
 a21910a <=( A232  and  a21909a );
 a21914a <=( A299  and  (not A298) );
 a21915a <=( A266  and  a21914a );
 a21916a <=( a21915a  and  a21910a );
 a21920a <=( (not A167)  and  (not A168) );
 a21921a <=( (not A170)  and  a21920a );
 a21925a <=( A200  and  (not A199) );
 a21926a <=( A166  and  a21925a );
 a21927a <=( a21926a  and  a21921a );
 a21931a <=( (not A265)  and  A233 );
 a21932a <=( A232  and  a21931a );
 a21936a <=( A299  and  (not A298) );
 a21937a <=( (not A266)  and  a21936a );
 a21938a <=( a21937a  and  a21932a );
 a21942a <=( (not A167)  and  (not A168) );
 a21943a <=( (not A170)  and  a21942a );
 a21947a <=( A200  and  (not A199) );
 a21948a <=( A166  and  a21947a );
 a21949a <=( a21948a  and  a21943a );
 a21953a <=( A265  and  A233 );
 a21954a <=( (not A232)  and  a21953a );
 a21958a <=( A268  and  A267 );
 a21959a <=( (not A266)  and  a21958a );
 a21960a <=( a21959a  and  a21954a );
 a21964a <=( (not A167)  and  (not A168) );
 a21965a <=( (not A170)  and  a21964a );
 a21969a <=( A200  and  (not A199) );
 a21970a <=( A166  and  a21969a );
 a21971a <=( a21970a  and  a21965a );
 a21975a <=( A265  and  A233 );
 a21976a <=( (not A232)  and  a21975a );
 a21980a <=( A269  and  A267 );
 a21981a <=( (not A266)  and  a21980a );
 a21982a <=( a21981a  and  a21976a );
 a21986a <=( (not A167)  and  (not A168) );
 a21987a <=( (not A170)  and  a21986a );
 a21991a <=( A200  and  (not A199) );
 a21992a <=( A166  and  a21991a );
 a21993a <=( a21992a  and  a21987a );
 a21997a <=( A265  and  (not A234) );
 a21998a <=( (not A233)  and  a21997a );
 a22002a <=( A299  and  (not A298) );
 a22003a <=( A266  and  a22002a );
 a22004a <=( a22003a  and  a21998a );
 a22008a <=( (not A167)  and  (not A168) );
 a22009a <=( (not A170)  and  a22008a );
 a22013a <=( A200  and  (not A199) );
 a22014a <=( A166  and  a22013a );
 a22015a <=( a22014a  and  a22009a );
 a22019a <=( (not A266)  and  (not A234) );
 a22020a <=( (not A233)  and  a22019a );
 a22024a <=( A299  and  (not A298) );
 a22025a <=( (not A267)  and  a22024a );
 a22026a <=( a22025a  and  a22020a );
 a22030a <=( (not A167)  and  (not A168) );
 a22031a <=( (not A170)  and  a22030a );
 a22035a <=( A200  and  (not A199) );
 a22036a <=( A166  and  a22035a );
 a22037a <=( a22036a  and  a22031a );
 a22041a <=( (not A265)  and  (not A234) );
 a22042a <=( (not A233)  and  a22041a );
 a22046a <=( A299  and  (not A298) );
 a22047a <=( (not A266)  and  a22046a );
 a22048a <=( a22047a  and  a22042a );
 a22052a <=( (not A167)  and  (not A168) );
 a22053a <=( (not A170)  and  a22052a );
 a22057a <=( A200  and  (not A199) );
 a22058a <=( A166  and  a22057a );
 a22059a <=( a22058a  and  a22053a );
 a22063a <=( A234  and  (not A233) );
 a22064a <=( A232  and  a22063a );
 a22068a <=( (not A300)  and  A298 );
 a22069a <=( A235  and  a22068a );
 a22070a <=( a22069a  and  a22064a );
 a22074a <=( (not A167)  and  (not A168) );
 a22075a <=( (not A170)  and  a22074a );
 a22079a <=( A200  and  (not A199) );
 a22080a <=( A166  and  a22079a );
 a22081a <=( a22080a  and  a22075a );
 a22085a <=( A234  and  (not A233) );
 a22086a <=( A232  and  a22085a );
 a22090a <=( A299  and  A298 );
 a22091a <=( A235  and  a22090a );
 a22092a <=( a22091a  and  a22086a );
 a22096a <=( (not A167)  and  (not A168) );
 a22097a <=( (not A170)  and  a22096a );
 a22101a <=( A200  and  (not A199) );
 a22102a <=( A166  and  a22101a );
 a22103a <=( a22102a  and  a22097a );
 a22107a <=( A234  and  (not A233) );
 a22108a <=( A232  and  a22107a );
 a22112a <=( (not A299)  and  (not A298) );
 a22113a <=( A235  and  a22112a );
 a22114a <=( a22113a  and  a22108a );
 a22118a <=( (not A167)  and  (not A168) );
 a22119a <=( (not A170)  and  a22118a );
 a22123a <=( A200  and  (not A199) );
 a22124a <=( A166  and  a22123a );
 a22125a <=( a22124a  and  a22119a );
 a22129a <=( A234  and  (not A233) );
 a22130a <=( A232  and  a22129a );
 a22134a <=( A266  and  (not A265) );
 a22135a <=( A235  and  a22134a );
 a22136a <=( a22135a  and  a22130a );
 a22140a <=( (not A167)  and  (not A168) );
 a22141a <=( (not A170)  and  a22140a );
 a22145a <=( A200  and  (not A199) );
 a22146a <=( A166  and  a22145a );
 a22147a <=( a22146a  and  a22141a );
 a22151a <=( A234  and  (not A233) );
 a22152a <=( A232  and  a22151a );
 a22156a <=( (not A300)  and  A298 );
 a22157a <=( A236  and  a22156a );
 a22158a <=( a22157a  and  a22152a );
 a22162a <=( (not A167)  and  (not A168) );
 a22163a <=( (not A170)  and  a22162a );
 a22167a <=( A200  and  (not A199) );
 a22168a <=( A166  and  a22167a );
 a22169a <=( a22168a  and  a22163a );
 a22173a <=( A234  and  (not A233) );
 a22174a <=( A232  and  a22173a );
 a22178a <=( A299  and  A298 );
 a22179a <=( A236  and  a22178a );
 a22180a <=( a22179a  and  a22174a );
 a22184a <=( (not A167)  and  (not A168) );
 a22185a <=( (not A170)  and  a22184a );
 a22189a <=( A200  and  (not A199) );
 a22190a <=( A166  and  a22189a );
 a22191a <=( a22190a  and  a22185a );
 a22195a <=( A234  and  (not A233) );
 a22196a <=( A232  and  a22195a );
 a22200a <=( (not A299)  and  (not A298) );
 a22201a <=( A236  and  a22200a );
 a22202a <=( a22201a  and  a22196a );
 a22206a <=( (not A167)  and  (not A168) );
 a22207a <=( (not A170)  and  a22206a );
 a22211a <=( A200  and  (not A199) );
 a22212a <=( A166  and  a22211a );
 a22213a <=( a22212a  and  a22207a );
 a22217a <=( A234  and  (not A233) );
 a22218a <=( A232  and  a22217a );
 a22222a <=( A266  and  (not A265) );
 a22223a <=( A236  and  a22222a );
 a22224a <=( a22223a  and  a22218a );
 a22228a <=( (not A167)  and  (not A168) );
 a22229a <=( (not A170)  and  a22228a );
 a22233a <=( A200  and  (not A199) );
 a22234a <=( A166  and  a22233a );
 a22235a <=( a22234a  and  a22229a );
 a22239a <=( A265  and  (not A233) );
 a22240a <=( (not A232)  and  a22239a );
 a22244a <=( A299  and  (not A298) );
 a22245a <=( A266  and  a22244a );
 a22246a <=( a22245a  and  a22240a );
 a22250a <=( (not A167)  and  (not A168) );
 a22251a <=( (not A170)  and  a22250a );
 a22255a <=( A200  and  (not A199) );
 a22256a <=( A166  and  a22255a );
 a22257a <=( a22256a  and  a22251a );
 a22261a <=( (not A266)  and  (not A233) );
 a22262a <=( (not A232)  and  a22261a );
 a22266a <=( A299  and  (not A298) );
 a22267a <=( (not A267)  and  a22266a );
 a22268a <=( a22267a  and  a22262a );
 a22272a <=( (not A167)  and  (not A168) );
 a22273a <=( (not A170)  and  a22272a );
 a22277a <=( A200  and  (not A199) );
 a22278a <=( A166  and  a22277a );
 a22279a <=( a22278a  and  a22273a );
 a22283a <=( (not A265)  and  (not A233) );
 a22284a <=( (not A232)  and  a22283a );
 a22288a <=( A299  and  (not A298) );
 a22289a <=( (not A266)  and  a22288a );
 a22290a <=( a22289a  and  a22284a );
 a22294a <=( A167  and  (not A168) );
 a22295a <=( A169  and  a22294a );
 a22299a <=( A200  and  (not A199) );
 a22300a <=( (not A166)  and  a22299a );
 a22301a <=( a22300a  and  a22295a );
 a22305a <=( A265  and  A233 );
 a22306a <=( A232  and  a22305a );
 a22310a <=( A299  and  (not A298) );
 a22311a <=( (not A267)  and  a22310a );
 a22312a <=( a22311a  and  a22306a );
 a22316a <=( A167  and  (not A168) );
 a22317a <=( A169  and  a22316a );
 a22321a <=( A200  and  (not A199) );
 a22322a <=( (not A166)  and  a22321a );
 a22323a <=( a22322a  and  a22317a );
 a22327a <=( A265  and  A233 );
 a22328a <=( A232  and  a22327a );
 a22332a <=( A299  and  (not A298) );
 a22333a <=( A266  and  a22332a );
 a22334a <=( a22333a  and  a22328a );
 a22338a <=( A167  and  (not A168) );
 a22339a <=( A169  and  a22338a );
 a22343a <=( A200  and  (not A199) );
 a22344a <=( (not A166)  and  a22343a );
 a22345a <=( a22344a  and  a22339a );
 a22349a <=( (not A265)  and  A233 );
 a22350a <=( A232  and  a22349a );
 a22354a <=( A299  and  (not A298) );
 a22355a <=( (not A266)  and  a22354a );
 a22356a <=( a22355a  and  a22350a );
 a22360a <=( A167  and  (not A168) );
 a22361a <=( A169  and  a22360a );
 a22365a <=( A200  and  (not A199) );
 a22366a <=( (not A166)  and  a22365a );
 a22367a <=( a22366a  and  a22361a );
 a22371a <=( A265  and  A233 );
 a22372a <=( (not A232)  and  a22371a );
 a22376a <=( A268  and  A267 );
 a22377a <=( (not A266)  and  a22376a );
 a22378a <=( a22377a  and  a22372a );
 a22382a <=( A167  and  (not A168) );
 a22383a <=( A169  and  a22382a );
 a22387a <=( A200  and  (not A199) );
 a22388a <=( (not A166)  and  a22387a );
 a22389a <=( a22388a  and  a22383a );
 a22393a <=( A265  and  A233 );
 a22394a <=( (not A232)  and  a22393a );
 a22398a <=( A269  and  A267 );
 a22399a <=( (not A266)  and  a22398a );
 a22400a <=( a22399a  and  a22394a );
 a22404a <=( A167  and  (not A168) );
 a22405a <=( A169  and  a22404a );
 a22409a <=( A200  and  (not A199) );
 a22410a <=( (not A166)  and  a22409a );
 a22411a <=( a22410a  and  a22405a );
 a22415a <=( A265  and  (not A234) );
 a22416a <=( (not A233)  and  a22415a );
 a22420a <=( A299  and  (not A298) );
 a22421a <=( A266  and  a22420a );
 a22422a <=( a22421a  and  a22416a );
 a22426a <=( A167  and  (not A168) );
 a22427a <=( A169  and  a22426a );
 a22431a <=( A200  and  (not A199) );
 a22432a <=( (not A166)  and  a22431a );
 a22433a <=( a22432a  and  a22427a );
 a22437a <=( (not A266)  and  (not A234) );
 a22438a <=( (not A233)  and  a22437a );
 a22442a <=( A299  and  (not A298) );
 a22443a <=( (not A267)  and  a22442a );
 a22444a <=( a22443a  and  a22438a );
 a22448a <=( A167  and  (not A168) );
 a22449a <=( A169  and  a22448a );
 a22453a <=( A200  and  (not A199) );
 a22454a <=( (not A166)  and  a22453a );
 a22455a <=( a22454a  and  a22449a );
 a22459a <=( (not A265)  and  (not A234) );
 a22460a <=( (not A233)  and  a22459a );
 a22464a <=( A299  and  (not A298) );
 a22465a <=( (not A266)  and  a22464a );
 a22466a <=( a22465a  and  a22460a );
 a22470a <=( A167  and  (not A168) );
 a22471a <=( A169  and  a22470a );
 a22475a <=( A200  and  (not A199) );
 a22476a <=( (not A166)  and  a22475a );
 a22477a <=( a22476a  and  a22471a );
 a22481a <=( A234  and  (not A233) );
 a22482a <=( A232  and  a22481a );
 a22486a <=( (not A300)  and  A298 );
 a22487a <=( A235  and  a22486a );
 a22488a <=( a22487a  and  a22482a );
 a22492a <=( A167  and  (not A168) );
 a22493a <=( A169  and  a22492a );
 a22497a <=( A200  and  (not A199) );
 a22498a <=( (not A166)  and  a22497a );
 a22499a <=( a22498a  and  a22493a );
 a22503a <=( A234  and  (not A233) );
 a22504a <=( A232  and  a22503a );
 a22508a <=( A299  and  A298 );
 a22509a <=( A235  and  a22508a );
 a22510a <=( a22509a  and  a22504a );
 a22514a <=( A167  and  (not A168) );
 a22515a <=( A169  and  a22514a );
 a22519a <=( A200  and  (not A199) );
 a22520a <=( (not A166)  and  a22519a );
 a22521a <=( a22520a  and  a22515a );
 a22525a <=( A234  and  (not A233) );
 a22526a <=( A232  and  a22525a );
 a22530a <=( (not A299)  and  (not A298) );
 a22531a <=( A235  and  a22530a );
 a22532a <=( a22531a  and  a22526a );
 a22536a <=( A167  and  (not A168) );
 a22537a <=( A169  and  a22536a );
 a22541a <=( A200  and  (not A199) );
 a22542a <=( (not A166)  and  a22541a );
 a22543a <=( a22542a  and  a22537a );
 a22547a <=( A234  and  (not A233) );
 a22548a <=( A232  and  a22547a );
 a22552a <=( A266  and  (not A265) );
 a22553a <=( A235  and  a22552a );
 a22554a <=( a22553a  and  a22548a );
 a22558a <=( A167  and  (not A168) );
 a22559a <=( A169  and  a22558a );
 a22563a <=( A200  and  (not A199) );
 a22564a <=( (not A166)  and  a22563a );
 a22565a <=( a22564a  and  a22559a );
 a22569a <=( A234  and  (not A233) );
 a22570a <=( A232  and  a22569a );
 a22574a <=( (not A300)  and  A298 );
 a22575a <=( A236  and  a22574a );
 a22576a <=( a22575a  and  a22570a );
 a22580a <=( A167  and  (not A168) );
 a22581a <=( A169  and  a22580a );
 a22585a <=( A200  and  (not A199) );
 a22586a <=( (not A166)  and  a22585a );
 a22587a <=( a22586a  and  a22581a );
 a22591a <=( A234  and  (not A233) );
 a22592a <=( A232  and  a22591a );
 a22596a <=( A299  and  A298 );
 a22597a <=( A236  and  a22596a );
 a22598a <=( a22597a  and  a22592a );
 a22602a <=( A167  and  (not A168) );
 a22603a <=( A169  and  a22602a );
 a22607a <=( A200  and  (not A199) );
 a22608a <=( (not A166)  and  a22607a );
 a22609a <=( a22608a  and  a22603a );
 a22613a <=( A234  and  (not A233) );
 a22614a <=( A232  and  a22613a );
 a22618a <=( (not A299)  and  (not A298) );
 a22619a <=( A236  and  a22618a );
 a22620a <=( a22619a  and  a22614a );
 a22624a <=( A167  and  (not A168) );
 a22625a <=( A169  and  a22624a );
 a22629a <=( A200  and  (not A199) );
 a22630a <=( (not A166)  and  a22629a );
 a22631a <=( a22630a  and  a22625a );
 a22635a <=( A234  and  (not A233) );
 a22636a <=( A232  and  a22635a );
 a22640a <=( A266  and  (not A265) );
 a22641a <=( A236  and  a22640a );
 a22642a <=( a22641a  and  a22636a );
 a22646a <=( A167  and  (not A168) );
 a22647a <=( A169  and  a22646a );
 a22651a <=( A200  and  (not A199) );
 a22652a <=( (not A166)  and  a22651a );
 a22653a <=( a22652a  and  a22647a );
 a22657a <=( A265  and  (not A233) );
 a22658a <=( (not A232)  and  a22657a );
 a22662a <=( A299  and  (not A298) );
 a22663a <=( A266  and  a22662a );
 a22664a <=( a22663a  and  a22658a );
 a22668a <=( A167  and  (not A168) );
 a22669a <=( A169  and  a22668a );
 a22673a <=( A200  and  (not A199) );
 a22674a <=( (not A166)  and  a22673a );
 a22675a <=( a22674a  and  a22669a );
 a22679a <=( (not A266)  and  (not A233) );
 a22680a <=( (not A232)  and  a22679a );
 a22684a <=( A299  and  (not A298) );
 a22685a <=( (not A267)  and  a22684a );
 a22686a <=( a22685a  and  a22680a );
 a22690a <=( A167  and  (not A168) );
 a22691a <=( A169  and  a22690a );
 a22695a <=( A200  and  (not A199) );
 a22696a <=( (not A166)  and  a22695a );
 a22697a <=( a22696a  and  a22691a );
 a22701a <=( (not A265)  and  (not A233) );
 a22702a <=( (not A232)  and  a22701a );
 a22706a <=( A299  and  (not A298) );
 a22707a <=( (not A266)  and  a22706a );
 a22708a <=( a22707a  and  a22702a );
 a22712a <=( A167  and  (not A168) );
 a22713a <=( A169  and  a22712a );
 a22717a <=( (not A200)  and  A199 );
 a22718a <=( (not A166)  and  a22717a );
 a22719a <=( a22718a  and  a22713a );
 a22723a <=( (not A232)  and  A202 );
 a22724a <=( A201  and  a22723a );
 a22728a <=( (not A300)  and  (not A299) );
 a22729a <=( A233  and  a22728a );
 a22730a <=( a22729a  and  a22724a );
 a22734a <=( A167  and  (not A168) );
 a22735a <=( A169  and  a22734a );
 a22739a <=( (not A200)  and  A199 );
 a22740a <=( (not A166)  and  a22739a );
 a22741a <=( a22740a  and  a22735a );
 a22745a <=( (not A232)  and  A202 );
 a22746a <=( A201  and  a22745a );
 a22750a <=( A299  and  A298 );
 a22751a <=( A233  and  a22750a );
 a22752a <=( a22751a  and  a22746a );
 a22756a <=( A167  and  (not A168) );
 a22757a <=( A169  and  a22756a );
 a22761a <=( (not A200)  and  A199 );
 a22762a <=( (not A166)  and  a22761a );
 a22763a <=( a22762a  and  a22757a );
 a22767a <=( (not A232)  and  A202 );
 a22768a <=( A201  and  a22767a );
 a22772a <=( (not A299)  and  (not A298) );
 a22773a <=( A233  and  a22772a );
 a22774a <=( a22773a  and  a22768a );
 a22778a <=( A167  and  (not A168) );
 a22779a <=( A169  and  a22778a );
 a22783a <=( (not A200)  and  A199 );
 a22784a <=( (not A166)  and  a22783a );
 a22785a <=( a22784a  and  a22779a );
 a22789a <=( (not A232)  and  A202 );
 a22790a <=( A201  and  a22789a );
 a22794a <=( A266  and  (not A265) );
 a22795a <=( A233  and  a22794a );
 a22796a <=( a22795a  and  a22790a );
 a22800a <=( A167  and  (not A168) );
 a22801a <=( A169  and  a22800a );
 a22805a <=( (not A200)  and  A199 );
 a22806a <=( (not A166)  and  a22805a );
 a22807a <=( a22806a  and  a22801a );
 a22811a <=( (not A232)  and  A203 );
 a22812a <=( A201  and  a22811a );
 a22816a <=( (not A300)  and  (not A299) );
 a22817a <=( A233  and  a22816a );
 a22818a <=( a22817a  and  a22812a );
 a22822a <=( A167  and  (not A168) );
 a22823a <=( A169  and  a22822a );
 a22827a <=( (not A200)  and  A199 );
 a22828a <=( (not A166)  and  a22827a );
 a22829a <=( a22828a  and  a22823a );
 a22833a <=( (not A232)  and  A203 );
 a22834a <=( A201  and  a22833a );
 a22838a <=( A299  and  A298 );
 a22839a <=( A233  and  a22838a );
 a22840a <=( a22839a  and  a22834a );
 a22844a <=( A167  and  (not A168) );
 a22845a <=( A169  and  a22844a );
 a22849a <=( (not A200)  and  A199 );
 a22850a <=( (not A166)  and  a22849a );
 a22851a <=( a22850a  and  a22845a );
 a22855a <=( (not A232)  and  A203 );
 a22856a <=( A201  and  a22855a );
 a22860a <=( (not A299)  and  (not A298) );
 a22861a <=( A233  and  a22860a );
 a22862a <=( a22861a  and  a22856a );
 a22866a <=( A167  and  (not A168) );
 a22867a <=( A169  and  a22866a );
 a22871a <=( (not A200)  and  A199 );
 a22872a <=( (not A166)  and  a22871a );
 a22873a <=( a22872a  and  a22867a );
 a22877a <=( (not A232)  and  A203 );
 a22878a <=( A201  and  a22877a );
 a22882a <=( A266  and  (not A265) );
 a22883a <=( A233  and  a22882a );
 a22884a <=( a22883a  and  a22878a );
 a22888a <=( (not A167)  and  (not A168) );
 a22889a <=( A169  and  a22888a );
 a22893a <=( A200  and  (not A199) );
 a22894a <=( A166  and  a22893a );
 a22895a <=( a22894a  and  a22889a );
 a22899a <=( A265  and  A233 );
 a22900a <=( A232  and  a22899a );
 a22904a <=( A299  and  (not A298) );
 a22905a <=( (not A267)  and  a22904a );
 a22906a <=( a22905a  and  a22900a );
 a22910a <=( (not A167)  and  (not A168) );
 a22911a <=( A169  and  a22910a );
 a22915a <=( A200  and  (not A199) );
 a22916a <=( A166  and  a22915a );
 a22917a <=( a22916a  and  a22911a );
 a22921a <=( A265  and  A233 );
 a22922a <=( A232  and  a22921a );
 a22926a <=( A299  and  (not A298) );
 a22927a <=( A266  and  a22926a );
 a22928a <=( a22927a  and  a22922a );
 a22932a <=( (not A167)  and  (not A168) );
 a22933a <=( A169  and  a22932a );
 a22937a <=( A200  and  (not A199) );
 a22938a <=( A166  and  a22937a );
 a22939a <=( a22938a  and  a22933a );
 a22943a <=( (not A265)  and  A233 );
 a22944a <=( A232  and  a22943a );
 a22948a <=( A299  and  (not A298) );
 a22949a <=( (not A266)  and  a22948a );
 a22950a <=( a22949a  and  a22944a );
 a22954a <=( (not A167)  and  (not A168) );
 a22955a <=( A169  and  a22954a );
 a22959a <=( A200  and  (not A199) );
 a22960a <=( A166  and  a22959a );
 a22961a <=( a22960a  and  a22955a );
 a22965a <=( A265  and  A233 );
 a22966a <=( (not A232)  and  a22965a );
 a22970a <=( A268  and  A267 );
 a22971a <=( (not A266)  and  a22970a );
 a22972a <=( a22971a  and  a22966a );
 a22976a <=( (not A167)  and  (not A168) );
 a22977a <=( A169  and  a22976a );
 a22981a <=( A200  and  (not A199) );
 a22982a <=( A166  and  a22981a );
 a22983a <=( a22982a  and  a22977a );
 a22987a <=( A265  and  A233 );
 a22988a <=( (not A232)  and  a22987a );
 a22992a <=( A269  and  A267 );
 a22993a <=( (not A266)  and  a22992a );
 a22994a <=( a22993a  and  a22988a );
 a22998a <=( (not A167)  and  (not A168) );
 a22999a <=( A169  and  a22998a );
 a23003a <=( A200  and  (not A199) );
 a23004a <=( A166  and  a23003a );
 a23005a <=( a23004a  and  a22999a );
 a23009a <=( A265  and  (not A234) );
 a23010a <=( (not A233)  and  a23009a );
 a23014a <=( A299  and  (not A298) );
 a23015a <=( A266  and  a23014a );
 a23016a <=( a23015a  and  a23010a );
 a23020a <=( (not A167)  and  (not A168) );
 a23021a <=( A169  and  a23020a );
 a23025a <=( A200  and  (not A199) );
 a23026a <=( A166  and  a23025a );
 a23027a <=( a23026a  and  a23021a );
 a23031a <=( (not A266)  and  (not A234) );
 a23032a <=( (not A233)  and  a23031a );
 a23036a <=( A299  and  (not A298) );
 a23037a <=( (not A267)  and  a23036a );
 a23038a <=( a23037a  and  a23032a );
 a23042a <=( (not A167)  and  (not A168) );
 a23043a <=( A169  and  a23042a );
 a23047a <=( A200  and  (not A199) );
 a23048a <=( A166  and  a23047a );
 a23049a <=( a23048a  and  a23043a );
 a23053a <=( (not A265)  and  (not A234) );
 a23054a <=( (not A233)  and  a23053a );
 a23058a <=( A299  and  (not A298) );
 a23059a <=( (not A266)  and  a23058a );
 a23060a <=( a23059a  and  a23054a );
 a23064a <=( (not A167)  and  (not A168) );
 a23065a <=( A169  and  a23064a );
 a23069a <=( A200  and  (not A199) );
 a23070a <=( A166  and  a23069a );
 a23071a <=( a23070a  and  a23065a );
 a23075a <=( A234  and  (not A233) );
 a23076a <=( A232  and  a23075a );
 a23080a <=( (not A300)  and  A298 );
 a23081a <=( A235  and  a23080a );
 a23082a <=( a23081a  and  a23076a );
 a23086a <=( (not A167)  and  (not A168) );
 a23087a <=( A169  and  a23086a );
 a23091a <=( A200  and  (not A199) );
 a23092a <=( A166  and  a23091a );
 a23093a <=( a23092a  and  a23087a );
 a23097a <=( A234  and  (not A233) );
 a23098a <=( A232  and  a23097a );
 a23102a <=( A299  and  A298 );
 a23103a <=( A235  and  a23102a );
 a23104a <=( a23103a  and  a23098a );
 a23108a <=( (not A167)  and  (not A168) );
 a23109a <=( A169  and  a23108a );
 a23113a <=( A200  and  (not A199) );
 a23114a <=( A166  and  a23113a );
 a23115a <=( a23114a  and  a23109a );
 a23119a <=( A234  and  (not A233) );
 a23120a <=( A232  and  a23119a );
 a23124a <=( (not A299)  and  (not A298) );
 a23125a <=( A235  and  a23124a );
 a23126a <=( a23125a  and  a23120a );
 a23130a <=( (not A167)  and  (not A168) );
 a23131a <=( A169  and  a23130a );
 a23135a <=( A200  and  (not A199) );
 a23136a <=( A166  and  a23135a );
 a23137a <=( a23136a  and  a23131a );
 a23141a <=( A234  and  (not A233) );
 a23142a <=( A232  and  a23141a );
 a23146a <=( A266  and  (not A265) );
 a23147a <=( A235  and  a23146a );
 a23148a <=( a23147a  and  a23142a );
 a23152a <=( (not A167)  and  (not A168) );
 a23153a <=( A169  and  a23152a );
 a23157a <=( A200  and  (not A199) );
 a23158a <=( A166  and  a23157a );
 a23159a <=( a23158a  and  a23153a );
 a23163a <=( A234  and  (not A233) );
 a23164a <=( A232  and  a23163a );
 a23168a <=( (not A300)  and  A298 );
 a23169a <=( A236  and  a23168a );
 a23170a <=( a23169a  and  a23164a );
 a23174a <=( (not A167)  and  (not A168) );
 a23175a <=( A169  and  a23174a );
 a23179a <=( A200  and  (not A199) );
 a23180a <=( A166  and  a23179a );
 a23181a <=( a23180a  and  a23175a );
 a23185a <=( A234  and  (not A233) );
 a23186a <=( A232  and  a23185a );
 a23190a <=( A299  and  A298 );
 a23191a <=( A236  and  a23190a );
 a23192a <=( a23191a  and  a23186a );
 a23196a <=( (not A167)  and  (not A168) );
 a23197a <=( A169  and  a23196a );
 a23201a <=( A200  and  (not A199) );
 a23202a <=( A166  and  a23201a );
 a23203a <=( a23202a  and  a23197a );
 a23207a <=( A234  and  (not A233) );
 a23208a <=( A232  and  a23207a );
 a23212a <=( (not A299)  and  (not A298) );
 a23213a <=( A236  and  a23212a );
 a23214a <=( a23213a  and  a23208a );
 a23218a <=( (not A167)  and  (not A168) );
 a23219a <=( A169  and  a23218a );
 a23223a <=( A200  and  (not A199) );
 a23224a <=( A166  and  a23223a );
 a23225a <=( a23224a  and  a23219a );
 a23229a <=( A234  and  (not A233) );
 a23230a <=( A232  and  a23229a );
 a23234a <=( A266  and  (not A265) );
 a23235a <=( A236  and  a23234a );
 a23236a <=( a23235a  and  a23230a );
 a23240a <=( (not A167)  and  (not A168) );
 a23241a <=( A169  and  a23240a );
 a23245a <=( A200  and  (not A199) );
 a23246a <=( A166  and  a23245a );
 a23247a <=( a23246a  and  a23241a );
 a23251a <=( A265  and  (not A233) );
 a23252a <=( (not A232)  and  a23251a );
 a23256a <=( A299  and  (not A298) );
 a23257a <=( A266  and  a23256a );
 a23258a <=( a23257a  and  a23252a );
 a23262a <=( (not A167)  and  (not A168) );
 a23263a <=( A169  and  a23262a );
 a23267a <=( A200  and  (not A199) );
 a23268a <=( A166  and  a23267a );
 a23269a <=( a23268a  and  a23263a );
 a23273a <=( (not A266)  and  (not A233) );
 a23274a <=( (not A232)  and  a23273a );
 a23278a <=( A299  and  (not A298) );
 a23279a <=( (not A267)  and  a23278a );
 a23280a <=( a23279a  and  a23274a );
 a23284a <=( (not A167)  and  (not A168) );
 a23285a <=( A169  and  a23284a );
 a23289a <=( A200  and  (not A199) );
 a23290a <=( A166  and  a23289a );
 a23291a <=( a23290a  and  a23285a );
 a23295a <=( (not A265)  and  (not A233) );
 a23296a <=( (not A232)  and  a23295a );
 a23300a <=( A299  and  (not A298) );
 a23301a <=( (not A266)  and  a23300a );
 a23302a <=( a23301a  and  a23296a );
 a23306a <=( (not A167)  and  (not A168) );
 a23307a <=( A169  and  a23306a );
 a23311a <=( (not A200)  and  A199 );
 a23312a <=( A166  and  a23311a );
 a23313a <=( a23312a  and  a23307a );
 a23317a <=( (not A232)  and  A202 );
 a23318a <=( A201  and  a23317a );
 a23322a <=( (not A300)  and  (not A299) );
 a23323a <=( A233  and  a23322a );
 a23324a <=( a23323a  and  a23318a );
 a23328a <=( (not A167)  and  (not A168) );
 a23329a <=( A169  and  a23328a );
 a23333a <=( (not A200)  and  A199 );
 a23334a <=( A166  and  a23333a );
 a23335a <=( a23334a  and  a23329a );
 a23339a <=( (not A232)  and  A202 );
 a23340a <=( A201  and  a23339a );
 a23344a <=( A299  and  A298 );
 a23345a <=( A233  and  a23344a );
 a23346a <=( a23345a  and  a23340a );
 a23350a <=( (not A167)  and  (not A168) );
 a23351a <=( A169  and  a23350a );
 a23355a <=( (not A200)  and  A199 );
 a23356a <=( A166  and  a23355a );
 a23357a <=( a23356a  and  a23351a );
 a23361a <=( (not A232)  and  A202 );
 a23362a <=( A201  and  a23361a );
 a23366a <=( (not A299)  and  (not A298) );
 a23367a <=( A233  and  a23366a );
 a23368a <=( a23367a  and  a23362a );
 a23372a <=( (not A167)  and  (not A168) );
 a23373a <=( A169  and  a23372a );
 a23377a <=( (not A200)  and  A199 );
 a23378a <=( A166  and  a23377a );
 a23379a <=( a23378a  and  a23373a );
 a23383a <=( (not A232)  and  A202 );
 a23384a <=( A201  and  a23383a );
 a23388a <=( A266  and  (not A265) );
 a23389a <=( A233  and  a23388a );
 a23390a <=( a23389a  and  a23384a );
 a23394a <=( (not A167)  and  (not A168) );
 a23395a <=( A169  and  a23394a );
 a23399a <=( (not A200)  and  A199 );
 a23400a <=( A166  and  a23399a );
 a23401a <=( a23400a  and  a23395a );
 a23405a <=( (not A232)  and  A203 );
 a23406a <=( A201  and  a23405a );
 a23410a <=( (not A300)  and  (not A299) );
 a23411a <=( A233  and  a23410a );
 a23412a <=( a23411a  and  a23406a );
 a23416a <=( (not A167)  and  (not A168) );
 a23417a <=( A169  and  a23416a );
 a23421a <=( (not A200)  and  A199 );
 a23422a <=( A166  and  a23421a );
 a23423a <=( a23422a  and  a23417a );
 a23427a <=( (not A232)  and  A203 );
 a23428a <=( A201  and  a23427a );
 a23432a <=( A299  and  A298 );
 a23433a <=( A233  and  a23432a );
 a23434a <=( a23433a  and  a23428a );
 a23438a <=( (not A167)  and  (not A168) );
 a23439a <=( A169  and  a23438a );
 a23443a <=( (not A200)  and  A199 );
 a23444a <=( A166  and  a23443a );
 a23445a <=( a23444a  and  a23439a );
 a23449a <=( (not A232)  and  A203 );
 a23450a <=( A201  and  a23449a );
 a23454a <=( (not A299)  and  (not A298) );
 a23455a <=( A233  and  a23454a );
 a23456a <=( a23455a  and  a23450a );
 a23460a <=( (not A167)  and  (not A168) );
 a23461a <=( A169  and  a23460a );
 a23465a <=( (not A200)  and  A199 );
 a23466a <=( A166  and  a23465a );
 a23467a <=( a23466a  and  a23461a );
 a23471a <=( (not A232)  and  A203 );
 a23472a <=( A201  and  a23471a );
 a23476a <=( A266  and  (not A265) );
 a23477a <=( A233  and  a23476a );
 a23478a <=( a23477a  and  a23472a );
 a23482a <=( (not A168)  and  A169 );
 a23483a <=( A170  and  a23482a );
 a23487a <=( A201  and  (not A200) );
 a23488a <=( A199  and  a23487a );
 a23489a <=( a23488a  and  a23483a );
 a23493a <=( A233  and  (not A232) );
 a23494a <=( A202  and  a23493a );
 a23498a <=( (not A302)  and  (not A301) );
 a23499a <=( (not A299)  and  a23498a );
 a23500a <=( a23499a  and  a23494a );
 a23504a <=( (not A168)  and  A169 );
 a23505a <=( A170  and  a23504a );
 a23509a <=( A201  and  (not A200) );
 a23510a <=( A199  and  a23509a );
 a23511a <=( a23510a  and  a23505a );
 a23515a <=( A233  and  (not A232) );
 a23516a <=( A203  and  a23515a );
 a23520a <=( (not A302)  and  (not A301) );
 a23521a <=( (not A299)  and  a23520a );
 a23522a <=( a23521a  and  a23516a );
 a23526a <=( A167  and  A169 );
 a23527a <=( (not A170)  and  a23526a );
 a23531a <=( A200  and  A199 );
 a23532a <=( A166  and  a23531a );
 a23533a <=( a23532a  and  a23527a );
 a23537a <=( A265  and  A233 );
 a23538a <=( A232  and  a23537a );
 a23542a <=( A299  and  (not A298) );
 a23543a <=( (not A267)  and  a23542a );
 a23544a <=( a23543a  and  a23538a );
 a23548a <=( A167  and  A169 );
 a23549a <=( (not A170)  and  a23548a );
 a23553a <=( A200  and  A199 );
 a23554a <=( A166  and  a23553a );
 a23555a <=( a23554a  and  a23549a );
 a23559a <=( A265  and  A233 );
 a23560a <=( A232  and  a23559a );
 a23564a <=( A299  and  (not A298) );
 a23565a <=( A266  and  a23564a );
 a23566a <=( a23565a  and  a23560a );
 a23570a <=( A167  and  A169 );
 a23571a <=( (not A170)  and  a23570a );
 a23575a <=( A200  and  A199 );
 a23576a <=( A166  and  a23575a );
 a23577a <=( a23576a  and  a23571a );
 a23581a <=( (not A265)  and  A233 );
 a23582a <=( A232  and  a23581a );
 a23586a <=( A299  and  (not A298) );
 a23587a <=( (not A266)  and  a23586a );
 a23588a <=( a23587a  and  a23582a );
 a23592a <=( A167  and  A169 );
 a23593a <=( (not A170)  and  a23592a );
 a23597a <=( A200  and  A199 );
 a23598a <=( A166  and  a23597a );
 a23599a <=( a23598a  and  a23593a );
 a23603a <=( A265  and  A233 );
 a23604a <=( (not A232)  and  a23603a );
 a23608a <=( A268  and  A267 );
 a23609a <=( (not A266)  and  a23608a );
 a23610a <=( a23609a  and  a23604a );
 a23614a <=( A167  and  A169 );
 a23615a <=( (not A170)  and  a23614a );
 a23619a <=( A200  and  A199 );
 a23620a <=( A166  and  a23619a );
 a23621a <=( a23620a  and  a23615a );
 a23625a <=( A265  and  A233 );
 a23626a <=( (not A232)  and  a23625a );
 a23630a <=( A269  and  A267 );
 a23631a <=( (not A266)  and  a23630a );
 a23632a <=( a23631a  and  a23626a );
 a23636a <=( A167  and  A169 );
 a23637a <=( (not A170)  and  a23636a );
 a23641a <=( A200  and  A199 );
 a23642a <=( A166  and  a23641a );
 a23643a <=( a23642a  and  a23637a );
 a23647a <=( A265  and  (not A234) );
 a23648a <=( (not A233)  and  a23647a );
 a23652a <=( A299  and  (not A298) );
 a23653a <=( A266  and  a23652a );
 a23654a <=( a23653a  and  a23648a );
 a23658a <=( A167  and  A169 );
 a23659a <=( (not A170)  and  a23658a );
 a23663a <=( A200  and  A199 );
 a23664a <=( A166  and  a23663a );
 a23665a <=( a23664a  and  a23659a );
 a23669a <=( (not A266)  and  (not A234) );
 a23670a <=( (not A233)  and  a23669a );
 a23674a <=( A299  and  (not A298) );
 a23675a <=( (not A267)  and  a23674a );
 a23676a <=( a23675a  and  a23670a );
 a23680a <=( A167  and  A169 );
 a23681a <=( (not A170)  and  a23680a );
 a23685a <=( A200  and  A199 );
 a23686a <=( A166  and  a23685a );
 a23687a <=( a23686a  and  a23681a );
 a23691a <=( (not A265)  and  (not A234) );
 a23692a <=( (not A233)  and  a23691a );
 a23696a <=( A299  and  (not A298) );
 a23697a <=( (not A266)  and  a23696a );
 a23698a <=( a23697a  and  a23692a );
 a23702a <=( A167  and  A169 );
 a23703a <=( (not A170)  and  a23702a );
 a23707a <=( A200  and  A199 );
 a23708a <=( A166  and  a23707a );
 a23709a <=( a23708a  and  a23703a );
 a23713a <=( A234  and  (not A233) );
 a23714a <=( A232  and  a23713a );
 a23718a <=( (not A300)  and  A298 );
 a23719a <=( A235  and  a23718a );
 a23720a <=( a23719a  and  a23714a );
 a23724a <=( A167  and  A169 );
 a23725a <=( (not A170)  and  a23724a );
 a23729a <=( A200  and  A199 );
 a23730a <=( A166  and  a23729a );
 a23731a <=( a23730a  and  a23725a );
 a23735a <=( A234  and  (not A233) );
 a23736a <=( A232  and  a23735a );
 a23740a <=( A299  and  A298 );
 a23741a <=( A235  and  a23740a );
 a23742a <=( a23741a  and  a23736a );
 a23746a <=( A167  and  A169 );
 a23747a <=( (not A170)  and  a23746a );
 a23751a <=( A200  and  A199 );
 a23752a <=( A166  and  a23751a );
 a23753a <=( a23752a  and  a23747a );
 a23757a <=( A234  and  (not A233) );
 a23758a <=( A232  and  a23757a );
 a23762a <=( (not A299)  and  (not A298) );
 a23763a <=( A235  and  a23762a );
 a23764a <=( a23763a  and  a23758a );
 a23768a <=( A167  and  A169 );
 a23769a <=( (not A170)  and  a23768a );
 a23773a <=( A200  and  A199 );
 a23774a <=( A166  and  a23773a );
 a23775a <=( a23774a  and  a23769a );
 a23779a <=( A234  and  (not A233) );
 a23780a <=( A232  and  a23779a );
 a23784a <=( A266  and  (not A265) );
 a23785a <=( A235  and  a23784a );
 a23786a <=( a23785a  and  a23780a );
 a23790a <=( A167  and  A169 );
 a23791a <=( (not A170)  and  a23790a );
 a23795a <=( A200  and  A199 );
 a23796a <=( A166  and  a23795a );
 a23797a <=( a23796a  and  a23791a );
 a23801a <=( A234  and  (not A233) );
 a23802a <=( A232  and  a23801a );
 a23806a <=( (not A300)  and  A298 );
 a23807a <=( A236  and  a23806a );
 a23808a <=( a23807a  and  a23802a );
 a23812a <=( A167  and  A169 );
 a23813a <=( (not A170)  and  a23812a );
 a23817a <=( A200  and  A199 );
 a23818a <=( A166  and  a23817a );
 a23819a <=( a23818a  and  a23813a );
 a23823a <=( A234  and  (not A233) );
 a23824a <=( A232  and  a23823a );
 a23828a <=( A299  and  A298 );
 a23829a <=( A236  and  a23828a );
 a23830a <=( a23829a  and  a23824a );
 a23834a <=( A167  and  A169 );
 a23835a <=( (not A170)  and  a23834a );
 a23839a <=( A200  and  A199 );
 a23840a <=( A166  and  a23839a );
 a23841a <=( a23840a  and  a23835a );
 a23845a <=( A234  and  (not A233) );
 a23846a <=( A232  and  a23845a );
 a23850a <=( (not A299)  and  (not A298) );
 a23851a <=( A236  and  a23850a );
 a23852a <=( a23851a  and  a23846a );
 a23856a <=( A167  and  A169 );
 a23857a <=( (not A170)  and  a23856a );
 a23861a <=( A200  and  A199 );
 a23862a <=( A166  and  a23861a );
 a23863a <=( a23862a  and  a23857a );
 a23867a <=( A234  and  (not A233) );
 a23868a <=( A232  and  a23867a );
 a23872a <=( A266  and  (not A265) );
 a23873a <=( A236  and  a23872a );
 a23874a <=( a23873a  and  a23868a );
 a23878a <=( A167  and  A169 );
 a23879a <=( (not A170)  and  a23878a );
 a23883a <=( A200  and  A199 );
 a23884a <=( A166  and  a23883a );
 a23885a <=( a23884a  and  a23879a );
 a23889a <=( A265  and  (not A233) );
 a23890a <=( (not A232)  and  a23889a );
 a23894a <=( A299  and  (not A298) );
 a23895a <=( A266  and  a23894a );
 a23896a <=( a23895a  and  a23890a );
 a23900a <=( A167  and  A169 );
 a23901a <=( (not A170)  and  a23900a );
 a23905a <=( A200  and  A199 );
 a23906a <=( A166  and  a23905a );
 a23907a <=( a23906a  and  a23901a );
 a23911a <=( (not A266)  and  (not A233) );
 a23912a <=( (not A232)  and  a23911a );
 a23916a <=( A299  and  (not A298) );
 a23917a <=( (not A267)  and  a23916a );
 a23918a <=( a23917a  and  a23912a );
 a23922a <=( A167  and  A169 );
 a23923a <=( (not A170)  and  a23922a );
 a23927a <=( A200  and  A199 );
 a23928a <=( A166  and  a23927a );
 a23929a <=( a23928a  and  a23923a );
 a23933a <=( (not A265)  and  (not A233) );
 a23934a <=( (not A232)  and  a23933a );
 a23938a <=( A299  and  (not A298) );
 a23939a <=( (not A266)  and  a23938a );
 a23940a <=( a23939a  and  a23934a );
 a23944a <=( A167  and  A169 );
 a23945a <=( (not A170)  and  a23944a );
 a23949a <=( (not A202)  and  (not A200) );
 a23950a <=( A166  and  a23949a );
 a23951a <=( a23950a  and  a23945a );
 a23955a <=( A233  and  (not A232) );
 a23956a <=( (not A203)  and  a23955a );
 a23960a <=( (not A302)  and  (not A301) );
 a23961a <=( (not A299)  and  a23960a );
 a23962a <=( a23961a  and  a23956a );
 a23966a <=( A167  and  A169 );
 a23967a <=( (not A170)  and  a23966a );
 a23971a <=( (not A201)  and  (not A200) );
 a23972a <=( A166  and  a23971a );
 a23973a <=( a23972a  and  a23967a );
 a23977a <=( A265  and  A233 );
 a23978a <=( A232  and  a23977a );
 a23982a <=( A299  and  (not A298) );
 a23983a <=( (not A267)  and  a23982a );
 a23984a <=( a23983a  and  a23978a );
 a23988a <=( A167  and  A169 );
 a23989a <=( (not A170)  and  a23988a );
 a23993a <=( (not A201)  and  (not A200) );
 a23994a <=( A166  and  a23993a );
 a23995a <=( a23994a  and  a23989a );
 a23999a <=( A265  and  A233 );
 a24000a <=( A232  and  a23999a );
 a24004a <=( A299  and  (not A298) );
 a24005a <=( A266  and  a24004a );
 a24006a <=( a24005a  and  a24000a );
 a24010a <=( A167  and  A169 );
 a24011a <=( (not A170)  and  a24010a );
 a24015a <=( (not A201)  and  (not A200) );
 a24016a <=( A166  and  a24015a );
 a24017a <=( a24016a  and  a24011a );
 a24021a <=( (not A265)  and  A233 );
 a24022a <=( A232  and  a24021a );
 a24026a <=( A299  and  (not A298) );
 a24027a <=( (not A266)  and  a24026a );
 a24028a <=( a24027a  and  a24022a );
 a24032a <=( A167  and  A169 );
 a24033a <=( (not A170)  and  a24032a );
 a24037a <=( (not A201)  and  (not A200) );
 a24038a <=( A166  and  a24037a );
 a24039a <=( a24038a  and  a24033a );
 a24043a <=( A265  and  A233 );
 a24044a <=( (not A232)  and  a24043a );
 a24048a <=( A268  and  A267 );
 a24049a <=( (not A266)  and  a24048a );
 a24050a <=( a24049a  and  a24044a );
 a24054a <=( A167  and  A169 );
 a24055a <=( (not A170)  and  a24054a );
 a24059a <=( (not A201)  and  (not A200) );
 a24060a <=( A166  and  a24059a );
 a24061a <=( a24060a  and  a24055a );
 a24065a <=( A265  and  A233 );
 a24066a <=( (not A232)  and  a24065a );
 a24070a <=( A269  and  A267 );
 a24071a <=( (not A266)  and  a24070a );
 a24072a <=( a24071a  and  a24066a );
 a24076a <=( A167  and  A169 );
 a24077a <=( (not A170)  and  a24076a );
 a24081a <=( (not A201)  and  (not A200) );
 a24082a <=( A166  and  a24081a );
 a24083a <=( a24082a  and  a24077a );
 a24087a <=( A265  and  (not A234) );
 a24088a <=( (not A233)  and  a24087a );
 a24092a <=( A299  and  (not A298) );
 a24093a <=( A266  and  a24092a );
 a24094a <=( a24093a  and  a24088a );
 a24098a <=( A167  and  A169 );
 a24099a <=( (not A170)  and  a24098a );
 a24103a <=( (not A201)  and  (not A200) );
 a24104a <=( A166  and  a24103a );
 a24105a <=( a24104a  and  a24099a );
 a24109a <=( (not A266)  and  (not A234) );
 a24110a <=( (not A233)  and  a24109a );
 a24114a <=( A299  and  (not A298) );
 a24115a <=( (not A267)  and  a24114a );
 a24116a <=( a24115a  and  a24110a );
 a24120a <=( A167  and  A169 );
 a24121a <=( (not A170)  and  a24120a );
 a24125a <=( (not A201)  and  (not A200) );
 a24126a <=( A166  and  a24125a );
 a24127a <=( a24126a  and  a24121a );
 a24131a <=( (not A265)  and  (not A234) );
 a24132a <=( (not A233)  and  a24131a );
 a24136a <=( A299  and  (not A298) );
 a24137a <=( (not A266)  and  a24136a );
 a24138a <=( a24137a  and  a24132a );
 a24142a <=( A167  and  A169 );
 a24143a <=( (not A170)  and  a24142a );
 a24147a <=( (not A201)  and  (not A200) );
 a24148a <=( A166  and  a24147a );
 a24149a <=( a24148a  and  a24143a );
 a24153a <=( A234  and  (not A233) );
 a24154a <=( A232  and  a24153a );
 a24158a <=( (not A300)  and  A298 );
 a24159a <=( A235  and  a24158a );
 a24160a <=( a24159a  and  a24154a );
 a24164a <=( A167  and  A169 );
 a24165a <=( (not A170)  and  a24164a );
 a24169a <=( (not A201)  and  (not A200) );
 a24170a <=( A166  and  a24169a );
 a24171a <=( a24170a  and  a24165a );
 a24175a <=( A234  and  (not A233) );
 a24176a <=( A232  and  a24175a );
 a24180a <=( A299  and  A298 );
 a24181a <=( A235  and  a24180a );
 a24182a <=( a24181a  and  a24176a );
 a24186a <=( A167  and  A169 );
 a24187a <=( (not A170)  and  a24186a );
 a24191a <=( (not A201)  and  (not A200) );
 a24192a <=( A166  and  a24191a );
 a24193a <=( a24192a  and  a24187a );
 a24197a <=( A234  and  (not A233) );
 a24198a <=( A232  and  a24197a );
 a24202a <=( (not A299)  and  (not A298) );
 a24203a <=( A235  and  a24202a );
 a24204a <=( a24203a  and  a24198a );
 a24208a <=( A167  and  A169 );
 a24209a <=( (not A170)  and  a24208a );
 a24213a <=( (not A201)  and  (not A200) );
 a24214a <=( A166  and  a24213a );
 a24215a <=( a24214a  and  a24209a );
 a24219a <=( A234  and  (not A233) );
 a24220a <=( A232  and  a24219a );
 a24224a <=( A266  and  (not A265) );
 a24225a <=( A235  and  a24224a );
 a24226a <=( a24225a  and  a24220a );
 a24230a <=( A167  and  A169 );
 a24231a <=( (not A170)  and  a24230a );
 a24235a <=( (not A201)  and  (not A200) );
 a24236a <=( A166  and  a24235a );
 a24237a <=( a24236a  and  a24231a );
 a24241a <=( A234  and  (not A233) );
 a24242a <=( A232  and  a24241a );
 a24246a <=( (not A300)  and  A298 );
 a24247a <=( A236  and  a24246a );
 a24248a <=( a24247a  and  a24242a );
 a24252a <=( A167  and  A169 );
 a24253a <=( (not A170)  and  a24252a );
 a24257a <=( (not A201)  and  (not A200) );
 a24258a <=( A166  and  a24257a );
 a24259a <=( a24258a  and  a24253a );
 a24263a <=( A234  and  (not A233) );
 a24264a <=( A232  and  a24263a );
 a24268a <=( A299  and  A298 );
 a24269a <=( A236  and  a24268a );
 a24270a <=( a24269a  and  a24264a );
 a24274a <=( A167  and  A169 );
 a24275a <=( (not A170)  and  a24274a );
 a24279a <=( (not A201)  and  (not A200) );
 a24280a <=( A166  and  a24279a );
 a24281a <=( a24280a  and  a24275a );
 a24285a <=( A234  and  (not A233) );
 a24286a <=( A232  and  a24285a );
 a24290a <=( (not A299)  and  (not A298) );
 a24291a <=( A236  and  a24290a );
 a24292a <=( a24291a  and  a24286a );
 a24296a <=( A167  and  A169 );
 a24297a <=( (not A170)  and  a24296a );
 a24301a <=( (not A201)  and  (not A200) );
 a24302a <=( A166  and  a24301a );
 a24303a <=( a24302a  and  a24297a );
 a24307a <=( A234  and  (not A233) );
 a24308a <=( A232  and  a24307a );
 a24312a <=( A266  and  (not A265) );
 a24313a <=( A236  and  a24312a );
 a24314a <=( a24313a  and  a24308a );
 a24318a <=( A167  and  A169 );
 a24319a <=( (not A170)  and  a24318a );
 a24323a <=( (not A201)  and  (not A200) );
 a24324a <=( A166  and  a24323a );
 a24325a <=( a24324a  and  a24319a );
 a24329a <=( A265  and  (not A233) );
 a24330a <=( (not A232)  and  a24329a );
 a24334a <=( A299  and  (not A298) );
 a24335a <=( A266  and  a24334a );
 a24336a <=( a24335a  and  a24330a );
 a24340a <=( A167  and  A169 );
 a24341a <=( (not A170)  and  a24340a );
 a24345a <=( (not A201)  and  (not A200) );
 a24346a <=( A166  and  a24345a );
 a24347a <=( a24346a  and  a24341a );
 a24351a <=( (not A266)  and  (not A233) );
 a24352a <=( (not A232)  and  a24351a );
 a24356a <=( A299  and  (not A298) );
 a24357a <=( (not A267)  and  a24356a );
 a24358a <=( a24357a  and  a24352a );
 a24362a <=( A167  and  A169 );
 a24363a <=( (not A170)  and  a24362a );
 a24367a <=( (not A201)  and  (not A200) );
 a24368a <=( A166  and  a24367a );
 a24369a <=( a24368a  and  a24363a );
 a24373a <=( (not A265)  and  (not A233) );
 a24374a <=( (not A232)  and  a24373a );
 a24378a <=( A299  and  (not A298) );
 a24379a <=( (not A266)  and  a24378a );
 a24380a <=( a24379a  and  a24374a );
 a24384a <=( A167  and  A169 );
 a24385a <=( (not A170)  and  a24384a );
 a24389a <=( (not A200)  and  (not A199) );
 a24390a <=( A166  and  a24389a );
 a24391a <=( a24390a  and  a24385a );
 a24395a <=( A265  and  A233 );
 a24396a <=( A232  and  a24395a );
 a24400a <=( A299  and  (not A298) );
 a24401a <=( (not A267)  and  a24400a );
 a24402a <=( a24401a  and  a24396a );
 a24406a <=( A167  and  A169 );
 a24407a <=( (not A170)  and  a24406a );
 a24411a <=( (not A200)  and  (not A199) );
 a24412a <=( A166  and  a24411a );
 a24413a <=( a24412a  and  a24407a );
 a24417a <=( A265  and  A233 );
 a24418a <=( A232  and  a24417a );
 a24422a <=( A299  and  (not A298) );
 a24423a <=( A266  and  a24422a );
 a24424a <=( a24423a  and  a24418a );
 a24428a <=( A167  and  A169 );
 a24429a <=( (not A170)  and  a24428a );
 a24433a <=( (not A200)  and  (not A199) );
 a24434a <=( A166  and  a24433a );
 a24435a <=( a24434a  and  a24429a );
 a24439a <=( (not A265)  and  A233 );
 a24440a <=( A232  and  a24439a );
 a24444a <=( A299  and  (not A298) );
 a24445a <=( (not A266)  and  a24444a );
 a24446a <=( a24445a  and  a24440a );
 a24450a <=( A167  and  A169 );
 a24451a <=( (not A170)  and  a24450a );
 a24455a <=( (not A200)  and  (not A199) );
 a24456a <=( A166  and  a24455a );
 a24457a <=( a24456a  and  a24451a );
 a24461a <=( A265  and  A233 );
 a24462a <=( (not A232)  and  a24461a );
 a24466a <=( A268  and  A267 );
 a24467a <=( (not A266)  and  a24466a );
 a24468a <=( a24467a  and  a24462a );
 a24472a <=( A167  and  A169 );
 a24473a <=( (not A170)  and  a24472a );
 a24477a <=( (not A200)  and  (not A199) );
 a24478a <=( A166  and  a24477a );
 a24479a <=( a24478a  and  a24473a );
 a24483a <=( A265  and  A233 );
 a24484a <=( (not A232)  and  a24483a );
 a24488a <=( A269  and  A267 );
 a24489a <=( (not A266)  and  a24488a );
 a24490a <=( a24489a  and  a24484a );
 a24494a <=( A167  and  A169 );
 a24495a <=( (not A170)  and  a24494a );
 a24499a <=( (not A200)  and  (not A199) );
 a24500a <=( A166  and  a24499a );
 a24501a <=( a24500a  and  a24495a );
 a24505a <=( A265  and  (not A234) );
 a24506a <=( (not A233)  and  a24505a );
 a24510a <=( A299  and  (not A298) );
 a24511a <=( A266  and  a24510a );
 a24512a <=( a24511a  and  a24506a );
 a24516a <=( A167  and  A169 );
 a24517a <=( (not A170)  and  a24516a );
 a24521a <=( (not A200)  and  (not A199) );
 a24522a <=( A166  and  a24521a );
 a24523a <=( a24522a  and  a24517a );
 a24527a <=( (not A266)  and  (not A234) );
 a24528a <=( (not A233)  and  a24527a );
 a24532a <=( A299  and  (not A298) );
 a24533a <=( (not A267)  and  a24532a );
 a24534a <=( a24533a  and  a24528a );
 a24538a <=( A167  and  A169 );
 a24539a <=( (not A170)  and  a24538a );
 a24543a <=( (not A200)  and  (not A199) );
 a24544a <=( A166  and  a24543a );
 a24545a <=( a24544a  and  a24539a );
 a24549a <=( (not A265)  and  (not A234) );
 a24550a <=( (not A233)  and  a24549a );
 a24554a <=( A299  and  (not A298) );
 a24555a <=( (not A266)  and  a24554a );
 a24556a <=( a24555a  and  a24550a );
 a24560a <=( A167  and  A169 );
 a24561a <=( (not A170)  and  a24560a );
 a24565a <=( (not A200)  and  (not A199) );
 a24566a <=( A166  and  a24565a );
 a24567a <=( a24566a  and  a24561a );
 a24571a <=( A234  and  (not A233) );
 a24572a <=( A232  and  a24571a );
 a24576a <=( (not A300)  and  A298 );
 a24577a <=( A235  and  a24576a );
 a24578a <=( a24577a  and  a24572a );
 a24582a <=( A167  and  A169 );
 a24583a <=( (not A170)  and  a24582a );
 a24587a <=( (not A200)  and  (not A199) );
 a24588a <=( A166  and  a24587a );
 a24589a <=( a24588a  and  a24583a );
 a24593a <=( A234  and  (not A233) );
 a24594a <=( A232  and  a24593a );
 a24598a <=( A299  and  A298 );
 a24599a <=( A235  and  a24598a );
 a24600a <=( a24599a  and  a24594a );
 a24604a <=( A167  and  A169 );
 a24605a <=( (not A170)  and  a24604a );
 a24609a <=( (not A200)  and  (not A199) );
 a24610a <=( A166  and  a24609a );
 a24611a <=( a24610a  and  a24605a );
 a24615a <=( A234  and  (not A233) );
 a24616a <=( A232  and  a24615a );
 a24620a <=( (not A299)  and  (not A298) );
 a24621a <=( A235  and  a24620a );
 a24622a <=( a24621a  and  a24616a );
 a24626a <=( A167  and  A169 );
 a24627a <=( (not A170)  and  a24626a );
 a24631a <=( (not A200)  and  (not A199) );
 a24632a <=( A166  and  a24631a );
 a24633a <=( a24632a  and  a24627a );
 a24637a <=( A234  and  (not A233) );
 a24638a <=( A232  and  a24637a );
 a24642a <=( A266  and  (not A265) );
 a24643a <=( A235  and  a24642a );
 a24644a <=( a24643a  and  a24638a );
 a24648a <=( A167  and  A169 );
 a24649a <=( (not A170)  and  a24648a );
 a24653a <=( (not A200)  and  (not A199) );
 a24654a <=( A166  and  a24653a );
 a24655a <=( a24654a  and  a24649a );
 a24659a <=( A234  and  (not A233) );
 a24660a <=( A232  and  a24659a );
 a24664a <=( (not A300)  and  A298 );
 a24665a <=( A236  and  a24664a );
 a24666a <=( a24665a  and  a24660a );
 a24670a <=( A167  and  A169 );
 a24671a <=( (not A170)  and  a24670a );
 a24675a <=( (not A200)  and  (not A199) );
 a24676a <=( A166  and  a24675a );
 a24677a <=( a24676a  and  a24671a );
 a24681a <=( A234  and  (not A233) );
 a24682a <=( A232  and  a24681a );
 a24686a <=( A299  and  A298 );
 a24687a <=( A236  and  a24686a );
 a24688a <=( a24687a  and  a24682a );
 a24692a <=( A167  and  A169 );
 a24693a <=( (not A170)  and  a24692a );
 a24697a <=( (not A200)  and  (not A199) );
 a24698a <=( A166  and  a24697a );
 a24699a <=( a24698a  and  a24693a );
 a24703a <=( A234  and  (not A233) );
 a24704a <=( A232  and  a24703a );
 a24708a <=( (not A299)  and  (not A298) );
 a24709a <=( A236  and  a24708a );
 a24710a <=( a24709a  and  a24704a );
 a24714a <=( A167  and  A169 );
 a24715a <=( (not A170)  and  a24714a );
 a24719a <=( (not A200)  and  (not A199) );
 a24720a <=( A166  and  a24719a );
 a24721a <=( a24720a  and  a24715a );
 a24725a <=( A234  and  (not A233) );
 a24726a <=( A232  and  a24725a );
 a24730a <=( A266  and  (not A265) );
 a24731a <=( A236  and  a24730a );
 a24732a <=( a24731a  and  a24726a );
 a24736a <=( A167  and  A169 );
 a24737a <=( (not A170)  and  a24736a );
 a24741a <=( (not A200)  and  (not A199) );
 a24742a <=( A166  and  a24741a );
 a24743a <=( a24742a  and  a24737a );
 a24747a <=( A265  and  (not A233) );
 a24748a <=( (not A232)  and  a24747a );
 a24752a <=( A299  and  (not A298) );
 a24753a <=( A266  and  a24752a );
 a24754a <=( a24753a  and  a24748a );
 a24758a <=( A167  and  A169 );
 a24759a <=( (not A170)  and  a24758a );
 a24763a <=( (not A200)  and  (not A199) );
 a24764a <=( A166  and  a24763a );
 a24765a <=( a24764a  and  a24759a );
 a24769a <=( (not A266)  and  (not A233) );
 a24770a <=( (not A232)  and  a24769a );
 a24774a <=( A299  and  (not A298) );
 a24775a <=( (not A267)  and  a24774a );
 a24776a <=( a24775a  and  a24770a );
 a24780a <=( A167  and  A169 );
 a24781a <=( (not A170)  and  a24780a );
 a24785a <=( (not A200)  and  (not A199) );
 a24786a <=( A166  and  a24785a );
 a24787a <=( a24786a  and  a24781a );
 a24791a <=( (not A265)  and  (not A233) );
 a24792a <=( (not A232)  and  a24791a );
 a24796a <=( A299  and  (not A298) );
 a24797a <=( (not A266)  and  a24796a );
 a24798a <=( a24797a  and  a24792a );
 a24802a <=( (not A167)  and  A169 );
 a24803a <=( (not A170)  and  a24802a );
 a24807a <=( A200  and  A199 );
 a24808a <=( (not A166)  and  a24807a );
 a24809a <=( a24808a  and  a24803a );
 a24813a <=( A265  and  A233 );
 a24814a <=( A232  and  a24813a );
 a24818a <=( A299  and  (not A298) );
 a24819a <=( (not A267)  and  a24818a );
 a24820a <=( a24819a  and  a24814a );
 a24824a <=( (not A167)  and  A169 );
 a24825a <=( (not A170)  and  a24824a );
 a24829a <=( A200  and  A199 );
 a24830a <=( (not A166)  and  a24829a );
 a24831a <=( a24830a  and  a24825a );
 a24835a <=( A265  and  A233 );
 a24836a <=( A232  and  a24835a );
 a24840a <=( A299  and  (not A298) );
 a24841a <=( A266  and  a24840a );
 a24842a <=( a24841a  and  a24836a );
 a24846a <=( (not A167)  and  A169 );
 a24847a <=( (not A170)  and  a24846a );
 a24851a <=( A200  and  A199 );
 a24852a <=( (not A166)  and  a24851a );
 a24853a <=( a24852a  and  a24847a );
 a24857a <=( (not A265)  and  A233 );
 a24858a <=( A232  and  a24857a );
 a24862a <=( A299  and  (not A298) );
 a24863a <=( (not A266)  and  a24862a );
 a24864a <=( a24863a  and  a24858a );
 a24868a <=( (not A167)  and  A169 );
 a24869a <=( (not A170)  and  a24868a );
 a24873a <=( A200  and  A199 );
 a24874a <=( (not A166)  and  a24873a );
 a24875a <=( a24874a  and  a24869a );
 a24879a <=( A265  and  A233 );
 a24880a <=( (not A232)  and  a24879a );
 a24884a <=( A268  and  A267 );
 a24885a <=( (not A266)  and  a24884a );
 a24886a <=( a24885a  and  a24880a );
 a24890a <=( (not A167)  and  A169 );
 a24891a <=( (not A170)  and  a24890a );
 a24895a <=( A200  and  A199 );
 a24896a <=( (not A166)  and  a24895a );
 a24897a <=( a24896a  and  a24891a );
 a24901a <=( A265  and  A233 );
 a24902a <=( (not A232)  and  a24901a );
 a24906a <=( A269  and  A267 );
 a24907a <=( (not A266)  and  a24906a );
 a24908a <=( a24907a  and  a24902a );
 a24912a <=( (not A167)  and  A169 );
 a24913a <=( (not A170)  and  a24912a );
 a24917a <=( A200  and  A199 );
 a24918a <=( (not A166)  and  a24917a );
 a24919a <=( a24918a  and  a24913a );
 a24923a <=( A265  and  (not A234) );
 a24924a <=( (not A233)  and  a24923a );
 a24928a <=( A299  and  (not A298) );
 a24929a <=( A266  and  a24928a );
 a24930a <=( a24929a  and  a24924a );
 a24934a <=( (not A167)  and  A169 );
 a24935a <=( (not A170)  and  a24934a );
 a24939a <=( A200  and  A199 );
 a24940a <=( (not A166)  and  a24939a );
 a24941a <=( a24940a  and  a24935a );
 a24945a <=( (not A266)  and  (not A234) );
 a24946a <=( (not A233)  and  a24945a );
 a24950a <=( A299  and  (not A298) );
 a24951a <=( (not A267)  and  a24950a );
 a24952a <=( a24951a  and  a24946a );
 a24956a <=( (not A167)  and  A169 );
 a24957a <=( (not A170)  and  a24956a );
 a24961a <=( A200  and  A199 );
 a24962a <=( (not A166)  and  a24961a );
 a24963a <=( a24962a  and  a24957a );
 a24967a <=( (not A265)  and  (not A234) );
 a24968a <=( (not A233)  and  a24967a );
 a24972a <=( A299  and  (not A298) );
 a24973a <=( (not A266)  and  a24972a );
 a24974a <=( a24973a  and  a24968a );
 a24978a <=( (not A167)  and  A169 );
 a24979a <=( (not A170)  and  a24978a );
 a24983a <=( A200  and  A199 );
 a24984a <=( (not A166)  and  a24983a );
 a24985a <=( a24984a  and  a24979a );
 a24989a <=( A234  and  (not A233) );
 a24990a <=( A232  and  a24989a );
 a24994a <=( (not A300)  and  A298 );
 a24995a <=( A235  and  a24994a );
 a24996a <=( a24995a  and  a24990a );
 a25000a <=( (not A167)  and  A169 );
 a25001a <=( (not A170)  and  a25000a );
 a25005a <=( A200  and  A199 );
 a25006a <=( (not A166)  and  a25005a );
 a25007a <=( a25006a  and  a25001a );
 a25011a <=( A234  and  (not A233) );
 a25012a <=( A232  and  a25011a );
 a25016a <=( A299  and  A298 );
 a25017a <=( A235  and  a25016a );
 a25018a <=( a25017a  and  a25012a );
 a25022a <=( (not A167)  and  A169 );
 a25023a <=( (not A170)  and  a25022a );
 a25027a <=( A200  and  A199 );
 a25028a <=( (not A166)  and  a25027a );
 a25029a <=( a25028a  and  a25023a );
 a25033a <=( A234  and  (not A233) );
 a25034a <=( A232  and  a25033a );
 a25038a <=( (not A299)  and  (not A298) );
 a25039a <=( A235  and  a25038a );
 a25040a <=( a25039a  and  a25034a );
 a25044a <=( (not A167)  and  A169 );
 a25045a <=( (not A170)  and  a25044a );
 a25049a <=( A200  and  A199 );
 a25050a <=( (not A166)  and  a25049a );
 a25051a <=( a25050a  and  a25045a );
 a25055a <=( A234  and  (not A233) );
 a25056a <=( A232  and  a25055a );
 a25060a <=( A266  and  (not A265) );
 a25061a <=( A235  and  a25060a );
 a25062a <=( a25061a  and  a25056a );
 a25066a <=( (not A167)  and  A169 );
 a25067a <=( (not A170)  and  a25066a );
 a25071a <=( A200  and  A199 );
 a25072a <=( (not A166)  and  a25071a );
 a25073a <=( a25072a  and  a25067a );
 a25077a <=( A234  and  (not A233) );
 a25078a <=( A232  and  a25077a );
 a25082a <=( (not A300)  and  A298 );
 a25083a <=( A236  and  a25082a );
 a25084a <=( a25083a  and  a25078a );
 a25088a <=( (not A167)  and  A169 );
 a25089a <=( (not A170)  and  a25088a );
 a25093a <=( A200  and  A199 );
 a25094a <=( (not A166)  and  a25093a );
 a25095a <=( a25094a  and  a25089a );
 a25099a <=( A234  and  (not A233) );
 a25100a <=( A232  and  a25099a );
 a25104a <=( A299  and  A298 );
 a25105a <=( A236  and  a25104a );
 a25106a <=( a25105a  and  a25100a );
 a25110a <=( (not A167)  and  A169 );
 a25111a <=( (not A170)  and  a25110a );
 a25115a <=( A200  and  A199 );
 a25116a <=( (not A166)  and  a25115a );
 a25117a <=( a25116a  and  a25111a );
 a25121a <=( A234  and  (not A233) );
 a25122a <=( A232  and  a25121a );
 a25126a <=( (not A299)  and  (not A298) );
 a25127a <=( A236  and  a25126a );
 a25128a <=( a25127a  and  a25122a );
 a25132a <=( (not A167)  and  A169 );
 a25133a <=( (not A170)  and  a25132a );
 a25137a <=( A200  and  A199 );
 a25138a <=( (not A166)  and  a25137a );
 a25139a <=( a25138a  and  a25133a );
 a25143a <=( A234  and  (not A233) );
 a25144a <=( A232  and  a25143a );
 a25148a <=( A266  and  (not A265) );
 a25149a <=( A236  and  a25148a );
 a25150a <=( a25149a  and  a25144a );
 a25154a <=( (not A167)  and  A169 );
 a25155a <=( (not A170)  and  a25154a );
 a25159a <=( A200  and  A199 );
 a25160a <=( (not A166)  and  a25159a );
 a25161a <=( a25160a  and  a25155a );
 a25165a <=( A265  and  (not A233) );
 a25166a <=( (not A232)  and  a25165a );
 a25170a <=( A299  and  (not A298) );
 a25171a <=( A266  and  a25170a );
 a25172a <=( a25171a  and  a25166a );
 a25176a <=( (not A167)  and  A169 );
 a25177a <=( (not A170)  and  a25176a );
 a25181a <=( A200  and  A199 );
 a25182a <=( (not A166)  and  a25181a );
 a25183a <=( a25182a  and  a25177a );
 a25187a <=( (not A266)  and  (not A233) );
 a25188a <=( (not A232)  and  a25187a );
 a25192a <=( A299  and  (not A298) );
 a25193a <=( (not A267)  and  a25192a );
 a25194a <=( a25193a  and  a25188a );
 a25198a <=( (not A167)  and  A169 );
 a25199a <=( (not A170)  and  a25198a );
 a25203a <=( A200  and  A199 );
 a25204a <=( (not A166)  and  a25203a );
 a25205a <=( a25204a  and  a25199a );
 a25209a <=( (not A265)  and  (not A233) );
 a25210a <=( (not A232)  and  a25209a );
 a25214a <=( A299  and  (not A298) );
 a25215a <=( (not A266)  and  a25214a );
 a25216a <=( a25215a  and  a25210a );
 a25220a <=( (not A167)  and  A169 );
 a25221a <=( (not A170)  and  a25220a );
 a25225a <=( (not A202)  and  (not A200) );
 a25226a <=( (not A166)  and  a25225a );
 a25227a <=( a25226a  and  a25221a );
 a25231a <=( A233  and  (not A232) );
 a25232a <=( (not A203)  and  a25231a );
 a25236a <=( (not A302)  and  (not A301) );
 a25237a <=( (not A299)  and  a25236a );
 a25238a <=( a25237a  and  a25232a );
 a25242a <=( (not A167)  and  A169 );
 a25243a <=( (not A170)  and  a25242a );
 a25247a <=( (not A201)  and  (not A200) );
 a25248a <=( (not A166)  and  a25247a );
 a25249a <=( a25248a  and  a25243a );
 a25253a <=( A265  and  A233 );
 a25254a <=( A232  and  a25253a );
 a25258a <=( A299  and  (not A298) );
 a25259a <=( (not A267)  and  a25258a );
 a25260a <=( a25259a  and  a25254a );
 a25264a <=( (not A167)  and  A169 );
 a25265a <=( (not A170)  and  a25264a );
 a25269a <=( (not A201)  and  (not A200) );
 a25270a <=( (not A166)  and  a25269a );
 a25271a <=( a25270a  and  a25265a );
 a25275a <=( A265  and  A233 );
 a25276a <=( A232  and  a25275a );
 a25280a <=( A299  and  (not A298) );
 a25281a <=( A266  and  a25280a );
 a25282a <=( a25281a  and  a25276a );
 a25286a <=( (not A167)  and  A169 );
 a25287a <=( (not A170)  and  a25286a );
 a25291a <=( (not A201)  and  (not A200) );
 a25292a <=( (not A166)  and  a25291a );
 a25293a <=( a25292a  and  a25287a );
 a25297a <=( (not A265)  and  A233 );
 a25298a <=( A232  and  a25297a );
 a25302a <=( A299  and  (not A298) );
 a25303a <=( (not A266)  and  a25302a );
 a25304a <=( a25303a  and  a25298a );
 a25308a <=( (not A167)  and  A169 );
 a25309a <=( (not A170)  and  a25308a );
 a25313a <=( (not A201)  and  (not A200) );
 a25314a <=( (not A166)  and  a25313a );
 a25315a <=( a25314a  and  a25309a );
 a25319a <=( A265  and  A233 );
 a25320a <=( (not A232)  and  a25319a );
 a25324a <=( A268  and  A267 );
 a25325a <=( (not A266)  and  a25324a );
 a25326a <=( a25325a  and  a25320a );
 a25330a <=( (not A167)  and  A169 );
 a25331a <=( (not A170)  and  a25330a );
 a25335a <=( (not A201)  and  (not A200) );
 a25336a <=( (not A166)  and  a25335a );
 a25337a <=( a25336a  and  a25331a );
 a25341a <=( A265  and  A233 );
 a25342a <=( (not A232)  and  a25341a );
 a25346a <=( A269  and  A267 );
 a25347a <=( (not A266)  and  a25346a );
 a25348a <=( a25347a  and  a25342a );
 a25352a <=( (not A167)  and  A169 );
 a25353a <=( (not A170)  and  a25352a );
 a25357a <=( (not A201)  and  (not A200) );
 a25358a <=( (not A166)  and  a25357a );
 a25359a <=( a25358a  and  a25353a );
 a25363a <=( A265  and  (not A234) );
 a25364a <=( (not A233)  and  a25363a );
 a25368a <=( A299  and  (not A298) );
 a25369a <=( A266  and  a25368a );
 a25370a <=( a25369a  and  a25364a );
 a25374a <=( (not A167)  and  A169 );
 a25375a <=( (not A170)  and  a25374a );
 a25379a <=( (not A201)  and  (not A200) );
 a25380a <=( (not A166)  and  a25379a );
 a25381a <=( a25380a  and  a25375a );
 a25385a <=( (not A266)  and  (not A234) );
 a25386a <=( (not A233)  and  a25385a );
 a25390a <=( A299  and  (not A298) );
 a25391a <=( (not A267)  and  a25390a );
 a25392a <=( a25391a  and  a25386a );
 a25396a <=( (not A167)  and  A169 );
 a25397a <=( (not A170)  and  a25396a );
 a25401a <=( (not A201)  and  (not A200) );
 a25402a <=( (not A166)  and  a25401a );
 a25403a <=( a25402a  and  a25397a );
 a25407a <=( (not A265)  and  (not A234) );
 a25408a <=( (not A233)  and  a25407a );
 a25412a <=( A299  and  (not A298) );
 a25413a <=( (not A266)  and  a25412a );
 a25414a <=( a25413a  and  a25408a );
 a25418a <=( (not A167)  and  A169 );
 a25419a <=( (not A170)  and  a25418a );
 a25423a <=( (not A201)  and  (not A200) );
 a25424a <=( (not A166)  and  a25423a );
 a25425a <=( a25424a  and  a25419a );
 a25429a <=( A234  and  (not A233) );
 a25430a <=( A232  and  a25429a );
 a25434a <=( (not A300)  and  A298 );
 a25435a <=( A235  and  a25434a );
 a25436a <=( a25435a  and  a25430a );
 a25440a <=( (not A167)  and  A169 );
 a25441a <=( (not A170)  and  a25440a );
 a25445a <=( (not A201)  and  (not A200) );
 a25446a <=( (not A166)  and  a25445a );
 a25447a <=( a25446a  and  a25441a );
 a25451a <=( A234  and  (not A233) );
 a25452a <=( A232  and  a25451a );
 a25456a <=( A299  and  A298 );
 a25457a <=( A235  and  a25456a );
 a25458a <=( a25457a  and  a25452a );
 a25462a <=( (not A167)  and  A169 );
 a25463a <=( (not A170)  and  a25462a );
 a25467a <=( (not A201)  and  (not A200) );
 a25468a <=( (not A166)  and  a25467a );
 a25469a <=( a25468a  and  a25463a );
 a25473a <=( A234  and  (not A233) );
 a25474a <=( A232  and  a25473a );
 a25478a <=( (not A299)  and  (not A298) );
 a25479a <=( A235  and  a25478a );
 a25480a <=( a25479a  and  a25474a );
 a25484a <=( (not A167)  and  A169 );
 a25485a <=( (not A170)  and  a25484a );
 a25489a <=( (not A201)  and  (not A200) );
 a25490a <=( (not A166)  and  a25489a );
 a25491a <=( a25490a  and  a25485a );
 a25495a <=( A234  and  (not A233) );
 a25496a <=( A232  and  a25495a );
 a25500a <=( A266  and  (not A265) );
 a25501a <=( A235  and  a25500a );
 a25502a <=( a25501a  and  a25496a );
 a25506a <=( (not A167)  and  A169 );
 a25507a <=( (not A170)  and  a25506a );
 a25511a <=( (not A201)  and  (not A200) );
 a25512a <=( (not A166)  and  a25511a );
 a25513a <=( a25512a  and  a25507a );
 a25517a <=( A234  and  (not A233) );
 a25518a <=( A232  and  a25517a );
 a25522a <=( (not A300)  and  A298 );
 a25523a <=( A236  and  a25522a );
 a25524a <=( a25523a  and  a25518a );
 a25528a <=( (not A167)  and  A169 );
 a25529a <=( (not A170)  and  a25528a );
 a25533a <=( (not A201)  and  (not A200) );
 a25534a <=( (not A166)  and  a25533a );
 a25535a <=( a25534a  and  a25529a );
 a25539a <=( A234  and  (not A233) );
 a25540a <=( A232  and  a25539a );
 a25544a <=( A299  and  A298 );
 a25545a <=( A236  and  a25544a );
 a25546a <=( a25545a  and  a25540a );
 a25550a <=( (not A167)  and  A169 );
 a25551a <=( (not A170)  and  a25550a );
 a25555a <=( (not A201)  and  (not A200) );
 a25556a <=( (not A166)  and  a25555a );
 a25557a <=( a25556a  and  a25551a );
 a25561a <=( A234  and  (not A233) );
 a25562a <=( A232  and  a25561a );
 a25566a <=( (not A299)  and  (not A298) );
 a25567a <=( A236  and  a25566a );
 a25568a <=( a25567a  and  a25562a );
 a25572a <=( (not A167)  and  A169 );
 a25573a <=( (not A170)  and  a25572a );
 a25577a <=( (not A201)  and  (not A200) );
 a25578a <=( (not A166)  and  a25577a );
 a25579a <=( a25578a  and  a25573a );
 a25583a <=( A234  and  (not A233) );
 a25584a <=( A232  and  a25583a );
 a25588a <=( A266  and  (not A265) );
 a25589a <=( A236  and  a25588a );
 a25590a <=( a25589a  and  a25584a );
 a25594a <=( (not A167)  and  A169 );
 a25595a <=( (not A170)  and  a25594a );
 a25599a <=( (not A201)  and  (not A200) );
 a25600a <=( (not A166)  and  a25599a );
 a25601a <=( a25600a  and  a25595a );
 a25605a <=( A265  and  (not A233) );
 a25606a <=( (not A232)  and  a25605a );
 a25610a <=( A299  and  (not A298) );
 a25611a <=( A266  and  a25610a );
 a25612a <=( a25611a  and  a25606a );
 a25616a <=( (not A167)  and  A169 );
 a25617a <=( (not A170)  and  a25616a );
 a25621a <=( (not A201)  and  (not A200) );
 a25622a <=( (not A166)  and  a25621a );
 a25623a <=( a25622a  and  a25617a );
 a25627a <=( (not A266)  and  (not A233) );
 a25628a <=( (not A232)  and  a25627a );
 a25632a <=( A299  and  (not A298) );
 a25633a <=( (not A267)  and  a25632a );
 a25634a <=( a25633a  and  a25628a );
 a25638a <=( (not A167)  and  A169 );
 a25639a <=( (not A170)  and  a25638a );
 a25643a <=( (not A201)  and  (not A200) );
 a25644a <=( (not A166)  and  a25643a );
 a25645a <=( a25644a  and  a25639a );
 a25649a <=( (not A265)  and  (not A233) );
 a25650a <=( (not A232)  and  a25649a );
 a25654a <=( A299  and  (not A298) );
 a25655a <=( (not A266)  and  a25654a );
 a25656a <=( a25655a  and  a25650a );
 a25660a <=( (not A167)  and  A169 );
 a25661a <=( (not A170)  and  a25660a );
 a25665a <=( (not A200)  and  (not A199) );
 a25666a <=( (not A166)  and  a25665a );
 a25667a <=( a25666a  and  a25661a );
 a25671a <=( A265  and  A233 );
 a25672a <=( A232  and  a25671a );
 a25676a <=( A299  and  (not A298) );
 a25677a <=( (not A267)  and  a25676a );
 a25678a <=( a25677a  and  a25672a );
 a25682a <=( (not A167)  and  A169 );
 a25683a <=( (not A170)  and  a25682a );
 a25687a <=( (not A200)  and  (not A199) );
 a25688a <=( (not A166)  and  a25687a );
 a25689a <=( a25688a  and  a25683a );
 a25693a <=( A265  and  A233 );
 a25694a <=( A232  and  a25693a );
 a25698a <=( A299  and  (not A298) );
 a25699a <=( A266  and  a25698a );
 a25700a <=( a25699a  and  a25694a );
 a25704a <=( (not A167)  and  A169 );
 a25705a <=( (not A170)  and  a25704a );
 a25709a <=( (not A200)  and  (not A199) );
 a25710a <=( (not A166)  and  a25709a );
 a25711a <=( a25710a  and  a25705a );
 a25715a <=( (not A265)  and  A233 );
 a25716a <=( A232  and  a25715a );
 a25720a <=( A299  and  (not A298) );
 a25721a <=( (not A266)  and  a25720a );
 a25722a <=( a25721a  and  a25716a );
 a25726a <=( (not A167)  and  A169 );
 a25727a <=( (not A170)  and  a25726a );
 a25731a <=( (not A200)  and  (not A199) );
 a25732a <=( (not A166)  and  a25731a );
 a25733a <=( a25732a  and  a25727a );
 a25737a <=( A265  and  A233 );
 a25738a <=( (not A232)  and  a25737a );
 a25742a <=( A268  and  A267 );
 a25743a <=( (not A266)  and  a25742a );
 a25744a <=( a25743a  and  a25738a );
 a25748a <=( (not A167)  and  A169 );
 a25749a <=( (not A170)  and  a25748a );
 a25753a <=( (not A200)  and  (not A199) );
 a25754a <=( (not A166)  and  a25753a );
 a25755a <=( a25754a  and  a25749a );
 a25759a <=( A265  and  A233 );
 a25760a <=( (not A232)  and  a25759a );
 a25764a <=( A269  and  A267 );
 a25765a <=( (not A266)  and  a25764a );
 a25766a <=( a25765a  and  a25760a );
 a25770a <=( (not A167)  and  A169 );
 a25771a <=( (not A170)  and  a25770a );
 a25775a <=( (not A200)  and  (not A199) );
 a25776a <=( (not A166)  and  a25775a );
 a25777a <=( a25776a  and  a25771a );
 a25781a <=( A265  and  (not A234) );
 a25782a <=( (not A233)  and  a25781a );
 a25786a <=( A299  and  (not A298) );
 a25787a <=( A266  and  a25786a );
 a25788a <=( a25787a  and  a25782a );
 a25792a <=( (not A167)  and  A169 );
 a25793a <=( (not A170)  and  a25792a );
 a25797a <=( (not A200)  and  (not A199) );
 a25798a <=( (not A166)  and  a25797a );
 a25799a <=( a25798a  and  a25793a );
 a25803a <=( (not A266)  and  (not A234) );
 a25804a <=( (not A233)  and  a25803a );
 a25808a <=( A299  and  (not A298) );
 a25809a <=( (not A267)  and  a25808a );
 a25810a <=( a25809a  and  a25804a );
 a25814a <=( (not A167)  and  A169 );
 a25815a <=( (not A170)  and  a25814a );
 a25819a <=( (not A200)  and  (not A199) );
 a25820a <=( (not A166)  and  a25819a );
 a25821a <=( a25820a  and  a25815a );
 a25825a <=( (not A265)  and  (not A234) );
 a25826a <=( (not A233)  and  a25825a );
 a25830a <=( A299  and  (not A298) );
 a25831a <=( (not A266)  and  a25830a );
 a25832a <=( a25831a  and  a25826a );
 a25836a <=( (not A167)  and  A169 );
 a25837a <=( (not A170)  and  a25836a );
 a25841a <=( (not A200)  and  (not A199) );
 a25842a <=( (not A166)  and  a25841a );
 a25843a <=( a25842a  and  a25837a );
 a25847a <=( A234  and  (not A233) );
 a25848a <=( A232  and  a25847a );
 a25852a <=( (not A300)  and  A298 );
 a25853a <=( A235  and  a25852a );
 a25854a <=( a25853a  and  a25848a );
 a25858a <=( (not A167)  and  A169 );
 a25859a <=( (not A170)  and  a25858a );
 a25863a <=( (not A200)  and  (not A199) );
 a25864a <=( (not A166)  and  a25863a );
 a25865a <=( a25864a  and  a25859a );
 a25869a <=( A234  and  (not A233) );
 a25870a <=( A232  and  a25869a );
 a25874a <=( A299  and  A298 );
 a25875a <=( A235  and  a25874a );
 a25876a <=( a25875a  and  a25870a );
 a25880a <=( (not A167)  and  A169 );
 a25881a <=( (not A170)  and  a25880a );
 a25885a <=( (not A200)  and  (not A199) );
 a25886a <=( (not A166)  and  a25885a );
 a25887a <=( a25886a  and  a25881a );
 a25891a <=( A234  and  (not A233) );
 a25892a <=( A232  and  a25891a );
 a25896a <=( (not A299)  and  (not A298) );
 a25897a <=( A235  and  a25896a );
 a25898a <=( a25897a  and  a25892a );
 a25902a <=( (not A167)  and  A169 );
 a25903a <=( (not A170)  and  a25902a );
 a25907a <=( (not A200)  and  (not A199) );
 a25908a <=( (not A166)  and  a25907a );
 a25909a <=( a25908a  and  a25903a );
 a25913a <=( A234  and  (not A233) );
 a25914a <=( A232  and  a25913a );
 a25918a <=( A266  and  (not A265) );
 a25919a <=( A235  and  a25918a );
 a25920a <=( a25919a  and  a25914a );
 a25924a <=( (not A167)  and  A169 );
 a25925a <=( (not A170)  and  a25924a );
 a25929a <=( (not A200)  and  (not A199) );
 a25930a <=( (not A166)  and  a25929a );
 a25931a <=( a25930a  and  a25925a );
 a25935a <=( A234  and  (not A233) );
 a25936a <=( A232  and  a25935a );
 a25940a <=( (not A300)  and  A298 );
 a25941a <=( A236  and  a25940a );
 a25942a <=( a25941a  and  a25936a );
 a25946a <=( (not A167)  and  A169 );
 a25947a <=( (not A170)  and  a25946a );
 a25951a <=( (not A200)  and  (not A199) );
 a25952a <=( (not A166)  and  a25951a );
 a25953a <=( a25952a  and  a25947a );
 a25957a <=( A234  and  (not A233) );
 a25958a <=( A232  and  a25957a );
 a25962a <=( A299  and  A298 );
 a25963a <=( A236  and  a25962a );
 a25964a <=( a25963a  and  a25958a );
 a25968a <=( (not A167)  and  A169 );
 a25969a <=( (not A170)  and  a25968a );
 a25973a <=( (not A200)  and  (not A199) );
 a25974a <=( (not A166)  and  a25973a );
 a25975a <=( a25974a  and  a25969a );
 a25979a <=( A234  and  (not A233) );
 a25980a <=( A232  and  a25979a );
 a25984a <=( (not A299)  and  (not A298) );
 a25985a <=( A236  and  a25984a );
 a25986a <=( a25985a  and  a25980a );
 a25990a <=( (not A167)  and  A169 );
 a25991a <=( (not A170)  and  a25990a );
 a25995a <=( (not A200)  and  (not A199) );
 a25996a <=( (not A166)  and  a25995a );
 a25997a <=( a25996a  and  a25991a );
 a26001a <=( A234  and  (not A233) );
 a26002a <=( A232  and  a26001a );
 a26006a <=( A266  and  (not A265) );
 a26007a <=( A236  and  a26006a );
 a26008a <=( a26007a  and  a26002a );
 a26012a <=( (not A167)  and  A169 );
 a26013a <=( (not A170)  and  a26012a );
 a26017a <=( (not A200)  and  (not A199) );
 a26018a <=( (not A166)  and  a26017a );
 a26019a <=( a26018a  and  a26013a );
 a26023a <=( A265  and  (not A233) );
 a26024a <=( (not A232)  and  a26023a );
 a26028a <=( A299  and  (not A298) );
 a26029a <=( A266  and  a26028a );
 a26030a <=( a26029a  and  a26024a );
 a26034a <=( (not A167)  and  A169 );
 a26035a <=( (not A170)  and  a26034a );
 a26039a <=( (not A200)  and  (not A199) );
 a26040a <=( (not A166)  and  a26039a );
 a26041a <=( a26040a  and  a26035a );
 a26045a <=( (not A266)  and  (not A233) );
 a26046a <=( (not A232)  and  a26045a );
 a26050a <=( A299  and  (not A298) );
 a26051a <=( (not A267)  and  a26050a );
 a26052a <=( a26051a  and  a26046a );
 a26056a <=( (not A167)  and  A169 );
 a26057a <=( (not A170)  and  a26056a );
 a26061a <=( (not A200)  and  (not A199) );
 a26062a <=( (not A166)  and  a26061a );
 a26063a <=( a26062a  and  a26057a );
 a26067a <=( (not A265)  and  (not A233) );
 a26068a <=( (not A232)  and  a26067a );
 a26072a <=( A299  and  (not A298) );
 a26073a <=( (not A266)  and  a26072a );
 a26074a <=( a26073a  and  a26068a );
 a26078a <=( (not A166)  and  (not A167) );
 a26079a <=( (not A169)  and  a26078a );
 a26083a <=( A232  and  A200 );
 a26084a <=( (not A199)  and  a26083a );
 a26085a <=( a26084a  and  a26079a );
 a26089a <=( (not A268)  and  A265 );
 a26090a <=( A233  and  a26089a );
 a26094a <=( A299  and  (not A298) );
 a26095a <=( (not A269)  and  a26094a );
 a26096a <=( a26095a  and  a26090a );
 a26100a <=( (not A166)  and  (not A167) );
 a26101a <=( (not A169)  and  a26100a );
 a26105a <=( (not A233)  and  A200 );
 a26106a <=( (not A199)  and  a26105a );
 a26107a <=( a26106a  and  a26101a );
 a26111a <=( A265  and  (not A236) );
 a26112a <=( (not A235)  and  a26111a );
 a26116a <=( A299  and  (not A298) );
 a26117a <=( A266  and  a26116a );
 a26118a <=( a26117a  and  a26112a );
 a26122a <=( (not A166)  and  (not A167) );
 a26123a <=( (not A169)  and  a26122a );
 a26127a <=( (not A233)  and  A200 );
 a26128a <=( (not A199)  and  a26127a );
 a26129a <=( a26128a  and  a26123a );
 a26133a <=( (not A266)  and  (not A236) );
 a26134a <=( (not A235)  and  a26133a );
 a26138a <=( A299  and  (not A298) );
 a26139a <=( (not A267)  and  a26138a );
 a26140a <=( a26139a  and  a26134a );
 a26144a <=( (not A166)  and  (not A167) );
 a26145a <=( (not A169)  and  a26144a );
 a26149a <=( (not A233)  and  A200 );
 a26150a <=( (not A199)  and  a26149a );
 a26151a <=( a26150a  and  a26145a );
 a26155a <=( (not A265)  and  (not A236) );
 a26156a <=( (not A235)  and  a26155a );
 a26160a <=( A299  and  (not A298) );
 a26161a <=( (not A266)  and  a26160a );
 a26162a <=( a26161a  and  a26156a );
 a26166a <=( (not A166)  and  (not A167) );
 a26167a <=( (not A169)  and  a26166a );
 a26171a <=( (not A233)  and  A200 );
 a26172a <=( (not A199)  and  a26171a );
 a26173a <=( a26172a  and  a26167a );
 a26177a <=( (not A268)  and  (not A266) );
 a26178a <=( (not A234)  and  a26177a );
 a26182a <=( A299  and  (not A298) );
 a26183a <=( (not A269)  and  a26182a );
 a26184a <=( a26183a  and  a26178a );
 a26188a <=( (not A166)  and  (not A167) );
 a26189a <=( (not A169)  and  a26188a );
 a26193a <=( A232  and  A200 );
 a26194a <=( (not A199)  and  a26193a );
 a26195a <=( a26194a  and  a26189a );
 a26199a <=( A235  and  A234 );
 a26200a <=( (not A233)  and  a26199a );
 a26204a <=( (not A302)  and  (not A301) );
 a26205a <=( A298  and  a26204a );
 a26206a <=( a26205a  and  a26200a );
 a26210a <=( (not A166)  and  (not A167) );
 a26211a <=( (not A169)  and  a26210a );
 a26215a <=( A232  and  A200 );
 a26216a <=( (not A199)  and  a26215a );
 a26217a <=( a26216a  and  a26211a );
 a26221a <=( A236  and  A234 );
 a26222a <=( (not A233)  and  a26221a );
 a26226a <=( (not A302)  and  (not A301) );
 a26227a <=( A298  and  a26226a );
 a26228a <=( a26227a  and  a26222a );
 a26232a <=( (not A166)  and  (not A167) );
 a26233a <=( (not A169)  and  a26232a );
 a26237a <=( (not A232)  and  A200 );
 a26238a <=( (not A199)  and  a26237a );
 a26239a <=( a26238a  and  a26233a );
 a26243a <=( (not A268)  and  (not A266) );
 a26244a <=( (not A233)  and  a26243a );
 a26248a <=( A299  and  (not A298) );
 a26249a <=( (not A269)  and  a26248a );
 a26250a <=( a26249a  and  a26244a );
 a26254a <=( (not A166)  and  (not A167) );
 a26255a <=( (not A169)  and  a26254a );
 a26259a <=( A201  and  (not A200) );
 a26260a <=( A199  and  a26259a );
 a26261a <=( a26260a  and  a26255a );
 a26265a <=( A233  and  (not A232) );
 a26266a <=( A202  and  a26265a );
 a26270a <=( (not A302)  and  (not A301) );
 a26271a <=( (not A299)  and  a26270a );
 a26272a <=( a26271a  and  a26266a );
 a26276a <=( (not A166)  and  (not A167) );
 a26277a <=( (not A169)  and  a26276a );
 a26281a <=( A201  and  (not A200) );
 a26282a <=( A199  and  a26281a );
 a26283a <=( a26282a  and  a26277a );
 a26287a <=( A233  and  (not A232) );
 a26288a <=( A203  and  a26287a );
 a26292a <=( (not A302)  and  (not A301) );
 a26293a <=( (not A299)  and  a26292a );
 a26294a <=( a26293a  and  a26288a );
 a26298a <=( A167  and  (not A168) );
 a26299a <=( (not A169)  and  a26298a );
 a26303a <=( A200  and  (not A199) );
 a26304a <=( A166  and  a26303a );
 a26305a <=( a26304a  and  a26299a );
 a26309a <=( A265  and  A233 );
 a26310a <=( A232  and  a26309a );
 a26314a <=( A299  and  (not A298) );
 a26315a <=( (not A267)  and  a26314a );
 a26316a <=( a26315a  and  a26310a );
 a26320a <=( A167  and  (not A168) );
 a26321a <=( (not A169)  and  a26320a );
 a26325a <=( A200  and  (not A199) );
 a26326a <=( A166  and  a26325a );
 a26327a <=( a26326a  and  a26321a );
 a26331a <=( A265  and  A233 );
 a26332a <=( A232  and  a26331a );
 a26336a <=( A299  and  (not A298) );
 a26337a <=( A266  and  a26336a );
 a26338a <=( a26337a  and  a26332a );
 a26342a <=( A167  and  (not A168) );
 a26343a <=( (not A169)  and  a26342a );
 a26347a <=( A200  and  (not A199) );
 a26348a <=( A166  and  a26347a );
 a26349a <=( a26348a  and  a26343a );
 a26353a <=( (not A265)  and  A233 );
 a26354a <=( A232  and  a26353a );
 a26358a <=( A299  and  (not A298) );
 a26359a <=( (not A266)  and  a26358a );
 a26360a <=( a26359a  and  a26354a );
 a26364a <=( A167  and  (not A168) );
 a26365a <=( (not A169)  and  a26364a );
 a26369a <=( A200  and  (not A199) );
 a26370a <=( A166  and  a26369a );
 a26371a <=( a26370a  and  a26365a );
 a26375a <=( A265  and  A233 );
 a26376a <=( (not A232)  and  a26375a );
 a26380a <=( A268  and  A267 );
 a26381a <=( (not A266)  and  a26380a );
 a26382a <=( a26381a  and  a26376a );
 a26386a <=( A167  and  (not A168) );
 a26387a <=( (not A169)  and  a26386a );
 a26391a <=( A200  and  (not A199) );
 a26392a <=( A166  and  a26391a );
 a26393a <=( a26392a  and  a26387a );
 a26397a <=( A265  and  A233 );
 a26398a <=( (not A232)  and  a26397a );
 a26402a <=( A269  and  A267 );
 a26403a <=( (not A266)  and  a26402a );
 a26404a <=( a26403a  and  a26398a );
 a26408a <=( A167  and  (not A168) );
 a26409a <=( (not A169)  and  a26408a );
 a26413a <=( A200  and  (not A199) );
 a26414a <=( A166  and  a26413a );
 a26415a <=( a26414a  and  a26409a );
 a26419a <=( A265  and  (not A234) );
 a26420a <=( (not A233)  and  a26419a );
 a26424a <=( A299  and  (not A298) );
 a26425a <=( A266  and  a26424a );
 a26426a <=( a26425a  and  a26420a );
 a26430a <=( A167  and  (not A168) );
 a26431a <=( (not A169)  and  a26430a );
 a26435a <=( A200  and  (not A199) );
 a26436a <=( A166  and  a26435a );
 a26437a <=( a26436a  and  a26431a );
 a26441a <=( (not A266)  and  (not A234) );
 a26442a <=( (not A233)  and  a26441a );
 a26446a <=( A299  and  (not A298) );
 a26447a <=( (not A267)  and  a26446a );
 a26448a <=( a26447a  and  a26442a );
 a26452a <=( A167  and  (not A168) );
 a26453a <=( (not A169)  and  a26452a );
 a26457a <=( A200  and  (not A199) );
 a26458a <=( A166  and  a26457a );
 a26459a <=( a26458a  and  a26453a );
 a26463a <=( (not A265)  and  (not A234) );
 a26464a <=( (not A233)  and  a26463a );
 a26468a <=( A299  and  (not A298) );
 a26469a <=( (not A266)  and  a26468a );
 a26470a <=( a26469a  and  a26464a );
 a26474a <=( A167  and  (not A168) );
 a26475a <=( (not A169)  and  a26474a );
 a26479a <=( A200  and  (not A199) );
 a26480a <=( A166  and  a26479a );
 a26481a <=( a26480a  and  a26475a );
 a26485a <=( A234  and  (not A233) );
 a26486a <=( A232  and  a26485a );
 a26490a <=( (not A300)  and  A298 );
 a26491a <=( A235  and  a26490a );
 a26492a <=( a26491a  and  a26486a );
 a26496a <=( A167  and  (not A168) );
 a26497a <=( (not A169)  and  a26496a );
 a26501a <=( A200  and  (not A199) );
 a26502a <=( A166  and  a26501a );
 a26503a <=( a26502a  and  a26497a );
 a26507a <=( A234  and  (not A233) );
 a26508a <=( A232  and  a26507a );
 a26512a <=( A299  and  A298 );
 a26513a <=( A235  and  a26512a );
 a26514a <=( a26513a  and  a26508a );
 a26518a <=( A167  and  (not A168) );
 a26519a <=( (not A169)  and  a26518a );
 a26523a <=( A200  and  (not A199) );
 a26524a <=( A166  and  a26523a );
 a26525a <=( a26524a  and  a26519a );
 a26529a <=( A234  and  (not A233) );
 a26530a <=( A232  and  a26529a );
 a26534a <=( (not A299)  and  (not A298) );
 a26535a <=( A235  and  a26534a );
 a26536a <=( a26535a  and  a26530a );
 a26540a <=( A167  and  (not A168) );
 a26541a <=( (not A169)  and  a26540a );
 a26545a <=( A200  and  (not A199) );
 a26546a <=( A166  and  a26545a );
 a26547a <=( a26546a  and  a26541a );
 a26551a <=( A234  and  (not A233) );
 a26552a <=( A232  and  a26551a );
 a26556a <=( A266  and  (not A265) );
 a26557a <=( A235  and  a26556a );
 a26558a <=( a26557a  and  a26552a );
 a26562a <=( A167  and  (not A168) );
 a26563a <=( (not A169)  and  a26562a );
 a26567a <=( A200  and  (not A199) );
 a26568a <=( A166  and  a26567a );
 a26569a <=( a26568a  and  a26563a );
 a26573a <=( A234  and  (not A233) );
 a26574a <=( A232  and  a26573a );
 a26578a <=( (not A300)  and  A298 );
 a26579a <=( A236  and  a26578a );
 a26580a <=( a26579a  and  a26574a );
 a26584a <=( A167  and  (not A168) );
 a26585a <=( (not A169)  and  a26584a );
 a26589a <=( A200  and  (not A199) );
 a26590a <=( A166  and  a26589a );
 a26591a <=( a26590a  and  a26585a );
 a26595a <=( A234  and  (not A233) );
 a26596a <=( A232  and  a26595a );
 a26600a <=( A299  and  A298 );
 a26601a <=( A236  and  a26600a );
 a26602a <=( a26601a  and  a26596a );
 a26606a <=( A167  and  (not A168) );
 a26607a <=( (not A169)  and  a26606a );
 a26611a <=( A200  and  (not A199) );
 a26612a <=( A166  and  a26611a );
 a26613a <=( a26612a  and  a26607a );
 a26617a <=( A234  and  (not A233) );
 a26618a <=( A232  and  a26617a );
 a26622a <=( (not A299)  and  (not A298) );
 a26623a <=( A236  and  a26622a );
 a26624a <=( a26623a  and  a26618a );
 a26628a <=( A167  and  (not A168) );
 a26629a <=( (not A169)  and  a26628a );
 a26633a <=( A200  and  (not A199) );
 a26634a <=( A166  and  a26633a );
 a26635a <=( a26634a  and  a26629a );
 a26639a <=( A234  and  (not A233) );
 a26640a <=( A232  and  a26639a );
 a26644a <=( A266  and  (not A265) );
 a26645a <=( A236  and  a26644a );
 a26646a <=( a26645a  and  a26640a );
 a26650a <=( A167  and  (not A168) );
 a26651a <=( (not A169)  and  a26650a );
 a26655a <=( A200  and  (not A199) );
 a26656a <=( A166  and  a26655a );
 a26657a <=( a26656a  and  a26651a );
 a26661a <=( A265  and  (not A233) );
 a26662a <=( (not A232)  and  a26661a );
 a26666a <=( A299  and  (not A298) );
 a26667a <=( A266  and  a26666a );
 a26668a <=( a26667a  and  a26662a );
 a26672a <=( A167  and  (not A168) );
 a26673a <=( (not A169)  and  a26672a );
 a26677a <=( A200  and  (not A199) );
 a26678a <=( A166  and  a26677a );
 a26679a <=( a26678a  and  a26673a );
 a26683a <=( (not A266)  and  (not A233) );
 a26684a <=( (not A232)  and  a26683a );
 a26688a <=( A299  and  (not A298) );
 a26689a <=( (not A267)  and  a26688a );
 a26690a <=( a26689a  and  a26684a );
 a26694a <=( A167  and  (not A168) );
 a26695a <=( (not A169)  and  a26694a );
 a26699a <=( A200  and  (not A199) );
 a26700a <=( A166  and  a26699a );
 a26701a <=( a26700a  and  a26695a );
 a26705a <=( (not A265)  and  (not A233) );
 a26706a <=( (not A232)  and  a26705a );
 a26710a <=( A299  and  (not A298) );
 a26711a <=( (not A266)  and  a26710a );
 a26712a <=( a26711a  and  a26706a );
 a26716a <=( A167  and  (not A168) );
 a26717a <=( (not A169)  and  a26716a );
 a26721a <=( (not A200)  and  A199 );
 a26722a <=( A166  and  a26721a );
 a26723a <=( a26722a  and  a26717a );
 a26727a <=( (not A232)  and  A202 );
 a26728a <=( A201  and  a26727a );
 a26732a <=( (not A300)  and  (not A299) );
 a26733a <=( A233  and  a26732a );
 a26734a <=( a26733a  and  a26728a );
 a26738a <=( A167  and  (not A168) );
 a26739a <=( (not A169)  and  a26738a );
 a26743a <=( (not A200)  and  A199 );
 a26744a <=( A166  and  a26743a );
 a26745a <=( a26744a  and  a26739a );
 a26749a <=( (not A232)  and  A202 );
 a26750a <=( A201  and  a26749a );
 a26754a <=( A299  and  A298 );
 a26755a <=( A233  and  a26754a );
 a26756a <=( a26755a  and  a26750a );
 a26760a <=( A167  and  (not A168) );
 a26761a <=( (not A169)  and  a26760a );
 a26765a <=( (not A200)  and  A199 );
 a26766a <=( A166  and  a26765a );
 a26767a <=( a26766a  and  a26761a );
 a26771a <=( (not A232)  and  A202 );
 a26772a <=( A201  and  a26771a );
 a26776a <=( (not A299)  and  (not A298) );
 a26777a <=( A233  and  a26776a );
 a26778a <=( a26777a  and  a26772a );
 a26782a <=( A167  and  (not A168) );
 a26783a <=( (not A169)  and  a26782a );
 a26787a <=( (not A200)  and  A199 );
 a26788a <=( A166  and  a26787a );
 a26789a <=( a26788a  and  a26783a );
 a26793a <=( (not A232)  and  A202 );
 a26794a <=( A201  and  a26793a );
 a26798a <=( A266  and  (not A265) );
 a26799a <=( A233  and  a26798a );
 a26800a <=( a26799a  and  a26794a );
 a26804a <=( A167  and  (not A168) );
 a26805a <=( (not A169)  and  a26804a );
 a26809a <=( (not A200)  and  A199 );
 a26810a <=( A166  and  a26809a );
 a26811a <=( a26810a  and  a26805a );
 a26815a <=( (not A232)  and  A203 );
 a26816a <=( A201  and  a26815a );
 a26820a <=( (not A300)  and  (not A299) );
 a26821a <=( A233  and  a26820a );
 a26822a <=( a26821a  and  a26816a );
 a26826a <=( A167  and  (not A168) );
 a26827a <=( (not A169)  and  a26826a );
 a26831a <=( (not A200)  and  A199 );
 a26832a <=( A166  and  a26831a );
 a26833a <=( a26832a  and  a26827a );
 a26837a <=( (not A232)  and  A203 );
 a26838a <=( A201  and  a26837a );
 a26842a <=( A299  and  A298 );
 a26843a <=( A233  and  a26842a );
 a26844a <=( a26843a  and  a26838a );
 a26848a <=( A167  and  (not A168) );
 a26849a <=( (not A169)  and  a26848a );
 a26853a <=( (not A200)  and  A199 );
 a26854a <=( A166  and  a26853a );
 a26855a <=( a26854a  and  a26849a );
 a26859a <=( (not A232)  and  A203 );
 a26860a <=( A201  and  a26859a );
 a26864a <=( (not A299)  and  (not A298) );
 a26865a <=( A233  and  a26864a );
 a26866a <=( a26865a  and  a26860a );
 a26870a <=( A167  and  (not A168) );
 a26871a <=( (not A169)  and  a26870a );
 a26875a <=( (not A200)  and  A199 );
 a26876a <=( A166  and  a26875a );
 a26877a <=( a26876a  and  a26871a );
 a26881a <=( (not A232)  and  A203 );
 a26882a <=( A201  and  a26881a );
 a26886a <=( A266  and  (not A265) );
 a26887a <=( A233  and  a26886a );
 a26888a <=( a26887a  and  a26882a );
 a26892a <=( A167  and  (not A169) );
 a26893a <=( A170  and  a26892a );
 a26897a <=( A200  and  A199 );
 a26898a <=( (not A166)  and  a26897a );
 a26899a <=( a26898a  and  a26893a );
 a26903a <=( A265  and  A233 );
 a26904a <=( A232  and  a26903a );
 a26908a <=( A299  and  (not A298) );
 a26909a <=( (not A267)  and  a26908a );
 a26910a <=( a26909a  and  a26904a );
 a26914a <=( A167  and  (not A169) );
 a26915a <=( A170  and  a26914a );
 a26919a <=( A200  and  A199 );
 a26920a <=( (not A166)  and  a26919a );
 a26921a <=( a26920a  and  a26915a );
 a26925a <=( A265  and  A233 );
 a26926a <=( A232  and  a26925a );
 a26930a <=( A299  and  (not A298) );
 a26931a <=( A266  and  a26930a );
 a26932a <=( a26931a  and  a26926a );
 a26936a <=( A167  and  (not A169) );
 a26937a <=( A170  and  a26936a );
 a26941a <=( A200  and  A199 );
 a26942a <=( (not A166)  and  a26941a );
 a26943a <=( a26942a  and  a26937a );
 a26947a <=( (not A265)  and  A233 );
 a26948a <=( A232  and  a26947a );
 a26952a <=( A299  and  (not A298) );
 a26953a <=( (not A266)  and  a26952a );
 a26954a <=( a26953a  and  a26948a );
 a26958a <=( A167  and  (not A169) );
 a26959a <=( A170  and  a26958a );
 a26963a <=( A200  and  A199 );
 a26964a <=( (not A166)  and  a26963a );
 a26965a <=( a26964a  and  a26959a );
 a26969a <=( A265  and  A233 );
 a26970a <=( (not A232)  and  a26969a );
 a26974a <=( A268  and  A267 );
 a26975a <=( (not A266)  and  a26974a );
 a26976a <=( a26975a  and  a26970a );
 a26980a <=( A167  and  (not A169) );
 a26981a <=( A170  and  a26980a );
 a26985a <=( A200  and  A199 );
 a26986a <=( (not A166)  and  a26985a );
 a26987a <=( a26986a  and  a26981a );
 a26991a <=( A265  and  A233 );
 a26992a <=( (not A232)  and  a26991a );
 a26996a <=( A269  and  A267 );
 a26997a <=( (not A266)  and  a26996a );
 a26998a <=( a26997a  and  a26992a );
 a27002a <=( A167  and  (not A169) );
 a27003a <=( A170  and  a27002a );
 a27007a <=( A200  and  A199 );
 a27008a <=( (not A166)  and  a27007a );
 a27009a <=( a27008a  and  a27003a );
 a27013a <=( A265  and  (not A234) );
 a27014a <=( (not A233)  and  a27013a );
 a27018a <=( A299  and  (not A298) );
 a27019a <=( A266  and  a27018a );
 a27020a <=( a27019a  and  a27014a );
 a27024a <=( A167  and  (not A169) );
 a27025a <=( A170  and  a27024a );
 a27029a <=( A200  and  A199 );
 a27030a <=( (not A166)  and  a27029a );
 a27031a <=( a27030a  and  a27025a );
 a27035a <=( (not A266)  and  (not A234) );
 a27036a <=( (not A233)  and  a27035a );
 a27040a <=( A299  and  (not A298) );
 a27041a <=( (not A267)  and  a27040a );
 a27042a <=( a27041a  and  a27036a );
 a27046a <=( A167  and  (not A169) );
 a27047a <=( A170  and  a27046a );
 a27051a <=( A200  and  A199 );
 a27052a <=( (not A166)  and  a27051a );
 a27053a <=( a27052a  and  a27047a );
 a27057a <=( (not A265)  and  (not A234) );
 a27058a <=( (not A233)  and  a27057a );
 a27062a <=( A299  and  (not A298) );
 a27063a <=( (not A266)  and  a27062a );
 a27064a <=( a27063a  and  a27058a );
 a27068a <=( A167  and  (not A169) );
 a27069a <=( A170  and  a27068a );
 a27073a <=( A200  and  A199 );
 a27074a <=( (not A166)  and  a27073a );
 a27075a <=( a27074a  and  a27069a );
 a27079a <=( A234  and  (not A233) );
 a27080a <=( A232  and  a27079a );
 a27084a <=( (not A300)  and  A298 );
 a27085a <=( A235  and  a27084a );
 a27086a <=( a27085a  and  a27080a );
 a27090a <=( A167  and  (not A169) );
 a27091a <=( A170  and  a27090a );
 a27095a <=( A200  and  A199 );
 a27096a <=( (not A166)  and  a27095a );
 a27097a <=( a27096a  and  a27091a );
 a27101a <=( A234  and  (not A233) );
 a27102a <=( A232  and  a27101a );
 a27106a <=( A299  and  A298 );
 a27107a <=( A235  and  a27106a );
 a27108a <=( a27107a  and  a27102a );
 a27112a <=( A167  and  (not A169) );
 a27113a <=( A170  and  a27112a );
 a27117a <=( A200  and  A199 );
 a27118a <=( (not A166)  and  a27117a );
 a27119a <=( a27118a  and  a27113a );
 a27123a <=( A234  and  (not A233) );
 a27124a <=( A232  and  a27123a );
 a27128a <=( (not A299)  and  (not A298) );
 a27129a <=( A235  and  a27128a );
 a27130a <=( a27129a  and  a27124a );
 a27134a <=( A167  and  (not A169) );
 a27135a <=( A170  and  a27134a );
 a27139a <=( A200  and  A199 );
 a27140a <=( (not A166)  and  a27139a );
 a27141a <=( a27140a  and  a27135a );
 a27145a <=( A234  and  (not A233) );
 a27146a <=( A232  and  a27145a );
 a27150a <=( A266  and  (not A265) );
 a27151a <=( A235  and  a27150a );
 a27152a <=( a27151a  and  a27146a );
 a27156a <=( A167  and  (not A169) );
 a27157a <=( A170  and  a27156a );
 a27161a <=( A200  and  A199 );
 a27162a <=( (not A166)  and  a27161a );
 a27163a <=( a27162a  and  a27157a );
 a27167a <=( A234  and  (not A233) );
 a27168a <=( A232  and  a27167a );
 a27172a <=( (not A300)  and  A298 );
 a27173a <=( A236  and  a27172a );
 a27174a <=( a27173a  and  a27168a );
 a27178a <=( A167  and  (not A169) );
 a27179a <=( A170  and  a27178a );
 a27183a <=( A200  and  A199 );
 a27184a <=( (not A166)  and  a27183a );
 a27185a <=( a27184a  and  a27179a );
 a27189a <=( A234  and  (not A233) );
 a27190a <=( A232  and  a27189a );
 a27194a <=( A299  and  A298 );
 a27195a <=( A236  and  a27194a );
 a27196a <=( a27195a  and  a27190a );
 a27200a <=( A167  and  (not A169) );
 a27201a <=( A170  and  a27200a );
 a27205a <=( A200  and  A199 );
 a27206a <=( (not A166)  and  a27205a );
 a27207a <=( a27206a  and  a27201a );
 a27211a <=( A234  and  (not A233) );
 a27212a <=( A232  and  a27211a );
 a27216a <=( (not A299)  and  (not A298) );
 a27217a <=( A236  and  a27216a );
 a27218a <=( a27217a  and  a27212a );
 a27222a <=( A167  and  (not A169) );
 a27223a <=( A170  and  a27222a );
 a27227a <=( A200  and  A199 );
 a27228a <=( (not A166)  and  a27227a );
 a27229a <=( a27228a  and  a27223a );
 a27233a <=( A234  and  (not A233) );
 a27234a <=( A232  and  a27233a );
 a27238a <=( A266  and  (not A265) );
 a27239a <=( A236  and  a27238a );
 a27240a <=( a27239a  and  a27234a );
 a27244a <=( A167  and  (not A169) );
 a27245a <=( A170  and  a27244a );
 a27249a <=( A200  and  A199 );
 a27250a <=( (not A166)  and  a27249a );
 a27251a <=( a27250a  and  a27245a );
 a27255a <=( A265  and  (not A233) );
 a27256a <=( (not A232)  and  a27255a );
 a27260a <=( A299  and  (not A298) );
 a27261a <=( A266  and  a27260a );
 a27262a <=( a27261a  and  a27256a );
 a27266a <=( A167  and  (not A169) );
 a27267a <=( A170  and  a27266a );
 a27271a <=( A200  and  A199 );
 a27272a <=( (not A166)  and  a27271a );
 a27273a <=( a27272a  and  a27267a );
 a27277a <=( (not A266)  and  (not A233) );
 a27278a <=( (not A232)  and  a27277a );
 a27282a <=( A299  and  (not A298) );
 a27283a <=( (not A267)  and  a27282a );
 a27284a <=( a27283a  and  a27278a );
 a27288a <=( A167  and  (not A169) );
 a27289a <=( A170  and  a27288a );
 a27293a <=( A200  and  A199 );
 a27294a <=( (not A166)  and  a27293a );
 a27295a <=( a27294a  and  a27289a );
 a27299a <=( (not A265)  and  (not A233) );
 a27300a <=( (not A232)  and  a27299a );
 a27304a <=( A299  and  (not A298) );
 a27305a <=( (not A266)  and  a27304a );
 a27306a <=( a27305a  and  a27300a );
 a27310a <=( A167  and  (not A169) );
 a27311a <=( A170  and  a27310a );
 a27315a <=( (not A202)  and  (not A200) );
 a27316a <=( (not A166)  and  a27315a );
 a27317a <=( a27316a  and  a27311a );
 a27321a <=( A233  and  (not A232) );
 a27322a <=( (not A203)  and  a27321a );
 a27326a <=( (not A302)  and  (not A301) );
 a27327a <=( (not A299)  and  a27326a );
 a27328a <=( a27327a  and  a27322a );
 a27332a <=( A167  and  (not A169) );
 a27333a <=( A170  and  a27332a );
 a27337a <=( (not A201)  and  (not A200) );
 a27338a <=( (not A166)  and  a27337a );
 a27339a <=( a27338a  and  a27333a );
 a27343a <=( A265  and  A233 );
 a27344a <=( A232  and  a27343a );
 a27348a <=( A299  and  (not A298) );
 a27349a <=( (not A267)  and  a27348a );
 a27350a <=( a27349a  and  a27344a );
 a27354a <=( A167  and  (not A169) );
 a27355a <=( A170  and  a27354a );
 a27359a <=( (not A201)  and  (not A200) );
 a27360a <=( (not A166)  and  a27359a );
 a27361a <=( a27360a  and  a27355a );
 a27365a <=( A265  and  A233 );
 a27366a <=( A232  and  a27365a );
 a27370a <=( A299  and  (not A298) );
 a27371a <=( A266  and  a27370a );
 a27372a <=( a27371a  and  a27366a );
 a27376a <=( A167  and  (not A169) );
 a27377a <=( A170  and  a27376a );
 a27381a <=( (not A201)  and  (not A200) );
 a27382a <=( (not A166)  and  a27381a );
 a27383a <=( a27382a  and  a27377a );
 a27387a <=( (not A265)  and  A233 );
 a27388a <=( A232  and  a27387a );
 a27392a <=( A299  and  (not A298) );
 a27393a <=( (not A266)  and  a27392a );
 a27394a <=( a27393a  and  a27388a );
 a27398a <=( A167  and  (not A169) );
 a27399a <=( A170  and  a27398a );
 a27403a <=( (not A201)  and  (not A200) );
 a27404a <=( (not A166)  and  a27403a );
 a27405a <=( a27404a  and  a27399a );
 a27409a <=( A265  and  A233 );
 a27410a <=( (not A232)  and  a27409a );
 a27414a <=( A268  and  A267 );
 a27415a <=( (not A266)  and  a27414a );
 a27416a <=( a27415a  and  a27410a );
 a27420a <=( A167  and  (not A169) );
 a27421a <=( A170  and  a27420a );
 a27425a <=( (not A201)  and  (not A200) );
 a27426a <=( (not A166)  and  a27425a );
 a27427a <=( a27426a  and  a27421a );
 a27431a <=( A265  and  A233 );
 a27432a <=( (not A232)  and  a27431a );
 a27436a <=( A269  and  A267 );
 a27437a <=( (not A266)  and  a27436a );
 a27438a <=( a27437a  and  a27432a );
 a27442a <=( A167  and  (not A169) );
 a27443a <=( A170  and  a27442a );
 a27447a <=( (not A201)  and  (not A200) );
 a27448a <=( (not A166)  and  a27447a );
 a27449a <=( a27448a  and  a27443a );
 a27453a <=( A265  and  (not A234) );
 a27454a <=( (not A233)  and  a27453a );
 a27458a <=( A299  and  (not A298) );
 a27459a <=( A266  and  a27458a );
 a27460a <=( a27459a  and  a27454a );
 a27464a <=( A167  and  (not A169) );
 a27465a <=( A170  and  a27464a );
 a27469a <=( (not A201)  and  (not A200) );
 a27470a <=( (not A166)  and  a27469a );
 a27471a <=( a27470a  and  a27465a );
 a27475a <=( (not A266)  and  (not A234) );
 a27476a <=( (not A233)  and  a27475a );
 a27480a <=( A299  and  (not A298) );
 a27481a <=( (not A267)  and  a27480a );
 a27482a <=( a27481a  and  a27476a );
 a27486a <=( A167  and  (not A169) );
 a27487a <=( A170  and  a27486a );
 a27491a <=( (not A201)  and  (not A200) );
 a27492a <=( (not A166)  and  a27491a );
 a27493a <=( a27492a  and  a27487a );
 a27497a <=( (not A265)  and  (not A234) );
 a27498a <=( (not A233)  and  a27497a );
 a27502a <=( A299  and  (not A298) );
 a27503a <=( (not A266)  and  a27502a );
 a27504a <=( a27503a  and  a27498a );
 a27508a <=( A167  and  (not A169) );
 a27509a <=( A170  and  a27508a );
 a27513a <=( (not A201)  and  (not A200) );
 a27514a <=( (not A166)  and  a27513a );
 a27515a <=( a27514a  and  a27509a );
 a27519a <=( A234  and  (not A233) );
 a27520a <=( A232  and  a27519a );
 a27524a <=( (not A300)  and  A298 );
 a27525a <=( A235  and  a27524a );
 a27526a <=( a27525a  and  a27520a );
 a27530a <=( A167  and  (not A169) );
 a27531a <=( A170  and  a27530a );
 a27535a <=( (not A201)  and  (not A200) );
 a27536a <=( (not A166)  and  a27535a );
 a27537a <=( a27536a  and  a27531a );
 a27541a <=( A234  and  (not A233) );
 a27542a <=( A232  and  a27541a );
 a27546a <=( A299  and  A298 );
 a27547a <=( A235  and  a27546a );
 a27548a <=( a27547a  and  a27542a );
 a27552a <=( A167  and  (not A169) );
 a27553a <=( A170  and  a27552a );
 a27557a <=( (not A201)  and  (not A200) );
 a27558a <=( (not A166)  and  a27557a );
 a27559a <=( a27558a  and  a27553a );
 a27563a <=( A234  and  (not A233) );
 a27564a <=( A232  and  a27563a );
 a27568a <=( (not A299)  and  (not A298) );
 a27569a <=( A235  and  a27568a );
 a27570a <=( a27569a  and  a27564a );
 a27574a <=( A167  and  (not A169) );
 a27575a <=( A170  and  a27574a );
 a27579a <=( (not A201)  and  (not A200) );
 a27580a <=( (not A166)  and  a27579a );
 a27581a <=( a27580a  and  a27575a );
 a27585a <=( A234  and  (not A233) );
 a27586a <=( A232  and  a27585a );
 a27590a <=( A266  and  (not A265) );
 a27591a <=( A235  and  a27590a );
 a27592a <=( a27591a  and  a27586a );
 a27596a <=( A167  and  (not A169) );
 a27597a <=( A170  and  a27596a );
 a27601a <=( (not A201)  and  (not A200) );
 a27602a <=( (not A166)  and  a27601a );
 a27603a <=( a27602a  and  a27597a );
 a27607a <=( A234  and  (not A233) );
 a27608a <=( A232  and  a27607a );
 a27612a <=( (not A300)  and  A298 );
 a27613a <=( A236  and  a27612a );
 a27614a <=( a27613a  and  a27608a );
 a27618a <=( A167  and  (not A169) );
 a27619a <=( A170  and  a27618a );
 a27623a <=( (not A201)  and  (not A200) );
 a27624a <=( (not A166)  and  a27623a );
 a27625a <=( a27624a  and  a27619a );
 a27629a <=( A234  and  (not A233) );
 a27630a <=( A232  and  a27629a );
 a27634a <=( A299  and  A298 );
 a27635a <=( A236  and  a27634a );
 a27636a <=( a27635a  and  a27630a );
 a27640a <=( A167  and  (not A169) );
 a27641a <=( A170  and  a27640a );
 a27645a <=( (not A201)  and  (not A200) );
 a27646a <=( (not A166)  and  a27645a );
 a27647a <=( a27646a  and  a27641a );
 a27651a <=( A234  and  (not A233) );
 a27652a <=( A232  and  a27651a );
 a27656a <=( (not A299)  and  (not A298) );
 a27657a <=( A236  and  a27656a );
 a27658a <=( a27657a  and  a27652a );
 a27662a <=( A167  and  (not A169) );
 a27663a <=( A170  and  a27662a );
 a27667a <=( (not A201)  and  (not A200) );
 a27668a <=( (not A166)  and  a27667a );
 a27669a <=( a27668a  and  a27663a );
 a27673a <=( A234  and  (not A233) );
 a27674a <=( A232  and  a27673a );
 a27678a <=( A266  and  (not A265) );
 a27679a <=( A236  and  a27678a );
 a27680a <=( a27679a  and  a27674a );
 a27684a <=( A167  and  (not A169) );
 a27685a <=( A170  and  a27684a );
 a27689a <=( (not A201)  and  (not A200) );
 a27690a <=( (not A166)  and  a27689a );
 a27691a <=( a27690a  and  a27685a );
 a27695a <=( A265  and  (not A233) );
 a27696a <=( (not A232)  and  a27695a );
 a27700a <=( A299  and  (not A298) );
 a27701a <=( A266  and  a27700a );
 a27702a <=( a27701a  and  a27696a );
 a27706a <=( A167  and  (not A169) );
 a27707a <=( A170  and  a27706a );
 a27711a <=( (not A201)  and  (not A200) );
 a27712a <=( (not A166)  and  a27711a );
 a27713a <=( a27712a  and  a27707a );
 a27717a <=( (not A266)  and  (not A233) );
 a27718a <=( (not A232)  and  a27717a );
 a27722a <=( A299  and  (not A298) );
 a27723a <=( (not A267)  and  a27722a );
 a27724a <=( a27723a  and  a27718a );
 a27728a <=( A167  and  (not A169) );
 a27729a <=( A170  and  a27728a );
 a27733a <=( (not A201)  and  (not A200) );
 a27734a <=( (not A166)  and  a27733a );
 a27735a <=( a27734a  and  a27729a );
 a27739a <=( (not A265)  and  (not A233) );
 a27740a <=( (not A232)  and  a27739a );
 a27744a <=( A299  and  (not A298) );
 a27745a <=( (not A266)  and  a27744a );
 a27746a <=( a27745a  and  a27740a );
 a27750a <=( A167  and  (not A169) );
 a27751a <=( A170  and  a27750a );
 a27755a <=( (not A200)  and  (not A199) );
 a27756a <=( (not A166)  and  a27755a );
 a27757a <=( a27756a  and  a27751a );
 a27761a <=( A265  and  A233 );
 a27762a <=( A232  and  a27761a );
 a27766a <=( A299  and  (not A298) );
 a27767a <=( (not A267)  and  a27766a );
 a27768a <=( a27767a  and  a27762a );
 a27772a <=( A167  and  (not A169) );
 a27773a <=( A170  and  a27772a );
 a27777a <=( (not A200)  and  (not A199) );
 a27778a <=( (not A166)  and  a27777a );
 a27779a <=( a27778a  and  a27773a );
 a27783a <=( A265  and  A233 );
 a27784a <=( A232  and  a27783a );
 a27788a <=( A299  and  (not A298) );
 a27789a <=( A266  and  a27788a );
 a27790a <=( a27789a  and  a27784a );
 a27794a <=( A167  and  (not A169) );
 a27795a <=( A170  and  a27794a );
 a27799a <=( (not A200)  and  (not A199) );
 a27800a <=( (not A166)  and  a27799a );
 a27801a <=( a27800a  and  a27795a );
 a27805a <=( (not A265)  and  A233 );
 a27806a <=( A232  and  a27805a );
 a27810a <=( A299  and  (not A298) );
 a27811a <=( (not A266)  and  a27810a );
 a27812a <=( a27811a  and  a27806a );
 a27816a <=( A167  and  (not A169) );
 a27817a <=( A170  and  a27816a );
 a27821a <=( (not A200)  and  (not A199) );
 a27822a <=( (not A166)  and  a27821a );
 a27823a <=( a27822a  and  a27817a );
 a27827a <=( A265  and  A233 );
 a27828a <=( (not A232)  and  a27827a );
 a27832a <=( A268  and  A267 );
 a27833a <=( (not A266)  and  a27832a );
 a27834a <=( a27833a  and  a27828a );
 a27838a <=( A167  and  (not A169) );
 a27839a <=( A170  and  a27838a );
 a27843a <=( (not A200)  and  (not A199) );
 a27844a <=( (not A166)  and  a27843a );
 a27845a <=( a27844a  and  a27839a );
 a27849a <=( A265  and  A233 );
 a27850a <=( (not A232)  and  a27849a );
 a27854a <=( A269  and  A267 );
 a27855a <=( (not A266)  and  a27854a );
 a27856a <=( a27855a  and  a27850a );
 a27860a <=( A167  and  (not A169) );
 a27861a <=( A170  and  a27860a );
 a27865a <=( (not A200)  and  (not A199) );
 a27866a <=( (not A166)  and  a27865a );
 a27867a <=( a27866a  and  a27861a );
 a27871a <=( A265  and  (not A234) );
 a27872a <=( (not A233)  and  a27871a );
 a27876a <=( A299  and  (not A298) );
 a27877a <=( A266  and  a27876a );
 a27878a <=( a27877a  and  a27872a );
 a27882a <=( A167  and  (not A169) );
 a27883a <=( A170  and  a27882a );
 a27887a <=( (not A200)  and  (not A199) );
 a27888a <=( (not A166)  and  a27887a );
 a27889a <=( a27888a  and  a27883a );
 a27893a <=( (not A266)  and  (not A234) );
 a27894a <=( (not A233)  and  a27893a );
 a27898a <=( A299  and  (not A298) );
 a27899a <=( (not A267)  and  a27898a );
 a27900a <=( a27899a  and  a27894a );
 a27904a <=( A167  and  (not A169) );
 a27905a <=( A170  and  a27904a );
 a27909a <=( (not A200)  and  (not A199) );
 a27910a <=( (not A166)  and  a27909a );
 a27911a <=( a27910a  and  a27905a );
 a27915a <=( (not A265)  and  (not A234) );
 a27916a <=( (not A233)  and  a27915a );
 a27920a <=( A299  and  (not A298) );
 a27921a <=( (not A266)  and  a27920a );
 a27922a <=( a27921a  and  a27916a );
 a27926a <=( A167  and  (not A169) );
 a27927a <=( A170  and  a27926a );
 a27931a <=( (not A200)  and  (not A199) );
 a27932a <=( (not A166)  and  a27931a );
 a27933a <=( a27932a  and  a27927a );
 a27937a <=( A234  and  (not A233) );
 a27938a <=( A232  and  a27937a );
 a27942a <=( (not A300)  and  A298 );
 a27943a <=( A235  and  a27942a );
 a27944a <=( a27943a  and  a27938a );
 a27948a <=( A167  and  (not A169) );
 a27949a <=( A170  and  a27948a );
 a27953a <=( (not A200)  and  (not A199) );
 a27954a <=( (not A166)  and  a27953a );
 a27955a <=( a27954a  and  a27949a );
 a27959a <=( A234  and  (not A233) );
 a27960a <=( A232  and  a27959a );
 a27964a <=( A299  and  A298 );
 a27965a <=( A235  and  a27964a );
 a27966a <=( a27965a  and  a27960a );
 a27970a <=( A167  and  (not A169) );
 a27971a <=( A170  and  a27970a );
 a27975a <=( (not A200)  and  (not A199) );
 a27976a <=( (not A166)  and  a27975a );
 a27977a <=( a27976a  and  a27971a );
 a27981a <=( A234  and  (not A233) );
 a27982a <=( A232  and  a27981a );
 a27986a <=( (not A299)  and  (not A298) );
 a27987a <=( A235  and  a27986a );
 a27988a <=( a27987a  and  a27982a );
 a27992a <=( A167  and  (not A169) );
 a27993a <=( A170  and  a27992a );
 a27997a <=( (not A200)  and  (not A199) );
 a27998a <=( (not A166)  and  a27997a );
 a27999a <=( a27998a  and  a27993a );
 a28003a <=( A234  and  (not A233) );
 a28004a <=( A232  and  a28003a );
 a28008a <=( A266  and  (not A265) );
 a28009a <=( A235  and  a28008a );
 a28010a <=( a28009a  and  a28004a );
 a28014a <=( A167  and  (not A169) );
 a28015a <=( A170  and  a28014a );
 a28019a <=( (not A200)  and  (not A199) );
 a28020a <=( (not A166)  and  a28019a );
 a28021a <=( a28020a  and  a28015a );
 a28025a <=( A234  and  (not A233) );
 a28026a <=( A232  and  a28025a );
 a28030a <=( (not A300)  and  A298 );
 a28031a <=( A236  and  a28030a );
 a28032a <=( a28031a  and  a28026a );
 a28036a <=( A167  and  (not A169) );
 a28037a <=( A170  and  a28036a );
 a28041a <=( (not A200)  and  (not A199) );
 a28042a <=( (not A166)  and  a28041a );
 a28043a <=( a28042a  and  a28037a );
 a28047a <=( A234  and  (not A233) );
 a28048a <=( A232  and  a28047a );
 a28052a <=( A299  and  A298 );
 a28053a <=( A236  and  a28052a );
 a28054a <=( a28053a  and  a28048a );
 a28058a <=( A167  and  (not A169) );
 a28059a <=( A170  and  a28058a );
 a28063a <=( (not A200)  and  (not A199) );
 a28064a <=( (not A166)  and  a28063a );
 a28065a <=( a28064a  and  a28059a );
 a28069a <=( A234  and  (not A233) );
 a28070a <=( A232  and  a28069a );
 a28074a <=( (not A299)  and  (not A298) );
 a28075a <=( A236  and  a28074a );
 a28076a <=( a28075a  and  a28070a );
 a28080a <=( A167  and  (not A169) );
 a28081a <=( A170  and  a28080a );
 a28085a <=( (not A200)  and  (not A199) );
 a28086a <=( (not A166)  and  a28085a );
 a28087a <=( a28086a  and  a28081a );
 a28091a <=( A234  and  (not A233) );
 a28092a <=( A232  and  a28091a );
 a28096a <=( A266  and  (not A265) );
 a28097a <=( A236  and  a28096a );
 a28098a <=( a28097a  and  a28092a );
 a28102a <=( A167  and  (not A169) );
 a28103a <=( A170  and  a28102a );
 a28107a <=( (not A200)  and  (not A199) );
 a28108a <=( (not A166)  and  a28107a );
 a28109a <=( a28108a  and  a28103a );
 a28113a <=( A265  and  (not A233) );
 a28114a <=( (not A232)  and  a28113a );
 a28118a <=( A299  and  (not A298) );
 a28119a <=( A266  and  a28118a );
 a28120a <=( a28119a  and  a28114a );
 a28124a <=( A167  and  (not A169) );
 a28125a <=( A170  and  a28124a );
 a28129a <=( (not A200)  and  (not A199) );
 a28130a <=( (not A166)  and  a28129a );
 a28131a <=( a28130a  and  a28125a );
 a28135a <=( (not A266)  and  (not A233) );
 a28136a <=( (not A232)  and  a28135a );
 a28140a <=( A299  and  (not A298) );
 a28141a <=( (not A267)  and  a28140a );
 a28142a <=( a28141a  and  a28136a );
 a28146a <=( A167  and  (not A169) );
 a28147a <=( A170  and  a28146a );
 a28151a <=( (not A200)  and  (not A199) );
 a28152a <=( (not A166)  and  a28151a );
 a28153a <=( a28152a  and  a28147a );
 a28157a <=( (not A265)  and  (not A233) );
 a28158a <=( (not A232)  and  a28157a );
 a28162a <=( A299  and  (not A298) );
 a28163a <=( (not A266)  and  a28162a );
 a28164a <=( a28163a  and  a28158a );
 a28168a <=( (not A167)  and  (not A169) );
 a28169a <=( A170  and  a28168a );
 a28173a <=( A200  and  A199 );
 a28174a <=( A166  and  a28173a );
 a28175a <=( a28174a  and  a28169a );
 a28179a <=( A265  and  A233 );
 a28180a <=( A232  and  a28179a );
 a28184a <=( A299  and  (not A298) );
 a28185a <=( (not A267)  and  a28184a );
 a28186a <=( a28185a  and  a28180a );
 a28190a <=( (not A167)  and  (not A169) );
 a28191a <=( A170  and  a28190a );
 a28195a <=( A200  and  A199 );
 a28196a <=( A166  and  a28195a );
 a28197a <=( a28196a  and  a28191a );
 a28201a <=( A265  and  A233 );
 a28202a <=( A232  and  a28201a );
 a28206a <=( A299  and  (not A298) );
 a28207a <=( A266  and  a28206a );
 a28208a <=( a28207a  and  a28202a );
 a28212a <=( (not A167)  and  (not A169) );
 a28213a <=( A170  and  a28212a );
 a28217a <=( A200  and  A199 );
 a28218a <=( A166  and  a28217a );
 a28219a <=( a28218a  and  a28213a );
 a28223a <=( (not A265)  and  A233 );
 a28224a <=( A232  and  a28223a );
 a28228a <=( A299  and  (not A298) );
 a28229a <=( (not A266)  and  a28228a );
 a28230a <=( a28229a  and  a28224a );
 a28234a <=( (not A167)  and  (not A169) );
 a28235a <=( A170  and  a28234a );
 a28239a <=( A200  and  A199 );
 a28240a <=( A166  and  a28239a );
 a28241a <=( a28240a  and  a28235a );
 a28245a <=( A265  and  A233 );
 a28246a <=( (not A232)  and  a28245a );
 a28250a <=( A268  and  A267 );
 a28251a <=( (not A266)  and  a28250a );
 a28252a <=( a28251a  and  a28246a );
 a28256a <=( (not A167)  and  (not A169) );
 a28257a <=( A170  and  a28256a );
 a28261a <=( A200  and  A199 );
 a28262a <=( A166  and  a28261a );
 a28263a <=( a28262a  and  a28257a );
 a28267a <=( A265  and  A233 );
 a28268a <=( (not A232)  and  a28267a );
 a28272a <=( A269  and  A267 );
 a28273a <=( (not A266)  and  a28272a );
 a28274a <=( a28273a  and  a28268a );
 a28278a <=( (not A167)  and  (not A169) );
 a28279a <=( A170  and  a28278a );
 a28283a <=( A200  and  A199 );
 a28284a <=( A166  and  a28283a );
 a28285a <=( a28284a  and  a28279a );
 a28289a <=( A265  and  (not A234) );
 a28290a <=( (not A233)  and  a28289a );
 a28294a <=( A299  and  (not A298) );
 a28295a <=( A266  and  a28294a );
 a28296a <=( a28295a  and  a28290a );
 a28300a <=( (not A167)  and  (not A169) );
 a28301a <=( A170  and  a28300a );
 a28305a <=( A200  and  A199 );
 a28306a <=( A166  and  a28305a );
 a28307a <=( a28306a  and  a28301a );
 a28311a <=( (not A266)  and  (not A234) );
 a28312a <=( (not A233)  and  a28311a );
 a28316a <=( A299  and  (not A298) );
 a28317a <=( (not A267)  and  a28316a );
 a28318a <=( a28317a  and  a28312a );
 a28322a <=( (not A167)  and  (not A169) );
 a28323a <=( A170  and  a28322a );
 a28327a <=( A200  and  A199 );
 a28328a <=( A166  and  a28327a );
 a28329a <=( a28328a  and  a28323a );
 a28333a <=( (not A265)  and  (not A234) );
 a28334a <=( (not A233)  and  a28333a );
 a28338a <=( A299  and  (not A298) );
 a28339a <=( (not A266)  and  a28338a );
 a28340a <=( a28339a  and  a28334a );
 a28344a <=( (not A167)  and  (not A169) );
 a28345a <=( A170  and  a28344a );
 a28349a <=( A200  and  A199 );
 a28350a <=( A166  and  a28349a );
 a28351a <=( a28350a  and  a28345a );
 a28355a <=( A234  and  (not A233) );
 a28356a <=( A232  and  a28355a );
 a28360a <=( (not A300)  and  A298 );
 a28361a <=( A235  and  a28360a );
 a28362a <=( a28361a  and  a28356a );
 a28366a <=( (not A167)  and  (not A169) );
 a28367a <=( A170  and  a28366a );
 a28371a <=( A200  and  A199 );
 a28372a <=( A166  and  a28371a );
 a28373a <=( a28372a  and  a28367a );
 a28377a <=( A234  and  (not A233) );
 a28378a <=( A232  and  a28377a );
 a28382a <=( A299  and  A298 );
 a28383a <=( A235  and  a28382a );
 a28384a <=( a28383a  and  a28378a );
 a28388a <=( (not A167)  and  (not A169) );
 a28389a <=( A170  and  a28388a );
 a28393a <=( A200  and  A199 );
 a28394a <=( A166  and  a28393a );
 a28395a <=( a28394a  and  a28389a );
 a28399a <=( A234  and  (not A233) );
 a28400a <=( A232  and  a28399a );
 a28404a <=( (not A299)  and  (not A298) );
 a28405a <=( A235  and  a28404a );
 a28406a <=( a28405a  and  a28400a );
 a28410a <=( (not A167)  and  (not A169) );
 a28411a <=( A170  and  a28410a );
 a28415a <=( A200  and  A199 );
 a28416a <=( A166  and  a28415a );
 a28417a <=( a28416a  and  a28411a );
 a28421a <=( A234  and  (not A233) );
 a28422a <=( A232  and  a28421a );
 a28426a <=( A266  and  (not A265) );
 a28427a <=( A235  and  a28426a );
 a28428a <=( a28427a  and  a28422a );
 a28432a <=( (not A167)  and  (not A169) );
 a28433a <=( A170  and  a28432a );
 a28437a <=( A200  and  A199 );
 a28438a <=( A166  and  a28437a );
 a28439a <=( a28438a  and  a28433a );
 a28443a <=( A234  and  (not A233) );
 a28444a <=( A232  and  a28443a );
 a28448a <=( (not A300)  and  A298 );
 a28449a <=( A236  and  a28448a );
 a28450a <=( a28449a  and  a28444a );
 a28454a <=( (not A167)  and  (not A169) );
 a28455a <=( A170  and  a28454a );
 a28459a <=( A200  and  A199 );
 a28460a <=( A166  and  a28459a );
 a28461a <=( a28460a  and  a28455a );
 a28465a <=( A234  and  (not A233) );
 a28466a <=( A232  and  a28465a );
 a28470a <=( A299  and  A298 );
 a28471a <=( A236  and  a28470a );
 a28472a <=( a28471a  and  a28466a );
 a28476a <=( (not A167)  and  (not A169) );
 a28477a <=( A170  and  a28476a );
 a28481a <=( A200  and  A199 );
 a28482a <=( A166  and  a28481a );
 a28483a <=( a28482a  and  a28477a );
 a28487a <=( A234  and  (not A233) );
 a28488a <=( A232  and  a28487a );
 a28492a <=( (not A299)  and  (not A298) );
 a28493a <=( A236  and  a28492a );
 a28494a <=( a28493a  and  a28488a );
 a28498a <=( (not A167)  and  (not A169) );
 a28499a <=( A170  and  a28498a );
 a28503a <=( A200  and  A199 );
 a28504a <=( A166  and  a28503a );
 a28505a <=( a28504a  and  a28499a );
 a28509a <=( A234  and  (not A233) );
 a28510a <=( A232  and  a28509a );
 a28514a <=( A266  and  (not A265) );
 a28515a <=( A236  and  a28514a );
 a28516a <=( a28515a  and  a28510a );
 a28520a <=( (not A167)  and  (not A169) );
 a28521a <=( A170  and  a28520a );
 a28525a <=( A200  and  A199 );
 a28526a <=( A166  and  a28525a );
 a28527a <=( a28526a  and  a28521a );
 a28531a <=( A265  and  (not A233) );
 a28532a <=( (not A232)  and  a28531a );
 a28536a <=( A299  and  (not A298) );
 a28537a <=( A266  and  a28536a );
 a28538a <=( a28537a  and  a28532a );
 a28542a <=( (not A167)  and  (not A169) );
 a28543a <=( A170  and  a28542a );
 a28547a <=( A200  and  A199 );
 a28548a <=( A166  and  a28547a );
 a28549a <=( a28548a  and  a28543a );
 a28553a <=( (not A266)  and  (not A233) );
 a28554a <=( (not A232)  and  a28553a );
 a28558a <=( A299  and  (not A298) );
 a28559a <=( (not A267)  and  a28558a );
 a28560a <=( a28559a  and  a28554a );
 a28564a <=( (not A167)  and  (not A169) );
 a28565a <=( A170  and  a28564a );
 a28569a <=( A200  and  A199 );
 a28570a <=( A166  and  a28569a );
 a28571a <=( a28570a  and  a28565a );
 a28575a <=( (not A265)  and  (not A233) );
 a28576a <=( (not A232)  and  a28575a );
 a28580a <=( A299  and  (not A298) );
 a28581a <=( (not A266)  and  a28580a );
 a28582a <=( a28581a  and  a28576a );
 a28586a <=( (not A167)  and  (not A169) );
 a28587a <=( A170  and  a28586a );
 a28591a <=( (not A202)  and  (not A200) );
 a28592a <=( A166  and  a28591a );
 a28593a <=( a28592a  and  a28587a );
 a28597a <=( A233  and  (not A232) );
 a28598a <=( (not A203)  and  a28597a );
 a28602a <=( (not A302)  and  (not A301) );
 a28603a <=( (not A299)  and  a28602a );
 a28604a <=( a28603a  and  a28598a );
 a28608a <=( (not A167)  and  (not A169) );
 a28609a <=( A170  and  a28608a );
 a28613a <=( (not A201)  and  (not A200) );
 a28614a <=( A166  and  a28613a );
 a28615a <=( a28614a  and  a28609a );
 a28619a <=( A265  and  A233 );
 a28620a <=( A232  and  a28619a );
 a28624a <=( A299  and  (not A298) );
 a28625a <=( (not A267)  and  a28624a );
 a28626a <=( a28625a  and  a28620a );
 a28630a <=( (not A167)  and  (not A169) );
 a28631a <=( A170  and  a28630a );
 a28635a <=( (not A201)  and  (not A200) );
 a28636a <=( A166  and  a28635a );
 a28637a <=( a28636a  and  a28631a );
 a28641a <=( A265  and  A233 );
 a28642a <=( A232  and  a28641a );
 a28646a <=( A299  and  (not A298) );
 a28647a <=( A266  and  a28646a );
 a28648a <=( a28647a  and  a28642a );
 a28652a <=( (not A167)  and  (not A169) );
 a28653a <=( A170  and  a28652a );
 a28657a <=( (not A201)  and  (not A200) );
 a28658a <=( A166  and  a28657a );
 a28659a <=( a28658a  and  a28653a );
 a28663a <=( (not A265)  and  A233 );
 a28664a <=( A232  and  a28663a );
 a28668a <=( A299  and  (not A298) );
 a28669a <=( (not A266)  and  a28668a );
 a28670a <=( a28669a  and  a28664a );
 a28674a <=( (not A167)  and  (not A169) );
 a28675a <=( A170  and  a28674a );
 a28679a <=( (not A201)  and  (not A200) );
 a28680a <=( A166  and  a28679a );
 a28681a <=( a28680a  and  a28675a );
 a28685a <=( A265  and  A233 );
 a28686a <=( (not A232)  and  a28685a );
 a28690a <=( A268  and  A267 );
 a28691a <=( (not A266)  and  a28690a );
 a28692a <=( a28691a  and  a28686a );
 a28696a <=( (not A167)  and  (not A169) );
 a28697a <=( A170  and  a28696a );
 a28701a <=( (not A201)  and  (not A200) );
 a28702a <=( A166  and  a28701a );
 a28703a <=( a28702a  and  a28697a );
 a28707a <=( A265  and  A233 );
 a28708a <=( (not A232)  and  a28707a );
 a28712a <=( A269  and  A267 );
 a28713a <=( (not A266)  and  a28712a );
 a28714a <=( a28713a  and  a28708a );
 a28718a <=( (not A167)  and  (not A169) );
 a28719a <=( A170  and  a28718a );
 a28723a <=( (not A201)  and  (not A200) );
 a28724a <=( A166  and  a28723a );
 a28725a <=( a28724a  and  a28719a );
 a28729a <=( A265  and  (not A234) );
 a28730a <=( (not A233)  and  a28729a );
 a28734a <=( A299  and  (not A298) );
 a28735a <=( A266  and  a28734a );
 a28736a <=( a28735a  and  a28730a );
 a28740a <=( (not A167)  and  (not A169) );
 a28741a <=( A170  and  a28740a );
 a28745a <=( (not A201)  and  (not A200) );
 a28746a <=( A166  and  a28745a );
 a28747a <=( a28746a  and  a28741a );
 a28751a <=( (not A266)  and  (not A234) );
 a28752a <=( (not A233)  and  a28751a );
 a28756a <=( A299  and  (not A298) );
 a28757a <=( (not A267)  and  a28756a );
 a28758a <=( a28757a  and  a28752a );
 a28762a <=( (not A167)  and  (not A169) );
 a28763a <=( A170  and  a28762a );
 a28767a <=( (not A201)  and  (not A200) );
 a28768a <=( A166  and  a28767a );
 a28769a <=( a28768a  and  a28763a );
 a28773a <=( (not A265)  and  (not A234) );
 a28774a <=( (not A233)  and  a28773a );
 a28778a <=( A299  and  (not A298) );
 a28779a <=( (not A266)  and  a28778a );
 a28780a <=( a28779a  and  a28774a );
 a28784a <=( (not A167)  and  (not A169) );
 a28785a <=( A170  and  a28784a );
 a28789a <=( (not A201)  and  (not A200) );
 a28790a <=( A166  and  a28789a );
 a28791a <=( a28790a  and  a28785a );
 a28795a <=( A234  and  (not A233) );
 a28796a <=( A232  and  a28795a );
 a28800a <=( (not A300)  and  A298 );
 a28801a <=( A235  and  a28800a );
 a28802a <=( a28801a  and  a28796a );
 a28806a <=( (not A167)  and  (not A169) );
 a28807a <=( A170  and  a28806a );
 a28811a <=( (not A201)  and  (not A200) );
 a28812a <=( A166  and  a28811a );
 a28813a <=( a28812a  and  a28807a );
 a28817a <=( A234  and  (not A233) );
 a28818a <=( A232  and  a28817a );
 a28822a <=( A299  and  A298 );
 a28823a <=( A235  and  a28822a );
 a28824a <=( a28823a  and  a28818a );
 a28828a <=( (not A167)  and  (not A169) );
 a28829a <=( A170  and  a28828a );
 a28833a <=( (not A201)  and  (not A200) );
 a28834a <=( A166  and  a28833a );
 a28835a <=( a28834a  and  a28829a );
 a28839a <=( A234  and  (not A233) );
 a28840a <=( A232  and  a28839a );
 a28844a <=( (not A299)  and  (not A298) );
 a28845a <=( A235  and  a28844a );
 a28846a <=( a28845a  and  a28840a );
 a28850a <=( (not A167)  and  (not A169) );
 a28851a <=( A170  and  a28850a );
 a28855a <=( (not A201)  and  (not A200) );
 a28856a <=( A166  and  a28855a );
 a28857a <=( a28856a  and  a28851a );
 a28861a <=( A234  and  (not A233) );
 a28862a <=( A232  and  a28861a );
 a28866a <=( A266  and  (not A265) );
 a28867a <=( A235  and  a28866a );
 a28868a <=( a28867a  and  a28862a );
 a28872a <=( (not A167)  and  (not A169) );
 a28873a <=( A170  and  a28872a );
 a28877a <=( (not A201)  and  (not A200) );
 a28878a <=( A166  and  a28877a );
 a28879a <=( a28878a  and  a28873a );
 a28883a <=( A234  and  (not A233) );
 a28884a <=( A232  and  a28883a );
 a28888a <=( (not A300)  and  A298 );
 a28889a <=( A236  and  a28888a );
 a28890a <=( a28889a  and  a28884a );
 a28894a <=( (not A167)  and  (not A169) );
 a28895a <=( A170  and  a28894a );
 a28899a <=( (not A201)  and  (not A200) );
 a28900a <=( A166  and  a28899a );
 a28901a <=( a28900a  and  a28895a );
 a28905a <=( A234  and  (not A233) );
 a28906a <=( A232  and  a28905a );
 a28910a <=( A299  and  A298 );
 a28911a <=( A236  and  a28910a );
 a28912a <=( a28911a  and  a28906a );
 a28916a <=( (not A167)  and  (not A169) );
 a28917a <=( A170  and  a28916a );
 a28921a <=( (not A201)  and  (not A200) );
 a28922a <=( A166  and  a28921a );
 a28923a <=( a28922a  and  a28917a );
 a28927a <=( A234  and  (not A233) );
 a28928a <=( A232  and  a28927a );
 a28932a <=( (not A299)  and  (not A298) );
 a28933a <=( A236  and  a28932a );
 a28934a <=( a28933a  and  a28928a );
 a28938a <=( (not A167)  and  (not A169) );
 a28939a <=( A170  and  a28938a );
 a28943a <=( (not A201)  and  (not A200) );
 a28944a <=( A166  and  a28943a );
 a28945a <=( a28944a  and  a28939a );
 a28949a <=( A234  and  (not A233) );
 a28950a <=( A232  and  a28949a );
 a28954a <=( A266  and  (not A265) );
 a28955a <=( A236  and  a28954a );
 a28956a <=( a28955a  and  a28950a );
 a28960a <=( (not A167)  and  (not A169) );
 a28961a <=( A170  and  a28960a );
 a28965a <=( (not A201)  and  (not A200) );
 a28966a <=( A166  and  a28965a );
 a28967a <=( a28966a  and  a28961a );
 a28971a <=( A265  and  (not A233) );
 a28972a <=( (not A232)  and  a28971a );
 a28976a <=( A299  and  (not A298) );
 a28977a <=( A266  and  a28976a );
 a28978a <=( a28977a  and  a28972a );
 a28982a <=( (not A167)  and  (not A169) );
 a28983a <=( A170  and  a28982a );
 a28987a <=( (not A201)  and  (not A200) );
 a28988a <=( A166  and  a28987a );
 a28989a <=( a28988a  and  a28983a );
 a28993a <=( (not A266)  and  (not A233) );
 a28994a <=( (not A232)  and  a28993a );
 a28998a <=( A299  and  (not A298) );
 a28999a <=( (not A267)  and  a28998a );
 a29000a <=( a28999a  and  a28994a );
 a29004a <=( (not A167)  and  (not A169) );
 a29005a <=( A170  and  a29004a );
 a29009a <=( (not A201)  and  (not A200) );
 a29010a <=( A166  and  a29009a );
 a29011a <=( a29010a  and  a29005a );
 a29015a <=( (not A265)  and  (not A233) );
 a29016a <=( (not A232)  and  a29015a );
 a29020a <=( A299  and  (not A298) );
 a29021a <=( (not A266)  and  a29020a );
 a29022a <=( a29021a  and  a29016a );
 a29026a <=( (not A167)  and  (not A169) );
 a29027a <=( A170  and  a29026a );
 a29031a <=( (not A200)  and  (not A199) );
 a29032a <=( A166  and  a29031a );
 a29033a <=( a29032a  and  a29027a );
 a29037a <=( A265  and  A233 );
 a29038a <=( A232  and  a29037a );
 a29042a <=( A299  and  (not A298) );
 a29043a <=( (not A267)  and  a29042a );
 a29044a <=( a29043a  and  a29038a );
 a29048a <=( (not A167)  and  (not A169) );
 a29049a <=( A170  and  a29048a );
 a29053a <=( (not A200)  and  (not A199) );
 a29054a <=( A166  and  a29053a );
 a29055a <=( a29054a  and  a29049a );
 a29059a <=( A265  and  A233 );
 a29060a <=( A232  and  a29059a );
 a29064a <=( A299  and  (not A298) );
 a29065a <=( A266  and  a29064a );
 a29066a <=( a29065a  and  a29060a );
 a29070a <=( (not A167)  and  (not A169) );
 a29071a <=( A170  and  a29070a );
 a29075a <=( (not A200)  and  (not A199) );
 a29076a <=( A166  and  a29075a );
 a29077a <=( a29076a  and  a29071a );
 a29081a <=( (not A265)  and  A233 );
 a29082a <=( A232  and  a29081a );
 a29086a <=( A299  and  (not A298) );
 a29087a <=( (not A266)  and  a29086a );
 a29088a <=( a29087a  and  a29082a );
 a29092a <=( (not A167)  and  (not A169) );
 a29093a <=( A170  and  a29092a );
 a29097a <=( (not A200)  and  (not A199) );
 a29098a <=( A166  and  a29097a );
 a29099a <=( a29098a  and  a29093a );
 a29103a <=( A265  and  A233 );
 a29104a <=( (not A232)  and  a29103a );
 a29108a <=( A268  and  A267 );
 a29109a <=( (not A266)  and  a29108a );
 a29110a <=( a29109a  and  a29104a );
 a29114a <=( (not A167)  and  (not A169) );
 a29115a <=( A170  and  a29114a );
 a29119a <=( (not A200)  and  (not A199) );
 a29120a <=( A166  and  a29119a );
 a29121a <=( a29120a  and  a29115a );
 a29125a <=( A265  and  A233 );
 a29126a <=( (not A232)  and  a29125a );
 a29130a <=( A269  and  A267 );
 a29131a <=( (not A266)  and  a29130a );
 a29132a <=( a29131a  and  a29126a );
 a29136a <=( (not A167)  and  (not A169) );
 a29137a <=( A170  and  a29136a );
 a29141a <=( (not A200)  and  (not A199) );
 a29142a <=( A166  and  a29141a );
 a29143a <=( a29142a  and  a29137a );
 a29147a <=( A265  and  (not A234) );
 a29148a <=( (not A233)  and  a29147a );
 a29152a <=( A299  and  (not A298) );
 a29153a <=( A266  and  a29152a );
 a29154a <=( a29153a  and  a29148a );
 a29158a <=( (not A167)  and  (not A169) );
 a29159a <=( A170  and  a29158a );
 a29163a <=( (not A200)  and  (not A199) );
 a29164a <=( A166  and  a29163a );
 a29165a <=( a29164a  and  a29159a );
 a29169a <=( (not A266)  and  (not A234) );
 a29170a <=( (not A233)  and  a29169a );
 a29174a <=( A299  and  (not A298) );
 a29175a <=( (not A267)  and  a29174a );
 a29176a <=( a29175a  and  a29170a );
 a29180a <=( (not A167)  and  (not A169) );
 a29181a <=( A170  and  a29180a );
 a29185a <=( (not A200)  and  (not A199) );
 a29186a <=( A166  and  a29185a );
 a29187a <=( a29186a  and  a29181a );
 a29191a <=( (not A265)  and  (not A234) );
 a29192a <=( (not A233)  and  a29191a );
 a29196a <=( A299  and  (not A298) );
 a29197a <=( (not A266)  and  a29196a );
 a29198a <=( a29197a  and  a29192a );
 a29202a <=( (not A167)  and  (not A169) );
 a29203a <=( A170  and  a29202a );
 a29207a <=( (not A200)  and  (not A199) );
 a29208a <=( A166  and  a29207a );
 a29209a <=( a29208a  and  a29203a );
 a29213a <=( A234  and  (not A233) );
 a29214a <=( A232  and  a29213a );
 a29218a <=( (not A300)  and  A298 );
 a29219a <=( A235  and  a29218a );
 a29220a <=( a29219a  and  a29214a );
 a29224a <=( (not A167)  and  (not A169) );
 a29225a <=( A170  and  a29224a );
 a29229a <=( (not A200)  and  (not A199) );
 a29230a <=( A166  and  a29229a );
 a29231a <=( a29230a  and  a29225a );
 a29235a <=( A234  and  (not A233) );
 a29236a <=( A232  and  a29235a );
 a29240a <=( A299  and  A298 );
 a29241a <=( A235  and  a29240a );
 a29242a <=( a29241a  and  a29236a );
 a29246a <=( (not A167)  and  (not A169) );
 a29247a <=( A170  and  a29246a );
 a29251a <=( (not A200)  and  (not A199) );
 a29252a <=( A166  and  a29251a );
 a29253a <=( a29252a  and  a29247a );
 a29257a <=( A234  and  (not A233) );
 a29258a <=( A232  and  a29257a );
 a29262a <=( (not A299)  and  (not A298) );
 a29263a <=( A235  and  a29262a );
 a29264a <=( a29263a  and  a29258a );
 a29268a <=( (not A167)  and  (not A169) );
 a29269a <=( A170  and  a29268a );
 a29273a <=( (not A200)  and  (not A199) );
 a29274a <=( A166  and  a29273a );
 a29275a <=( a29274a  and  a29269a );
 a29279a <=( A234  and  (not A233) );
 a29280a <=( A232  and  a29279a );
 a29284a <=( A266  and  (not A265) );
 a29285a <=( A235  and  a29284a );
 a29286a <=( a29285a  and  a29280a );
 a29290a <=( (not A167)  and  (not A169) );
 a29291a <=( A170  and  a29290a );
 a29295a <=( (not A200)  and  (not A199) );
 a29296a <=( A166  and  a29295a );
 a29297a <=( a29296a  and  a29291a );
 a29301a <=( A234  and  (not A233) );
 a29302a <=( A232  and  a29301a );
 a29306a <=( (not A300)  and  A298 );
 a29307a <=( A236  and  a29306a );
 a29308a <=( a29307a  and  a29302a );
 a29312a <=( (not A167)  and  (not A169) );
 a29313a <=( A170  and  a29312a );
 a29317a <=( (not A200)  and  (not A199) );
 a29318a <=( A166  and  a29317a );
 a29319a <=( a29318a  and  a29313a );
 a29323a <=( A234  and  (not A233) );
 a29324a <=( A232  and  a29323a );
 a29328a <=( A299  and  A298 );
 a29329a <=( A236  and  a29328a );
 a29330a <=( a29329a  and  a29324a );
 a29334a <=( (not A167)  and  (not A169) );
 a29335a <=( A170  and  a29334a );
 a29339a <=( (not A200)  and  (not A199) );
 a29340a <=( A166  and  a29339a );
 a29341a <=( a29340a  and  a29335a );
 a29345a <=( A234  and  (not A233) );
 a29346a <=( A232  and  a29345a );
 a29350a <=( (not A299)  and  (not A298) );
 a29351a <=( A236  and  a29350a );
 a29352a <=( a29351a  and  a29346a );
 a29356a <=( (not A167)  and  (not A169) );
 a29357a <=( A170  and  a29356a );
 a29361a <=( (not A200)  and  (not A199) );
 a29362a <=( A166  and  a29361a );
 a29363a <=( a29362a  and  a29357a );
 a29367a <=( A234  and  (not A233) );
 a29368a <=( A232  and  a29367a );
 a29372a <=( A266  and  (not A265) );
 a29373a <=( A236  and  a29372a );
 a29374a <=( a29373a  and  a29368a );
 a29378a <=( (not A167)  and  (not A169) );
 a29379a <=( A170  and  a29378a );
 a29383a <=( (not A200)  and  (not A199) );
 a29384a <=( A166  and  a29383a );
 a29385a <=( a29384a  and  a29379a );
 a29389a <=( A265  and  (not A233) );
 a29390a <=( (not A232)  and  a29389a );
 a29394a <=( A299  and  (not A298) );
 a29395a <=( A266  and  a29394a );
 a29396a <=( a29395a  and  a29390a );
 a29400a <=( (not A167)  and  (not A169) );
 a29401a <=( A170  and  a29400a );
 a29405a <=( (not A200)  and  (not A199) );
 a29406a <=( A166  and  a29405a );
 a29407a <=( a29406a  and  a29401a );
 a29411a <=( (not A266)  and  (not A233) );
 a29412a <=( (not A232)  and  a29411a );
 a29416a <=( A299  and  (not A298) );
 a29417a <=( (not A267)  and  a29416a );
 a29418a <=( a29417a  and  a29412a );
 a29422a <=( (not A167)  and  (not A169) );
 a29423a <=( A170  and  a29422a );
 a29427a <=( (not A200)  and  (not A199) );
 a29428a <=( A166  and  a29427a );
 a29429a <=( a29428a  and  a29423a );
 a29433a <=( (not A265)  and  (not A233) );
 a29434a <=( (not A232)  and  a29433a );
 a29438a <=( A299  and  (not A298) );
 a29439a <=( (not A266)  and  a29438a );
 a29440a <=( a29439a  and  a29434a );
 a29444a <=( (not A168)  and  (not A169) );
 a29445a <=( (not A170)  and  a29444a );
 a29449a <=( A201  and  (not A200) );
 a29450a <=( A199  and  a29449a );
 a29451a <=( a29450a  and  a29445a );
 a29455a <=( A233  and  (not A232) );
 a29456a <=( A202  and  a29455a );
 a29460a <=( (not A302)  and  (not A301) );
 a29461a <=( (not A299)  and  a29460a );
 a29462a <=( a29461a  and  a29456a );
 a29466a <=( (not A168)  and  (not A169) );
 a29467a <=( (not A170)  and  a29466a );
 a29471a <=( A201  and  (not A200) );
 a29472a <=( A199  and  a29471a );
 a29473a <=( a29472a  and  a29467a );
 a29477a <=( A233  and  (not A232) );
 a29478a <=( A203  and  a29477a );
 a29482a <=( (not A302)  and  (not A301) );
 a29483a <=( (not A299)  and  a29482a );
 a29484a <=( a29483a  and  a29478a );
 a29488a <=( A199  and  A166 );
 a29489a <=( A168  and  a29488a );
 a29493a <=( A233  and  A232 );
 a29494a <=( A200  and  a29493a );
 a29495a <=( a29494a  and  a29489a );
 a29499a <=( (not A269)  and  (not A268) );
 a29500a <=( A265  and  a29499a );
 a29503a <=( (not A299)  and  A298 );
 a29506a <=( A301  and  A300 );
 a29507a <=( a29506a  and  a29503a );
 a29508a <=( a29507a  and  a29500a );
 a29512a <=( A199  and  A166 );
 a29513a <=( A168  and  a29512a );
 a29517a <=( A233  and  A232 );
 a29518a <=( A200  and  a29517a );
 a29519a <=( a29518a  and  a29513a );
 a29523a <=( (not A269)  and  (not A268) );
 a29524a <=( A265  and  a29523a );
 a29527a <=( (not A299)  and  A298 );
 a29530a <=( A302  and  A300 );
 a29531a <=( a29530a  and  a29527a );
 a29532a <=( a29531a  and  a29524a );
 a29536a <=( A199  and  A166 );
 a29537a <=( A168  and  a29536a );
 a29541a <=( (not A235)  and  (not A233) );
 a29542a <=( A200  and  a29541a );
 a29543a <=( a29542a  and  a29537a );
 a29547a <=( A266  and  A265 );
 a29548a <=( (not A236)  and  a29547a );
 a29551a <=( (not A299)  and  A298 );
 a29554a <=( A301  and  A300 );
 a29555a <=( a29554a  and  a29551a );
 a29556a <=( a29555a  and  a29548a );
 a29560a <=( A199  and  A166 );
 a29561a <=( A168  and  a29560a );
 a29565a <=( (not A235)  and  (not A233) );
 a29566a <=( A200  and  a29565a );
 a29567a <=( a29566a  and  a29561a );
 a29571a <=( A266  and  A265 );
 a29572a <=( (not A236)  and  a29571a );
 a29575a <=( (not A299)  and  A298 );
 a29578a <=( A302  and  A300 );
 a29579a <=( a29578a  and  a29575a );
 a29580a <=( a29579a  and  a29572a );
 a29584a <=( A199  and  A166 );
 a29585a <=( A168  and  a29584a );
 a29589a <=( (not A235)  and  (not A233) );
 a29590a <=( A200  and  a29589a );
 a29591a <=( a29590a  and  a29585a );
 a29595a <=( (not A267)  and  (not A266) );
 a29596a <=( (not A236)  and  a29595a );
 a29599a <=( (not A299)  and  A298 );
 a29602a <=( A301  and  A300 );
 a29603a <=( a29602a  and  a29599a );
 a29604a <=( a29603a  and  a29596a );
 a29608a <=( A199  and  A166 );
 a29609a <=( A168  and  a29608a );
 a29613a <=( (not A235)  and  (not A233) );
 a29614a <=( A200  and  a29613a );
 a29615a <=( a29614a  and  a29609a );
 a29619a <=( (not A267)  and  (not A266) );
 a29620a <=( (not A236)  and  a29619a );
 a29623a <=( (not A299)  and  A298 );
 a29626a <=( A302  and  A300 );
 a29627a <=( a29626a  and  a29623a );
 a29628a <=( a29627a  and  a29620a );
 a29632a <=( A199  and  A166 );
 a29633a <=( A168  and  a29632a );
 a29637a <=( (not A235)  and  (not A233) );
 a29638a <=( A200  and  a29637a );
 a29639a <=( a29638a  and  a29633a );
 a29643a <=( (not A266)  and  (not A265) );
 a29644a <=( (not A236)  and  a29643a );
 a29647a <=( (not A299)  and  A298 );
 a29650a <=( A301  and  A300 );
 a29651a <=( a29650a  and  a29647a );
 a29652a <=( a29651a  and  a29644a );
 a29656a <=( A199  and  A166 );
 a29657a <=( A168  and  a29656a );
 a29661a <=( (not A235)  and  (not A233) );
 a29662a <=( A200  and  a29661a );
 a29663a <=( a29662a  and  a29657a );
 a29667a <=( (not A266)  and  (not A265) );
 a29668a <=( (not A236)  and  a29667a );
 a29671a <=( (not A299)  and  A298 );
 a29674a <=( A302  and  A300 );
 a29675a <=( a29674a  and  a29671a );
 a29676a <=( a29675a  and  a29668a );
 a29680a <=( A199  and  A166 );
 a29681a <=( A168  and  a29680a );
 a29685a <=( (not A234)  and  (not A233) );
 a29686a <=( A200  and  a29685a );
 a29687a <=( a29686a  and  a29681a );
 a29691a <=( (not A269)  and  (not A268) );
 a29692a <=( (not A266)  and  a29691a );
 a29695a <=( (not A299)  and  A298 );
 a29698a <=( A301  and  A300 );
 a29699a <=( a29698a  and  a29695a );
 a29700a <=( a29699a  and  a29692a );
 a29704a <=( A199  and  A166 );
 a29705a <=( A168  and  a29704a );
 a29709a <=( (not A234)  and  (not A233) );
 a29710a <=( A200  and  a29709a );
 a29711a <=( a29710a  and  a29705a );
 a29715a <=( (not A269)  and  (not A268) );
 a29716a <=( (not A266)  and  a29715a );
 a29719a <=( (not A299)  and  A298 );
 a29722a <=( A302  and  A300 );
 a29723a <=( a29722a  and  a29719a );
 a29724a <=( a29723a  and  a29716a );
 a29728a <=( A199  and  A166 );
 a29729a <=( A168  and  a29728a );
 a29733a <=( (not A233)  and  (not A232) );
 a29734a <=( A200  and  a29733a );
 a29735a <=( a29734a  and  a29729a );
 a29739a <=( (not A269)  and  (not A268) );
 a29740a <=( (not A266)  and  a29739a );
 a29743a <=( (not A299)  and  A298 );
 a29746a <=( A301  and  A300 );
 a29747a <=( a29746a  and  a29743a );
 a29748a <=( a29747a  and  a29740a );
 a29752a <=( A199  and  A166 );
 a29753a <=( A168  and  a29752a );
 a29757a <=( (not A233)  and  (not A232) );
 a29758a <=( A200  and  a29757a );
 a29759a <=( a29758a  and  a29753a );
 a29763a <=( (not A269)  and  (not A268) );
 a29764a <=( (not A266)  and  a29763a );
 a29767a <=( (not A299)  and  A298 );
 a29770a <=( A302  and  A300 );
 a29771a <=( a29770a  and  a29767a );
 a29772a <=( a29771a  and  a29764a );
 a29776a <=( (not A200)  and  A166 );
 a29777a <=( A168  and  a29776a );
 a29781a <=( A232  and  (not A203) );
 a29782a <=( (not A202)  and  a29781a );
 a29783a <=( a29782a  and  a29777a );
 a29787a <=( (not A267)  and  A265 );
 a29788a <=( A233  and  a29787a );
 a29791a <=( (not A299)  and  A298 );
 a29794a <=( A301  and  A300 );
 a29795a <=( a29794a  and  a29791a );
 a29796a <=( a29795a  and  a29788a );
 a29800a <=( (not A200)  and  A166 );
 a29801a <=( A168  and  a29800a );
 a29805a <=( A232  and  (not A203) );
 a29806a <=( (not A202)  and  a29805a );
 a29807a <=( a29806a  and  a29801a );
 a29811a <=( (not A267)  and  A265 );
 a29812a <=( A233  and  a29811a );
 a29815a <=( (not A299)  and  A298 );
 a29818a <=( A302  and  A300 );
 a29819a <=( a29818a  and  a29815a );
 a29820a <=( a29819a  and  a29812a );
 a29824a <=( (not A200)  and  A166 );
 a29825a <=( A168  and  a29824a );
 a29829a <=( A232  and  (not A203) );
 a29830a <=( (not A202)  and  a29829a );
 a29831a <=( a29830a  and  a29825a );
 a29835a <=( A266  and  A265 );
 a29836a <=( A233  and  a29835a );
 a29839a <=( (not A299)  and  A298 );
 a29842a <=( A301  and  A300 );
 a29843a <=( a29842a  and  a29839a );
 a29844a <=( a29843a  and  a29836a );
 a29848a <=( (not A200)  and  A166 );
 a29849a <=( A168  and  a29848a );
 a29853a <=( A232  and  (not A203) );
 a29854a <=( (not A202)  and  a29853a );
 a29855a <=( a29854a  and  a29849a );
 a29859a <=( A266  and  A265 );
 a29860a <=( A233  and  a29859a );
 a29863a <=( (not A299)  and  A298 );
 a29866a <=( A302  and  A300 );
 a29867a <=( a29866a  and  a29863a );
 a29868a <=( a29867a  and  a29860a );
 a29872a <=( (not A200)  and  A166 );
 a29873a <=( A168  and  a29872a );
 a29877a <=( A232  and  (not A203) );
 a29878a <=( (not A202)  and  a29877a );
 a29879a <=( a29878a  and  a29873a );
 a29883a <=( (not A266)  and  (not A265) );
 a29884a <=( A233  and  a29883a );
 a29887a <=( (not A299)  and  A298 );
 a29890a <=( A301  and  A300 );
 a29891a <=( a29890a  and  a29887a );
 a29892a <=( a29891a  and  a29884a );
 a29896a <=( (not A200)  and  A166 );
 a29897a <=( A168  and  a29896a );
 a29901a <=( A232  and  (not A203) );
 a29902a <=( (not A202)  and  a29901a );
 a29903a <=( a29902a  and  a29897a );
 a29907a <=( (not A266)  and  (not A265) );
 a29908a <=( A233  and  a29907a );
 a29911a <=( (not A299)  and  A298 );
 a29914a <=( A302  and  A300 );
 a29915a <=( a29914a  and  a29911a );
 a29916a <=( a29915a  and  a29908a );
 a29920a <=( (not A200)  and  A166 );
 a29921a <=( A168  and  a29920a );
 a29925a <=( (not A233)  and  (not A203) );
 a29926a <=( (not A202)  and  a29925a );
 a29927a <=( a29926a  and  a29921a );
 a29931a <=( (not A266)  and  (not A236) );
 a29932a <=( (not A235)  and  a29931a );
 a29935a <=( (not A269)  and  (not A268) );
 a29938a <=( A299  and  (not A298) );
 a29939a <=( a29938a  and  a29935a );
 a29940a <=( a29939a  and  a29932a );
 a29944a <=( (not A200)  and  A166 );
 a29945a <=( A168  and  a29944a );
 a29949a <=( (not A233)  and  (not A203) );
 a29950a <=( (not A202)  and  a29949a );
 a29951a <=( a29950a  and  a29945a );
 a29955a <=( A266  and  A265 );
 a29956a <=( (not A234)  and  a29955a );
 a29959a <=( (not A299)  and  A298 );
 a29962a <=( A301  and  A300 );
 a29963a <=( a29962a  and  a29959a );
 a29964a <=( a29963a  and  a29956a );
 a29968a <=( (not A200)  and  A166 );
 a29969a <=( A168  and  a29968a );
 a29973a <=( (not A233)  and  (not A203) );
 a29974a <=( (not A202)  and  a29973a );
 a29975a <=( a29974a  and  a29969a );
 a29979a <=( A266  and  A265 );
 a29980a <=( (not A234)  and  a29979a );
 a29983a <=( (not A299)  and  A298 );
 a29986a <=( A302  and  A300 );
 a29987a <=( a29986a  and  a29983a );
 a29988a <=( a29987a  and  a29980a );
 a29992a <=( (not A200)  and  A166 );
 a29993a <=( A168  and  a29992a );
 a29997a <=( (not A233)  and  (not A203) );
 a29998a <=( (not A202)  and  a29997a );
 a29999a <=( a29998a  and  a29993a );
 a30003a <=( (not A267)  and  (not A266) );
 a30004a <=( (not A234)  and  a30003a );
 a30007a <=( (not A299)  and  A298 );
 a30010a <=( A301  and  A300 );
 a30011a <=( a30010a  and  a30007a );
 a30012a <=( a30011a  and  a30004a );
 a30016a <=( (not A200)  and  A166 );
 a30017a <=( A168  and  a30016a );
 a30021a <=( (not A233)  and  (not A203) );
 a30022a <=( (not A202)  and  a30021a );
 a30023a <=( a30022a  and  a30017a );
 a30027a <=( (not A267)  and  (not A266) );
 a30028a <=( (not A234)  and  a30027a );
 a30031a <=( (not A299)  and  A298 );
 a30034a <=( A302  and  A300 );
 a30035a <=( a30034a  and  a30031a );
 a30036a <=( a30035a  and  a30028a );
 a30040a <=( (not A200)  and  A166 );
 a30041a <=( A168  and  a30040a );
 a30045a <=( (not A233)  and  (not A203) );
 a30046a <=( (not A202)  and  a30045a );
 a30047a <=( a30046a  and  a30041a );
 a30051a <=( (not A266)  and  (not A265) );
 a30052a <=( (not A234)  and  a30051a );
 a30055a <=( (not A299)  and  A298 );
 a30058a <=( A301  and  A300 );
 a30059a <=( a30058a  and  a30055a );
 a30060a <=( a30059a  and  a30052a );
 a30064a <=( (not A200)  and  A166 );
 a30065a <=( A168  and  a30064a );
 a30069a <=( (not A233)  and  (not A203) );
 a30070a <=( (not A202)  and  a30069a );
 a30071a <=( a30070a  and  a30065a );
 a30075a <=( (not A266)  and  (not A265) );
 a30076a <=( (not A234)  and  a30075a );
 a30079a <=( (not A299)  and  A298 );
 a30082a <=( A302  and  A300 );
 a30083a <=( a30082a  and  a30079a );
 a30084a <=( a30083a  and  a30076a );
 a30088a <=( (not A200)  and  A166 );
 a30089a <=( A168  and  a30088a );
 a30093a <=( A232  and  (not A203) );
 a30094a <=( (not A202)  and  a30093a );
 a30095a <=( a30094a  and  a30089a );
 a30099a <=( A235  and  A234 );
 a30100a <=( (not A233)  and  a30099a );
 a30103a <=( (not A266)  and  A265 );
 a30106a <=( A268  and  A267 );
 a30107a <=( a30106a  and  a30103a );
 a30108a <=( a30107a  and  a30100a );
 a30112a <=( (not A200)  and  A166 );
 a30113a <=( A168  and  a30112a );
 a30117a <=( A232  and  (not A203) );
 a30118a <=( (not A202)  and  a30117a );
 a30119a <=( a30118a  and  a30113a );
 a30123a <=( A235  and  A234 );
 a30124a <=( (not A233)  and  a30123a );
 a30127a <=( (not A266)  and  A265 );
 a30130a <=( A269  and  A267 );
 a30131a <=( a30130a  and  a30127a );
 a30132a <=( a30131a  and  a30124a );
 a30136a <=( (not A200)  and  A166 );
 a30137a <=( A168  and  a30136a );
 a30141a <=( A232  and  (not A203) );
 a30142a <=( (not A202)  and  a30141a );
 a30143a <=( a30142a  and  a30137a );
 a30147a <=( A236  and  A234 );
 a30148a <=( (not A233)  and  a30147a );
 a30151a <=( (not A266)  and  A265 );
 a30154a <=( A268  and  A267 );
 a30155a <=( a30154a  and  a30151a );
 a30156a <=( a30155a  and  a30148a );
 a30160a <=( (not A200)  and  A166 );
 a30161a <=( A168  and  a30160a );
 a30165a <=( A232  and  (not A203) );
 a30166a <=( (not A202)  and  a30165a );
 a30167a <=( a30166a  and  a30161a );
 a30171a <=( A236  and  A234 );
 a30172a <=( (not A233)  and  a30171a );
 a30175a <=( (not A266)  and  A265 );
 a30178a <=( A269  and  A267 );
 a30179a <=( a30178a  and  a30175a );
 a30180a <=( a30179a  and  a30172a );
 a30184a <=( (not A200)  and  A166 );
 a30185a <=( A168  and  a30184a );
 a30189a <=( (not A232)  and  (not A203) );
 a30190a <=( (not A202)  and  a30189a );
 a30191a <=( a30190a  and  a30185a );
 a30195a <=( A266  and  A265 );
 a30196a <=( (not A233)  and  a30195a );
 a30199a <=( (not A299)  and  A298 );
 a30202a <=( A301  and  A300 );
 a30203a <=( a30202a  and  a30199a );
 a30204a <=( a30203a  and  a30196a );
 a30208a <=( (not A200)  and  A166 );
 a30209a <=( A168  and  a30208a );
 a30213a <=( (not A232)  and  (not A203) );
 a30214a <=( (not A202)  and  a30213a );
 a30215a <=( a30214a  and  a30209a );
 a30219a <=( A266  and  A265 );
 a30220a <=( (not A233)  and  a30219a );
 a30223a <=( (not A299)  and  A298 );
 a30226a <=( A302  and  A300 );
 a30227a <=( a30226a  and  a30223a );
 a30228a <=( a30227a  and  a30220a );
 a30232a <=( (not A200)  and  A166 );
 a30233a <=( A168  and  a30232a );
 a30237a <=( (not A232)  and  (not A203) );
 a30238a <=( (not A202)  and  a30237a );
 a30239a <=( a30238a  and  a30233a );
 a30243a <=( (not A267)  and  (not A266) );
 a30244a <=( (not A233)  and  a30243a );
 a30247a <=( (not A299)  and  A298 );
 a30250a <=( A301  and  A300 );
 a30251a <=( a30250a  and  a30247a );
 a30252a <=( a30251a  and  a30244a );
 a30256a <=( (not A200)  and  A166 );
 a30257a <=( A168  and  a30256a );
 a30261a <=( (not A232)  and  (not A203) );
 a30262a <=( (not A202)  and  a30261a );
 a30263a <=( a30262a  and  a30257a );
 a30267a <=( (not A267)  and  (not A266) );
 a30268a <=( (not A233)  and  a30267a );
 a30271a <=( (not A299)  and  A298 );
 a30274a <=( A302  and  A300 );
 a30275a <=( a30274a  and  a30271a );
 a30276a <=( a30275a  and  a30268a );
 a30280a <=( (not A200)  and  A166 );
 a30281a <=( A168  and  a30280a );
 a30285a <=( (not A232)  and  (not A203) );
 a30286a <=( (not A202)  and  a30285a );
 a30287a <=( a30286a  and  a30281a );
 a30291a <=( (not A266)  and  (not A265) );
 a30292a <=( (not A233)  and  a30291a );
 a30295a <=( (not A299)  and  A298 );
 a30298a <=( A301  and  A300 );
 a30299a <=( a30298a  and  a30295a );
 a30300a <=( a30299a  and  a30292a );
 a30304a <=( (not A200)  and  A166 );
 a30305a <=( A168  and  a30304a );
 a30309a <=( (not A232)  and  (not A203) );
 a30310a <=( (not A202)  and  a30309a );
 a30311a <=( a30310a  and  a30305a );
 a30315a <=( (not A266)  and  (not A265) );
 a30316a <=( (not A233)  and  a30315a );
 a30319a <=( (not A299)  and  A298 );
 a30322a <=( A302  and  A300 );
 a30323a <=( a30322a  and  a30319a );
 a30324a <=( a30323a  and  a30316a );
 a30328a <=( (not A200)  and  A166 );
 a30329a <=( A168  and  a30328a );
 a30333a <=( A233  and  A232 );
 a30334a <=( (not A201)  and  a30333a );
 a30335a <=( a30334a  and  a30329a );
 a30339a <=( (not A269)  and  (not A268) );
 a30340a <=( A265  and  a30339a );
 a30343a <=( (not A299)  and  A298 );
 a30346a <=( A301  and  A300 );
 a30347a <=( a30346a  and  a30343a );
 a30348a <=( a30347a  and  a30340a );
 a30352a <=( (not A200)  and  A166 );
 a30353a <=( A168  and  a30352a );
 a30357a <=( A233  and  A232 );
 a30358a <=( (not A201)  and  a30357a );
 a30359a <=( a30358a  and  a30353a );
 a30363a <=( (not A269)  and  (not A268) );
 a30364a <=( A265  and  a30363a );
 a30367a <=( (not A299)  and  A298 );
 a30370a <=( A302  and  A300 );
 a30371a <=( a30370a  and  a30367a );
 a30372a <=( a30371a  and  a30364a );
 a30376a <=( (not A200)  and  A166 );
 a30377a <=( A168  and  a30376a );
 a30381a <=( (not A235)  and  (not A233) );
 a30382a <=( (not A201)  and  a30381a );
 a30383a <=( a30382a  and  a30377a );
 a30387a <=( A266  and  A265 );
 a30388a <=( (not A236)  and  a30387a );
 a30391a <=( (not A299)  and  A298 );
 a30394a <=( A301  and  A300 );
 a30395a <=( a30394a  and  a30391a );
 a30396a <=( a30395a  and  a30388a );
 a30400a <=( (not A200)  and  A166 );
 a30401a <=( A168  and  a30400a );
 a30405a <=( (not A235)  and  (not A233) );
 a30406a <=( (not A201)  and  a30405a );
 a30407a <=( a30406a  and  a30401a );
 a30411a <=( A266  and  A265 );
 a30412a <=( (not A236)  and  a30411a );
 a30415a <=( (not A299)  and  A298 );
 a30418a <=( A302  and  A300 );
 a30419a <=( a30418a  and  a30415a );
 a30420a <=( a30419a  and  a30412a );
 a30424a <=( (not A200)  and  A166 );
 a30425a <=( A168  and  a30424a );
 a30429a <=( (not A235)  and  (not A233) );
 a30430a <=( (not A201)  and  a30429a );
 a30431a <=( a30430a  and  a30425a );
 a30435a <=( (not A267)  and  (not A266) );
 a30436a <=( (not A236)  and  a30435a );
 a30439a <=( (not A299)  and  A298 );
 a30442a <=( A301  and  A300 );
 a30443a <=( a30442a  and  a30439a );
 a30444a <=( a30443a  and  a30436a );
 a30448a <=( (not A200)  and  A166 );
 a30449a <=( A168  and  a30448a );
 a30453a <=( (not A235)  and  (not A233) );
 a30454a <=( (not A201)  and  a30453a );
 a30455a <=( a30454a  and  a30449a );
 a30459a <=( (not A267)  and  (not A266) );
 a30460a <=( (not A236)  and  a30459a );
 a30463a <=( (not A299)  and  A298 );
 a30466a <=( A302  and  A300 );
 a30467a <=( a30466a  and  a30463a );
 a30468a <=( a30467a  and  a30460a );
 a30472a <=( (not A200)  and  A166 );
 a30473a <=( A168  and  a30472a );
 a30477a <=( (not A235)  and  (not A233) );
 a30478a <=( (not A201)  and  a30477a );
 a30479a <=( a30478a  and  a30473a );
 a30483a <=( (not A266)  and  (not A265) );
 a30484a <=( (not A236)  and  a30483a );
 a30487a <=( (not A299)  and  A298 );
 a30490a <=( A301  and  A300 );
 a30491a <=( a30490a  and  a30487a );
 a30492a <=( a30491a  and  a30484a );
 a30496a <=( (not A200)  and  A166 );
 a30497a <=( A168  and  a30496a );
 a30501a <=( (not A235)  and  (not A233) );
 a30502a <=( (not A201)  and  a30501a );
 a30503a <=( a30502a  and  a30497a );
 a30507a <=( (not A266)  and  (not A265) );
 a30508a <=( (not A236)  and  a30507a );
 a30511a <=( (not A299)  and  A298 );
 a30514a <=( A302  and  A300 );
 a30515a <=( a30514a  and  a30511a );
 a30516a <=( a30515a  and  a30508a );
 a30520a <=( (not A200)  and  A166 );
 a30521a <=( A168  and  a30520a );
 a30525a <=( (not A234)  and  (not A233) );
 a30526a <=( (not A201)  and  a30525a );
 a30527a <=( a30526a  and  a30521a );
 a30531a <=( (not A269)  and  (not A268) );
 a30532a <=( (not A266)  and  a30531a );
 a30535a <=( (not A299)  and  A298 );
 a30538a <=( A301  and  A300 );
 a30539a <=( a30538a  and  a30535a );
 a30540a <=( a30539a  and  a30532a );
 a30544a <=( (not A200)  and  A166 );
 a30545a <=( A168  and  a30544a );
 a30549a <=( (not A234)  and  (not A233) );
 a30550a <=( (not A201)  and  a30549a );
 a30551a <=( a30550a  and  a30545a );
 a30555a <=( (not A269)  and  (not A268) );
 a30556a <=( (not A266)  and  a30555a );
 a30559a <=( (not A299)  and  A298 );
 a30562a <=( A302  and  A300 );
 a30563a <=( a30562a  and  a30559a );
 a30564a <=( a30563a  and  a30556a );
 a30568a <=( (not A200)  and  A166 );
 a30569a <=( A168  and  a30568a );
 a30573a <=( (not A233)  and  (not A232) );
 a30574a <=( (not A201)  and  a30573a );
 a30575a <=( a30574a  and  a30569a );
 a30579a <=( (not A269)  and  (not A268) );
 a30580a <=( (not A266)  and  a30579a );
 a30583a <=( (not A299)  and  A298 );
 a30586a <=( A301  and  A300 );
 a30587a <=( a30586a  and  a30583a );
 a30588a <=( a30587a  and  a30580a );
 a30592a <=( (not A200)  and  A166 );
 a30593a <=( A168  and  a30592a );
 a30597a <=( (not A233)  and  (not A232) );
 a30598a <=( (not A201)  and  a30597a );
 a30599a <=( a30598a  and  a30593a );
 a30603a <=( (not A269)  and  (not A268) );
 a30604a <=( (not A266)  and  a30603a );
 a30607a <=( (not A299)  and  A298 );
 a30610a <=( A302  and  A300 );
 a30611a <=( a30610a  and  a30607a );
 a30612a <=( a30611a  and  a30604a );
 a30616a <=( (not A199)  and  A166 );
 a30617a <=( A168  and  a30616a );
 a30621a <=( A233  and  A232 );
 a30622a <=( (not A200)  and  a30621a );
 a30623a <=( a30622a  and  a30617a );
 a30627a <=( (not A269)  and  (not A268) );
 a30628a <=( A265  and  a30627a );
 a30631a <=( (not A299)  and  A298 );
 a30634a <=( A301  and  A300 );
 a30635a <=( a30634a  and  a30631a );
 a30636a <=( a30635a  and  a30628a );
 a30640a <=( (not A199)  and  A166 );
 a30641a <=( A168  and  a30640a );
 a30645a <=( A233  and  A232 );
 a30646a <=( (not A200)  and  a30645a );
 a30647a <=( a30646a  and  a30641a );
 a30651a <=( (not A269)  and  (not A268) );
 a30652a <=( A265  and  a30651a );
 a30655a <=( (not A299)  and  A298 );
 a30658a <=( A302  and  A300 );
 a30659a <=( a30658a  and  a30655a );
 a30660a <=( a30659a  and  a30652a );
 a30664a <=( (not A199)  and  A166 );
 a30665a <=( A168  and  a30664a );
 a30669a <=( (not A235)  and  (not A233) );
 a30670a <=( (not A200)  and  a30669a );
 a30671a <=( a30670a  and  a30665a );
 a30675a <=( A266  and  A265 );
 a30676a <=( (not A236)  and  a30675a );
 a30679a <=( (not A299)  and  A298 );
 a30682a <=( A301  and  A300 );
 a30683a <=( a30682a  and  a30679a );
 a30684a <=( a30683a  and  a30676a );
 a30688a <=( (not A199)  and  A166 );
 a30689a <=( A168  and  a30688a );
 a30693a <=( (not A235)  and  (not A233) );
 a30694a <=( (not A200)  and  a30693a );
 a30695a <=( a30694a  and  a30689a );
 a30699a <=( A266  and  A265 );
 a30700a <=( (not A236)  and  a30699a );
 a30703a <=( (not A299)  and  A298 );
 a30706a <=( A302  and  A300 );
 a30707a <=( a30706a  and  a30703a );
 a30708a <=( a30707a  and  a30700a );
 a30712a <=( (not A199)  and  A166 );
 a30713a <=( A168  and  a30712a );
 a30717a <=( (not A235)  and  (not A233) );
 a30718a <=( (not A200)  and  a30717a );
 a30719a <=( a30718a  and  a30713a );
 a30723a <=( (not A267)  and  (not A266) );
 a30724a <=( (not A236)  and  a30723a );
 a30727a <=( (not A299)  and  A298 );
 a30730a <=( A301  and  A300 );
 a30731a <=( a30730a  and  a30727a );
 a30732a <=( a30731a  and  a30724a );
 a30736a <=( (not A199)  and  A166 );
 a30737a <=( A168  and  a30736a );
 a30741a <=( (not A235)  and  (not A233) );
 a30742a <=( (not A200)  and  a30741a );
 a30743a <=( a30742a  and  a30737a );
 a30747a <=( (not A267)  and  (not A266) );
 a30748a <=( (not A236)  and  a30747a );
 a30751a <=( (not A299)  and  A298 );
 a30754a <=( A302  and  A300 );
 a30755a <=( a30754a  and  a30751a );
 a30756a <=( a30755a  and  a30748a );
 a30760a <=( (not A199)  and  A166 );
 a30761a <=( A168  and  a30760a );
 a30765a <=( (not A235)  and  (not A233) );
 a30766a <=( (not A200)  and  a30765a );
 a30767a <=( a30766a  and  a30761a );
 a30771a <=( (not A266)  and  (not A265) );
 a30772a <=( (not A236)  and  a30771a );
 a30775a <=( (not A299)  and  A298 );
 a30778a <=( A301  and  A300 );
 a30779a <=( a30778a  and  a30775a );
 a30780a <=( a30779a  and  a30772a );
 a30784a <=( (not A199)  and  A166 );
 a30785a <=( A168  and  a30784a );
 a30789a <=( (not A235)  and  (not A233) );
 a30790a <=( (not A200)  and  a30789a );
 a30791a <=( a30790a  and  a30785a );
 a30795a <=( (not A266)  and  (not A265) );
 a30796a <=( (not A236)  and  a30795a );
 a30799a <=( (not A299)  and  A298 );
 a30802a <=( A302  and  A300 );
 a30803a <=( a30802a  and  a30799a );
 a30804a <=( a30803a  and  a30796a );
 a30808a <=( (not A199)  and  A166 );
 a30809a <=( A168  and  a30808a );
 a30813a <=( (not A234)  and  (not A233) );
 a30814a <=( (not A200)  and  a30813a );
 a30815a <=( a30814a  and  a30809a );
 a30819a <=( (not A269)  and  (not A268) );
 a30820a <=( (not A266)  and  a30819a );
 a30823a <=( (not A299)  and  A298 );
 a30826a <=( A301  and  A300 );
 a30827a <=( a30826a  and  a30823a );
 a30828a <=( a30827a  and  a30820a );
 a30832a <=( (not A199)  and  A166 );
 a30833a <=( A168  and  a30832a );
 a30837a <=( (not A234)  and  (not A233) );
 a30838a <=( (not A200)  and  a30837a );
 a30839a <=( a30838a  and  a30833a );
 a30843a <=( (not A269)  and  (not A268) );
 a30844a <=( (not A266)  and  a30843a );
 a30847a <=( (not A299)  and  A298 );
 a30850a <=( A302  and  A300 );
 a30851a <=( a30850a  and  a30847a );
 a30852a <=( a30851a  and  a30844a );
 a30856a <=( (not A199)  and  A166 );
 a30857a <=( A168  and  a30856a );
 a30861a <=( (not A233)  and  (not A232) );
 a30862a <=( (not A200)  and  a30861a );
 a30863a <=( a30862a  and  a30857a );
 a30867a <=( (not A269)  and  (not A268) );
 a30868a <=( (not A266)  and  a30867a );
 a30871a <=( (not A299)  and  A298 );
 a30874a <=( A301  and  A300 );
 a30875a <=( a30874a  and  a30871a );
 a30876a <=( a30875a  and  a30868a );
 a30880a <=( (not A199)  and  A166 );
 a30881a <=( A168  and  a30880a );
 a30885a <=( (not A233)  and  (not A232) );
 a30886a <=( (not A200)  and  a30885a );
 a30887a <=( a30886a  and  a30881a );
 a30891a <=( (not A269)  and  (not A268) );
 a30892a <=( (not A266)  and  a30891a );
 a30895a <=( (not A299)  and  A298 );
 a30898a <=( A302  and  A300 );
 a30899a <=( a30898a  and  a30895a );
 a30900a <=( a30899a  and  a30892a );
 a30904a <=( A199  and  A167 );
 a30905a <=( A168  and  a30904a );
 a30909a <=( A233  and  A232 );
 a30910a <=( A200  and  a30909a );
 a30911a <=( a30910a  and  a30905a );
 a30915a <=( (not A269)  and  (not A268) );
 a30916a <=( A265  and  a30915a );
 a30919a <=( (not A299)  and  A298 );
 a30922a <=( A301  and  A300 );
 a30923a <=( a30922a  and  a30919a );
 a30924a <=( a30923a  and  a30916a );
 a30928a <=( A199  and  A167 );
 a30929a <=( A168  and  a30928a );
 a30933a <=( A233  and  A232 );
 a30934a <=( A200  and  a30933a );
 a30935a <=( a30934a  and  a30929a );
 a30939a <=( (not A269)  and  (not A268) );
 a30940a <=( A265  and  a30939a );
 a30943a <=( (not A299)  and  A298 );
 a30946a <=( A302  and  A300 );
 a30947a <=( a30946a  and  a30943a );
 a30948a <=( a30947a  and  a30940a );
 a30952a <=( A199  and  A167 );
 a30953a <=( A168  and  a30952a );
 a30957a <=( (not A235)  and  (not A233) );
 a30958a <=( A200  and  a30957a );
 a30959a <=( a30958a  and  a30953a );
 a30963a <=( A266  and  A265 );
 a30964a <=( (not A236)  and  a30963a );
 a30967a <=( (not A299)  and  A298 );
 a30970a <=( A301  and  A300 );
 a30971a <=( a30970a  and  a30967a );
 a30972a <=( a30971a  and  a30964a );
 a30976a <=( A199  and  A167 );
 a30977a <=( A168  and  a30976a );
 a30981a <=( (not A235)  and  (not A233) );
 a30982a <=( A200  and  a30981a );
 a30983a <=( a30982a  and  a30977a );
 a30987a <=( A266  and  A265 );
 a30988a <=( (not A236)  and  a30987a );
 a30991a <=( (not A299)  and  A298 );
 a30994a <=( A302  and  A300 );
 a30995a <=( a30994a  and  a30991a );
 a30996a <=( a30995a  and  a30988a );
 a31000a <=( A199  and  A167 );
 a31001a <=( A168  and  a31000a );
 a31005a <=( (not A235)  and  (not A233) );
 a31006a <=( A200  and  a31005a );
 a31007a <=( a31006a  and  a31001a );
 a31011a <=( (not A267)  and  (not A266) );
 a31012a <=( (not A236)  and  a31011a );
 a31015a <=( (not A299)  and  A298 );
 a31018a <=( A301  and  A300 );
 a31019a <=( a31018a  and  a31015a );
 a31020a <=( a31019a  and  a31012a );
 a31024a <=( A199  and  A167 );
 a31025a <=( A168  and  a31024a );
 a31029a <=( (not A235)  and  (not A233) );
 a31030a <=( A200  and  a31029a );
 a31031a <=( a31030a  and  a31025a );
 a31035a <=( (not A267)  and  (not A266) );
 a31036a <=( (not A236)  and  a31035a );
 a31039a <=( (not A299)  and  A298 );
 a31042a <=( A302  and  A300 );
 a31043a <=( a31042a  and  a31039a );
 a31044a <=( a31043a  and  a31036a );
 a31048a <=( A199  and  A167 );
 a31049a <=( A168  and  a31048a );
 a31053a <=( (not A235)  and  (not A233) );
 a31054a <=( A200  and  a31053a );
 a31055a <=( a31054a  and  a31049a );
 a31059a <=( (not A266)  and  (not A265) );
 a31060a <=( (not A236)  and  a31059a );
 a31063a <=( (not A299)  and  A298 );
 a31066a <=( A301  and  A300 );
 a31067a <=( a31066a  and  a31063a );
 a31068a <=( a31067a  and  a31060a );
 a31072a <=( A199  and  A167 );
 a31073a <=( A168  and  a31072a );
 a31077a <=( (not A235)  and  (not A233) );
 a31078a <=( A200  and  a31077a );
 a31079a <=( a31078a  and  a31073a );
 a31083a <=( (not A266)  and  (not A265) );
 a31084a <=( (not A236)  and  a31083a );
 a31087a <=( (not A299)  and  A298 );
 a31090a <=( A302  and  A300 );
 a31091a <=( a31090a  and  a31087a );
 a31092a <=( a31091a  and  a31084a );
 a31096a <=( A199  and  A167 );
 a31097a <=( A168  and  a31096a );
 a31101a <=( (not A234)  and  (not A233) );
 a31102a <=( A200  and  a31101a );
 a31103a <=( a31102a  and  a31097a );
 a31107a <=( (not A269)  and  (not A268) );
 a31108a <=( (not A266)  and  a31107a );
 a31111a <=( (not A299)  and  A298 );
 a31114a <=( A301  and  A300 );
 a31115a <=( a31114a  and  a31111a );
 a31116a <=( a31115a  and  a31108a );
 a31120a <=( A199  and  A167 );
 a31121a <=( A168  and  a31120a );
 a31125a <=( (not A234)  and  (not A233) );
 a31126a <=( A200  and  a31125a );
 a31127a <=( a31126a  and  a31121a );
 a31131a <=( (not A269)  and  (not A268) );
 a31132a <=( (not A266)  and  a31131a );
 a31135a <=( (not A299)  and  A298 );
 a31138a <=( A302  and  A300 );
 a31139a <=( a31138a  and  a31135a );
 a31140a <=( a31139a  and  a31132a );
 a31144a <=( A199  and  A167 );
 a31145a <=( A168  and  a31144a );
 a31149a <=( (not A233)  and  (not A232) );
 a31150a <=( A200  and  a31149a );
 a31151a <=( a31150a  and  a31145a );
 a31155a <=( (not A269)  and  (not A268) );
 a31156a <=( (not A266)  and  a31155a );
 a31159a <=( (not A299)  and  A298 );
 a31162a <=( A301  and  A300 );
 a31163a <=( a31162a  and  a31159a );
 a31164a <=( a31163a  and  a31156a );
 a31168a <=( A199  and  A167 );
 a31169a <=( A168  and  a31168a );
 a31173a <=( (not A233)  and  (not A232) );
 a31174a <=( A200  and  a31173a );
 a31175a <=( a31174a  and  a31169a );
 a31179a <=( (not A269)  and  (not A268) );
 a31180a <=( (not A266)  and  a31179a );
 a31183a <=( (not A299)  and  A298 );
 a31186a <=( A302  and  A300 );
 a31187a <=( a31186a  and  a31183a );
 a31188a <=( a31187a  and  a31180a );
 a31192a <=( (not A200)  and  A167 );
 a31193a <=( A168  and  a31192a );
 a31197a <=( A232  and  (not A203) );
 a31198a <=( (not A202)  and  a31197a );
 a31199a <=( a31198a  and  a31193a );
 a31203a <=( (not A267)  and  A265 );
 a31204a <=( A233  and  a31203a );
 a31207a <=( (not A299)  and  A298 );
 a31210a <=( A301  and  A300 );
 a31211a <=( a31210a  and  a31207a );
 a31212a <=( a31211a  and  a31204a );
 a31216a <=( (not A200)  and  A167 );
 a31217a <=( A168  and  a31216a );
 a31221a <=( A232  and  (not A203) );
 a31222a <=( (not A202)  and  a31221a );
 a31223a <=( a31222a  and  a31217a );
 a31227a <=( (not A267)  and  A265 );
 a31228a <=( A233  and  a31227a );
 a31231a <=( (not A299)  and  A298 );
 a31234a <=( A302  and  A300 );
 a31235a <=( a31234a  and  a31231a );
 a31236a <=( a31235a  and  a31228a );
 a31240a <=( (not A200)  and  A167 );
 a31241a <=( A168  and  a31240a );
 a31245a <=( A232  and  (not A203) );
 a31246a <=( (not A202)  and  a31245a );
 a31247a <=( a31246a  and  a31241a );
 a31251a <=( A266  and  A265 );
 a31252a <=( A233  and  a31251a );
 a31255a <=( (not A299)  and  A298 );
 a31258a <=( A301  and  A300 );
 a31259a <=( a31258a  and  a31255a );
 a31260a <=( a31259a  and  a31252a );
 a31264a <=( (not A200)  and  A167 );
 a31265a <=( A168  and  a31264a );
 a31269a <=( A232  and  (not A203) );
 a31270a <=( (not A202)  and  a31269a );
 a31271a <=( a31270a  and  a31265a );
 a31275a <=( A266  and  A265 );
 a31276a <=( A233  and  a31275a );
 a31279a <=( (not A299)  and  A298 );
 a31282a <=( A302  and  A300 );
 a31283a <=( a31282a  and  a31279a );
 a31284a <=( a31283a  and  a31276a );
 a31288a <=( (not A200)  and  A167 );
 a31289a <=( A168  and  a31288a );
 a31293a <=( A232  and  (not A203) );
 a31294a <=( (not A202)  and  a31293a );
 a31295a <=( a31294a  and  a31289a );
 a31299a <=( (not A266)  and  (not A265) );
 a31300a <=( A233  and  a31299a );
 a31303a <=( (not A299)  and  A298 );
 a31306a <=( A301  and  A300 );
 a31307a <=( a31306a  and  a31303a );
 a31308a <=( a31307a  and  a31300a );
 a31312a <=( (not A200)  and  A167 );
 a31313a <=( A168  and  a31312a );
 a31317a <=( A232  and  (not A203) );
 a31318a <=( (not A202)  and  a31317a );
 a31319a <=( a31318a  and  a31313a );
 a31323a <=( (not A266)  and  (not A265) );
 a31324a <=( A233  and  a31323a );
 a31327a <=( (not A299)  and  A298 );
 a31330a <=( A302  and  A300 );
 a31331a <=( a31330a  and  a31327a );
 a31332a <=( a31331a  and  a31324a );
 a31336a <=( (not A200)  and  A167 );
 a31337a <=( A168  and  a31336a );
 a31341a <=( (not A233)  and  (not A203) );
 a31342a <=( (not A202)  and  a31341a );
 a31343a <=( a31342a  and  a31337a );
 a31347a <=( (not A266)  and  (not A236) );
 a31348a <=( (not A235)  and  a31347a );
 a31351a <=( (not A269)  and  (not A268) );
 a31354a <=( A299  and  (not A298) );
 a31355a <=( a31354a  and  a31351a );
 a31356a <=( a31355a  and  a31348a );
 a31360a <=( (not A200)  and  A167 );
 a31361a <=( A168  and  a31360a );
 a31365a <=( (not A233)  and  (not A203) );
 a31366a <=( (not A202)  and  a31365a );
 a31367a <=( a31366a  and  a31361a );
 a31371a <=( A266  and  A265 );
 a31372a <=( (not A234)  and  a31371a );
 a31375a <=( (not A299)  and  A298 );
 a31378a <=( A301  and  A300 );
 a31379a <=( a31378a  and  a31375a );
 a31380a <=( a31379a  and  a31372a );
 a31384a <=( (not A200)  and  A167 );
 a31385a <=( A168  and  a31384a );
 a31389a <=( (not A233)  and  (not A203) );
 a31390a <=( (not A202)  and  a31389a );
 a31391a <=( a31390a  and  a31385a );
 a31395a <=( A266  and  A265 );
 a31396a <=( (not A234)  and  a31395a );
 a31399a <=( (not A299)  and  A298 );
 a31402a <=( A302  and  A300 );
 a31403a <=( a31402a  and  a31399a );
 a31404a <=( a31403a  and  a31396a );
 a31408a <=( (not A200)  and  A167 );
 a31409a <=( A168  and  a31408a );
 a31413a <=( (not A233)  and  (not A203) );
 a31414a <=( (not A202)  and  a31413a );
 a31415a <=( a31414a  and  a31409a );
 a31419a <=( (not A267)  and  (not A266) );
 a31420a <=( (not A234)  and  a31419a );
 a31423a <=( (not A299)  and  A298 );
 a31426a <=( A301  and  A300 );
 a31427a <=( a31426a  and  a31423a );
 a31428a <=( a31427a  and  a31420a );
 a31432a <=( (not A200)  and  A167 );
 a31433a <=( A168  and  a31432a );
 a31437a <=( (not A233)  and  (not A203) );
 a31438a <=( (not A202)  and  a31437a );
 a31439a <=( a31438a  and  a31433a );
 a31443a <=( (not A267)  and  (not A266) );
 a31444a <=( (not A234)  and  a31443a );
 a31447a <=( (not A299)  and  A298 );
 a31450a <=( A302  and  A300 );
 a31451a <=( a31450a  and  a31447a );
 a31452a <=( a31451a  and  a31444a );
 a31456a <=( (not A200)  and  A167 );
 a31457a <=( A168  and  a31456a );
 a31461a <=( (not A233)  and  (not A203) );
 a31462a <=( (not A202)  and  a31461a );
 a31463a <=( a31462a  and  a31457a );
 a31467a <=( (not A266)  and  (not A265) );
 a31468a <=( (not A234)  and  a31467a );
 a31471a <=( (not A299)  and  A298 );
 a31474a <=( A301  and  A300 );
 a31475a <=( a31474a  and  a31471a );
 a31476a <=( a31475a  and  a31468a );
 a31480a <=( (not A200)  and  A167 );
 a31481a <=( A168  and  a31480a );
 a31485a <=( (not A233)  and  (not A203) );
 a31486a <=( (not A202)  and  a31485a );
 a31487a <=( a31486a  and  a31481a );
 a31491a <=( (not A266)  and  (not A265) );
 a31492a <=( (not A234)  and  a31491a );
 a31495a <=( (not A299)  and  A298 );
 a31498a <=( A302  and  A300 );
 a31499a <=( a31498a  and  a31495a );
 a31500a <=( a31499a  and  a31492a );
 a31504a <=( (not A200)  and  A167 );
 a31505a <=( A168  and  a31504a );
 a31509a <=( A232  and  (not A203) );
 a31510a <=( (not A202)  and  a31509a );
 a31511a <=( a31510a  and  a31505a );
 a31515a <=( A235  and  A234 );
 a31516a <=( (not A233)  and  a31515a );
 a31519a <=( (not A266)  and  A265 );
 a31522a <=( A268  and  A267 );
 a31523a <=( a31522a  and  a31519a );
 a31524a <=( a31523a  and  a31516a );
 a31528a <=( (not A200)  and  A167 );
 a31529a <=( A168  and  a31528a );
 a31533a <=( A232  and  (not A203) );
 a31534a <=( (not A202)  and  a31533a );
 a31535a <=( a31534a  and  a31529a );
 a31539a <=( A235  and  A234 );
 a31540a <=( (not A233)  and  a31539a );
 a31543a <=( (not A266)  and  A265 );
 a31546a <=( A269  and  A267 );
 a31547a <=( a31546a  and  a31543a );
 a31548a <=( a31547a  and  a31540a );
 a31552a <=( (not A200)  and  A167 );
 a31553a <=( A168  and  a31552a );
 a31557a <=( A232  and  (not A203) );
 a31558a <=( (not A202)  and  a31557a );
 a31559a <=( a31558a  and  a31553a );
 a31563a <=( A236  and  A234 );
 a31564a <=( (not A233)  and  a31563a );
 a31567a <=( (not A266)  and  A265 );
 a31570a <=( A268  and  A267 );
 a31571a <=( a31570a  and  a31567a );
 a31572a <=( a31571a  and  a31564a );
 a31576a <=( (not A200)  and  A167 );
 a31577a <=( A168  and  a31576a );
 a31581a <=( A232  and  (not A203) );
 a31582a <=( (not A202)  and  a31581a );
 a31583a <=( a31582a  and  a31577a );
 a31587a <=( A236  and  A234 );
 a31588a <=( (not A233)  and  a31587a );
 a31591a <=( (not A266)  and  A265 );
 a31594a <=( A269  and  A267 );
 a31595a <=( a31594a  and  a31591a );
 a31596a <=( a31595a  and  a31588a );
 a31600a <=( (not A200)  and  A167 );
 a31601a <=( A168  and  a31600a );
 a31605a <=( (not A232)  and  (not A203) );
 a31606a <=( (not A202)  and  a31605a );
 a31607a <=( a31606a  and  a31601a );
 a31611a <=( A266  and  A265 );
 a31612a <=( (not A233)  and  a31611a );
 a31615a <=( (not A299)  and  A298 );
 a31618a <=( A301  and  A300 );
 a31619a <=( a31618a  and  a31615a );
 a31620a <=( a31619a  and  a31612a );
 a31624a <=( (not A200)  and  A167 );
 a31625a <=( A168  and  a31624a );
 a31629a <=( (not A232)  and  (not A203) );
 a31630a <=( (not A202)  and  a31629a );
 a31631a <=( a31630a  and  a31625a );
 a31635a <=( A266  and  A265 );
 a31636a <=( (not A233)  and  a31635a );
 a31639a <=( (not A299)  and  A298 );
 a31642a <=( A302  and  A300 );
 a31643a <=( a31642a  and  a31639a );
 a31644a <=( a31643a  and  a31636a );
 a31648a <=( (not A200)  and  A167 );
 a31649a <=( A168  and  a31648a );
 a31653a <=( (not A232)  and  (not A203) );
 a31654a <=( (not A202)  and  a31653a );
 a31655a <=( a31654a  and  a31649a );
 a31659a <=( (not A267)  and  (not A266) );
 a31660a <=( (not A233)  and  a31659a );
 a31663a <=( (not A299)  and  A298 );
 a31666a <=( A301  and  A300 );
 a31667a <=( a31666a  and  a31663a );
 a31668a <=( a31667a  and  a31660a );
 a31672a <=( (not A200)  and  A167 );
 a31673a <=( A168  and  a31672a );
 a31677a <=( (not A232)  and  (not A203) );
 a31678a <=( (not A202)  and  a31677a );
 a31679a <=( a31678a  and  a31673a );
 a31683a <=( (not A267)  and  (not A266) );
 a31684a <=( (not A233)  and  a31683a );
 a31687a <=( (not A299)  and  A298 );
 a31690a <=( A302  and  A300 );
 a31691a <=( a31690a  and  a31687a );
 a31692a <=( a31691a  and  a31684a );
 a31696a <=( (not A200)  and  A167 );
 a31697a <=( A168  and  a31696a );
 a31701a <=( (not A232)  and  (not A203) );
 a31702a <=( (not A202)  and  a31701a );
 a31703a <=( a31702a  and  a31697a );
 a31707a <=( (not A266)  and  (not A265) );
 a31708a <=( (not A233)  and  a31707a );
 a31711a <=( (not A299)  and  A298 );
 a31714a <=( A301  and  A300 );
 a31715a <=( a31714a  and  a31711a );
 a31716a <=( a31715a  and  a31708a );
 a31720a <=( (not A200)  and  A167 );
 a31721a <=( A168  and  a31720a );
 a31725a <=( (not A232)  and  (not A203) );
 a31726a <=( (not A202)  and  a31725a );
 a31727a <=( a31726a  and  a31721a );
 a31731a <=( (not A266)  and  (not A265) );
 a31732a <=( (not A233)  and  a31731a );
 a31735a <=( (not A299)  and  A298 );
 a31738a <=( A302  and  A300 );
 a31739a <=( a31738a  and  a31735a );
 a31740a <=( a31739a  and  a31732a );
 a31744a <=( (not A200)  and  A167 );
 a31745a <=( A168  and  a31744a );
 a31749a <=( A233  and  A232 );
 a31750a <=( (not A201)  and  a31749a );
 a31751a <=( a31750a  and  a31745a );
 a31755a <=( (not A269)  and  (not A268) );
 a31756a <=( A265  and  a31755a );
 a31759a <=( (not A299)  and  A298 );
 a31762a <=( A301  and  A300 );
 a31763a <=( a31762a  and  a31759a );
 a31764a <=( a31763a  and  a31756a );
 a31768a <=( (not A200)  and  A167 );
 a31769a <=( A168  and  a31768a );
 a31773a <=( A233  and  A232 );
 a31774a <=( (not A201)  and  a31773a );
 a31775a <=( a31774a  and  a31769a );
 a31779a <=( (not A269)  and  (not A268) );
 a31780a <=( A265  and  a31779a );
 a31783a <=( (not A299)  and  A298 );
 a31786a <=( A302  and  A300 );
 a31787a <=( a31786a  and  a31783a );
 a31788a <=( a31787a  and  a31780a );
 a31792a <=( (not A200)  and  A167 );
 a31793a <=( A168  and  a31792a );
 a31797a <=( (not A235)  and  (not A233) );
 a31798a <=( (not A201)  and  a31797a );
 a31799a <=( a31798a  and  a31793a );
 a31803a <=( A266  and  A265 );
 a31804a <=( (not A236)  and  a31803a );
 a31807a <=( (not A299)  and  A298 );
 a31810a <=( A301  and  A300 );
 a31811a <=( a31810a  and  a31807a );
 a31812a <=( a31811a  and  a31804a );
 a31816a <=( (not A200)  and  A167 );
 a31817a <=( A168  and  a31816a );
 a31821a <=( (not A235)  and  (not A233) );
 a31822a <=( (not A201)  and  a31821a );
 a31823a <=( a31822a  and  a31817a );
 a31827a <=( A266  and  A265 );
 a31828a <=( (not A236)  and  a31827a );
 a31831a <=( (not A299)  and  A298 );
 a31834a <=( A302  and  A300 );
 a31835a <=( a31834a  and  a31831a );
 a31836a <=( a31835a  and  a31828a );
 a31840a <=( (not A200)  and  A167 );
 a31841a <=( A168  and  a31840a );
 a31845a <=( (not A235)  and  (not A233) );
 a31846a <=( (not A201)  and  a31845a );
 a31847a <=( a31846a  and  a31841a );
 a31851a <=( (not A267)  and  (not A266) );
 a31852a <=( (not A236)  and  a31851a );
 a31855a <=( (not A299)  and  A298 );
 a31858a <=( A301  and  A300 );
 a31859a <=( a31858a  and  a31855a );
 a31860a <=( a31859a  and  a31852a );
 a31864a <=( (not A200)  and  A167 );
 a31865a <=( A168  and  a31864a );
 a31869a <=( (not A235)  and  (not A233) );
 a31870a <=( (not A201)  and  a31869a );
 a31871a <=( a31870a  and  a31865a );
 a31875a <=( (not A267)  and  (not A266) );
 a31876a <=( (not A236)  and  a31875a );
 a31879a <=( (not A299)  and  A298 );
 a31882a <=( A302  and  A300 );
 a31883a <=( a31882a  and  a31879a );
 a31884a <=( a31883a  and  a31876a );
 a31888a <=( (not A200)  and  A167 );
 a31889a <=( A168  and  a31888a );
 a31893a <=( (not A235)  and  (not A233) );
 a31894a <=( (not A201)  and  a31893a );
 a31895a <=( a31894a  and  a31889a );
 a31899a <=( (not A266)  and  (not A265) );
 a31900a <=( (not A236)  and  a31899a );
 a31903a <=( (not A299)  and  A298 );
 a31906a <=( A301  and  A300 );
 a31907a <=( a31906a  and  a31903a );
 a31908a <=( a31907a  and  a31900a );
 a31912a <=( (not A200)  and  A167 );
 a31913a <=( A168  and  a31912a );
 a31917a <=( (not A235)  and  (not A233) );
 a31918a <=( (not A201)  and  a31917a );
 a31919a <=( a31918a  and  a31913a );
 a31923a <=( (not A266)  and  (not A265) );
 a31924a <=( (not A236)  and  a31923a );
 a31927a <=( (not A299)  and  A298 );
 a31930a <=( A302  and  A300 );
 a31931a <=( a31930a  and  a31927a );
 a31932a <=( a31931a  and  a31924a );
 a31936a <=( (not A200)  and  A167 );
 a31937a <=( A168  and  a31936a );
 a31941a <=( (not A234)  and  (not A233) );
 a31942a <=( (not A201)  and  a31941a );
 a31943a <=( a31942a  and  a31937a );
 a31947a <=( (not A269)  and  (not A268) );
 a31948a <=( (not A266)  and  a31947a );
 a31951a <=( (not A299)  and  A298 );
 a31954a <=( A301  and  A300 );
 a31955a <=( a31954a  and  a31951a );
 a31956a <=( a31955a  and  a31948a );
 a31960a <=( (not A200)  and  A167 );
 a31961a <=( A168  and  a31960a );
 a31965a <=( (not A234)  and  (not A233) );
 a31966a <=( (not A201)  and  a31965a );
 a31967a <=( a31966a  and  a31961a );
 a31971a <=( (not A269)  and  (not A268) );
 a31972a <=( (not A266)  and  a31971a );
 a31975a <=( (not A299)  and  A298 );
 a31978a <=( A302  and  A300 );
 a31979a <=( a31978a  and  a31975a );
 a31980a <=( a31979a  and  a31972a );
 a31984a <=( (not A200)  and  A167 );
 a31985a <=( A168  and  a31984a );
 a31989a <=( (not A233)  and  (not A232) );
 a31990a <=( (not A201)  and  a31989a );
 a31991a <=( a31990a  and  a31985a );
 a31995a <=( (not A269)  and  (not A268) );
 a31996a <=( (not A266)  and  a31995a );
 a31999a <=( (not A299)  and  A298 );
 a32002a <=( A301  and  A300 );
 a32003a <=( a32002a  and  a31999a );
 a32004a <=( a32003a  and  a31996a );
 a32008a <=( (not A200)  and  A167 );
 a32009a <=( A168  and  a32008a );
 a32013a <=( (not A233)  and  (not A232) );
 a32014a <=( (not A201)  and  a32013a );
 a32015a <=( a32014a  and  a32009a );
 a32019a <=( (not A269)  and  (not A268) );
 a32020a <=( (not A266)  and  a32019a );
 a32023a <=( (not A299)  and  A298 );
 a32026a <=( A302  and  A300 );
 a32027a <=( a32026a  and  a32023a );
 a32028a <=( a32027a  and  a32020a );
 a32032a <=( (not A199)  and  A167 );
 a32033a <=( A168  and  a32032a );
 a32037a <=( A233  and  A232 );
 a32038a <=( (not A200)  and  a32037a );
 a32039a <=( a32038a  and  a32033a );
 a32043a <=( (not A269)  and  (not A268) );
 a32044a <=( A265  and  a32043a );
 a32047a <=( (not A299)  and  A298 );
 a32050a <=( A301  and  A300 );
 a32051a <=( a32050a  and  a32047a );
 a32052a <=( a32051a  and  a32044a );
 a32056a <=( (not A199)  and  A167 );
 a32057a <=( A168  and  a32056a );
 a32061a <=( A233  and  A232 );
 a32062a <=( (not A200)  and  a32061a );
 a32063a <=( a32062a  and  a32057a );
 a32067a <=( (not A269)  and  (not A268) );
 a32068a <=( A265  and  a32067a );
 a32071a <=( (not A299)  and  A298 );
 a32074a <=( A302  and  A300 );
 a32075a <=( a32074a  and  a32071a );
 a32076a <=( a32075a  and  a32068a );
 a32080a <=( (not A199)  and  A167 );
 a32081a <=( A168  and  a32080a );
 a32085a <=( (not A235)  and  (not A233) );
 a32086a <=( (not A200)  and  a32085a );
 a32087a <=( a32086a  and  a32081a );
 a32091a <=( A266  and  A265 );
 a32092a <=( (not A236)  and  a32091a );
 a32095a <=( (not A299)  and  A298 );
 a32098a <=( A301  and  A300 );
 a32099a <=( a32098a  and  a32095a );
 a32100a <=( a32099a  and  a32092a );
 a32104a <=( (not A199)  and  A167 );
 a32105a <=( A168  and  a32104a );
 a32109a <=( (not A235)  and  (not A233) );
 a32110a <=( (not A200)  and  a32109a );
 a32111a <=( a32110a  and  a32105a );
 a32115a <=( A266  and  A265 );
 a32116a <=( (not A236)  and  a32115a );
 a32119a <=( (not A299)  and  A298 );
 a32122a <=( A302  and  A300 );
 a32123a <=( a32122a  and  a32119a );
 a32124a <=( a32123a  and  a32116a );
 a32128a <=( (not A199)  and  A167 );
 a32129a <=( A168  and  a32128a );
 a32133a <=( (not A235)  and  (not A233) );
 a32134a <=( (not A200)  and  a32133a );
 a32135a <=( a32134a  and  a32129a );
 a32139a <=( (not A267)  and  (not A266) );
 a32140a <=( (not A236)  and  a32139a );
 a32143a <=( (not A299)  and  A298 );
 a32146a <=( A301  and  A300 );
 a32147a <=( a32146a  and  a32143a );
 a32148a <=( a32147a  and  a32140a );
 a32152a <=( (not A199)  and  A167 );
 a32153a <=( A168  and  a32152a );
 a32157a <=( (not A235)  and  (not A233) );
 a32158a <=( (not A200)  and  a32157a );
 a32159a <=( a32158a  and  a32153a );
 a32163a <=( (not A267)  and  (not A266) );
 a32164a <=( (not A236)  and  a32163a );
 a32167a <=( (not A299)  and  A298 );
 a32170a <=( A302  and  A300 );
 a32171a <=( a32170a  and  a32167a );
 a32172a <=( a32171a  and  a32164a );
 a32176a <=( (not A199)  and  A167 );
 a32177a <=( A168  and  a32176a );
 a32181a <=( (not A235)  and  (not A233) );
 a32182a <=( (not A200)  and  a32181a );
 a32183a <=( a32182a  and  a32177a );
 a32187a <=( (not A266)  and  (not A265) );
 a32188a <=( (not A236)  and  a32187a );
 a32191a <=( (not A299)  and  A298 );
 a32194a <=( A301  and  A300 );
 a32195a <=( a32194a  and  a32191a );
 a32196a <=( a32195a  and  a32188a );
 a32200a <=( (not A199)  and  A167 );
 a32201a <=( A168  and  a32200a );
 a32205a <=( (not A235)  and  (not A233) );
 a32206a <=( (not A200)  and  a32205a );
 a32207a <=( a32206a  and  a32201a );
 a32211a <=( (not A266)  and  (not A265) );
 a32212a <=( (not A236)  and  a32211a );
 a32215a <=( (not A299)  and  A298 );
 a32218a <=( A302  and  A300 );
 a32219a <=( a32218a  and  a32215a );
 a32220a <=( a32219a  and  a32212a );
 a32224a <=( (not A199)  and  A167 );
 a32225a <=( A168  and  a32224a );
 a32229a <=( (not A234)  and  (not A233) );
 a32230a <=( (not A200)  and  a32229a );
 a32231a <=( a32230a  and  a32225a );
 a32235a <=( (not A269)  and  (not A268) );
 a32236a <=( (not A266)  and  a32235a );
 a32239a <=( (not A299)  and  A298 );
 a32242a <=( A301  and  A300 );
 a32243a <=( a32242a  and  a32239a );
 a32244a <=( a32243a  and  a32236a );
 a32248a <=( (not A199)  and  A167 );
 a32249a <=( A168  and  a32248a );
 a32253a <=( (not A234)  and  (not A233) );
 a32254a <=( (not A200)  and  a32253a );
 a32255a <=( a32254a  and  a32249a );
 a32259a <=( (not A269)  and  (not A268) );
 a32260a <=( (not A266)  and  a32259a );
 a32263a <=( (not A299)  and  A298 );
 a32266a <=( A302  and  A300 );
 a32267a <=( a32266a  and  a32263a );
 a32268a <=( a32267a  and  a32260a );
 a32272a <=( (not A199)  and  A167 );
 a32273a <=( A168  and  a32272a );
 a32277a <=( (not A233)  and  (not A232) );
 a32278a <=( (not A200)  and  a32277a );
 a32279a <=( a32278a  and  a32273a );
 a32283a <=( (not A269)  and  (not A268) );
 a32284a <=( (not A266)  and  a32283a );
 a32287a <=( (not A299)  and  A298 );
 a32290a <=( A301  and  A300 );
 a32291a <=( a32290a  and  a32287a );
 a32292a <=( a32291a  and  a32284a );
 a32296a <=( (not A199)  and  A167 );
 a32297a <=( A168  and  a32296a );
 a32301a <=( (not A233)  and  (not A232) );
 a32302a <=( (not A200)  and  a32301a );
 a32303a <=( a32302a  and  a32297a );
 a32307a <=( (not A269)  and  (not A268) );
 a32308a <=( (not A266)  and  a32307a );
 a32311a <=( (not A299)  and  A298 );
 a32314a <=( A302  and  A300 );
 a32315a <=( a32314a  and  a32311a );
 a32316a <=( a32315a  and  a32308a );
 a32320a <=( (not A166)  and  (not A167) );
 a32321a <=( A170  and  a32320a );
 a32325a <=( A232  and  A200 );
 a32326a <=( (not A199)  and  a32325a );
 a32327a <=( a32326a  and  a32321a );
 a32331a <=( (not A267)  and  A265 );
 a32332a <=( A233  and  a32331a );
 a32335a <=( (not A299)  and  A298 );
 a32338a <=( A301  and  A300 );
 a32339a <=( a32338a  and  a32335a );
 a32340a <=( a32339a  and  a32332a );
 a32344a <=( (not A166)  and  (not A167) );
 a32345a <=( A170  and  a32344a );
 a32349a <=( A232  and  A200 );
 a32350a <=( (not A199)  and  a32349a );
 a32351a <=( a32350a  and  a32345a );
 a32355a <=( (not A267)  and  A265 );
 a32356a <=( A233  and  a32355a );
 a32359a <=( (not A299)  and  A298 );
 a32362a <=( A302  and  A300 );
 a32363a <=( a32362a  and  a32359a );
 a32364a <=( a32363a  and  a32356a );
 a32368a <=( (not A166)  and  (not A167) );
 a32369a <=( A170  and  a32368a );
 a32373a <=( A232  and  A200 );
 a32374a <=( (not A199)  and  a32373a );
 a32375a <=( a32374a  and  a32369a );
 a32379a <=( A266  and  A265 );
 a32380a <=( A233  and  a32379a );
 a32383a <=( (not A299)  and  A298 );
 a32386a <=( A301  and  A300 );
 a32387a <=( a32386a  and  a32383a );
 a32388a <=( a32387a  and  a32380a );
 a32392a <=( (not A166)  and  (not A167) );
 a32393a <=( A170  and  a32392a );
 a32397a <=( A232  and  A200 );
 a32398a <=( (not A199)  and  a32397a );
 a32399a <=( a32398a  and  a32393a );
 a32403a <=( A266  and  A265 );
 a32404a <=( A233  and  a32403a );
 a32407a <=( (not A299)  and  A298 );
 a32410a <=( A302  and  A300 );
 a32411a <=( a32410a  and  a32407a );
 a32412a <=( a32411a  and  a32404a );
 a32416a <=( (not A166)  and  (not A167) );
 a32417a <=( A170  and  a32416a );
 a32421a <=( A232  and  A200 );
 a32422a <=( (not A199)  and  a32421a );
 a32423a <=( a32422a  and  a32417a );
 a32427a <=( (not A266)  and  (not A265) );
 a32428a <=( A233  and  a32427a );
 a32431a <=( (not A299)  and  A298 );
 a32434a <=( A301  and  A300 );
 a32435a <=( a32434a  and  a32431a );
 a32436a <=( a32435a  and  a32428a );
 a32440a <=( (not A166)  and  (not A167) );
 a32441a <=( A170  and  a32440a );
 a32445a <=( A232  and  A200 );
 a32446a <=( (not A199)  and  a32445a );
 a32447a <=( a32446a  and  a32441a );
 a32451a <=( (not A266)  and  (not A265) );
 a32452a <=( A233  and  a32451a );
 a32455a <=( (not A299)  and  A298 );
 a32458a <=( A302  and  A300 );
 a32459a <=( a32458a  and  a32455a );
 a32460a <=( a32459a  and  a32452a );
 a32464a <=( (not A166)  and  (not A167) );
 a32465a <=( A170  and  a32464a );
 a32469a <=( (not A233)  and  A200 );
 a32470a <=( (not A199)  and  a32469a );
 a32471a <=( a32470a  and  a32465a );
 a32475a <=( (not A266)  and  (not A236) );
 a32476a <=( (not A235)  and  a32475a );
 a32479a <=( (not A269)  and  (not A268) );
 a32482a <=( A299  and  (not A298) );
 a32483a <=( a32482a  and  a32479a );
 a32484a <=( a32483a  and  a32476a );
 a32488a <=( (not A166)  and  (not A167) );
 a32489a <=( A170  and  a32488a );
 a32493a <=( (not A233)  and  A200 );
 a32494a <=( (not A199)  and  a32493a );
 a32495a <=( a32494a  and  a32489a );
 a32499a <=( A266  and  A265 );
 a32500a <=( (not A234)  and  a32499a );
 a32503a <=( (not A299)  and  A298 );
 a32506a <=( A301  and  A300 );
 a32507a <=( a32506a  and  a32503a );
 a32508a <=( a32507a  and  a32500a );
 a32512a <=( (not A166)  and  (not A167) );
 a32513a <=( A170  and  a32512a );
 a32517a <=( (not A233)  and  A200 );
 a32518a <=( (not A199)  and  a32517a );
 a32519a <=( a32518a  and  a32513a );
 a32523a <=( A266  and  A265 );
 a32524a <=( (not A234)  and  a32523a );
 a32527a <=( (not A299)  and  A298 );
 a32530a <=( A302  and  A300 );
 a32531a <=( a32530a  and  a32527a );
 a32532a <=( a32531a  and  a32524a );
 a32536a <=( (not A166)  and  (not A167) );
 a32537a <=( A170  and  a32536a );
 a32541a <=( (not A233)  and  A200 );
 a32542a <=( (not A199)  and  a32541a );
 a32543a <=( a32542a  and  a32537a );
 a32547a <=( (not A267)  and  (not A266) );
 a32548a <=( (not A234)  and  a32547a );
 a32551a <=( (not A299)  and  A298 );
 a32554a <=( A301  and  A300 );
 a32555a <=( a32554a  and  a32551a );
 a32556a <=( a32555a  and  a32548a );
 a32560a <=( (not A166)  and  (not A167) );
 a32561a <=( A170  and  a32560a );
 a32565a <=( (not A233)  and  A200 );
 a32566a <=( (not A199)  and  a32565a );
 a32567a <=( a32566a  and  a32561a );
 a32571a <=( (not A267)  and  (not A266) );
 a32572a <=( (not A234)  and  a32571a );
 a32575a <=( (not A299)  and  A298 );
 a32578a <=( A302  and  A300 );
 a32579a <=( a32578a  and  a32575a );
 a32580a <=( a32579a  and  a32572a );
 a32584a <=( (not A166)  and  (not A167) );
 a32585a <=( A170  and  a32584a );
 a32589a <=( (not A233)  and  A200 );
 a32590a <=( (not A199)  and  a32589a );
 a32591a <=( a32590a  and  a32585a );
 a32595a <=( (not A266)  and  (not A265) );
 a32596a <=( (not A234)  and  a32595a );
 a32599a <=( (not A299)  and  A298 );
 a32602a <=( A301  and  A300 );
 a32603a <=( a32602a  and  a32599a );
 a32604a <=( a32603a  and  a32596a );
 a32608a <=( (not A166)  and  (not A167) );
 a32609a <=( A170  and  a32608a );
 a32613a <=( (not A233)  and  A200 );
 a32614a <=( (not A199)  and  a32613a );
 a32615a <=( a32614a  and  a32609a );
 a32619a <=( (not A266)  and  (not A265) );
 a32620a <=( (not A234)  and  a32619a );
 a32623a <=( (not A299)  and  A298 );
 a32626a <=( A302  and  A300 );
 a32627a <=( a32626a  and  a32623a );
 a32628a <=( a32627a  and  a32620a );
 a32632a <=( (not A166)  and  (not A167) );
 a32633a <=( A170  and  a32632a );
 a32637a <=( A232  and  A200 );
 a32638a <=( (not A199)  and  a32637a );
 a32639a <=( a32638a  and  a32633a );
 a32643a <=( A235  and  A234 );
 a32644a <=( (not A233)  and  a32643a );
 a32647a <=( (not A266)  and  A265 );
 a32650a <=( A268  and  A267 );
 a32651a <=( a32650a  and  a32647a );
 a32652a <=( a32651a  and  a32644a );
 a32656a <=( (not A166)  and  (not A167) );
 a32657a <=( A170  and  a32656a );
 a32661a <=( A232  and  A200 );
 a32662a <=( (not A199)  and  a32661a );
 a32663a <=( a32662a  and  a32657a );
 a32667a <=( A235  and  A234 );
 a32668a <=( (not A233)  and  a32667a );
 a32671a <=( (not A266)  and  A265 );
 a32674a <=( A269  and  A267 );
 a32675a <=( a32674a  and  a32671a );
 a32676a <=( a32675a  and  a32668a );
 a32680a <=( (not A166)  and  (not A167) );
 a32681a <=( A170  and  a32680a );
 a32685a <=( A232  and  A200 );
 a32686a <=( (not A199)  and  a32685a );
 a32687a <=( a32686a  and  a32681a );
 a32691a <=( A236  and  A234 );
 a32692a <=( (not A233)  and  a32691a );
 a32695a <=( (not A266)  and  A265 );
 a32698a <=( A268  and  A267 );
 a32699a <=( a32698a  and  a32695a );
 a32700a <=( a32699a  and  a32692a );
 a32704a <=( (not A166)  and  (not A167) );
 a32705a <=( A170  and  a32704a );
 a32709a <=( A232  and  A200 );
 a32710a <=( (not A199)  and  a32709a );
 a32711a <=( a32710a  and  a32705a );
 a32715a <=( A236  and  A234 );
 a32716a <=( (not A233)  and  a32715a );
 a32719a <=( (not A266)  and  A265 );
 a32722a <=( A269  and  A267 );
 a32723a <=( a32722a  and  a32719a );
 a32724a <=( a32723a  and  a32716a );
 a32728a <=( (not A166)  and  (not A167) );
 a32729a <=( A170  and  a32728a );
 a32733a <=( (not A232)  and  A200 );
 a32734a <=( (not A199)  and  a32733a );
 a32735a <=( a32734a  and  a32729a );
 a32739a <=( A266  and  A265 );
 a32740a <=( (not A233)  and  a32739a );
 a32743a <=( (not A299)  and  A298 );
 a32746a <=( A301  and  A300 );
 a32747a <=( a32746a  and  a32743a );
 a32748a <=( a32747a  and  a32740a );
 a32752a <=( (not A166)  and  (not A167) );
 a32753a <=( A170  and  a32752a );
 a32757a <=( (not A232)  and  A200 );
 a32758a <=( (not A199)  and  a32757a );
 a32759a <=( a32758a  and  a32753a );
 a32763a <=( A266  and  A265 );
 a32764a <=( (not A233)  and  a32763a );
 a32767a <=( (not A299)  and  A298 );
 a32770a <=( A302  and  A300 );
 a32771a <=( a32770a  and  a32767a );
 a32772a <=( a32771a  and  a32764a );
 a32776a <=( (not A166)  and  (not A167) );
 a32777a <=( A170  and  a32776a );
 a32781a <=( (not A232)  and  A200 );
 a32782a <=( (not A199)  and  a32781a );
 a32783a <=( a32782a  and  a32777a );
 a32787a <=( (not A267)  and  (not A266) );
 a32788a <=( (not A233)  and  a32787a );
 a32791a <=( (not A299)  and  A298 );
 a32794a <=( A301  and  A300 );
 a32795a <=( a32794a  and  a32791a );
 a32796a <=( a32795a  and  a32788a );
 a32800a <=( (not A166)  and  (not A167) );
 a32801a <=( A170  and  a32800a );
 a32805a <=( (not A232)  and  A200 );
 a32806a <=( (not A199)  and  a32805a );
 a32807a <=( a32806a  and  a32801a );
 a32811a <=( (not A267)  and  (not A266) );
 a32812a <=( (not A233)  and  a32811a );
 a32815a <=( (not A299)  and  A298 );
 a32818a <=( A302  and  A300 );
 a32819a <=( a32818a  and  a32815a );
 a32820a <=( a32819a  and  a32812a );
 a32824a <=( (not A166)  and  (not A167) );
 a32825a <=( A170  and  a32824a );
 a32829a <=( (not A232)  and  A200 );
 a32830a <=( (not A199)  and  a32829a );
 a32831a <=( a32830a  and  a32825a );
 a32835a <=( (not A266)  and  (not A265) );
 a32836a <=( (not A233)  and  a32835a );
 a32839a <=( (not A299)  and  A298 );
 a32842a <=( A301  and  A300 );
 a32843a <=( a32842a  and  a32839a );
 a32844a <=( a32843a  and  a32836a );
 a32848a <=( (not A166)  and  (not A167) );
 a32849a <=( A170  and  a32848a );
 a32853a <=( (not A232)  and  A200 );
 a32854a <=( (not A199)  and  a32853a );
 a32855a <=( a32854a  and  a32849a );
 a32859a <=( (not A266)  and  (not A265) );
 a32860a <=( (not A233)  and  a32859a );
 a32863a <=( (not A299)  and  A298 );
 a32866a <=( A302  and  A300 );
 a32867a <=( a32866a  and  a32863a );
 a32868a <=( a32867a  and  a32860a );
 a32872a <=( (not A166)  and  (not A167) );
 a32873a <=( A170  and  a32872a );
 a32877a <=( A201  and  (not A200) );
 a32878a <=( A199  and  a32877a );
 a32879a <=( a32878a  and  a32873a );
 a32883a <=( A233  and  A232 );
 a32884a <=( A202  and  a32883a );
 a32887a <=( (not A267)  and  A265 );
 a32890a <=( A299  and  (not A298) );
 a32891a <=( a32890a  and  a32887a );
 a32892a <=( a32891a  and  a32884a );
 a32896a <=( (not A166)  and  (not A167) );
 a32897a <=( A170  and  a32896a );
 a32901a <=( A201  and  (not A200) );
 a32902a <=( A199  and  a32901a );
 a32903a <=( a32902a  and  a32897a );
 a32907a <=( A233  and  A232 );
 a32908a <=( A202  and  a32907a );
 a32911a <=( A266  and  A265 );
 a32914a <=( A299  and  (not A298) );
 a32915a <=( a32914a  and  a32911a );
 a32916a <=( a32915a  and  a32908a );
 a32920a <=( (not A166)  and  (not A167) );
 a32921a <=( A170  and  a32920a );
 a32925a <=( A201  and  (not A200) );
 a32926a <=( A199  and  a32925a );
 a32927a <=( a32926a  and  a32921a );
 a32931a <=( A233  and  A232 );
 a32932a <=( A202  and  a32931a );
 a32935a <=( (not A266)  and  (not A265) );
 a32938a <=( A299  and  (not A298) );
 a32939a <=( a32938a  and  a32935a );
 a32940a <=( a32939a  and  a32932a );
 a32944a <=( (not A166)  and  (not A167) );
 a32945a <=( A170  and  a32944a );
 a32949a <=( A201  and  (not A200) );
 a32950a <=( A199  and  a32949a );
 a32951a <=( a32950a  and  a32945a );
 a32955a <=( A233  and  (not A232) );
 a32956a <=( A202  and  a32955a );
 a32959a <=( (not A266)  and  A265 );
 a32962a <=( A268  and  A267 );
 a32963a <=( a32962a  and  a32959a );
 a32964a <=( a32963a  and  a32956a );
 a32968a <=( (not A166)  and  (not A167) );
 a32969a <=( A170  and  a32968a );
 a32973a <=( A201  and  (not A200) );
 a32974a <=( A199  and  a32973a );
 a32975a <=( a32974a  and  a32969a );
 a32979a <=( A233  and  (not A232) );
 a32980a <=( A202  and  a32979a );
 a32983a <=( (not A266)  and  A265 );
 a32986a <=( A269  and  A267 );
 a32987a <=( a32986a  and  a32983a );
 a32988a <=( a32987a  and  a32980a );
 a32992a <=( (not A166)  and  (not A167) );
 a32993a <=( A170  and  a32992a );
 a32997a <=( A201  and  (not A200) );
 a32998a <=( A199  and  a32997a );
 a32999a <=( a32998a  and  a32993a );
 a33003a <=( (not A234)  and  (not A233) );
 a33004a <=( A202  and  a33003a );
 a33007a <=( A266  and  A265 );
 a33010a <=( A299  and  (not A298) );
 a33011a <=( a33010a  and  a33007a );
 a33012a <=( a33011a  and  a33004a );
 a33016a <=( (not A166)  and  (not A167) );
 a33017a <=( A170  and  a33016a );
 a33021a <=( A201  and  (not A200) );
 a33022a <=( A199  and  a33021a );
 a33023a <=( a33022a  and  a33017a );
 a33027a <=( (not A234)  and  (not A233) );
 a33028a <=( A202  and  a33027a );
 a33031a <=( (not A267)  and  (not A266) );
 a33034a <=( A299  and  (not A298) );
 a33035a <=( a33034a  and  a33031a );
 a33036a <=( a33035a  and  a33028a );
 a33040a <=( (not A166)  and  (not A167) );
 a33041a <=( A170  and  a33040a );
 a33045a <=( A201  and  (not A200) );
 a33046a <=( A199  and  a33045a );
 a33047a <=( a33046a  and  a33041a );
 a33051a <=( (not A234)  and  (not A233) );
 a33052a <=( A202  and  a33051a );
 a33055a <=( (not A266)  and  (not A265) );
 a33058a <=( A299  and  (not A298) );
 a33059a <=( a33058a  and  a33055a );
 a33060a <=( a33059a  and  a33052a );
 a33064a <=( (not A166)  and  (not A167) );
 a33065a <=( A170  and  a33064a );
 a33069a <=( A201  and  (not A200) );
 a33070a <=( A199  and  a33069a );
 a33071a <=( a33070a  and  a33065a );
 a33075a <=( (not A233)  and  A232 );
 a33076a <=( A202  and  a33075a );
 a33079a <=( A235  and  A234 );
 a33082a <=( (not A300)  and  A298 );
 a33083a <=( a33082a  and  a33079a );
 a33084a <=( a33083a  and  a33076a );
 a33088a <=( (not A166)  and  (not A167) );
 a33089a <=( A170  and  a33088a );
 a33093a <=( A201  and  (not A200) );
 a33094a <=( A199  and  a33093a );
 a33095a <=( a33094a  and  a33089a );
 a33099a <=( (not A233)  and  A232 );
 a33100a <=( A202  and  a33099a );
 a33103a <=( A235  and  A234 );
 a33106a <=( A299  and  A298 );
 a33107a <=( a33106a  and  a33103a );
 a33108a <=( a33107a  and  a33100a );
 a33112a <=( (not A166)  and  (not A167) );
 a33113a <=( A170  and  a33112a );
 a33117a <=( A201  and  (not A200) );
 a33118a <=( A199  and  a33117a );
 a33119a <=( a33118a  and  a33113a );
 a33123a <=( (not A233)  and  A232 );
 a33124a <=( A202  and  a33123a );
 a33127a <=( A235  and  A234 );
 a33130a <=( (not A299)  and  (not A298) );
 a33131a <=( a33130a  and  a33127a );
 a33132a <=( a33131a  and  a33124a );
 a33136a <=( (not A166)  and  (not A167) );
 a33137a <=( A170  and  a33136a );
 a33141a <=( A201  and  (not A200) );
 a33142a <=( A199  and  a33141a );
 a33143a <=( a33142a  and  a33137a );
 a33147a <=( (not A233)  and  A232 );
 a33148a <=( A202  and  a33147a );
 a33151a <=( A235  and  A234 );
 a33154a <=( A266  and  (not A265) );
 a33155a <=( a33154a  and  a33151a );
 a33156a <=( a33155a  and  a33148a );
 a33160a <=( (not A166)  and  (not A167) );
 a33161a <=( A170  and  a33160a );
 a33165a <=( A201  and  (not A200) );
 a33166a <=( A199  and  a33165a );
 a33167a <=( a33166a  and  a33161a );
 a33171a <=( (not A233)  and  A232 );
 a33172a <=( A202  and  a33171a );
 a33175a <=( A236  and  A234 );
 a33178a <=( (not A300)  and  A298 );
 a33179a <=( a33178a  and  a33175a );
 a33180a <=( a33179a  and  a33172a );
 a33184a <=( (not A166)  and  (not A167) );
 a33185a <=( A170  and  a33184a );
 a33189a <=( A201  and  (not A200) );
 a33190a <=( A199  and  a33189a );
 a33191a <=( a33190a  and  a33185a );
 a33195a <=( (not A233)  and  A232 );
 a33196a <=( A202  and  a33195a );
 a33199a <=( A236  and  A234 );
 a33202a <=( A299  and  A298 );
 a33203a <=( a33202a  and  a33199a );
 a33204a <=( a33203a  and  a33196a );
 a33208a <=( (not A166)  and  (not A167) );
 a33209a <=( A170  and  a33208a );
 a33213a <=( A201  and  (not A200) );
 a33214a <=( A199  and  a33213a );
 a33215a <=( a33214a  and  a33209a );
 a33219a <=( (not A233)  and  A232 );
 a33220a <=( A202  and  a33219a );
 a33223a <=( A236  and  A234 );
 a33226a <=( (not A299)  and  (not A298) );
 a33227a <=( a33226a  and  a33223a );
 a33228a <=( a33227a  and  a33220a );
 a33232a <=( (not A166)  and  (not A167) );
 a33233a <=( A170  and  a33232a );
 a33237a <=( A201  and  (not A200) );
 a33238a <=( A199  and  a33237a );
 a33239a <=( a33238a  and  a33233a );
 a33243a <=( (not A233)  and  A232 );
 a33244a <=( A202  and  a33243a );
 a33247a <=( A236  and  A234 );
 a33250a <=( A266  and  (not A265) );
 a33251a <=( a33250a  and  a33247a );
 a33252a <=( a33251a  and  a33244a );
 a33256a <=( (not A166)  and  (not A167) );
 a33257a <=( A170  and  a33256a );
 a33261a <=( A201  and  (not A200) );
 a33262a <=( A199  and  a33261a );
 a33263a <=( a33262a  and  a33257a );
 a33267a <=( (not A233)  and  (not A232) );
 a33268a <=( A202  and  a33267a );
 a33271a <=( A266  and  A265 );
 a33274a <=( A299  and  (not A298) );
 a33275a <=( a33274a  and  a33271a );
 a33276a <=( a33275a  and  a33268a );
 a33280a <=( (not A166)  and  (not A167) );
 a33281a <=( A170  and  a33280a );
 a33285a <=( A201  and  (not A200) );
 a33286a <=( A199  and  a33285a );
 a33287a <=( a33286a  and  a33281a );
 a33291a <=( (not A233)  and  (not A232) );
 a33292a <=( A202  and  a33291a );
 a33295a <=( (not A267)  and  (not A266) );
 a33298a <=( A299  and  (not A298) );
 a33299a <=( a33298a  and  a33295a );
 a33300a <=( a33299a  and  a33292a );
 a33304a <=( (not A166)  and  (not A167) );
 a33305a <=( A170  and  a33304a );
 a33309a <=( A201  and  (not A200) );
 a33310a <=( A199  and  a33309a );
 a33311a <=( a33310a  and  a33305a );
 a33315a <=( (not A233)  and  (not A232) );
 a33316a <=( A202  and  a33315a );
 a33319a <=( (not A266)  and  (not A265) );
 a33322a <=( A299  and  (not A298) );
 a33323a <=( a33322a  and  a33319a );
 a33324a <=( a33323a  and  a33316a );
 a33328a <=( (not A166)  and  (not A167) );
 a33329a <=( A170  and  a33328a );
 a33333a <=( A201  and  (not A200) );
 a33334a <=( A199  and  a33333a );
 a33335a <=( a33334a  and  a33329a );
 a33339a <=( A233  and  A232 );
 a33340a <=( A203  and  a33339a );
 a33343a <=( (not A267)  and  A265 );
 a33346a <=( A299  and  (not A298) );
 a33347a <=( a33346a  and  a33343a );
 a33348a <=( a33347a  and  a33340a );
 a33352a <=( (not A166)  and  (not A167) );
 a33353a <=( A170  and  a33352a );
 a33357a <=( A201  and  (not A200) );
 a33358a <=( A199  and  a33357a );
 a33359a <=( a33358a  and  a33353a );
 a33363a <=( A233  and  A232 );
 a33364a <=( A203  and  a33363a );
 a33367a <=( A266  and  A265 );
 a33370a <=( A299  and  (not A298) );
 a33371a <=( a33370a  and  a33367a );
 a33372a <=( a33371a  and  a33364a );
 a33376a <=( (not A166)  and  (not A167) );
 a33377a <=( A170  and  a33376a );
 a33381a <=( A201  and  (not A200) );
 a33382a <=( A199  and  a33381a );
 a33383a <=( a33382a  and  a33377a );
 a33387a <=( A233  and  A232 );
 a33388a <=( A203  and  a33387a );
 a33391a <=( (not A266)  and  (not A265) );
 a33394a <=( A299  and  (not A298) );
 a33395a <=( a33394a  and  a33391a );
 a33396a <=( a33395a  and  a33388a );
 a33400a <=( (not A166)  and  (not A167) );
 a33401a <=( A170  and  a33400a );
 a33405a <=( A201  and  (not A200) );
 a33406a <=( A199  and  a33405a );
 a33407a <=( a33406a  and  a33401a );
 a33411a <=( A233  and  (not A232) );
 a33412a <=( A203  and  a33411a );
 a33415a <=( (not A266)  and  A265 );
 a33418a <=( A268  and  A267 );
 a33419a <=( a33418a  and  a33415a );
 a33420a <=( a33419a  and  a33412a );
 a33424a <=( (not A166)  and  (not A167) );
 a33425a <=( A170  and  a33424a );
 a33429a <=( A201  and  (not A200) );
 a33430a <=( A199  and  a33429a );
 a33431a <=( a33430a  and  a33425a );
 a33435a <=( A233  and  (not A232) );
 a33436a <=( A203  and  a33435a );
 a33439a <=( (not A266)  and  A265 );
 a33442a <=( A269  and  A267 );
 a33443a <=( a33442a  and  a33439a );
 a33444a <=( a33443a  and  a33436a );
 a33448a <=( (not A166)  and  (not A167) );
 a33449a <=( A170  and  a33448a );
 a33453a <=( A201  and  (not A200) );
 a33454a <=( A199  and  a33453a );
 a33455a <=( a33454a  and  a33449a );
 a33459a <=( (not A234)  and  (not A233) );
 a33460a <=( A203  and  a33459a );
 a33463a <=( A266  and  A265 );
 a33466a <=( A299  and  (not A298) );
 a33467a <=( a33466a  and  a33463a );
 a33468a <=( a33467a  and  a33460a );
 a33472a <=( (not A166)  and  (not A167) );
 a33473a <=( A170  and  a33472a );
 a33477a <=( A201  and  (not A200) );
 a33478a <=( A199  and  a33477a );
 a33479a <=( a33478a  and  a33473a );
 a33483a <=( (not A234)  and  (not A233) );
 a33484a <=( A203  and  a33483a );
 a33487a <=( (not A267)  and  (not A266) );
 a33490a <=( A299  and  (not A298) );
 a33491a <=( a33490a  and  a33487a );
 a33492a <=( a33491a  and  a33484a );
 a33496a <=( (not A166)  and  (not A167) );
 a33497a <=( A170  and  a33496a );
 a33501a <=( A201  and  (not A200) );
 a33502a <=( A199  and  a33501a );
 a33503a <=( a33502a  and  a33497a );
 a33507a <=( (not A234)  and  (not A233) );
 a33508a <=( A203  and  a33507a );
 a33511a <=( (not A266)  and  (not A265) );
 a33514a <=( A299  and  (not A298) );
 a33515a <=( a33514a  and  a33511a );
 a33516a <=( a33515a  and  a33508a );
 a33520a <=( (not A166)  and  (not A167) );
 a33521a <=( A170  and  a33520a );
 a33525a <=( A201  and  (not A200) );
 a33526a <=( A199  and  a33525a );
 a33527a <=( a33526a  and  a33521a );
 a33531a <=( (not A233)  and  A232 );
 a33532a <=( A203  and  a33531a );
 a33535a <=( A235  and  A234 );
 a33538a <=( (not A300)  and  A298 );
 a33539a <=( a33538a  and  a33535a );
 a33540a <=( a33539a  and  a33532a );
 a33544a <=( (not A166)  and  (not A167) );
 a33545a <=( A170  and  a33544a );
 a33549a <=( A201  and  (not A200) );
 a33550a <=( A199  and  a33549a );
 a33551a <=( a33550a  and  a33545a );
 a33555a <=( (not A233)  and  A232 );
 a33556a <=( A203  and  a33555a );
 a33559a <=( A235  and  A234 );
 a33562a <=( A299  and  A298 );
 a33563a <=( a33562a  and  a33559a );
 a33564a <=( a33563a  and  a33556a );
 a33568a <=( (not A166)  and  (not A167) );
 a33569a <=( A170  and  a33568a );
 a33573a <=( A201  and  (not A200) );
 a33574a <=( A199  and  a33573a );
 a33575a <=( a33574a  and  a33569a );
 a33579a <=( (not A233)  and  A232 );
 a33580a <=( A203  and  a33579a );
 a33583a <=( A235  and  A234 );
 a33586a <=( (not A299)  and  (not A298) );
 a33587a <=( a33586a  and  a33583a );
 a33588a <=( a33587a  and  a33580a );
 a33592a <=( (not A166)  and  (not A167) );
 a33593a <=( A170  and  a33592a );
 a33597a <=( A201  and  (not A200) );
 a33598a <=( A199  and  a33597a );
 a33599a <=( a33598a  and  a33593a );
 a33603a <=( (not A233)  and  A232 );
 a33604a <=( A203  and  a33603a );
 a33607a <=( A235  and  A234 );
 a33610a <=( A266  and  (not A265) );
 a33611a <=( a33610a  and  a33607a );
 a33612a <=( a33611a  and  a33604a );
 a33616a <=( (not A166)  and  (not A167) );
 a33617a <=( A170  and  a33616a );
 a33621a <=( A201  and  (not A200) );
 a33622a <=( A199  and  a33621a );
 a33623a <=( a33622a  and  a33617a );
 a33627a <=( (not A233)  and  A232 );
 a33628a <=( A203  and  a33627a );
 a33631a <=( A236  and  A234 );
 a33634a <=( (not A300)  and  A298 );
 a33635a <=( a33634a  and  a33631a );
 a33636a <=( a33635a  and  a33628a );
 a33640a <=( (not A166)  and  (not A167) );
 a33641a <=( A170  and  a33640a );
 a33645a <=( A201  and  (not A200) );
 a33646a <=( A199  and  a33645a );
 a33647a <=( a33646a  and  a33641a );
 a33651a <=( (not A233)  and  A232 );
 a33652a <=( A203  and  a33651a );
 a33655a <=( A236  and  A234 );
 a33658a <=( A299  and  A298 );
 a33659a <=( a33658a  and  a33655a );
 a33660a <=( a33659a  and  a33652a );
 a33664a <=( (not A166)  and  (not A167) );
 a33665a <=( A170  and  a33664a );
 a33669a <=( A201  and  (not A200) );
 a33670a <=( A199  and  a33669a );
 a33671a <=( a33670a  and  a33665a );
 a33675a <=( (not A233)  and  A232 );
 a33676a <=( A203  and  a33675a );
 a33679a <=( A236  and  A234 );
 a33682a <=( (not A299)  and  (not A298) );
 a33683a <=( a33682a  and  a33679a );
 a33684a <=( a33683a  and  a33676a );
 a33688a <=( (not A166)  and  (not A167) );
 a33689a <=( A170  and  a33688a );
 a33693a <=( A201  and  (not A200) );
 a33694a <=( A199  and  a33693a );
 a33695a <=( a33694a  and  a33689a );
 a33699a <=( (not A233)  and  A232 );
 a33700a <=( A203  and  a33699a );
 a33703a <=( A236  and  A234 );
 a33706a <=( A266  and  (not A265) );
 a33707a <=( a33706a  and  a33703a );
 a33708a <=( a33707a  and  a33700a );
 a33712a <=( (not A166)  and  (not A167) );
 a33713a <=( A170  and  a33712a );
 a33717a <=( A201  and  (not A200) );
 a33718a <=( A199  and  a33717a );
 a33719a <=( a33718a  and  a33713a );
 a33723a <=( (not A233)  and  (not A232) );
 a33724a <=( A203  and  a33723a );
 a33727a <=( A266  and  A265 );
 a33730a <=( A299  and  (not A298) );
 a33731a <=( a33730a  and  a33727a );
 a33732a <=( a33731a  and  a33724a );
 a33736a <=( (not A166)  and  (not A167) );
 a33737a <=( A170  and  a33736a );
 a33741a <=( A201  and  (not A200) );
 a33742a <=( A199  and  a33741a );
 a33743a <=( a33742a  and  a33737a );
 a33747a <=( (not A233)  and  (not A232) );
 a33748a <=( A203  and  a33747a );
 a33751a <=( (not A267)  and  (not A266) );
 a33754a <=( A299  and  (not A298) );
 a33755a <=( a33754a  and  a33751a );
 a33756a <=( a33755a  and  a33748a );
 a33760a <=( (not A166)  and  (not A167) );
 a33761a <=( A170  and  a33760a );
 a33765a <=( A201  and  (not A200) );
 a33766a <=( A199  and  a33765a );
 a33767a <=( a33766a  and  a33761a );
 a33771a <=( (not A233)  and  (not A232) );
 a33772a <=( A203  and  a33771a );
 a33775a <=( (not A266)  and  (not A265) );
 a33778a <=( A299  and  (not A298) );
 a33779a <=( a33778a  and  a33775a );
 a33780a <=( a33779a  and  a33772a );
 a33784a <=( A167  and  (not A168) );
 a33785a <=( A170  and  a33784a );
 a33789a <=( A200  and  (not A199) );
 a33790a <=( A166  and  a33789a );
 a33791a <=( a33790a  and  a33785a );
 a33795a <=( A265  and  A233 );
 a33796a <=( A232  and  a33795a );
 a33799a <=( (not A269)  and  (not A268) );
 a33802a <=( A299  and  (not A298) );
 a33803a <=( a33802a  and  a33799a );
 a33804a <=( a33803a  and  a33796a );
 a33808a <=( A167  and  (not A168) );
 a33809a <=( A170  and  a33808a );
 a33813a <=( A200  and  (not A199) );
 a33814a <=( A166  and  a33813a );
 a33815a <=( a33814a  and  a33809a );
 a33819a <=( (not A236)  and  (not A235) );
 a33820a <=( (not A233)  and  a33819a );
 a33823a <=( A266  and  A265 );
 a33826a <=( A299  and  (not A298) );
 a33827a <=( a33826a  and  a33823a );
 a33828a <=( a33827a  and  a33820a );
 a33832a <=( A167  and  (not A168) );
 a33833a <=( A170  and  a33832a );
 a33837a <=( A200  and  (not A199) );
 a33838a <=( A166  and  a33837a );
 a33839a <=( a33838a  and  a33833a );
 a33843a <=( (not A236)  and  (not A235) );
 a33844a <=( (not A233)  and  a33843a );
 a33847a <=( (not A267)  and  (not A266) );
 a33850a <=( A299  and  (not A298) );
 a33851a <=( a33850a  and  a33847a );
 a33852a <=( a33851a  and  a33844a );
 a33856a <=( A167  and  (not A168) );
 a33857a <=( A170  and  a33856a );
 a33861a <=( A200  and  (not A199) );
 a33862a <=( A166  and  a33861a );
 a33863a <=( a33862a  and  a33857a );
 a33867a <=( (not A236)  and  (not A235) );
 a33868a <=( (not A233)  and  a33867a );
 a33871a <=( (not A266)  and  (not A265) );
 a33874a <=( A299  and  (not A298) );
 a33875a <=( a33874a  and  a33871a );
 a33876a <=( a33875a  and  a33868a );
 a33880a <=( A167  and  (not A168) );
 a33881a <=( A170  and  a33880a );
 a33885a <=( A200  and  (not A199) );
 a33886a <=( A166  and  a33885a );
 a33887a <=( a33886a  and  a33881a );
 a33891a <=( (not A266)  and  (not A234) );
 a33892a <=( (not A233)  and  a33891a );
 a33895a <=( (not A269)  and  (not A268) );
 a33898a <=( A299  and  (not A298) );
 a33899a <=( a33898a  and  a33895a );
 a33900a <=( a33899a  and  a33892a );
 a33904a <=( A167  and  (not A168) );
 a33905a <=( A170  and  a33904a );
 a33909a <=( A200  and  (not A199) );
 a33910a <=( A166  and  a33909a );
 a33911a <=( a33910a  and  a33905a );
 a33915a <=( A234  and  (not A233) );
 a33916a <=( A232  and  a33915a );
 a33919a <=( A298  and  A235 );
 a33922a <=( (not A302)  and  (not A301) );
 a33923a <=( a33922a  and  a33919a );
 a33924a <=( a33923a  and  a33916a );
 a33928a <=( A167  and  (not A168) );
 a33929a <=( A170  and  a33928a );
 a33933a <=( A200  and  (not A199) );
 a33934a <=( A166  and  a33933a );
 a33935a <=( a33934a  and  a33929a );
 a33939a <=( A234  and  (not A233) );
 a33940a <=( A232  and  a33939a );
 a33943a <=( A298  and  A236 );
 a33946a <=( (not A302)  and  (not A301) );
 a33947a <=( a33946a  and  a33943a );
 a33948a <=( a33947a  and  a33940a );
 a33952a <=( A167  and  (not A168) );
 a33953a <=( A170  and  a33952a );
 a33957a <=( A200  and  (not A199) );
 a33958a <=( A166  and  a33957a );
 a33959a <=( a33958a  and  a33953a );
 a33963a <=( (not A266)  and  (not A233) );
 a33964a <=( (not A232)  and  a33963a );
 a33967a <=( (not A269)  and  (not A268) );
 a33970a <=( A299  and  (not A298) );
 a33971a <=( a33970a  and  a33967a );
 a33972a <=( a33971a  and  a33964a );
 a33976a <=( A167  and  (not A168) );
 a33977a <=( (not A170)  and  a33976a );
 a33981a <=( A200  and  (not A199) );
 a33982a <=( (not A166)  and  a33981a );
 a33983a <=( a33982a  and  a33977a );
 a33987a <=( A265  and  A233 );
 a33988a <=( A232  and  a33987a );
 a33991a <=( (not A269)  and  (not A268) );
 a33994a <=( A299  and  (not A298) );
 a33995a <=( a33994a  and  a33991a );
 a33996a <=( a33995a  and  a33988a );
 a34000a <=( A167  and  (not A168) );
 a34001a <=( (not A170)  and  a34000a );
 a34005a <=( A200  and  (not A199) );
 a34006a <=( (not A166)  and  a34005a );
 a34007a <=( a34006a  and  a34001a );
 a34011a <=( (not A236)  and  (not A235) );
 a34012a <=( (not A233)  and  a34011a );
 a34015a <=( A266  and  A265 );
 a34018a <=( A299  and  (not A298) );
 a34019a <=( a34018a  and  a34015a );
 a34020a <=( a34019a  and  a34012a );
 a34024a <=( A167  and  (not A168) );
 a34025a <=( (not A170)  and  a34024a );
 a34029a <=( A200  and  (not A199) );
 a34030a <=( (not A166)  and  a34029a );
 a34031a <=( a34030a  and  a34025a );
 a34035a <=( (not A236)  and  (not A235) );
 a34036a <=( (not A233)  and  a34035a );
 a34039a <=( (not A267)  and  (not A266) );
 a34042a <=( A299  and  (not A298) );
 a34043a <=( a34042a  and  a34039a );
 a34044a <=( a34043a  and  a34036a );
 a34048a <=( A167  and  (not A168) );
 a34049a <=( (not A170)  and  a34048a );
 a34053a <=( A200  and  (not A199) );
 a34054a <=( (not A166)  and  a34053a );
 a34055a <=( a34054a  and  a34049a );
 a34059a <=( (not A236)  and  (not A235) );
 a34060a <=( (not A233)  and  a34059a );
 a34063a <=( (not A266)  and  (not A265) );
 a34066a <=( A299  and  (not A298) );
 a34067a <=( a34066a  and  a34063a );
 a34068a <=( a34067a  and  a34060a );
 a34072a <=( A167  and  (not A168) );
 a34073a <=( (not A170)  and  a34072a );
 a34077a <=( A200  and  (not A199) );
 a34078a <=( (not A166)  and  a34077a );
 a34079a <=( a34078a  and  a34073a );
 a34083a <=( (not A266)  and  (not A234) );
 a34084a <=( (not A233)  and  a34083a );
 a34087a <=( (not A269)  and  (not A268) );
 a34090a <=( A299  and  (not A298) );
 a34091a <=( a34090a  and  a34087a );
 a34092a <=( a34091a  and  a34084a );
 a34096a <=( A167  and  (not A168) );
 a34097a <=( (not A170)  and  a34096a );
 a34101a <=( A200  and  (not A199) );
 a34102a <=( (not A166)  and  a34101a );
 a34103a <=( a34102a  and  a34097a );
 a34107a <=( A234  and  (not A233) );
 a34108a <=( A232  and  a34107a );
 a34111a <=( A298  and  A235 );
 a34114a <=( (not A302)  and  (not A301) );
 a34115a <=( a34114a  and  a34111a );
 a34116a <=( a34115a  and  a34108a );
 a34120a <=( A167  and  (not A168) );
 a34121a <=( (not A170)  and  a34120a );
 a34125a <=( A200  and  (not A199) );
 a34126a <=( (not A166)  and  a34125a );
 a34127a <=( a34126a  and  a34121a );
 a34131a <=( A234  and  (not A233) );
 a34132a <=( A232  and  a34131a );
 a34135a <=( A298  and  A236 );
 a34138a <=( (not A302)  and  (not A301) );
 a34139a <=( a34138a  and  a34135a );
 a34140a <=( a34139a  and  a34132a );
 a34144a <=( A167  and  (not A168) );
 a34145a <=( (not A170)  and  a34144a );
 a34149a <=( A200  and  (not A199) );
 a34150a <=( (not A166)  and  a34149a );
 a34151a <=( a34150a  and  a34145a );
 a34155a <=( (not A266)  and  (not A233) );
 a34156a <=( (not A232)  and  a34155a );
 a34159a <=( (not A269)  and  (not A268) );
 a34162a <=( A299  and  (not A298) );
 a34163a <=( a34162a  and  a34159a );
 a34164a <=( a34163a  and  a34156a );
 a34168a <=( (not A167)  and  (not A168) );
 a34169a <=( (not A170)  and  a34168a );
 a34173a <=( A200  and  (not A199) );
 a34174a <=( A166  and  a34173a );
 a34175a <=( a34174a  and  a34169a );
 a34179a <=( A265  and  A233 );
 a34180a <=( A232  and  a34179a );
 a34183a <=( (not A269)  and  (not A268) );
 a34186a <=( A299  and  (not A298) );
 a34187a <=( a34186a  and  a34183a );
 a34188a <=( a34187a  and  a34180a );
 a34192a <=( (not A167)  and  (not A168) );
 a34193a <=( (not A170)  and  a34192a );
 a34197a <=( A200  and  (not A199) );
 a34198a <=( A166  and  a34197a );
 a34199a <=( a34198a  and  a34193a );
 a34203a <=( (not A236)  and  (not A235) );
 a34204a <=( (not A233)  and  a34203a );
 a34207a <=( A266  and  A265 );
 a34210a <=( A299  and  (not A298) );
 a34211a <=( a34210a  and  a34207a );
 a34212a <=( a34211a  and  a34204a );
 a34216a <=( (not A167)  and  (not A168) );
 a34217a <=( (not A170)  and  a34216a );
 a34221a <=( A200  and  (not A199) );
 a34222a <=( A166  and  a34221a );
 a34223a <=( a34222a  and  a34217a );
 a34227a <=( (not A236)  and  (not A235) );
 a34228a <=( (not A233)  and  a34227a );
 a34231a <=( (not A267)  and  (not A266) );
 a34234a <=( A299  and  (not A298) );
 a34235a <=( a34234a  and  a34231a );
 a34236a <=( a34235a  and  a34228a );
 a34240a <=( (not A167)  and  (not A168) );
 a34241a <=( (not A170)  and  a34240a );
 a34245a <=( A200  and  (not A199) );
 a34246a <=( A166  and  a34245a );
 a34247a <=( a34246a  and  a34241a );
 a34251a <=( (not A236)  and  (not A235) );
 a34252a <=( (not A233)  and  a34251a );
 a34255a <=( (not A266)  and  (not A265) );
 a34258a <=( A299  and  (not A298) );
 a34259a <=( a34258a  and  a34255a );
 a34260a <=( a34259a  and  a34252a );
 a34264a <=( (not A167)  and  (not A168) );
 a34265a <=( (not A170)  and  a34264a );
 a34269a <=( A200  and  (not A199) );
 a34270a <=( A166  and  a34269a );
 a34271a <=( a34270a  and  a34265a );
 a34275a <=( (not A266)  and  (not A234) );
 a34276a <=( (not A233)  and  a34275a );
 a34279a <=( (not A269)  and  (not A268) );
 a34282a <=( A299  and  (not A298) );
 a34283a <=( a34282a  and  a34279a );
 a34284a <=( a34283a  and  a34276a );
 a34288a <=( (not A167)  and  (not A168) );
 a34289a <=( (not A170)  and  a34288a );
 a34293a <=( A200  and  (not A199) );
 a34294a <=( A166  and  a34293a );
 a34295a <=( a34294a  and  a34289a );
 a34299a <=( A234  and  (not A233) );
 a34300a <=( A232  and  a34299a );
 a34303a <=( A298  and  A235 );
 a34306a <=( (not A302)  and  (not A301) );
 a34307a <=( a34306a  and  a34303a );
 a34308a <=( a34307a  and  a34300a );
 a34312a <=( (not A167)  and  (not A168) );
 a34313a <=( (not A170)  and  a34312a );
 a34317a <=( A200  and  (not A199) );
 a34318a <=( A166  and  a34317a );
 a34319a <=( a34318a  and  a34313a );
 a34323a <=( A234  and  (not A233) );
 a34324a <=( A232  and  a34323a );
 a34327a <=( A298  and  A236 );
 a34330a <=( (not A302)  and  (not A301) );
 a34331a <=( a34330a  and  a34327a );
 a34332a <=( a34331a  and  a34324a );
 a34336a <=( (not A167)  and  (not A168) );
 a34337a <=( (not A170)  and  a34336a );
 a34341a <=( A200  and  (not A199) );
 a34342a <=( A166  and  a34341a );
 a34343a <=( a34342a  and  a34337a );
 a34347a <=( (not A266)  and  (not A233) );
 a34348a <=( (not A232)  and  a34347a );
 a34351a <=( (not A269)  and  (not A268) );
 a34354a <=( A299  and  (not A298) );
 a34355a <=( a34354a  and  a34351a );
 a34356a <=( a34355a  and  a34348a );
 a34360a <=( A167  and  (not A168) );
 a34361a <=( A169  and  a34360a );
 a34365a <=( A200  and  (not A199) );
 a34366a <=( (not A166)  and  a34365a );
 a34367a <=( a34366a  and  a34361a );
 a34371a <=( A265  and  A233 );
 a34372a <=( A232  and  a34371a );
 a34375a <=( (not A269)  and  (not A268) );
 a34378a <=( A299  and  (not A298) );
 a34379a <=( a34378a  and  a34375a );
 a34380a <=( a34379a  and  a34372a );
 a34384a <=( A167  and  (not A168) );
 a34385a <=( A169  and  a34384a );
 a34389a <=( A200  and  (not A199) );
 a34390a <=( (not A166)  and  a34389a );
 a34391a <=( a34390a  and  a34385a );
 a34395a <=( (not A236)  and  (not A235) );
 a34396a <=( (not A233)  and  a34395a );
 a34399a <=( A266  and  A265 );
 a34402a <=( A299  and  (not A298) );
 a34403a <=( a34402a  and  a34399a );
 a34404a <=( a34403a  and  a34396a );
 a34408a <=( A167  and  (not A168) );
 a34409a <=( A169  and  a34408a );
 a34413a <=( A200  and  (not A199) );
 a34414a <=( (not A166)  and  a34413a );
 a34415a <=( a34414a  and  a34409a );
 a34419a <=( (not A236)  and  (not A235) );
 a34420a <=( (not A233)  and  a34419a );
 a34423a <=( (not A267)  and  (not A266) );
 a34426a <=( A299  and  (not A298) );
 a34427a <=( a34426a  and  a34423a );
 a34428a <=( a34427a  and  a34420a );
 a34432a <=( A167  and  (not A168) );
 a34433a <=( A169  and  a34432a );
 a34437a <=( A200  and  (not A199) );
 a34438a <=( (not A166)  and  a34437a );
 a34439a <=( a34438a  and  a34433a );
 a34443a <=( (not A236)  and  (not A235) );
 a34444a <=( (not A233)  and  a34443a );
 a34447a <=( (not A266)  and  (not A265) );
 a34450a <=( A299  and  (not A298) );
 a34451a <=( a34450a  and  a34447a );
 a34452a <=( a34451a  and  a34444a );
 a34456a <=( A167  and  (not A168) );
 a34457a <=( A169  and  a34456a );
 a34461a <=( A200  and  (not A199) );
 a34462a <=( (not A166)  and  a34461a );
 a34463a <=( a34462a  and  a34457a );
 a34467a <=( (not A266)  and  (not A234) );
 a34468a <=( (not A233)  and  a34467a );
 a34471a <=( (not A269)  and  (not A268) );
 a34474a <=( A299  and  (not A298) );
 a34475a <=( a34474a  and  a34471a );
 a34476a <=( a34475a  and  a34468a );
 a34480a <=( A167  and  (not A168) );
 a34481a <=( A169  and  a34480a );
 a34485a <=( A200  and  (not A199) );
 a34486a <=( (not A166)  and  a34485a );
 a34487a <=( a34486a  and  a34481a );
 a34491a <=( A234  and  (not A233) );
 a34492a <=( A232  and  a34491a );
 a34495a <=( A298  and  A235 );
 a34498a <=( (not A302)  and  (not A301) );
 a34499a <=( a34498a  and  a34495a );
 a34500a <=( a34499a  and  a34492a );
 a34504a <=( A167  and  (not A168) );
 a34505a <=( A169  and  a34504a );
 a34509a <=( A200  and  (not A199) );
 a34510a <=( (not A166)  and  a34509a );
 a34511a <=( a34510a  and  a34505a );
 a34515a <=( A234  and  (not A233) );
 a34516a <=( A232  and  a34515a );
 a34519a <=( A298  and  A236 );
 a34522a <=( (not A302)  and  (not A301) );
 a34523a <=( a34522a  and  a34519a );
 a34524a <=( a34523a  and  a34516a );
 a34528a <=( A167  and  (not A168) );
 a34529a <=( A169  and  a34528a );
 a34533a <=( A200  and  (not A199) );
 a34534a <=( (not A166)  and  a34533a );
 a34535a <=( a34534a  and  a34529a );
 a34539a <=( (not A266)  and  (not A233) );
 a34540a <=( (not A232)  and  a34539a );
 a34543a <=( (not A269)  and  (not A268) );
 a34546a <=( A299  and  (not A298) );
 a34547a <=( a34546a  and  a34543a );
 a34548a <=( a34547a  and  a34540a );
 a34552a <=( A167  and  (not A168) );
 a34553a <=( A169  and  a34552a );
 a34557a <=( (not A200)  and  A199 );
 a34558a <=( (not A166)  and  a34557a );
 a34559a <=( a34558a  and  a34553a );
 a34563a <=( (not A232)  and  A202 );
 a34564a <=( A201  and  a34563a );
 a34567a <=( (not A299)  and  A233 );
 a34570a <=( (not A302)  and  (not A301) );
 a34571a <=( a34570a  and  a34567a );
 a34572a <=( a34571a  and  a34564a );
 a34576a <=( A167  and  (not A168) );
 a34577a <=( A169  and  a34576a );
 a34581a <=( (not A200)  and  A199 );
 a34582a <=( (not A166)  and  a34581a );
 a34583a <=( a34582a  and  a34577a );
 a34587a <=( (not A232)  and  A203 );
 a34588a <=( A201  and  a34587a );
 a34591a <=( (not A299)  and  A233 );
 a34594a <=( (not A302)  and  (not A301) );
 a34595a <=( a34594a  and  a34591a );
 a34596a <=( a34595a  and  a34588a );
 a34600a <=( (not A167)  and  (not A168) );
 a34601a <=( A169  and  a34600a );
 a34605a <=( A200  and  (not A199) );
 a34606a <=( A166  and  a34605a );
 a34607a <=( a34606a  and  a34601a );
 a34611a <=( A265  and  A233 );
 a34612a <=( A232  and  a34611a );
 a34615a <=( (not A269)  and  (not A268) );
 a34618a <=( A299  and  (not A298) );
 a34619a <=( a34618a  and  a34615a );
 a34620a <=( a34619a  and  a34612a );
 a34624a <=( (not A167)  and  (not A168) );
 a34625a <=( A169  and  a34624a );
 a34629a <=( A200  and  (not A199) );
 a34630a <=( A166  and  a34629a );
 a34631a <=( a34630a  and  a34625a );
 a34635a <=( (not A236)  and  (not A235) );
 a34636a <=( (not A233)  and  a34635a );
 a34639a <=( A266  and  A265 );
 a34642a <=( A299  and  (not A298) );
 a34643a <=( a34642a  and  a34639a );
 a34644a <=( a34643a  and  a34636a );
 a34648a <=( (not A167)  and  (not A168) );
 a34649a <=( A169  and  a34648a );
 a34653a <=( A200  and  (not A199) );
 a34654a <=( A166  and  a34653a );
 a34655a <=( a34654a  and  a34649a );
 a34659a <=( (not A236)  and  (not A235) );
 a34660a <=( (not A233)  and  a34659a );
 a34663a <=( (not A267)  and  (not A266) );
 a34666a <=( A299  and  (not A298) );
 a34667a <=( a34666a  and  a34663a );
 a34668a <=( a34667a  and  a34660a );
 a34672a <=( (not A167)  and  (not A168) );
 a34673a <=( A169  and  a34672a );
 a34677a <=( A200  and  (not A199) );
 a34678a <=( A166  and  a34677a );
 a34679a <=( a34678a  and  a34673a );
 a34683a <=( (not A236)  and  (not A235) );
 a34684a <=( (not A233)  and  a34683a );
 a34687a <=( (not A266)  and  (not A265) );
 a34690a <=( A299  and  (not A298) );
 a34691a <=( a34690a  and  a34687a );
 a34692a <=( a34691a  and  a34684a );
 a34696a <=( (not A167)  and  (not A168) );
 a34697a <=( A169  and  a34696a );
 a34701a <=( A200  and  (not A199) );
 a34702a <=( A166  and  a34701a );
 a34703a <=( a34702a  and  a34697a );
 a34707a <=( (not A266)  and  (not A234) );
 a34708a <=( (not A233)  and  a34707a );
 a34711a <=( (not A269)  and  (not A268) );
 a34714a <=( A299  and  (not A298) );
 a34715a <=( a34714a  and  a34711a );
 a34716a <=( a34715a  and  a34708a );
 a34720a <=( (not A167)  and  (not A168) );
 a34721a <=( A169  and  a34720a );
 a34725a <=( A200  and  (not A199) );
 a34726a <=( A166  and  a34725a );
 a34727a <=( a34726a  and  a34721a );
 a34731a <=( A234  and  (not A233) );
 a34732a <=( A232  and  a34731a );
 a34735a <=( A298  and  A235 );
 a34738a <=( (not A302)  and  (not A301) );
 a34739a <=( a34738a  and  a34735a );
 a34740a <=( a34739a  and  a34732a );
 a34744a <=( (not A167)  and  (not A168) );
 a34745a <=( A169  and  a34744a );
 a34749a <=( A200  and  (not A199) );
 a34750a <=( A166  and  a34749a );
 a34751a <=( a34750a  and  a34745a );
 a34755a <=( A234  and  (not A233) );
 a34756a <=( A232  and  a34755a );
 a34759a <=( A298  and  A236 );
 a34762a <=( (not A302)  and  (not A301) );
 a34763a <=( a34762a  and  a34759a );
 a34764a <=( a34763a  and  a34756a );
 a34768a <=( (not A167)  and  (not A168) );
 a34769a <=( A169  and  a34768a );
 a34773a <=( A200  and  (not A199) );
 a34774a <=( A166  and  a34773a );
 a34775a <=( a34774a  and  a34769a );
 a34779a <=( (not A266)  and  (not A233) );
 a34780a <=( (not A232)  and  a34779a );
 a34783a <=( (not A269)  and  (not A268) );
 a34786a <=( A299  and  (not A298) );
 a34787a <=( a34786a  and  a34783a );
 a34788a <=( a34787a  and  a34780a );
 a34792a <=( (not A167)  and  (not A168) );
 a34793a <=( A169  and  a34792a );
 a34797a <=( (not A200)  and  A199 );
 a34798a <=( A166  and  a34797a );
 a34799a <=( a34798a  and  a34793a );
 a34803a <=( (not A232)  and  A202 );
 a34804a <=( A201  and  a34803a );
 a34807a <=( (not A299)  and  A233 );
 a34810a <=( (not A302)  and  (not A301) );
 a34811a <=( a34810a  and  a34807a );
 a34812a <=( a34811a  and  a34804a );
 a34816a <=( (not A167)  and  (not A168) );
 a34817a <=( A169  and  a34816a );
 a34821a <=( (not A200)  and  A199 );
 a34822a <=( A166  and  a34821a );
 a34823a <=( a34822a  and  a34817a );
 a34827a <=( (not A232)  and  A203 );
 a34828a <=( A201  and  a34827a );
 a34831a <=( (not A299)  and  A233 );
 a34834a <=( (not A302)  and  (not A301) );
 a34835a <=( a34834a  and  a34831a );
 a34836a <=( a34835a  and  a34828a );
 a34840a <=( (not A168)  and  A169 );
 a34841a <=( A170  and  a34840a );
 a34845a <=( A201  and  (not A200) );
 a34846a <=( A199  and  a34845a );
 a34847a <=( a34846a  and  a34841a );
 a34851a <=( A233  and  A232 );
 a34852a <=( A202  and  a34851a );
 a34855a <=( (not A267)  and  A265 );
 a34858a <=( A299  and  (not A298) );
 a34859a <=( a34858a  and  a34855a );
 a34860a <=( a34859a  and  a34852a );
 a34864a <=( (not A168)  and  A169 );
 a34865a <=( A170  and  a34864a );
 a34869a <=( A201  and  (not A200) );
 a34870a <=( A199  and  a34869a );
 a34871a <=( a34870a  and  a34865a );
 a34875a <=( A233  and  A232 );
 a34876a <=( A202  and  a34875a );
 a34879a <=( A266  and  A265 );
 a34882a <=( A299  and  (not A298) );
 a34883a <=( a34882a  and  a34879a );
 a34884a <=( a34883a  and  a34876a );
 a34888a <=( (not A168)  and  A169 );
 a34889a <=( A170  and  a34888a );
 a34893a <=( A201  and  (not A200) );
 a34894a <=( A199  and  a34893a );
 a34895a <=( a34894a  and  a34889a );
 a34899a <=( A233  and  A232 );
 a34900a <=( A202  and  a34899a );
 a34903a <=( (not A266)  and  (not A265) );
 a34906a <=( A299  and  (not A298) );
 a34907a <=( a34906a  and  a34903a );
 a34908a <=( a34907a  and  a34900a );
 a34912a <=( (not A168)  and  A169 );
 a34913a <=( A170  and  a34912a );
 a34917a <=( A201  and  (not A200) );
 a34918a <=( A199  and  a34917a );
 a34919a <=( a34918a  and  a34913a );
 a34923a <=( A233  and  (not A232) );
 a34924a <=( A202  and  a34923a );
 a34927a <=( (not A266)  and  A265 );
 a34930a <=( A268  and  A267 );
 a34931a <=( a34930a  and  a34927a );
 a34932a <=( a34931a  and  a34924a );
 a34936a <=( (not A168)  and  A169 );
 a34937a <=( A170  and  a34936a );
 a34941a <=( A201  and  (not A200) );
 a34942a <=( A199  and  a34941a );
 a34943a <=( a34942a  and  a34937a );
 a34947a <=( A233  and  (not A232) );
 a34948a <=( A202  and  a34947a );
 a34951a <=( (not A266)  and  A265 );
 a34954a <=( A269  and  A267 );
 a34955a <=( a34954a  and  a34951a );
 a34956a <=( a34955a  and  a34948a );
 a34960a <=( (not A168)  and  A169 );
 a34961a <=( A170  and  a34960a );
 a34965a <=( A201  and  (not A200) );
 a34966a <=( A199  and  a34965a );
 a34967a <=( a34966a  and  a34961a );
 a34971a <=( (not A234)  and  (not A233) );
 a34972a <=( A202  and  a34971a );
 a34975a <=( A266  and  A265 );
 a34978a <=( A299  and  (not A298) );
 a34979a <=( a34978a  and  a34975a );
 a34980a <=( a34979a  and  a34972a );
 a34984a <=( (not A168)  and  A169 );
 a34985a <=( A170  and  a34984a );
 a34989a <=( A201  and  (not A200) );
 a34990a <=( A199  and  a34989a );
 a34991a <=( a34990a  and  a34985a );
 a34995a <=( (not A234)  and  (not A233) );
 a34996a <=( A202  and  a34995a );
 a34999a <=( (not A267)  and  (not A266) );
 a35002a <=( A299  and  (not A298) );
 a35003a <=( a35002a  and  a34999a );
 a35004a <=( a35003a  and  a34996a );
 a35008a <=( (not A168)  and  A169 );
 a35009a <=( A170  and  a35008a );
 a35013a <=( A201  and  (not A200) );
 a35014a <=( A199  and  a35013a );
 a35015a <=( a35014a  and  a35009a );
 a35019a <=( (not A234)  and  (not A233) );
 a35020a <=( A202  and  a35019a );
 a35023a <=( (not A266)  and  (not A265) );
 a35026a <=( A299  and  (not A298) );
 a35027a <=( a35026a  and  a35023a );
 a35028a <=( a35027a  and  a35020a );
 a35032a <=( (not A168)  and  A169 );
 a35033a <=( A170  and  a35032a );
 a35037a <=( A201  and  (not A200) );
 a35038a <=( A199  and  a35037a );
 a35039a <=( a35038a  and  a35033a );
 a35043a <=( (not A233)  and  A232 );
 a35044a <=( A202  and  a35043a );
 a35047a <=( A235  and  A234 );
 a35050a <=( (not A300)  and  A298 );
 a35051a <=( a35050a  and  a35047a );
 a35052a <=( a35051a  and  a35044a );
 a35056a <=( (not A168)  and  A169 );
 a35057a <=( A170  and  a35056a );
 a35061a <=( A201  and  (not A200) );
 a35062a <=( A199  and  a35061a );
 a35063a <=( a35062a  and  a35057a );
 a35067a <=( (not A233)  and  A232 );
 a35068a <=( A202  and  a35067a );
 a35071a <=( A235  and  A234 );
 a35074a <=( A299  and  A298 );
 a35075a <=( a35074a  and  a35071a );
 a35076a <=( a35075a  and  a35068a );
 a35080a <=( (not A168)  and  A169 );
 a35081a <=( A170  and  a35080a );
 a35085a <=( A201  and  (not A200) );
 a35086a <=( A199  and  a35085a );
 a35087a <=( a35086a  and  a35081a );
 a35091a <=( (not A233)  and  A232 );
 a35092a <=( A202  and  a35091a );
 a35095a <=( A235  and  A234 );
 a35098a <=( (not A299)  and  (not A298) );
 a35099a <=( a35098a  and  a35095a );
 a35100a <=( a35099a  and  a35092a );
 a35104a <=( (not A168)  and  A169 );
 a35105a <=( A170  and  a35104a );
 a35109a <=( A201  and  (not A200) );
 a35110a <=( A199  and  a35109a );
 a35111a <=( a35110a  and  a35105a );
 a35115a <=( (not A233)  and  A232 );
 a35116a <=( A202  and  a35115a );
 a35119a <=( A235  and  A234 );
 a35122a <=( A266  and  (not A265) );
 a35123a <=( a35122a  and  a35119a );
 a35124a <=( a35123a  and  a35116a );
 a35128a <=( (not A168)  and  A169 );
 a35129a <=( A170  and  a35128a );
 a35133a <=( A201  and  (not A200) );
 a35134a <=( A199  and  a35133a );
 a35135a <=( a35134a  and  a35129a );
 a35139a <=( (not A233)  and  A232 );
 a35140a <=( A202  and  a35139a );
 a35143a <=( A236  and  A234 );
 a35146a <=( (not A300)  and  A298 );
 a35147a <=( a35146a  and  a35143a );
 a35148a <=( a35147a  and  a35140a );
 a35152a <=( (not A168)  and  A169 );
 a35153a <=( A170  and  a35152a );
 a35157a <=( A201  and  (not A200) );
 a35158a <=( A199  and  a35157a );
 a35159a <=( a35158a  and  a35153a );
 a35163a <=( (not A233)  and  A232 );
 a35164a <=( A202  and  a35163a );
 a35167a <=( A236  and  A234 );
 a35170a <=( A299  and  A298 );
 a35171a <=( a35170a  and  a35167a );
 a35172a <=( a35171a  and  a35164a );
 a35176a <=( (not A168)  and  A169 );
 a35177a <=( A170  and  a35176a );
 a35181a <=( A201  and  (not A200) );
 a35182a <=( A199  and  a35181a );
 a35183a <=( a35182a  and  a35177a );
 a35187a <=( (not A233)  and  A232 );
 a35188a <=( A202  and  a35187a );
 a35191a <=( A236  and  A234 );
 a35194a <=( (not A299)  and  (not A298) );
 a35195a <=( a35194a  and  a35191a );
 a35196a <=( a35195a  and  a35188a );
 a35200a <=( (not A168)  and  A169 );
 a35201a <=( A170  and  a35200a );
 a35205a <=( A201  and  (not A200) );
 a35206a <=( A199  and  a35205a );
 a35207a <=( a35206a  and  a35201a );
 a35211a <=( (not A233)  and  A232 );
 a35212a <=( A202  and  a35211a );
 a35215a <=( A236  and  A234 );
 a35218a <=( A266  and  (not A265) );
 a35219a <=( a35218a  and  a35215a );
 a35220a <=( a35219a  and  a35212a );
 a35224a <=( (not A168)  and  A169 );
 a35225a <=( A170  and  a35224a );
 a35229a <=( A201  and  (not A200) );
 a35230a <=( A199  and  a35229a );
 a35231a <=( a35230a  and  a35225a );
 a35235a <=( (not A233)  and  (not A232) );
 a35236a <=( A202  and  a35235a );
 a35239a <=( A266  and  A265 );
 a35242a <=( A299  and  (not A298) );
 a35243a <=( a35242a  and  a35239a );
 a35244a <=( a35243a  and  a35236a );
 a35248a <=( (not A168)  and  A169 );
 a35249a <=( A170  and  a35248a );
 a35253a <=( A201  and  (not A200) );
 a35254a <=( A199  and  a35253a );
 a35255a <=( a35254a  and  a35249a );
 a35259a <=( (not A233)  and  (not A232) );
 a35260a <=( A202  and  a35259a );
 a35263a <=( (not A267)  and  (not A266) );
 a35266a <=( A299  and  (not A298) );
 a35267a <=( a35266a  and  a35263a );
 a35268a <=( a35267a  and  a35260a );
 a35272a <=( (not A168)  and  A169 );
 a35273a <=( A170  and  a35272a );
 a35277a <=( A201  and  (not A200) );
 a35278a <=( A199  and  a35277a );
 a35279a <=( a35278a  and  a35273a );
 a35283a <=( (not A233)  and  (not A232) );
 a35284a <=( A202  and  a35283a );
 a35287a <=( (not A266)  and  (not A265) );
 a35290a <=( A299  and  (not A298) );
 a35291a <=( a35290a  and  a35287a );
 a35292a <=( a35291a  and  a35284a );
 a35296a <=( (not A168)  and  A169 );
 a35297a <=( A170  and  a35296a );
 a35301a <=( A201  and  (not A200) );
 a35302a <=( A199  and  a35301a );
 a35303a <=( a35302a  and  a35297a );
 a35307a <=( A233  and  A232 );
 a35308a <=( A203  and  a35307a );
 a35311a <=( (not A267)  and  A265 );
 a35314a <=( A299  and  (not A298) );
 a35315a <=( a35314a  and  a35311a );
 a35316a <=( a35315a  and  a35308a );
 a35320a <=( (not A168)  and  A169 );
 a35321a <=( A170  and  a35320a );
 a35325a <=( A201  and  (not A200) );
 a35326a <=( A199  and  a35325a );
 a35327a <=( a35326a  and  a35321a );
 a35331a <=( A233  and  A232 );
 a35332a <=( A203  and  a35331a );
 a35335a <=( A266  and  A265 );
 a35338a <=( A299  and  (not A298) );
 a35339a <=( a35338a  and  a35335a );
 a35340a <=( a35339a  and  a35332a );
 a35344a <=( (not A168)  and  A169 );
 a35345a <=( A170  and  a35344a );
 a35349a <=( A201  and  (not A200) );
 a35350a <=( A199  and  a35349a );
 a35351a <=( a35350a  and  a35345a );
 a35355a <=( A233  and  A232 );
 a35356a <=( A203  and  a35355a );
 a35359a <=( (not A266)  and  (not A265) );
 a35362a <=( A299  and  (not A298) );
 a35363a <=( a35362a  and  a35359a );
 a35364a <=( a35363a  and  a35356a );
 a35368a <=( (not A168)  and  A169 );
 a35369a <=( A170  and  a35368a );
 a35373a <=( A201  and  (not A200) );
 a35374a <=( A199  and  a35373a );
 a35375a <=( a35374a  and  a35369a );
 a35379a <=( A233  and  (not A232) );
 a35380a <=( A203  and  a35379a );
 a35383a <=( (not A266)  and  A265 );
 a35386a <=( A268  and  A267 );
 a35387a <=( a35386a  and  a35383a );
 a35388a <=( a35387a  and  a35380a );
 a35392a <=( (not A168)  and  A169 );
 a35393a <=( A170  and  a35392a );
 a35397a <=( A201  and  (not A200) );
 a35398a <=( A199  and  a35397a );
 a35399a <=( a35398a  and  a35393a );
 a35403a <=( A233  and  (not A232) );
 a35404a <=( A203  and  a35403a );
 a35407a <=( (not A266)  and  A265 );
 a35410a <=( A269  and  A267 );
 a35411a <=( a35410a  and  a35407a );
 a35412a <=( a35411a  and  a35404a );
 a35416a <=( (not A168)  and  A169 );
 a35417a <=( A170  and  a35416a );
 a35421a <=( A201  and  (not A200) );
 a35422a <=( A199  and  a35421a );
 a35423a <=( a35422a  and  a35417a );
 a35427a <=( (not A234)  and  (not A233) );
 a35428a <=( A203  and  a35427a );
 a35431a <=( A266  and  A265 );
 a35434a <=( A299  and  (not A298) );
 a35435a <=( a35434a  and  a35431a );
 a35436a <=( a35435a  and  a35428a );
 a35440a <=( (not A168)  and  A169 );
 a35441a <=( A170  and  a35440a );
 a35445a <=( A201  and  (not A200) );
 a35446a <=( A199  and  a35445a );
 a35447a <=( a35446a  and  a35441a );
 a35451a <=( (not A234)  and  (not A233) );
 a35452a <=( A203  and  a35451a );
 a35455a <=( (not A267)  and  (not A266) );
 a35458a <=( A299  and  (not A298) );
 a35459a <=( a35458a  and  a35455a );
 a35460a <=( a35459a  and  a35452a );
 a35464a <=( (not A168)  and  A169 );
 a35465a <=( A170  and  a35464a );
 a35469a <=( A201  and  (not A200) );
 a35470a <=( A199  and  a35469a );
 a35471a <=( a35470a  and  a35465a );
 a35475a <=( (not A234)  and  (not A233) );
 a35476a <=( A203  and  a35475a );
 a35479a <=( (not A266)  and  (not A265) );
 a35482a <=( A299  and  (not A298) );
 a35483a <=( a35482a  and  a35479a );
 a35484a <=( a35483a  and  a35476a );
 a35488a <=( (not A168)  and  A169 );
 a35489a <=( A170  and  a35488a );
 a35493a <=( A201  and  (not A200) );
 a35494a <=( A199  and  a35493a );
 a35495a <=( a35494a  and  a35489a );
 a35499a <=( (not A233)  and  A232 );
 a35500a <=( A203  and  a35499a );
 a35503a <=( A235  and  A234 );
 a35506a <=( (not A300)  and  A298 );
 a35507a <=( a35506a  and  a35503a );
 a35508a <=( a35507a  and  a35500a );
 a35512a <=( (not A168)  and  A169 );
 a35513a <=( A170  and  a35512a );
 a35517a <=( A201  and  (not A200) );
 a35518a <=( A199  and  a35517a );
 a35519a <=( a35518a  and  a35513a );
 a35523a <=( (not A233)  and  A232 );
 a35524a <=( A203  and  a35523a );
 a35527a <=( A235  and  A234 );
 a35530a <=( A299  and  A298 );
 a35531a <=( a35530a  and  a35527a );
 a35532a <=( a35531a  and  a35524a );
 a35536a <=( (not A168)  and  A169 );
 a35537a <=( A170  and  a35536a );
 a35541a <=( A201  and  (not A200) );
 a35542a <=( A199  and  a35541a );
 a35543a <=( a35542a  and  a35537a );
 a35547a <=( (not A233)  and  A232 );
 a35548a <=( A203  and  a35547a );
 a35551a <=( A235  and  A234 );
 a35554a <=( (not A299)  and  (not A298) );
 a35555a <=( a35554a  and  a35551a );
 a35556a <=( a35555a  and  a35548a );
 a35560a <=( (not A168)  and  A169 );
 a35561a <=( A170  and  a35560a );
 a35565a <=( A201  and  (not A200) );
 a35566a <=( A199  and  a35565a );
 a35567a <=( a35566a  and  a35561a );
 a35571a <=( (not A233)  and  A232 );
 a35572a <=( A203  and  a35571a );
 a35575a <=( A235  and  A234 );
 a35578a <=( A266  and  (not A265) );
 a35579a <=( a35578a  and  a35575a );
 a35580a <=( a35579a  and  a35572a );
 a35584a <=( (not A168)  and  A169 );
 a35585a <=( A170  and  a35584a );
 a35589a <=( A201  and  (not A200) );
 a35590a <=( A199  and  a35589a );
 a35591a <=( a35590a  and  a35585a );
 a35595a <=( (not A233)  and  A232 );
 a35596a <=( A203  and  a35595a );
 a35599a <=( A236  and  A234 );
 a35602a <=( (not A300)  and  A298 );
 a35603a <=( a35602a  and  a35599a );
 a35604a <=( a35603a  and  a35596a );
 a35608a <=( (not A168)  and  A169 );
 a35609a <=( A170  and  a35608a );
 a35613a <=( A201  and  (not A200) );
 a35614a <=( A199  and  a35613a );
 a35615a <=( a35614a  and  a35609a );
 a35619a <=( (not A233)  and  A232 );
 a35620a <=( A203  and  a35619a );
 a35623a <=( A236  and  A234 );
 a35626a <=( A299  and  A298 );
 a35627a <=( a35626a  and  a35623a );
 a35628a <=( a35627a  and  a35620a );
 a35632a <=( (not A168)  and  A169 );
 a35633a <=( A170  and  a35632a );
 a35637a <=( A201  and  (not A200) );
 a35638a <=( A199  and  a35637a );
 a35639a <=( a35638a  and  a35633a );
 a35643a <=( (not A233)  and  A232 );
 a35644a <=( A203  and  a35643a );
 a35647a <=( A236  and  A234 );
 a35650a <=( (not A299)  and  (not A298) );
 a35651a <=( a35650a  and  a35647a );
 a35652a <=( a35651a  and  a35644a );
 a35656a <=( (not A168)  and  A169 );
 a35657a <=( A170  and  a35656a );
 a35661a <=( A201  and  (not A200) );
 a35662a <=( A199  and  a35661a );
 a35663a <=( a35662a  and  a35657a );
 a35667a <=( (not A233)  and  A232 );
 a35668a <=( A203  and  a35667a );
 a35671a <=( A236  and  A234 );
 a35674a <=( A266  and  (not A265) );
 a35675a <=( a35674a  and  a35671a );
 a35676a <=( a35675a  and  a35668a );
 a35680a <=( (not A168)  and  A169 );
 a35681a <=( A170  and  a35680a );
 a35685a <=( A201  and  (not A200) );
 a35686a <=( A199  and  a35685a );
 a35687a <=( a35686a  and  a35681a );
 a35691a <=( (not A233)  and  (not A232) );
 a35692a <=( A203  and  a35691a );
 a35695a <=( A266  and  A265 );
 a35698a <=( A299  and  (not A298) );
 a35699a <=( a35698a  and  a35695a );
 a35700a <=( a35699a  and  a35692a );
 a35704a <=( (not A168)  and  A169 );
 a35705a <=( A170  and  a35704a );
 a35709a <=( A201  and  (not A200) );
 a35710a <=( A199  and  a35709a );
 a35711a <=( a35710a  and  a35705a );
 a35715a <=( (not A233)  and  (not A232) );
 a35716a <=( A203  and  a35715a );
 a35719a <=( (not A267)  and  (not A266) );
 a35722a <=( A299  and  (not A298) );
 a35723a <=( a35722a  and  a35719a );
 a35724a <=( a35723a  and  a35716a );
 a35728a <=( (not A168)  and  A169 );
 a35729a <=( A170  and  a35728a );
 a35733a <=( A201  and  (not A200) );
 a35734a <=( A199  and  a35733a );
 a35735a <=( a35734a  and  a35729a );
 a35739a <=( (not A233)  and  (not A232) );
 a35740a <=( A203  and  a35739a );
 a35743a <=( (not A266)  and  (not A265) );
 a35746a <=( A299  and  (not A298) );
 a35747a <=( a35746a  and  a35743a );
 a35748a <=( a35747a  and  a35740a );
 a35752a <=( A167  and  A169 );
 a35753a <=( (not A170)  and  a35752a );
 a35757a <=( A200  and  A199 );
 a35758a <=( A166  and  a35757a );
 a35759a <=( a35758a  and  a35753a );
 a35763a <=( A265  and  A233 );
 a35764a <=( A232  and  a35763a );
 a35767a <=( (not A269)  and  (not A268) );
 a35770a <=( A299  and  (not A298) );
 a35771a <=( a35770a  and  a35767a );
 a35772a <=( a35771a  and  a35764a );
 a35776a <=( A167  and  A169 );
 a35777a <=( (not A170)  and  a35776a );
 a35781a <=( A200  and  A199 );
 a35782a <=( A166  and  a35781a );
 a35783a <=( a35782a  and  a35777a );
 a35787a <=( (not A236)  and  (not A235) );
 a35788a <=( (not A233)  and  a35787a );
 a35791a <=( A266  and  A265 );
 a35794a <=( A299  and  (not A298) );
 a35795a <=( a35794a  and  a35791a );
 a35796a <=( a35795a  and  a35788a );
 a35800a <=( A167  and  A169 );
 a35801a <=( (not A170)  and  a35800a );
 a35805a <=( A200  and  A199 );
 a35806a <=( A166  and  a35805a );
 a35807a <=( a35806a  and  a35801a );
 a35811a <=( (not A236)  and  (not A235) );
 a35812a <=( (not A233)  and  a35811a );
 a35815a <=( (not A267)  and  (not A266) );
 a35818a <=( A299  and  (not A298) );
 a35819a <=( a35818a  and  a35815a );
 a35820a <=( a35819a  and  a35812a );
 a35824a <=( A167  and  A169 );
 a35825a <=( (not A170)  and  a35824a );
 a35829a <=( A200  and  A199 );
 a35830a <=( A166  and  a35829a );
 a35831a <=( a35830a  and  a35825a );
 a35835a <=( (not A236)  and  (not A235) );
 a35836a <=( (not A233)  and  a35835a );
 a35839a <=( (not A266)  and  (not A265) );
 a35842a <=( A299  and  (not A298) );
 a35843a <=( a35842a  and  a35839a );
 a35844a <=( a35843a  and  a35836a );
 a35848a <=( A167  and  A169 );
 a35849a <=( (not A170)  and  a35848a );
 a35853a <=( A200  and  A199 );
 a35854a <=( A166  and  a35853a );
 a35855a <=( a35854a  and  a35849a );
 a35859a <=( (not A266)  and  (not A234) );
 a35860a <=( (not A233)  and  a35859a );
 a35863a <=( (not A269)  and  (not A268) );
 a35866a <=( A299  and  (not A298) );
 a35867a <=( a35866a  and  a35863a );
 a35868a <=( a35867a  and  a35860a );
 a35872a <=( A167  and  A169 );
 a35873a <=( (not A170)  and  a35872a );
 a35877a <=( A200  and  A199 );
 a35878a <=( A166  and  a35877a );
 a35879a <=( a35878a  and  a35873a );
 a35883a <=( A234  and  (not A233) );
 a35884a <=( A232  and  a35883a );
 a35887a <=( A298  and  A235 );
 a35890a <=( (not A302)  and  (not A301) );
 a35891a <=( a35890a  and  a35887a );
 a35892a <=( a35891a  and  a35884a );
 a35896a <=( A167  and  A169 );
 a35897a <=( (not A170)  and  a35896a );
 a35901a <=( A200  and  A199 );
 a35902a <=( A166  and  a35901a );
 a35903a <=( a35902a  and  a35897a );
 a35907a <=( A234  and  (not A233) );
 a35908a <=( A232  and  a35907a );
 a35911a <=( A298  and  A236 );
 a35914a <=( (not A302)  and  (not A301) );
 a35915a <=( a35914a  and  a35911a );
 a35916a <=( a35915a  and  a35908a );
 a35920a <=( A167  and  A169 );
 a35921a <=( (not A170)  and  a35920a );
 a35925a <=( A200  and  A199 );
 a35926a <=( A166  and  a35925a );
 a35927a <=( a35926a  and  a35921a );
 a35931a <=( (not A266)  and  (not A233) );
 a35932a <=( (not A232)  and  a35931a );
 a35935a <=( (not A269)  and  (not A268) );
 a35938a <=( A299  and  (not A298) );
 a35939a <=( a35938a  and  a35935a );
 a35940a <=( a35939a  and  a35932a );
 a35944a <=( A167  and  A169 );
 a35945a <=( (not A170)  and  a35944a );
 a35949a <=( (not A202)  and  (not A200) );
 a35950a <=( A166  and  a35949a );
 a35951a <=( a35950a  and  a35945a );
 a35955a <=( A233  and  A232 );
 a35956a <=( (not A203)  and  a35955a );
 a35959a <=( (not A267)  and  A265 );
 a35962a <=( A299  and  (not A298) );
 a35963a <=( a35962a  and  a35959a );
 a35964a <=( a35963a  and  a35956a );
 a35968a <=( A167  and  A169 );
 a35969a <=( (not A170)  and  a35968a );
 a35973a <=( (not A202)  and  (not A200) );
 a35974a <=( A166  and  a35973a );
 a35975a <=( a35974a  and  a35969a );
 a35979a <=( A233  and  A232 );
 a35980a <=( (not A203)  and  a35979a );
 a35983a <=( A266  and  A265 );
 a35986a <=( A299  and  (not A298) );
 a35987a <=( a35986a  and  a35983a );
 a35988a <=( a35987a  and  a35980a );
 a35992a <=( A167  and  A169 );
 a35993a <=( (not A170)  and  a35992a );
 a35997a <=( (not A202)  and  (not A200) );
 a35998a <=( A166  and  a35997a );
 a35999a <=( a35998a  and  a35993a );
 a36003a <=( A233  and  A232 );
 a36004a <=( (not A203)  and  a36003a );
 a36007a <=( (not A266)  and  (not A265) );
 a36010a <=( A299  and  (not A298) );
 a36011a <=( a36010a  and  a36007a );
 a36012a <=( a36011a  and  a36004a );
 a36016a <=( A167  and  A169 );
 a36017a <=( (not A170)  and  a36016a );
 a36021a <=( (not A202)  and  (not A200) );
 a36022a <=( A166  and  a36021a );
 a36023a <=( a36022a  and  a36017a );
 a36027a <=( A233  and  (not A232) );
 a36028a <=( (not A203)  and  a36027a );
 a36031a <=( (not A266)  and  A265 );
 a36034a <=( A268  and  A267 );
 a36035a <=( a36034a  and  a36031a );
 a36036a <=( a36035a  and  a36028a );
 a36040a <=( A167  and  A169 );
 a36041a <=( (not A170)  and  a36040a );
 a36045a <=( (not A202)  and  (not A200) );
 a36046a <=( A166  and  a36045a );
 a36047a <=( a36046a  and  a36041a );
 a36051a <=( A233  and  (not A232) );
 a36052a <=( (not A203)  and  a36051a );
 a36055a <=( (not A266)  and  A265 );
 a36058a <=( A269  and  A267 );
 a36059a <=( a36058a  and  a36055a );
 a36060a <=( a36059a  and  a36052a );
 a36064a <=( A167  and  A169 );
 a36065a <=( (not A170)  and  a36064a );
 a36069a <=( (not A202)  and  (not A200) );
 a36070a <=( A166  and  a36069a );
 a36071a <=( a36070a  and  a36065a );
 a36075a <=( (not A234)  and  (not A233) );
 a36076a <=( (not A203)  and  a36075a );
 a36079a <=( A266  and  A265 );
 a36082a <=( A299  and  (not A298) );
 a36083a <=( a36082a  and  a36079a );
 a36084a <=( a36083a  and  a36076a );
 a36088a <=( A167  and  A169 );
 a36089a <=( (not A170)  and  a36088a );
 a36093a <=( (not A202)  and  (not A200) );
 a36094a <=( A166  and  a36093a );
 a36095a <=( a36094a  and  a36089a );
 a36099a <=( (not A234)  and  (not A233) );
 a36100a <=( (not A203)  and  a36099a );
 a36103a <=( (not A267)  and  (not A266) );
 a36106a <=( A299  and  (not A298) );
 a36107a <=( a36106a  and  a36103a );
 a36108a <=( a36107a  and  a36100a );
 a36112a <=( A167  and  A169 );
 a36113a <=( (not A170)  and  a36112a );
 a36117a <=( (not A202)  and  (not A200) );
 a36118a <=( A166  and  a36117a );
 a36119a <=( a36118a  and  a36113a );
 a36123a <=( (not A234)  and  (not A233) );
 a36124a <=( (not A203)  and  a36123a );
 a36127a <=( (not A266)  and  (not A265) );
 a36130a <=( A299  and  (not A298) );
 a36131a <=( a36130a  and  a36127a );
 a36132a <=( a36131a  and  a36124a );
 a36136a <=( A167  and  A169 );
 a36137a <=( (not A170)  and  a36136a );
 a36141a <=( (not A202)  and  (not A200) );
 a36142a <=( A166  and  a36141a );
 a36143a <=( a36142a  and  a36137a );
 a36147a <=( (not A233)  and  A232 );
 a36148a <=( (not A203)  and  a36147a );
 a36151a <=( A235  and  A234 );
 a36154a <=( (not A300)  and  A298 );
 a36155a <=( a36154a  and  a36151a );
 a36156a <=( a36155a  and  a36148a );
 a36160a <=( A167  and  A169 );
 a36161a <=( (not A170)  and  a36160a );
 a36165a <=( (not A202)  and  (not A200) );
 a36166a <=( A166  and  a36165a );
 a36167a <=( a36166a  and  a36161a );
 a36171a <=( (not A233)  and  A232 );
 a36172a <=( (not A203)  and  a36171a );
 a36175a <=( A235  and  A234 );
 a36178a <=( A299  and  A298 );
 a36179a <=( a36178a  and  a36175a );
 a36180a <=( a36179a  and  a36172a );
 a36184a <=( A167  and  A169 );
 a36185a <=( (not A170)  and  a36184a );
 a36189a <=( (not A202)  and  (not A200) );
 a36190a <=( A166  and  a36189a );
 a36191a <=( a36190a  and  a36185a );
 a36195a <=( (not A233)  and  A232 );
 a36196a <=( (not A203)  and  a36195a );
 a36199a <=( A235  and  A234 );
 a36202a <=( (not A299)  and  (not A298) );
 a36203a <=( a36202a  and  a36199a );
 a36204a <=( a36203a  and  a36196a );
 a36208a <=( A167  and  A169 );
 a36209a <=( (not A170)  and  a36208a );
 a36213a <=( (not A202)  and  (not A200) );
 a36214a <=( A166  and  a36213a );
 a36215a <=( a36214a  and  a36209a );
 a36219a <=( (not A233)  and  A232 );
 a36220a <=( (not A203)  and  a36219a );
 a36223a <=( A235  and  A234 );
 a36226a <=( A266  and  (not A265) );
 a36227a <=( a36226a  and  a36223a );
 a36228a <=( a36227a  and  a36220a );
 a36232a <=( A167  and  A169 );
 a36233a <=( (not A170)  and  a36232a );
 a36237a <=( (not A202)  and  (not A200) );
 a36238a <=( A166  and  a36237a );
 a36239a <=( a36238a  and  a36233a );
 a36243a <=( (not A233)  and  A232 );
 a36244a <=( (not A203)  and  a36243a );
 a36247a <=( A236  and  A234 );
 a36250a <=( (not A300)  and  A298 );
 a36251a <=( a36250a  and  a36247a );
 a36252a <=( a36251a  and  a36244a );
 a36256a <=( A167  and  A169 );
 a36257a <=( (not A170)  and  a36256a );
 a36261a <=( (not A202)  and  (not A200) );
 a36262a <=( A166  and  a36261a );
 a36263a <=( a36262a  and  a36257a );
 a36267a <=( (not A233)  and  A232 );
 a36268a <=( (not A203)  and  a36267a );
 a36271a <=( A236  and  A234 );
 a36274a <=( A299  and  A298 );
 a36275a <=( a36274a  and  a36271a );
 a36276a <=( a36275a  and  a36268a );
 a36280a <=( A167  and  A169 );
 a36281a <=( (not A170)  and  a36280a );
 a36285a <=( (not A202)  and  (not A200) );
 a36286a <=( A166  and  a36285a );
 a36287a <=( a36286a  and  a36281a );
 a36291a <=( (not A233)  and  A232 );
 a36292a <=( (not A203)  and  a36291a );
 a36295a <=( A236  and  A234 );
 a36298a <=( (not A299)  and  (not A298) );
 a36299a <=( a36298a  and  a36295a );
 a36300a <=( a36299a  and  a36292a );
 a36304a <=( A167  and  A169 );
 a36305a <=( (not A170)  and  a36304a );
 a36309a <=( (not A202)  and  (not A200) );
 a36310a <=( A166  and  a36309a );
 a36311a <=( a36310a  and  a36305a );
 a36315a <=( (not A233)  and  A232 );
 a36316a <=( (not A203)  and  a36315a );
 a36319a <=( A236  and  A234 );
 a36322a <=( A266  and  (not A265) );
 a36323a <=( a36322a  and  a36319a );
 a36324a <=( a36323a  and  a36316a );
 a36328a <=( A167  and  A169 );
 a36329a <=( (not A170)  and  a36328a );
 a36333a <=( (not A202)  and  (not A200) );
 a36334a <=( A166  and  a36333a );
 a36335a <=( a36334a  and  a36329a );
 a36339a <=( (not A233)  and  (not A232) );
 a36340a <=( (not A203)  and  a36339a );
 a36343a <=( A266  and  A265 );
 a36346a <=( A299  and  (not A298) );
 a36347a <=( a36346a  and  a36343a );
 a36348a <=( a36347a  and  a36340a );
 a36352a <=( A167  and  A169 );
 a36353a <=( (not A170)  and  a36352a );
 a36357a <=( (not A202)  and  (not A200) );
 a36358a <=( A166  and  a36357a );
 a36359a <=( a36358a  and  a36353a );
 a36363a <=( (not A233)  and  (not A232) );
 a36364a <=( (not A203)  and  a36363a );
 a36367a <=( (not A267)  and  (not A266) );
 a36370a <=( A299  and  (not A298) );
 a36371a <=( a36370a  and  a36367a );
 a36372a <=( a36371a  and  a36364a );
 a36376a <=( A167  and  A169 );
 a36377a <=( (not A170)  and  a36376a );
 a36381a <=( (not A202)  and  (not A200) );
 a36382a <=( A166  and  a36381a );
 a36383a <=( a36382a  and  a36377a );
 a36387a <=( (not A233)  and  (not A232) );
 a36388a <=( (not A203)  and  a36387a );
 a36391a <=( (not A266)  and  (not A265) );
 a36394a <=( A299  and  (not A298) );
 a36395a <=( a36394a  and  a36391a );
 a36396a <=( a36395a  and  a36388a );
 a36400a <=( A167  and  A169 );
 a36401a <=( (not A170)  and  a36400a );
 a36405a <=( (not A201)  and  (not A200) );
 a36406a <=( A166  and  a36405a );
 a36407a <=( a36406a  and  a36401a );
 a36411a <=( A265  and  A233 );
 a36412a <=( A232  and  a36411a );
 a36415a <=( (not A269)  and  (not A268) );
 a36418a <=( A299  and  (not A298) );
 a36419a <=( a36418a  and  a36415a );
 a36420a <=( a36419a  and  a36412a );
 a36424a <=( A167  and  A169 );
 a36425a <=( (not A170)  and  a36424a );
 a36429a <=( (not A201)  and  (not A200) );
 a36430a <=( A166  and  a36429a );
 a36431a <=( a36430a  and  a36425a );
 a36435a <=( (not A236)  and  (not A235) );
 a36436a <=( (not A233)  and  a36435a );
 a36439a <=( A266  and  A265 );
 a36442a <=( A299  and  (not A298) );
 a36443a <=( a36442a  and  a36439a );
 a36444a <=( a36443a  and  a36436a );
 a36448a <=( A167  and  A169 );
 a36449a <=( (not A170)  and  a36448a );
 a36453a <=( (not A201)  and  (not A200) );
 a36454a <=( A166  and  a36453a );
 a36455a <=( a36454a  and  a36449a );
 a36459a <=( (not A236)  and  (not A235) );
 a36460a <=( (not A233)  and  a36459a );
 a36463a <=( (not A267)  and  (not A266) );
 a36466a <=( A299  and  (not A298) );
 a36467a <=( a36466a  and  a36463a );
 a36468a <=( a36467a  and  a36460a );
 a36472a <=( A167  and  A169 );
 a36473a <=( (not A170)  and  a36472a );
 a36477a <=( (not A201)  and  (not A200) );
 a36478a <=( A166  and  a36477a );
 a36479a <=( a36478a  and  a36473a );
 a36483a <=( (not A236)  and  (not A235) );
 a36484a <=( (not A233)  and  a36483a );
 a36487a <=( (not A266)  and  (not A265) );
 a36490a <=( A299  and  (not A298) );
 a36491a <=( a36490a  and  a36487a );
 a36492a <=( a36491a  and  a36484a );
 a36496a <=( A167  and  A169 );
 a36497a <=( (not A170)  and  a36496a );
 a36501a <=( (not A201)  and  (not A200) );
 a36502a <=( A166  and  a36501a );
 a36503a <=( a36502a  and  a36497a );
 a36507a <=( (not A266)  and  (not A234) );
 a36508a <=( (not A233)  and  a36507a );
 a36511a <=( (not A269)  and  (not A268) );
 a36514a <=( A299  and  (not A298) );
 a36515a <=( a36514a  and  a36511a );
 a36516a <=( a36515a  and  a36508a );
 a36520a <=( A167  and  A169 );
 a36521a <=( (not A170)  and  a36520a );
 a36525a <=( (not A201)  and  (not A200) );
 a36526a <=( A166  and  a36525a );
 a36527a <=( a36526a  and  a36521a );
 a36531a <=( A234  and  (not A233) );
 a36532a <=( A232  and  a36531a );
 a36535a <=( A298  and  A235 );
 a36538a <=( (not A302)  and  (not A301) );
 a36539a <=( a36538a  and  a36535a );
 a36540a <=( a36539a  and  a36532a );
 a36544a <=( A167  and  A169 );
 a36545a <=( (not A170)  and  a36544a );
 a36549a <=( (not A201)  and  (not A200) );
 a36550a <=( A166  and  a36549a );
 a36551a <=( a36550a  and  a36545a );
 a36555a <=( A234  and  (not A233) );
 a36556a <=( A232  and  a36555a );
 a36559a <=( A298  and  A236 );
 a36562a <=( (not A302)  and  (not A301) );
 a36563a <=( a36562a  and  a36559a );
 a36564a <=( a36563a  and  a36556a );
 a36568a <=( A167  and  A169 );
 a36569a <=( (not A170)  and  a36568a );
 a36573a <=( (not A201)  and  (not A200) );
 a36574a <=( A166  and  a36573a );
 a36575a <=( a36574a  and  a36569a );
 a36579a <=( (not A266)  and  (not A233) );
 a36580a <=( (not A232)  and  a36579a );
 a36583a <=( (not A269)  and  (not A268) );
 a36586a <=( A299  and  (not A298) );
 a36587a <=( a36586a  and  a36583a );
 a36588a <=( a36587a  and  a36580a );
 a36592a <=( A167  and  A169 );
 a36593a <=( (not A170)  and  a36592a );
 a36597a <=( (not A200)  and  (not A199) );
 a36598a <=( A166  and  a36597a );
 a36599a <=( a36598a  and  a36593a );
 a36603a <=( A265  and  A233 );
 a36604a <=( A232  and  a36603a );
 a36607a <=( (not A269)  and  (not A268) );
 a36610a <=( A299  and  (not A298) );
 a36611a <=( a36610a  and  a36607a );
 a36612a <=( a36611a  and  a36604a );
 a36616a <=( A167  and  A169 );
 a36617a <=( (not A170)  and  a36616a );
 a36621a <=( (not A200)  and  (not A199) );
 a36622a <=( A166  and  a36621a );
 a36623a <=( a36622a  and  a36617a );
 a36627a <=( (not A236)  and  (not A235) );
 a36628a <=( (not A233)  and  a36627a );
 a36631a <=( A266  and  A265 );
 a36634a <=( A299  and  (not A298) );
 a36635a <=( a36634a  and  a36631a );
 a36636a <=( a36635a  and  a36628a );
 a36640a <=( A167  and  A169 );
 a36641a <=( (not A170)  and  a36640a );
 a36645a <=( (not A200)  and  (not A199) );
 a36646a <=( A166  and  a36645a );
 a36647a <=( a36646a  and  a36641a );
 a36651a <=( (not A236)  and  (not A235) );
 a36652a <=( (not A233)  and  a36651a );
 a36655a <=( (not A267)  and  (not A266) );
 a36658a <=( A299  and  (not A298) );
 a36659a <=( a36658a  and  a36655a );
 a36660a <=( a36659a  and  a36652a );
 a36664a <=( A167  and  A169 );
 a36665a <=( (not A170)  and  a36664a );
 a36669a <=( (not A200)  and  (not A199) );
 a36670a <=( A166  and  a36669a );
 a36671a <=( a36670a  and  a36665a );
 a36675a <=( (not A236)  and  (not A235) );
 a36676a <=( (not A233)  and  a36675a );
 a36679a <=( (not A266)  and  (not A265) );
 a36682a <=( A299  and  (not A298) );
 a36683a <=( a36682a  and  a36679a );
 a36684a <=( a36683a  and  a36676a );
 a36688a <=( A167  and  A169 );
 a36689a <=( (not A170)  and  a36688a );
 a36693a <=( (not A200)  and  (not A199) );
 a36694a <=( A166  and  a36693a );
 a36695a <=( a36694a  and  a36689a );
 a36699a <=( (not A266)  and  (not A234) );
 a36700a <=( (not A233)  and  a36699a );
 a36703a <=( (not A269)  and  (not A268) );
 a36706a <=( A299  and  (not A298) );
 a36707a <=( a36706a  and  a36703a );
 a36708a <=( a36707a  and  a36700a );
 a36712a <=( A167  and  A169 );
 a36713a <=( (not A170)  and  a36712a );
 a36717a <=( (not A200)  and  (not A199) );
 a36718a <=( A166  and  a36717a );
 a36719a <=( a36718a  and  a36713a );
 a36723a <=( A234  and  (not A233) );
 a36724a <=( A232  and  a36723a );
 a36727a <=( A298  and  A235 );
 a36730a <=( (not A302)  and  (not A301) );
 a36731a <=( a36730a  and  a36727a );
 a36732a <=( a36731a  and  a36724a );
 a36736a <=( A167  and  A169 );
 a36737a <=( (not A170)  and  a36736a );
 a36741a <=( (not A200)  and  (not A199) );
 a36742a <=( A166  and  a36741a );
 a36743a <=( a36742a  and  a36737a );
 a36747a <=( A234  and  (not A233) );
 a36748a <=( A232  and  a36747a );
 a36751a <=( A298  and  A236 );
 a36754a <=( (not A302)  and  (not A301) );
 a36755a <=( a36754a  and  a36751a );
 a36756a <=( a36755a  and  a36748a );
 a36760a <=( A167  and  A169 );
 a36761a <=( (not A170)  and  a36760a );
 a36765a <=( (not A200)  and  (not A199) );
 a36766a <=( A166  and  a36765a );
 a36767a <=( a36766a  and  a36761a );
 a36771a <=( (not A266)  and  (not A233) );
 a36772a <=( (not A232)  and  a36771a );
 a36775a <=( (not A269)  and  (not A268) );
 a36778a <=( A299  and  (not A298) );
 a36779a <=( a36778a  and  a36775a );
 a36780a <=( a36779a  and  a36772a );
 a36784a <=( (not A167)  and  A169 );
 a36785a <=( (not A170)  and  a36784a );
 a36789a <=( A200  and  A199 );
 a36790a <=( (not A166)  and  a36789a );
 a36791a <=( a36790a  and  a36785a );
 a36795a <=( A265  and  A233 );
 a36796a <=( A232  and  a36795a );
 a36799a <=( (not A269)  and  (not A268) );
 a36802a <=( A299  and  (not A298) );
 a36803a <=( a36802a  and  a36799a );
 a36804a <=( a36803a  and  a36796a );
 a36808a <=( (not A167)  and  A169 );
 a36809a <=( (not A170)  and  a36808a );
 a36813a <=( A200  and  A199 );
 a36814a <=( (not A166)  and  a36813a );
 a36815a <=( a36814a  and  a36809a );
 a36819a <=( (not A236)  and  (not A235) );
 a36820a <=( (not A233)  and  a36819a );
 a36823a <=( A266  and  A265 );
 a36826a <=( A299  and  (not A298) );
 a36827a <=( a36826a  and  a36823a );
 a36828a <=( a36827a  and  a36820a );
 a36832a <=( (not A167)  and  A169 );
 a36833a <=( (not A170)  and  a36832a );
 a36837a <=( A200  and  A199 );
 a36838a <=( (not A166)  and  a36837a );
 a36839a <=( a36838a  and  a36833a );
 a36843a <=( (not A236)  and  (not A235) );
 a36844a <=( (not A233)  and  a36843a );
 a36847a <=( (not A267)  and  (not A266) );
 a36850a <=( A299  and  (not A298) );
 a36851a <=( a36850a  and  a36847a );
 a36852a <=( a36851a  and  a36844a );
 a36856a <=( (not A167)  and  A169 );
 a36857a <=( (not A170)  and  a36856a );
 a36861a <=( A200  and  A199 );
 a36862a <=( (not A166)  and  a36861a );
 a36863a <=( a36862a  and  a36857a );
 a36867a <=( (not A236)  and  (not A235) );
 a36868a <=( (not A233)  and  a36867a );
 a36871a <=( (not A266)  and  (not A265) );
 a36874a <=( A299  and  (not A298) );
 a36875a <=( a36874a  and  a36871a );
 a36876a <=( a36875a  and  a36868a );
 a36880a <=( (not A167)  and  A169 );
 a36881a <=( (not A170)  and  a36880a );
 a36885a <=( A200  and  A199 );
 a36886a <=( (not A166)  and  a36885a );
 a36887a <=( a36886a  and  a36881a );
 a36891a <=( (not A266)  and  (not A234) );
 a36892a <=( (not A233)  and  a36891a );
 a36895a <=( (not A269)  and  (not A268) );
 a36898a <=( A299  and  (not A298) );
 a36899a <=( a36898a  and  a36895a );
 a36900a <=( a36899a  and  a36892a );
 a36904a <=( (not A167)  and  A169 );
 a36905a <=( (not A170)  and  a36904a );
 a36909a <=( A200  and  A199 );
 a36910a <=( (not A166)  and  a36909a );
 a36911a <=( a36910a  and  a36905a );
 a36915a <=( A234  and  (not A233) );
 a36916a <=( A232  and  a36915a );
 a36919a <=( A298  and  A235 );
 a36922a <=( (not A302)  and  (not A301) );
 a36923a <=( a36922a  and  a36919a );
 a36924a <=( a36923a  and  a36916a );
 a36928a <=( (not A167)  and  A169 );
 a36929a <=( (not A170)  and  a36928a );
 a36933a <=( A200  and  A199 );
 a36934a <=( (not A166)  and  a36933a );
 a36935a <=( a36934a  and  a36929a );
 a36939a <=( A234  and  (not A233) );
 a36940a <=( A232  and  a36939a );
 a36943a <=( A298  and  A236 );
 a36946a <=( (not A302)  and  (not A301) );
 a36947a <=( a36946a  and  a36943a );
 a36948a <=( a36947a  and  a36940a );
 a36952a <=( (not A167)  and  A169 );
 a36953a <=( (not A170)  and  a36952a );
 a36957a <=( A200  and  A199 );
 a36958a <=( (not A166)  and  a36957a );
 a36959a <=( a36958a  and  a36953a );
 a36963a <=( (not A266)  and  (not A233) );
 a36964a <=( (not A232)  and  a36963a );
 a36967a <=( (not A269)  and  (not A268) );
 a36970a <=( A299  and  (not A298) );
 a36971a <=( a36970a  and  a36967a );
 a36972a <=( a36971a  and  a36964a );
 a36976a <=( (not A167)  and  A169 );
 a36977a <=( (not A170)  and  a36976a );
 a36981a <=( (not A202)  and  (not A200) );
 a36982a <=( (not A166)  and  a36981a );
 a36983a <=( a36982a  and  a36977a );
 a36987a <=( A233  and  A232 );
 a36988a <=( (not A203)  and  a36987a );
 a36991a <=( (not A267)  and  A265 );
 a36994a <=( A299  and  (not A298) );
 a36995a <=( a36994a  and  a36991a );
 a36996a <=( a36995a  and  a36988a );
 a37000a <=( (not A167)  and  A169 );
 a37001a <=( (not A170)  and  a37000a );
 a37005a <=( (not A202)  and  (not A200) );
 a37006a <=( (not A166)  and  a37005a );
 a37007a <=( a37006a  and  a37001a );
 a37011a <=( A233  and  A232 );
 a37012a <=( (not A203)  and  a37011a );
 a37015a <=( A266  and  A265 );
 a37018a <=( A299  and  (not A298) );
 a37019a <=( a37018a  and  a37015a );
 a37020a <=( a37019a  and  a37012a );
 a37024a <=( (not A167)  and  A169 );
 a37025a <=( (not A170)  and  a37024a );
 a37029a <=( (not A202)  and  (not A200) );
 a37030a <=( (not A166)  and  a37029a );
 a37031a <=( a37030a  and  a37025a );
 a37035a <=( A233  and  A232 );
 a37036a <=( (not A203)  and  a37035a );
 a37039a <=( (not A266)  and  (not A265) );
 a37042a <=( A299  and  (not A298) );
 a37043a <=( a37042a  and  a37039a );
 a37044a <=( a37043a  and  a37036a );
 a37048a <=( (not A167)  and  A169 );
 a37049a <=( (not A170)  and  a37048a );
 a37053a <=( (not A202)  and  (not A200) );
 a37054a <=( (not A166)  and  a37053a );
 a37055a <=( a37054a  and  a37049a );
 a37059a <=( A233  and  (not A232) );
 a37060a <=( (not A203)  and  a37059a );
 a37063a <=( (not A266)  and  A265 );
 a37066a <=( A268  and  A267 );
 a37067a <=( a37066a  and  a37063a );
 a37068a <=( a37067a  and  a37060a );
 a37072a <=( (not A167)  and  A169 );
 a37073a <=( (not A170)  and  a37072a );
 a37077a <=( (not A202)  and  (not A200) );
 a37078a <=( (not A166)  and  a37077a );
 a37079a <=( a37078a  and  a37073a );
 a37083a <=( A233  and  (not A232) );
 a37084a <=( (not A203)  and  a37083a );
 a37087a <=( (not A266)  and  A265 );
 a37090a <=( A269  and  A267 );
 a37091a <=( a37090a  and  a37087a );
 a37092a <=( a37091a  and  a37084a );
 a37096a <=( (not A167)  and  A169 );
 a37097a <=( (not A170)  and  a37096a );
 a37101a <=( (not A202)  and  (not A200) );
 a37102a <=( (not A166)  and  a37101a );
 a37103a <=( a37102a  and  a37097a );
 a37107a <=( (not A234)  and  (not A233) );
 a37108a <=( (not A203)  and  a37107a );
 a37111a <=( A266  and  A265 );
 a37114a <=( A299  and  (not A298) );
 a37115a <=( a37114a  and  a37111a );
 a37116a <=( a37115a  and  a37108a );
 a37120a <=( (not A167)  and  A169 );
 a37121a <=( (not A170)  and  a37120a );
 a37125a <=( (not A202)  and  (not A200) );
 a37126a <=( (not A166)  and  a37125a );
 a37127a <=( a37126a  and  a37121a );
 a37131a <=( (not A234)  and  (not A233) );
 a37132a <=( (not A203)  and  a37131a );
 a37135a <=( (not A267)  and  (not A266) );
 a37138a <=( A299  and  (not A298) );
 a37139a <=( a37138a  and  a37135a );
 a37140a <=( a37139a  and  a37132a );
 a37144a <=( (not A167)  and  A169 );
 a37145a <=( (not A170)  and  a37144a );
 a37149a <=( (not A202)  and  (not A200) );
 a37150a <=( (not A166)  and  a37149a );
 a37151a <=( a37150a  and  a37145a );
 a37155a <=( (not A234)  and  (not A233) );
 a37156a <=( (not A203)  and  a37155a );
 a37159a <=( (not A266)  and  (not A265) );
 a37162a <=( A299  and  (not A298) );
 a37163a <=( a37162a  and  a37159a );
 a37164a <=( a37163a  and  a37156a );
 a37168a <=( (not A167)  and  A169 );
 a37169a <=( (not A170)  and  a37168a );
 a37173a <=( (not A202)  and  (not A200) );
 a37174a <=( (not A166)  and  a37173a );
 a37175a <=( a37174a  and  a37169a );
 a37179a <=( (not A233)  and  A232 );
 a37180a <=( (not A203)  and  a37179a );
 a37183a <=( A235  and  A234 );
 a37186a <=( (not A300)  and  A298 );
 a37187a <=( a37186a  and  a37183a );
 a37188a <=( a37187a  and  a37180a );
 a37192a <=( (not A167)  and  A169 );
 a37193a <=( (not A170)  and  a37192a );
 a37197a <=( (not A202)  and  (not A200) );
 a37198a <=( (not A166)  and  a37197a );
 a37199a <=( a37198a  and  a37193a );
 a37203a <=( (not A233)  and  A232 );
 a37204a <=( (not A203)  and  a37203a );
 a37207a <=( A235  and  A234 );
 a37210a <=( A299  and  A298 );
 a37211a <=( a37210a  and  a37207a );
 a37212a <=( a37211a  and  a37204a );
 a37216a <=( (not A167)  and  A169 );
 a37217a <=( (not A170)  and  a37216a );
 a37221a <=( (not A202)  and  (not A200) );
 a37222a <=( (not A166)  and  a37221a );
 a37223a <=( a37222a  and  a37217a );
 a37227a <=( (not A233)  and  A232 );
 a37228a <=( (not A203)  and  a37227a );
 a37231a <=( A235  and  A234 );
 a37234a <=( (not A299)  and  (not A298) );
 a37235a <=( a37234a  and  a37231a );
 a37236a <=( a37235a  and  a37228a );
 a37240a <=( (not A167)  and  A169 );
 a37241a <=( (not A170)  and  a37240a );
 a37245a <=( (not A202)  and  (not A200) );
 a37246a <=( (not A166)  and  a37245a );
 a37247a <=( a37246a  and  a37241a );
 a37251a <=( (not A233)  and  A232 );
 a37252a <=( (not A203)  and  a37251a );
 a37255a <=( A235  and  A234 );
 a37258a <=( A266  and  (not A265) );
 a37259a <=( a37258a  and  a37255a );
 a37260a <=( a37259a  and  a37252a );
 a37264a <=( (not A167)  and  A169 );
 a37265a <=( (not A170)  and  a37264a );
 a37269a <=( (not A202)  and  (not A200) );
 a37270a <=( (not A166)  and  a37269a );
 a37271a <=( a37270a  and  a37265a );
 a37275a <=( (not A233)  and  A232 );
 a37276a <=( (not A203)  and  a37275a );
 a37279a <=( A236  and  A234 );
 a37282a <=( (not A300)  and  A298 );
 a37283a <=( a37282a  and  a37279a );
 a37284a <=( a37283a  and  a37276a );
 a37288a <=( (not A167)  and  A169 );
 a37289a <=( (not A170)  and  a37288a );
 a37293a <=( (not A202)  and  (not A200) );
 a37294a <=( (not A166)  and  a37293a );
 a37295a <=( a37294a  and  a37289a );
 a37299a <=( (not A233)  and  A232 );
 a37300a <=( (not A203)  and  a37299a );
 a37303a <=( A236  and  A234 );
 a37306a <=( A299  and  A298 );
 a37307a <=( a37306a  and  a37303a );
 a37308a <=( a37307a  and  a37300a );
 a37312a <=( (not A167)  and  A169 );
 a37313a <=( (not A170)  and  a37312a );
 a37317a <=( (not A202)  and  (not A200) );
 a37318a <=( (not A166)  and  a37317a );
 a37319a <=( a37318a  and  a37313a );
 a37323a <=( (not A233)  and  A232 );
 a37324a <=( (not A203)  and  a37323a );
 a37327a <=( A236  and  A234 );
 a37330a <=( (not A299)  and  (not A298) );
 a37331a <=( a37330a  and  a37327a );
 a37332a <=( a37331a  and  a37324a );
 a37336a <=( (not A167)  and  A169 );
 a37337a <=( (not A170)  and  a37336a );
 a37341a <=( (not A202)  and  (not A200) );
 a37342a <=( (not A166)  and  a37341a );
 a37343a <=( a37342a  and  a37337a );
 a37347a <=( (not A233)  and  A232 );
 a37348a <=( (not A203)  and  a37347a );
 a37351a <=( A236  and  A234 );
 a37354a <=( A266  and  (not A265) );
 a37355a <=( a37354a  and  a37351a );
 a37356a <=( a37355a  and  a37348a );
 a37360a <=( (not A167)  and  A169 );
 a37361a <=( (not A170)  and  a37360a );
 a37365a <=( (not A202)  and  (not A200) );
 a37366a <=( (not A166)  and  a37365a );
 a37367a <=( a37366a  and  a37361a );
 a37371a <=( (not A233)  and  (not A232) );
 a37372a <=( (not A203)  and  a37371a );
 a37375a <=( A266  and  A265 );
 a37378a <=( A299  and  (not A298) );
 a37379a <=( a37378a  and  a37375a );
 a37380a <=( a37379a  and  a37372a );
 a37384a <=( (not A167)  and  A169 );
 a37385a <=( (not A170)  and  a37384a );
 a37389a <=( (not A202)  and  (not A200) );
 a37390a <=( (not A166)  and  a37389a );
 a37391a <=( a37390a  and  a37385a );
 a37395a <=( (not A233)  and  (not A232) );
 a37396a <=( (not A203)  and  a37395a );
 a37399a <=( (not A267)  and  (not A266) );
 a37402a <=( A299  and  (not A298) );
 a37403a <=( a37402a  and  a37399a );
 a37404a <=( a37403a  and  a37396a );
 a37408a <=( (not A167)  and  A169 );
 a37409a <=( (not A170)  and  a37408a );
 a37413a <=( (not A202)  and  (not A200) );
 a37414a <=( (not A166)  and  a37413a );
 a37415a <=( a37414a  and  a37409a );
 a37419a <=( (not A233)  and  (not A232) );
 a37420a <=( (not A203)  and  a37419a );
 a37423a <=( (not A266)  and  (not A265) );
 a37426a <=( A299  and  (not A298) );
 a37427a <=( a37426a  and  a37423a );
 a37428a <=( a37427a  and  a37420a );
 a37432a <=( (not A167)  and  A169 );
 a37433a <=( (not A170)  and  a37432a );
 a37437a <=( (not A201)  and  (not A200) );
 a37438a <=( (not A166)  and  a37437a );
 a37439a <=( a37438a  and  a37433a );
 a37443a <=( A265  and  A233 );
 a37444a <=( A232  and  a37443a );
 a37447a <=( (not A269)  and  (not A268) );
 a37450a <=( A299  and  (not A298) );
 a37451a <=( a37450a  and  a37447a );
 a37452a <=( a37451a  and  a37444a );
 a37456a <=( (not A167)  and  A169 );
 a37457a <=( (not A170)  and  a37456a );
 a37461a <=( (not A201)  and  (not A200) );
 a37462a <=( (not A166)  and  a37461a );
 a37463a <=( a37462a  and  a37457a );
 a37467a <=( (not A236)  and  (not A235) );
 a37468a <=( (not A233)  and  a37467a );
 a37471a <=( A266  and  A265 );
 a37474a <=( A299  and  (not A298) );
 a37475a <=( a37474a  and  a37471a );
 a37476a <=( a37475a  and  a37468a );
 a37480a <=( (not A167)  and  A169 );
 a37481a <=( (not A170)  and  a37480a );
 a37485a <=( (not A201)  and  (not A200) );
 a37486a <=( (not A166)  and  a37485a );
 a37487a <=( a37486a  and  a37481a );
 a37491a <=( (not A236)  and  (not A235) );
 a37492a <=( (not A233)  and  a37491a );
 a37495a <=( (not A267)  and  (not A266) );
 a37498a <=( A299  and  (not A298) );
 a37499a <=( a37498a  and  a37495a );
 a37500a <=( a37499a  and  a37492a );
 a37504a <=( (not A167)  and  A169 );
 a37505a <=( (not A170)  and  a37504a );
 a37509a <=( (not A201)  and  (not A200) );
 a37510a <=( (not A166)  and  a37509a );
 a37511a <=( a37510a  and  a37505a );
 a37515a <=( (not A236)  and  (not A235) );
 a37516a <=( (not A233)  and  a37515a );
 a37519a <=( (not A266)  and  (not A265) );
 a37522a <=( A299  and  (not A298) );
 a37523a <=( a37522a  and  a37519a );
 a37524a <=( a37523a  and  a37516a );
 a37528a <=( (not A167)  and  A169 );
 a37529a <=( (not A170)  and  a37528a );
 a37533a <=( (not A201)  and  (not A200) );
 a37534a <=( (not A166)  and  a37533a );
 a37535a <=( a37534a  and  a37529a );
 a37539a <=( (not A266)  and  (not A234) );
 a37540a <=( (not A233)  and  a37539a );
 a37543a <=( (not A269)  and  (not A268) );
 a37546a <=( A299  and  (not A298) );
 a37547a <=( a37546a  and  a37543a );
 a37548a <=( a37547a  and  a37540a );
 a37552a <=( (not A167)  and  A169 );
 a37553a <=( (not A170)  and  a37552a );
 a37557a <=( (not A201)  and  (not A200) );
 a37558a <=( (not A166)  and  a37557a );
 a37559a <=( a37558a  and  a37553a );
 a37563a <=( A234  and  (not A233) );
 a37564a <=( A232  and  a37563a );
 a37567a <=( A298  and  A235 );
 a37570a <=( (not A302)  and  (not A301) );
 a37571a <=( a37570a  and  a37567a );
 a37572a <=( a37571a  and  a37564a );
 a37576a <=( (not A167)  and  A169 );
 a37577a <=( (not A170)  and  a37576a );
 a37581a <=( (not A201)  and  (not A200) );
 a37582a <=( (not A166)  and  a37581a );
 a37583a <=( a37582a  and  a37577a );
 a37587a <=( A234  and  (not A233) );
 a37588a <=( A232  and  a37587a );
 a37591a <=( A298  and  A236 );
 a37594a <=( (not A302)  and  (not A301) );
 a37595a <=( a37594a  and  a37591a );
 a37596a <=( a37595a  and  a37588a );
 a37600a <=( (not A167)  and  A169 );
 a37601a <=( (not A170)  and  a37600a );
 a37605a <=( (not A201)  and  (not A200) );
 a37606a <=( (not A166)  and  a37605a );
 a37607a <=( a37606a  and  a37601a );
 a37611a <=( (not A266)  and  (not A233) );
 a37612a <=( (not A232)  and  a37611a );
 a37615a <=( (not A269)  and  (not A268) );
 a37618a <=( A299  and  (not A298) );
 a37619a <=( a37618a  and  a37615a );
 a37620a <=( a37619a  and  a37612a );
 a37624a <=( (not A167)  and  A169 );
 a37625a <=( (not A170)  and  a37624a );
 a37629a <=( (not A200)  and  (not A199) );
 a37630a <=( (not A166)  and  a37629a );
 a37631a <=( a37630a  and  a37625a );
 a37635a <=( A265  and  A233 );
 a37636a <=( A232  and  a37635a );
 a37639a <=( (not A269)  and  (not A268) );
 a37642a <=( A299  and  (not A298) );
 a37643a <=( a37642a  and  a37639a );
 a37644a <=( a37643a  and  a37636a );
 a37648a <=( (not A167)  and  A169 );
 a37649a <=( (not A170)  and  a37648a );
 a37653a <=( (not A200)  and  (not A199) );
 a37654a <=( (not A166)  and  a37653a );
 a37655a <=( a37654a  and  a37649a );
 a37659a <=( (not A236)  and  (not A235) );
 a37660a <=( (not A233)  and  a37659a );
 a37663a <=( A266  and  A265 );
 a37666a <=( A299  and  (not A298) );
 a37667a <=( a37666a  and  a37663a );
 a37668a <=( a37667a  and  a37660a );
 a37672a <=( (not A167)  and  A169 );
 a37673a <=( (not A170)  and  a37672a );
 a37677a <=( (not A200)  and  (not A199) );
 a37678a <=( (not A166)  and  a37677a );
 a37679a <=( a37678a  and  a37673a );
 a37683a <=( (not A236)  and  (not A235) );
 a37684a <=( (not A233)  and  a37683a );
 a37687a <=( (not A267)  and  (not A266) );
 a37690a <=( A299  and  (not A298) );
 a37691a <=( a37690a  and  a37687a );
 a37692a <=( a37691a  and  a37684a );
 a37696a <=( (not A167)  and  A169 );
 a37697a <=( (not A170)  and  a37696a );
 a37701a <=( (not A200)  and  (not A199) );
 a37702a <=( (not A166)  and  a37701a );
 a37703a <=( a37702a  and  a37697a );
 a37707a <=( (not A236)  and  (not A235) );
 a37708a <=( (not A233)  and  a37707a );
 a37711a <=( (not A266)  and  (not A265) );
 a37714a <=( A299  and  (not A298) );
 a37715a <=( a37714a  and  a37711a );
 a37716a <=( a37715a  and  a37708a );
 a37720a <=( (not A167)  and  A169 );
 a37721a <=( (not A170)  and  a37720a );
 a37725a <=( (not A200)  and  (not A199) );
 a37726a <=( (not A166)  and  a37725a );
 a37727a <=( a37726a  and  a37721a );
 a37731a <=( (not A266)  and  (not A234) );
 a37732a <=( (not A233)  and  a37731a );
 a37735a <=( (not A269)  and  (not A268) );
 a37738a <=( A299  and  (not A298) );
 a37739a <=( a37738a  and  a37735a );
 a37740a <=( a37739a  and  a37732a );
 a37744a <=( (not A167)  and  A169 );
 a37745a <=( (not A170)  and  a37744a );
 a37749a <=( (not A200)  and  (not A199) );
 a37750a <=( (not A166)  and  a37749a );
 a37751a <=( a37750a  and  a37745a );
 a37755a <=( A234  and  (not A233) );
 a37756a <=( A232  and  a37755a );
 a37759a <=( A298  and  A235 );
 a37762a <=( (not A302)  and  (not A301) );
 a37763a <=( a37762a  and  a37759a );
 a37764a <=( a37763a  and  a37756a );
 a37768a <=( (not A167)  and  A169 );
 a37769a <=( (not A170)  and  a37768a );
 a37773a <=( (not A200)  and  (not A199) );
 a37774a <=( (not A166)  and  a37773a );
 a37775a <=( a37774a  and  a37769a );
 a37779a <=( A234  and  (not A233) );
 a37780a <=( A232  and  a37779a );
 a37783a <=( A298  and  A236 );
 a37786a <=( (not A302)  and  (not A301) );
 a37787a <=( a37786a  and  a37783a );
 a37788a <=( a37787a  and  a37780a );
 a37792a <=( (not A167)  and  A169 );
 a37793a <=( (not A170)  and  a37792a );
 a37797a <=( (not A200)  and  (not A199) );
 a37798a <=( (not A166)  and  a37797a );
 a37799a <=( a37798a  and  a37793a );
 a37803a <=( (not A266)  and  (not A233) );
 a37804a <=( (not A232)  and  a37803a );
 a37807a <=( (not A269)  and  (not A268) );
 a37810a <=( A299  and  (not A298) );
 a37811a <=( a37810a  and  a37807a );
 a37812a <=( a37811a  and  a37804a );
 a37816a <=( (not A166)  and  (not A167) );
 a37817a <=( (not A169)  and  a37816a );
 a37821a <=( A232  and  A200 );
 a37822a <=( (not A199)  and  a37821a );
 a37823a <=( a37822a  and  a37817a );
 a37827a <=( (not A267)  and  A265 );
 a37828a <=( A233  and  a37827a );
 a37831a <=( (not A299)  and  A298 );
 a37834a <=( A301  and  A300 );
 a37835a <=( a37834a  and  a37831a );
 a37836a <=( a37835a  and  a37828a );
 a37840a <=( (not A166)  and  (not A167) );
 a37841a <=( (not A169)  and  a37840a );
 a37845a <=( A232  and  A200 );
 a37846a <=( (not A199)  and  a37845a );
 a37847a <=( a37846a  and  a37841a );
 a37851a <=( (not A267)  and  A265 );
 a37852a <=( A233  and  a37851a );
 a37855a <=( (not A299)  and  A298 );
 a37858a <=( A302  and  A300 );
 a37859a <=( a37858a  and  a37855a );
 a37860a <=( a37859a  and  a37852a );
 a37864a <=( (not A166)  and  (not A167) );
 a37865a <=( (not A169)  and  a37864a );
 a37869a <=( A232  and  A200 );
 a37870a <=( (not A199)  and  a37869a );
 a37871a <=( a37870a  and  a37865a );
 a37875a <=( A266  and  A265 );
 a37876a <=( A233  and  a37875a );
 a37879a <=( (not A299)  and  A298 );
 a37882a <=( A301  and  A300 );
 a37883a <=( a37882a  and  a37879a );
 a37884a <=( a37883a  and  a37876a );
 a37888a <=( (not A166)  and  (not A167) );
 a37889a <=( (not A169)  and  a37888a );
 a37893a <=( A232  and  A200 );
 a37894a <=( (not A199)  and  a37893a );
 a37895a <=( a37894a  and  a37889a );
 a37899a <=( A266  and  A265 );
 a37900a <=( A233  and  a37899a );
 a37903a <=( (not A299)  and  A298 );
 a37906a <=( A302  and  A300 );
 a37907a <=( a37906a  and  a37903a );
 a37908a <=( a37907a  and  a37900a );
 a37912a <=( (not A166)  and  (not A167) );
 a37913a <=( (not A169)  and  a37912a );
 a37917a <=( A232  and  A200 );
 a37918a <=( (not A199)  and  a37917a );
 a37919a <=( a37918a  and  a37913a );
 a37923a <=( (not A266)  and  (not A265) );
 a37924a <=( A233  and  a37923a );
 a37927a <=( (not A299)  and  A298 );
 a37930a <=( A301  and  A300 );
 a37931a <=( a37930a  and  a37927a );
 a37932a <=( a37931a  and  a37924a );
 a37936a <=( (not A166)  and  (not A167) );
 a37937a <=( (not A169)  and  a37936a );
 a37941a <=( A232  and  A200 );
 a37942a <=( (not A199)  and  a37941a );
 a37943a <=( a37942a  and  a37937a );
 a37947a <=( (not A266)  and  (not A265) );
 a37948a <=( A233  and  a37947a );
 a37951a <=( (not A299)  and  A298 );
 a37954a <=( A302  and  A300 );
 a37955a <=( a37954a  and  a37951a );
 a37956a <=( a37955a  and  a37948a );
 a37960a <=( (not A166)  and  (not A167) );
 a37961a <=( (not A169)  and  a37960a );
 a37965a <=( (not A233)  and  A200 );
 a37966a <=( (not A199)  and  a37965a );
 a37967a <=( a37966a  and  a37961a );
 a37971a <=( (not A266)  and  (not A236) );
 a37972a <=( (not A235)  and  a37971a );
 a37975a <=( (not A269)  and  (not A268) );
 a37978a <=( A299  and  (not A298) );
 a37979a <=( a37978a  and  a37975a );
 a37980a <=( a37979a  and  a37972a );
 a37984a <=( (not A166)  and  (not A167) );
 a37985a <=( (not A169)  and  a37984a );
 a37989a <=( (not A233)  and  A200 );
 a37990a <=( (not A199)  and  a37989a );
 a37991a <=( a37990a  and  a37985a );
 a37995a <=( A266  and  A265 );
 a37996a <=( (not A234)  and  a37995a );
 a37999a <=( (not A299)  and  A298 );
 a38002a <=( A301  and  A300 );
 a38003a <=( a38002a  and  a37999a );
 a38004a <=( a38003a  and  a37996a );
 a38008a <=( (not A166)  and  (not A167) );
 a38009a <=( (not A169)  and  a38008a );
 a38013a <=( (not A233)  and  A200 );
 a38014a <=( (not A199)  and  a38013a );
 a38015a <=( a38014a  and  a38009a );
 a38019a <=( A266  and  A265 );
 a38020a <=( (not A234)  and  a38019a );
 a38023a <=( (not A299)  and  A298 );
 a38026a <=( A302  and  A300 );
 a38027a <=( a38026a  and  a38023a );
 a38028a <=( a38027a  and  a38020a );
 a38032a <=( (not A166)  and  (not A167) );
 a38033a <=( (not A169)  and  a38032a );
 a38037a <=( (not A233)  and  A200 );
 a38038a <=( (not A199)  and  a38037a );
 a38039a <=( a38038a  and  a38033a );
 a38043a <=( (not A267)  and  (not A266) );
 a38044a <=( (not A234)  and  a38043a );
 a38047a <=( (not A299)  and  A298 );
 a38050a <=( A301  and  A300 );
 a38051a <=( a38050a  and  a38047a );
 a38052a <=( a38051a  and  a38044a );
 a38056a <=( (not A166)  and  (not A167) );
 a38057a <=( (not A169)  and  a38056a );
 a38061a <=( (not A233)  and  A200 );
 a38062a <=( (not A199)  and  a38061a );
 a38063a <=( a38062a  and  a38057a );
 a38067a <=( (not A267)  and  (not A266) );
 a38068a <=( (not A234)  and  a38067a );
 a38071a <=( (not A299)  and  A298 );
 a38074a <=( A302  and  A300 );
 a38075a <=( a38074a  and  a38071a );
 a38076a <=( a38075a  and  a38068a );
 a38080a <=( (not A166)  and  (not A167) );
 a38081a <=( (not A169)  and  a38080a );
 a38085a <=( (not A233)  and  A200 );
 a38086a <=( (not A199)  and  a38085a );
 a38087a <=( a38086a  and  a38081a );
 a38091a <=( (not A266)  and  (not A265) );
 a38092a <=( (not A234)  and  a38091a );
 a38095a <=( (not A299)  and  A298 );
 a38098a <=( A301  and  A300 );
 a38099a <=( a38098a  and  a38095a );
 a38100a <=( a38099a  and  a38092a );
 a38104a <=( (not A166)  and  (not A167) );
 a38105a <=( (not A169)  and  a38104a );
 a38109a <=( (not A233)  and  A200 );
 a38110a <=( (not A199)  and  a38109a );
 a38111a <=( a38110a  and  a38105a );
 a38115a <=( (not A266)  and  (not A265) );
 a38116a <=( (not A234)  and  a38115a );
 a38119a <=( (not A299)  and  A298 );
 a38122a <=( A302  and  A300 );
 a38123a <=( a38122a  and  a38119a );
 a38124a <=( a38123a  and  a38116a );
 a38128a <=( (not A166)  and  (not A167) );
 a38129a <=( (not A169)  and  a38128a );
 a38133a <=( A232  and  A200 );
 a38134a <=( (not A199)  and  a38133a );
 a38135a <=( a38134a  and  a38129a );
 a38139a <=( A235  and  A234 );
 a38140a <=( (not A233)  and  a38139a );
 a38143a <=( (not A266)  and  A265 );
 a38146a <=( A268  and  A267 );
 a38147a <=( a38146a  and  a38143a );
 a38148a <=( a38147a  and  a38140a );
 a38152a <=( (not A166)  and  (not A167) );
 a38153a <=( (not A169)  and  a38152a );
 a38157a <=( A232  and  A200 );
 a38158a <=( (not A199)  and  a38157a );
 a38159a <=( a38158a  and  a38153a );
 a38163a <=( A235  and  A234 );
 a38164a <=( (not A233)  and  a38163a );
 a38167a <=( (not A266)  and  A265 );
 a38170a <=( A269  and  A267 );
 a38171a <=( a38170a  and  a38167a );
 a38172a <=( a38171a  and  a38164a );
 a38176a <=( (not A166)  and  (not A167) );
 a38177a <=( (not A169)  and  a38176a );
 a38181a <=( A232  and  A200 );
 a38182a <=( (not A199)  and  a38181a );
 a38183a <=( a38182a  and  a38177a );
 a38187a <=( A236  and  A234 );
 a38188a <=( (not A233)  and  a38187a );
 a38191a <=( (not A266)  and  A265 );
 a38194a <=( A268  and  A267 );
 a38195a <=( a38194a  and  a38191a );
 a38196a <=( a38195a  and  a38188a );
 a38200a <=( (not A166)  and  (not A167) );
 a38201a <=( (not A169)  and  a38200a );
 a38205a <=( A232  and  A200 );
 a38206a <=( (not A199)  and  a38205a );
 a38207a <=( a38206a  and  a38201a );
 a38211a <=( A236  and  A234 );
 a38212a <=( (not A233)  and  a38211a );
 a38215a <=( (not A266)  and  A265 );
 a38218a <=( A269  and  A267 );
 a38219a <=( a38218a  and  a38215a );
 a38220a <=( a38219a  and  a38212a );
 a38224a <=( (not A166)  and  (not A167) );
 a38225a <=( (not A169)  and  a38224a );
 a38229a <=( (not A232)  and  A200 );
 a38230a <=( (not A199)  and  a38229a );
 a38231a <=( a38230a  and  a38225a );
 a38235a <=( A266  and  A265 );
 a38236a <=( (not A233)  and  a38235a );
 a38239a <=( (not A299)  and  A298 );
 a38242a <=( A301  and  A300 );
 a38243a <=( a38242a  and  a38239a );
 a38244a <=( a38243a  and  a38236a );
 a38248a <=( (not A166)  and  (not A167) );
 a38249a <=( (not A169)  and  a38248a );
 a38253a <=( (not A232)  and  A200 );
 a38254a <=( (not A199)  and  a38253a );
 a38255a <=( a38254a  and  a38249a );
 a38259a <=( A266  and  A265 );
 a38260a <=( (not A233)  and  a38259a );
 a38263a <=( (not A299)  and  A298 );
 a38266a <=( A302  and  A300 );
 a38267a <=( a38266a  and  a38263a );
 a38268a <=( a38267a  and  a38260a );
 a38272a <=( (not A166)  and  (not A167) );
 a38273a <=( (not A169)  and  a38272a );
 a38277a <=( (not A232)  and  A200 );
 a38278a <=( (not A199)  and  a38277a );
 a38279a <=( a38278a  and  a38273a );
 a38283a <=( (not A267)  and  (not A266) );
 a38284a <=( (not A233)  and  a38283a );
 a38287a <=( (not A299)  and  A298 );
 a38290a <=( A301  and  A300 );
 a38291a <=( a38290a  and  a38287a );
 a38292a <=( a38291a  and  a38284a );
 a38296a <=( (not A166)  and  (not A167) );
 a38297a <=( (not A169)  and  a38296a );
 a38301a <=( (not A232)  and  A200 );
 a38302a <=( (not A199)  and  a38301a );
 a38303a <=( a38302a  and  a38297a );
 a38307a <=( (not A267)  and  (not A266) );
 a38308a <=( (not A233)  and  a38307a );
 a38311a <=( (not A299)  and  A298 );
 a38314a <=( A302  and  A300 );
 a38315a <=( a38314a  and  a38311a );
 a38316a <=( a38315a  and  a38308a );
 a38320a <=( (not A166)  and  (not A167) );
 a38321a <=( (not A169)  and  a38320a );
 a38325a <=( (not A232)  and  A200 );
 a38326a <=( (not A199)  and  a38325a );
 a38327a <=( a38326a  and  a38321a );
 a38331a <=( (not A266)  and  (not A265) );
 a38332a <=( (not A233)  and  a38331a );
 a38335a <=( (not A299)  and  A298 );
 a38338a <=( A301  and  A300 );
 a38339a <=( a38338a  and  a38335a );
 a38340a <=( a38339a  and  a38332a );
 a38344a <=( (not A166)  and  (not A167) );
 a38345a <=( (not A169)  and  a38344a );
 a38349a <=( (not A232)  and  A200 );
 a38350a <=( (not A199)  and  a38349a );
 a38351a <=( a38350a  and  a38345a );
 a38355a <=( (not A266)  and  (not A265) );
 a38356a <=( (not A233)  and  a38355a );
 a38359a <=( (not A299)  and  A298 );
 a38362a <=( A302  and  A300 );
 a38363a <=( a38362a  and  a38359a );
 a38364a <=( a38363a  and  a38356a );
 a38368a <=( (not A166)  and  (not A167) );
 a38369a <=( (not A169)  and  a38368a );
 a38373a <=( A201  and  (not A200) );
 a38374a <=( A199  and  a38373a );
 a38375a <=( a38374a  and  a38369a );
 a38379a <=( A233  and  A232 );
 a38380a <=( A202  and  a38379a );
 a38383a <=( (not A267)  and  A265 );
 a38386a <=( A299  and  (not A298) );
 a38387a <=( a38386a  and  a38383a );
 a38388a <=( a38387a  and  a38380a );
 a38392a <=( (not A166)  and  (not A167) );
 a38393a <=( (not A169)  and  a38392a );
 a38397a <=( A201  and  (not A200) );
 a38398a <=( A199  and  a38397a );
 a38399a <=( a38398a  and  a38393a );
 a38403a <=( A233  and  A232 );
 a38404a <=( A202  and  a38403a );
 a38407a <=( A266  and  A265 );
 a38410a <=( A299  and  (not A298) );
 a38411a <=( a38410a  and  a38407a );
 a38412a <=( a38411a  and  a38404a );
 a38416a <=( (not A166)  and  (not A167) );
 a38417a <=( (not A169)  and  a38416a );
 a38421a <=( A201  and  (not A200) );
 a38422a <=( A199  and  a38421a );
 a38423a <=( a38422a  and  a38417a );
 a38427a <=( A233  and  A232 );
 a38428a <=( A202  and  a38427a );
 a38431a <=( (not A266)  and  (not A265) );
 a38434a <=( A299  and  (not A298) );
 a38435a <=( a38434a  and  a38431a );
 a38436a <=( a38435a  and  a38428a );
 a38440a <=( (not A166)  and  (not A167) );
 a38441a <=( (not A169)  and  a38440a );
 a38445a <=( A201  and  (not A200) );
 a38446a <=( A199  and  a38445a );
 a38447a <=( a38446a  and  a38441a );
 a38451a <=( A233  and  (not A232) );
 a38452a <=( A202  and  a38451a );
 a38455a <=( (not A266)  and  A265 );
 a38458a <=( A268  and  A267 );
 a38459a <=( a38458a  and  a38455a );
 a38460a <=( a38459a  and  a38452a );
 a38464a <=( (not A166)  and  (not A167) );
 a38465a <=( (not A169)  and  a38464a );
 a38469a <=( A201  and  (not A200) );
 a38470a <=( A199  and  a38469a );
 a38471a <=( a38470a  and  a38465a );
 a38475a <=( A233  and  (not A232) );
 a38476a <=( A202  and  a38475a );
 a38479a <=( (not A266)  and  A265 );
 a38482a <=( A269  and  A267 );
 a38483a <=( a38482a  and  a38479a );
 a38484a <=( a38483a  and  a38476a );
 a38488a <=( (not A166)  and  (not A167) );
 a38489a <=( (not A169)  and  a38488a );
 a38493a <=( A201  and  (not A200) );
 a38494a <=( A199  and  a38493a );
 a38495a <=( a38494a  and  a38489a );
 a38499a <=( (not A234)  and  (not A233) );
 a38500a <=( A202  and  a38499a );
 a38503a <=( A266  and  A265 );
 a38506a <=( A299  and  (not A298) );
 a38507a <=( a38506a  and  a38503a );
 a38508a <=( a38507a  and  a38500a );
 a38512a <=( (not A166)  and  (not A167) );
 a38513a <=( (not A169)  and  a38512a );
 a38517a <=( A201  and  (not A200) );
 a38518a <=( A199  and  a38517a );
 a38519a <=( a38518a  and  a38513a );
 a38523a <=( (not A234)  and  (not A233) );
 a38524a <=( A202  and  a38523a );
 a38527a <=( (not A267)  and  (not A266) );
 a38530a <=( A299  and  (not A298) );
 a38531a <=( a38530a  and  a38527a );
 a38532a <=( a38531a  and  a38524a );
 a38536a <=( (not A166)  and  (not A167) );
 a38537a <=( (not A169)  and  a38536a );
 a38541a <=( A201  and  (not A200) );
 a38542a <=( A199  and  a38541a );
 a38543a <=( a38542a  and  a38537a );
 a38547a <=( (not A234)  and  (not A233) );
 a38548a <=( A202  and  a38547a );
 a38551a <=( (not A266)  and  (not A265) );
 a38554a <=( A299  and  (not A298) );
 a38555a <=( a38554a  and  a38551a );
 a38556a <=( a38555a  and  a38548a );
 a38560a <=( (not A166)  and  (not A167) );
 a38561a <=( (not A169)  and  a38560a );
 a38565a <=( A201  and  (not A200) );
 a38566a <=( A199  and  a38565a );
 a38567a <=( a38566a  and  a38561a );
 a38571a <=( (not A233)  and  A232 );
 a38572a <=( A202  and  a38571a );
 a38575a <=( A235  and  A234 );
 a38578a <=( (not A300)  and  A298 );
 a38579a <=( a38578a  and  a38575a );
 a38580a <=( a38579a  and  a38572a );
 a38584a <=( (not A166)  and  (not A167) );
 a38585a <=( (not A169)  and  a38584a );
 a38589a <=( A201  and  (not A200) );
 a38590a <=( A199  and  a38589a );
 a38591a <=( a38590a  and  a38585a );
 a38595a <=( (not A233)  and  A232 );
 a38596a <=( A202  and  a38595a );
 a38599a <=( A235  and  A234 );
 a38602a <=( A299  and  A298 );
 a38603a <=( a38602a  and  a38599a );
 a38604a <=( a38603a  and  a38596a );
 a38608a <=( (not A166)  and  (not A167) );
 a38609a <=( (not A169)  and  a38608a );
 a38613a <=( A201  and  (not A200) );
 a38614a <=( A199  and  a38613a );
 a38615a <=( a38614a  and  a38609a );
 a38619a <=( (not A233)  and  A232 );
 a38620a <=( A202  and  a38619a );
 a38623a <=( A235  and  A234 );
 a38626a <=( (not A299)  and  (not A298) );
 a38627a <=( a38626a  and  a38623a );
 a38628a <=( a38627a  and  a38620a );
 a38632a <=( (not A166)  and  (not A167) );
 a38633a <=( (not A169)  and  a38632a );
 a38637a <=( A201  and  (not A200) );
 a38638a <=( A199  and  a38637a );
 a38639a <=( a38638a  and  a38633a );
 a38643a <=( (not A233)  and  A232 );
 a38644a <=( A202  and  a38643a );
 a38647a <=( A235  and  A234 );
 a38650a <=( A266  and  (not A265) );
 a38651a <=( a38650a  and  a38647a );
 a38652a <=( a38651a  and  a38644a );
 a38656a <=( (not A166)  and  (not A167) );
 a38657a <=( (not A169)  and  a38656a );
 a38661a <=( A201  and  (not A200) );
 a38662a <=( A199  and  a38661a );
 a38663a <=( a38662a  and  a38657a );
 a38667a <=( (not A233)  and  A232 );
 a38668a <=( A202  and  a38667a );
 a38671a <=( A236  and  A234 );
 a38674a <=( (not A300)  and  A298 );
 a38675a <=( a38674a  and  a38671a );
 a38676a <=( a38675a  and  a38668a );
 a38680a <=( (not A166)  and  (not A167) );
 a38681a <=( (not A169)  and  a38680a );
 a38685a <=( A201  and  (not A200) );
 a38686a <=( A199  and  a38685a );
 a38687a <=( a38686a  and  a38681a );
 a38691a <=( (not A233)  and  A232 );
 a38692a <=( A202  and  a38691a );
 a38695a <=( A236  and  A234 );
 a38698a <=( A299  and  A298 );
 a38699a <=( a38698a  and  a38695a );
 a38700a <=( a38699a  and  a38692a );
 a38704a <=( (not A166)  and  (not A167) );
 a38705a <=( (not A169)  and  a38704a );
 a38709a <=( A201  and  (not A200) );
 a38710a <=( A199  and  a38709a );
 a38711a <=( a38710a  and  a38705a );
 a38715a <=( (not A233)  and  A232 );
 a38716a <=( A202  and  a38715a );
 a38719a <=( A236  and  A234 );
 a38722a <=( (not A299)  and  (not A298) );
 a38723a <=( a38722a  and  a38719a );
 a38724a <=( a38723a  and  a38716a );
 a38728a <=( (not A166)  and  (not A167) );
 a38729a <=( (not A169)  and  a38728a );
 a38733a <=( A201  and  (not A200) );
 a38734a <=( A199  and  a38733a );
 a38735a <=( a38734a  and  a38729a );
 a38739a <=( (not A233)  and  A232 );
 a38740a <=( A202  and  a38739a );
 a38743a <=( A236  and  A234 );
 a38746a <=( A266  and  (not A265) );
 a38747a <=( a38746a  and  a38743a );
 a38748a <=( a38747a  and  a38740a );
 a38752a <=( (not A166)  and  (not A167) );
 a38753a <=( (not A169)  and  a38752a );
 a38757a <=( A201  and  (not A200) );
 a38758a <=( A199  and  a38757a );
 a38759a <=( a38758a  and  a38753a );
 a38763a <=( (not A233)  and  (not A232) );
 a38764a <=( A202  and  a38763a );
 a38767a <=( A266  and  A265 );
 a38770a <=( A299  and  (not A298) );
 a38771a <=( a38770a  and  a38767a );
 a38772a <=( a38771a  and  a38764a );
 a38776a <=( (not A166)  and  (not A167) );
 a38777a <=( (not A169)  and  a38776a );
 a38781a <=( A201  and  (not A200) );
 a38782a <=( A199  and  a38781a );
 a38783a <=( a38782a  and  a38777a );
 a38787a <=( (not A233)  and  (not A232) );
 a38788a <=( A202  and  a38787a );
 a38791a <=( (not A267)  and  (not A266) );
 a38794a <=( A299  and  (not A298) );
 a38795a <=( a38794a  and  a38791a );
 a38796a <=( a38795a  and  a38788a );
 a38800a <=( (not A166)  and  (not A167) );
 a38801a <=( (not A169)  and  a38800a );
 a38805a <=( A201  and  (not A200) );
 a38806a <=( A199  and  a38805a );
 a38807a <=( a38806a  and  a38801a );
 a38811a <=( (not A233)  and  (not A232) );
 a38812a <=( A202  and  a38811a );
 a38815a <=( (not A266)  and  (not A265) );
 a38818a <=( A299  and  (not A298) );
 a38819a <=( a38818a  and  a38815a );
 a38820a <=( a38819a  and  a38812a );
 a38824a <=( (not A166)  and  (not A167) );
 a38825a <=( (not A169)  and  a38824a );
 a38829a <=( A201  and  (not A200) );
 a38830a <=( A199  and  a38829a );
 a38831a <=( a38830a  and  a38825a );
 a38835a <=( A233  and  A232 );
 a38836a <=( A203  and  a38835a );
 a38839a <=( (not A267)  and  A265 );
 a38842a <=( A299  and  (not A298) );
 a38843a <=( a38842a  and  a38839a );
 a38844a <=( a38843a  and  a38836a );
 a38848a <=( (not A166)  and  (not A167) );
 a38849a <=( (not A169)  and  a38848a );
 a38853a <=( A201  and  (not A200) );
 a38854a <=( A199  and  a38853a );
 a38855a <=( a38854a  and  a38849a );
 a38859a <=( A233  and  A232 );
 a38860a <=( A203  and  a38859a );
 a38863a <=( A266  and  A265 );
 a38866a <=( A299  and  (not A298) );
 a38867a <=( a38866a  and  a38863a );
 a38868a <=( a38867a  and  a38860a );
 a38872a <=( (not A166)  and  (not A167) );
 a38873a <=( (not A169)  and  a38872a );
 a38877a <=( A201  and  (not A200) );
 a38878a <=( A199  and  a38877a );
 a38879a <=( a38878a  and  a38873a );
 a38883a <=( A233  and  A232 );
 a38884a <=( A203  and  a38883a );
 a38887a <=( (not A266)  and  (not A265) );
 a38890a <=( A299  and  (not A298) );
 a38891a <=( a38890a  and  a38887a );
 a38892a <=( a38891a  and  a38884a );
 a38896a <=( (not A166)  and  (not A167) );
 a38897a <=( (not A169)  and  a38896a );
 a38901a <=( A201  and  (not A200) );
 a38902a <=( A199  and  a38901a );
 a38903a <=( a38902a  and  a38897a );
 a38907a <=( A233  and  (not A232) );
 a38908a <=( A203  and  a38907a );
 a38911a <=( (not A266)  and  A265 );
 a38914a <=( A268  and  A267 );
 a38915a <=( a38914a  and  a38911a );
 a38916a <=( a38915a  and  a38908a );
 a38920a <=( (not A166)  and  (not A167) );
 a38921a <=( (not A169)  and  a38920a );
 a38925a <=( A201  and  (not A200) );
 a38926a <=( A199  and  a38925a );
 a38927a <=( a38926a  and  a38921a );
 a38931a <=( A233  and  (not A232) );
 a38932a <=( A203  and  a38931a );
 a38935a <=( (not A266)  and  A265 );
 a38938a <=( A269  and  A267 );
 a38939a <=( a38938a  and  a38935a );
 a38940a <=( a38939a  and  a38932a );
 a38944a <=( (not A166)  and  (not A167) );
 a38945a <=( (not A169)  and  a38944a );
 a38949a <=( A201  and  (not A200) );
 a38950a <=( A199  and  a38949a );
 a38951a <=( a38950a  and  a38945a );
 a38955a <=( (not A234)  and  (not A233) );
 a38956a <=( A203  and  a38955a );
 a38959a <=( A266  and  A265 );
 a38962a <=( A299  and  (not A298) );
 a38963a <=( a38962a  and  a38959a );
 a38964a <=( a38963a  and  a38956a );
 a38968a <=( (not A166)  and  (not A167) );
 a38969a <=( (not A169)  and  a38968a );
 a38973a <=( A201  and  (not A200) );
 a38974a <=( A199  and  a38973a );
 a38975a <=( a38974a  and  a38969a );
 a38979a <=( (not A234)  and  (not A233) );
 a38980a <=( A203  and  a38979a );
 a38983a <=( (not A267)  and  (not A266) );
 a38986a <=( A299  and  (not A298) );
 a38987a <=( a38986a  and  a38983a );
 a38988a <=( a38987a  and  a38980a );
 a38992a <=( (not A166)  and  (not A167) );
 a38993a <=( (not A169)  and  a38992a );
 a38997a <=( A201  and  (not A200) );
 a38998a <=( A199  and  a38997a );
 a38999a <=( a38998a  and  a38993a );
 a39003a <=( (not A234)  and  (not A233) );
 a39004a <=( A203  and  a39003a );
 a39007a <=( (not A266)  and  (not A265) );
 a39010a <=( A299  and  (not A298) );
 a39011a <=( a39010a  and  a39007a );
 a39012a <=( a39011a  and  a39004a );
 a39016a <=( (not A166)  and  (not A167) );
 a39017a <=( (not A169)  and  a39016a );
 a39021a <=( A201  and  (not A200) );
 a39022a <=( A199  and  a39021a );
 a39023a <=( a39022a  and  a39017a );
 a39027a <=( (not A233)  and  A232 );
 a39028a <=( A203  and  a39027a );
 a39031a <=( A235  and  A234 );
 a39034a <=( (not A300)  and  A298 );
 a39035a <=( a39034a  and  a39031a );
 a39036a <=( a39035a  and  a39028a );
 a39040a <=( (not A166)  and  (not A167) );
 a39041a <=( (not A169)  and  a39040a );
 a39045a <=( A201  and  (not A200) );
 a39046a <=( A199  and  a39045a );
 a39047a <=( a39046a  and  a39041a );
 a39051a <=( (not A233)  and  A232 );
 a39052a <=( A203  and  a39051a );
 a39055a <=( A235  and  A234 );
 a39058a <=( A299  and  A298 );
 a39059a <=( a39058a  and  a39055a );
 a39060a <=( a39059a  and  a39052a );
 a39064a <=( (not A166)  and  (not A167) );
 a39065a <=( (not A169)  and  a39064a );
 a39069a <=( A201  and  (not A200) );
 a39070a <=( A199  and  a39069a );
 a39071a <=( a39070a  and  a39065a );
 a39075a <=( (not A233)  and  A232 );
 a39076a <=( A203  and  a39075a );
 a39079a <=( A235  and  A234 );
 a39082a <=( (not A299)  and  (not A298) );
 a39083a <=( a39082a  and  a39079a );
 a39084a <=( a39083a  and  a39076a );
 a39088a <=( (not A166)  and  (not A167) );
 a39089a <=( (not A169)  and  a39088a );
 a39093a <=( A201  and  (not A200) );
 a39094a <=( A199  and  a39093a );
 a39095a <=( a39094a  and  a39089a );
 a39099a <=( (not A233)  and  A232 );
 a39100a <=( A203  and  a39099a );
 a39103a <=( A235  and  A234 );
 a39106a <=( A266  and  (not A265) );
 a39107a <=( a39106a  and  a39103a );
 a39108a <=( a39107a  and  a39100a );
 a39112a <=( (not A166)  and  (not A167) );
 a39113a <=( (not A169)  and  a39112a );
 a39117a <=( A201  and  (not A200) );
 a39118a <=( A199  and  a39117a );
 a39119a <=( a39118a  and  a39113a );
 a39123a <=( (not A233)  and  A232 );
 a39124a <=( A203  and  a39123a );
 a39127a <=( A236  and  A234 );
 a39130a <=( (not A300)  and  A298 );
 a39131a <=( a39130a  and  a39127a );
 a39132a <=( a39131a  and  a39124a );
 a39136a <=( (not A166)  and  (not A167) );
 a39137a <=( (not A169)  and  a39136a );
 a39141a <=( A201  and  (not A200) );
 a39142a <=( A199  and  a39141a );
 a39143a <=( a39142a  and  a39137a );
 a39147a <=( (not A233)  and  A232 );
 a39148a <=( A203  and  a39147a );
 a39151a <=( A236  and  A234 );
 a39154a <=( A299  and  A298 );
 a39155a <=( a39154a  and  a39151a );
 a39156a <=( a39155a  and  a39148a );
 a39160a <=( (not A166)  and  (not A167) );
 a39161a <=( (not A169)  and  a39160a );
 a39165a <=( A201  and  (not A200) );
 a39166a <=( A199  and  a39165a );
 a39167a <=( a39166a  and  a39161a );
 a39171a <=( (not A233)  and  A232 );
 a39172a <=( A203  and  a39171a );
 a39175a <=( A236  and  A234 );
 a39178a <=( (not A299)  and  (not A298) );
 a39179a <=( a39178a  and  a39175a );
 a39180a <=( a39179a  and  a39172a );
 a39184a <=( (not A166)  and  (not A167) );
 a39185a <=( (not A169)  and  a39184a );
 a39189a <=( A201  and  (not A200) );
 a39190a <=( A199  and  a39189a );
 a39191a <=( a39190a  and  a39185a );
 a39195a <=( (not A233)  and  A232 );
 a39196a <=( A203  and  a39195a );
 a39199a <=( A236  and  A234 );
 a39202a <=( A266  and  (not A265) );
 a39203a <=( a39202a  and  a39199a );
 a39204a <=( a39203a  and  a39196a );
 a39208a <=( (not A166)  and  (not A167) );
 a39209a <=( (not A169)  and  a39208a );
 a39213a <=( A201  and  (not A200) );
 a39214a <=( A199  and  a39213a );
 a39215a <=( a39214a  and  a39209a );
 a39219a <=( (not A233)  and  (not A232) );
 a39220a <=( A203  and  a39219a );
 a39223a <=( A266  and  A265 );
 a39226a <=( A299  and  (not A298) );
 a39227a <=( a39226a  and  a39223a );
 a39228a <=( a39227a  and  a39220a );
 a39232a <=( (not A166)  and  (not A167) );
 a39233a <=( (not A169)  and  a39232a );
 a39237a <=( A201  and  (not A200) );
 a39238a <=( A199  and  a39237a );
 a39239a <=( a39238a  and  a39233a );
 a39243a <=( (not A233)  and  (not A232) );
 a39244a <=( A203  and  a39243a );
 a39247a <=( (not A267)  and  (not A266) );
 a39250a <=( A299  and  (not A298) );
 a39251a <=( a39250a  and  a39247a );
 a39252a <=( a39251a  and  a39244a );
 a39256a <=( (not A166)  and  (not A167) );
 a39257a <=( (not A169)  and  a39256a );
 a39261a <=( A201  and  (not A200) );
 a39262a <=( A199  and  a39261a );
 a39263a <=( a39262a  and  a39257a );
 a39267a <=( (not A233)  and  (not A232) );
 a39268a <=( A203  and  a39267a );
 a39271a <=( (not A266)  and  (not A265) );
 a39274a <=( A299  and  (not A298) );
 a39275a <=( a39274a  and  a39271a );
 a39276a <=( a39275a  and  a39268a );
 a39280a <=( A167  and  (not A168) );
 a39281a <=( (not A169)  and  a39280a );
 a39285a <=( A200  and  (not A199) );
 a39286a <=( A166  and  a39285a );
 a39287a <=( a39286a  and  a39281a );
 a39291a <=( A265  and  A233 );
 a39292a <=( A232  and  a39291a );
 a39295a <=( (not A269)  and  (not A268) );
 a39298a <=( A299  and  (not A298) );
 a39299a <=( a39298a  and  a39295a );
 a39300a <=( a39299a  and  a39292a );
 a39304a <=( A167  and  (not A168) );
 a39305a <=( (not A169)  and  a39304a );
 a39309a <=( A200  and  (not A199) );
 a39310a <=( A166  and  a39309a );
 a39311a <=( a39310a  and  a39305a );
 a39315a <=( (not A236)  and  (not A235) );
 a39316a <=( (not A233)  and  a39315a );
 a39319a <=( A266  and  A265 );
 a39322a <=( A299  and  (not A298) );
 a39323a <=( a39322a  and  a39319a );
 a39324a <=( a39323a  and  a39316a );
 a39328a <=( A167  and  (not A168) );
 a39329a <=( (not A169)  and  a39328a );
 a39333a <=( A200  and  (not A199) );
 a39334a <=( A166  and  a39333a );
 a39335a <=( a39334a  and  a39329a );
 a39339a <=( (not A236)  and  (not A235) );
 a39340a <=( (not A233)  and  a39339a );
 a39343a <=( (not A267)  and  (not A266) );
 a39346a <=( A299  and  (not A298) );
 a39347a <=( a39346a  and  a39343a );
 a39348a <=( a39347a  and  a39340a );
 a39352a <=( A167  and  (not A168) );
 a39353a <=( (not A169)  and  a39352a );
 a39357a <=( A200  and  (not A199) );
 a39358a <=( A166  and  a39357a );
 a39359a <=( a39358a  and  a39353a );
 a39363a <=( (not A236)  and  (not A235) );
 a39364a <=( (not A233)  and  a39363a );
 a39367a <=( (not A266)  and  (not A265) );
 a39370a <=( A299  and  (not A298) );
 a39371a <=( a39370a  and  a39367a );
 a39372a <=( a39371a  and  a39364a );
 a39376a <=( A167  and  (not A168) );
 a39377a <=( (not A169)  and  a39376a );
 a39381a <=( A200  and  (not A199) );
 a39382a <=( A166  and  a39381a );
 a39383a <=( a39382a  and  a39377a );
 a39387a <=( (not A266)  and  (not A234) );
 a39388a <=( (not A233)  and  a39387a );
 a39391a <=( (not A269)  and  (not A268) );
 a39394a <=( A299  and  (not A298) );
 a39395a <=( a39394a  and  a39391a );
 a39396a <=( a39395a  and  a39388a );
 a39400a <=( A167  and  (not A168) );
 a39401a <=( (not A169)  and  a39400a );
 a39405a <=( A200  and  (not A199) );
 a39406a <=( A166  and  a39405a );
 a39407a <=( a39406a  and  a39401a );
 a39411a <=( A234  and  (not A233) );
 a39412a <=( A232  and  a39411a );
 a39415a <=( A298  and  A235 );
 a39418a <=( (not A302)  and  (not A301) );
 a39419a <=( a39418a  and  a39415a );
 a39420a <=( a39419a  and  a39412a );
 a39424a <=( A167  and  (not A168) );
 a39425a <=( (not A169)  and  a39424a );
 a39429a <=( A200  and  (not A199) );
 a39430a <=( A166  and  a39429a );
 a39431a <=( a39430a  and  a39425a );
 a39435a <=( A234  and  (not A233) );
 a39436a <=( A232  and  a39435a );
 a39439a <=( A298  and  A236 );
 a39442a <=( (not A302)  and  (not A301) );
 a39443a <=( a39442a  and  a39439a );
 a39444a <=( a39443a  and  a39436a );
 a39448a <=( A167  and  (not A168) );
 a39449a <=( (not A169)  and  a39448a );
 a39453a <=( A200  and  (not A199) );
 a39454a <=( A166  and  a39453a );
 a39455a <=( a39454a  and  a39449a );
 a39459a <=( (not A266)  and  (not A233) );
 a39460a <=( (not A232)  and  a39459a );
 a39463a <=( (not A269)  and  (not A268) );
 a39466a <=( A299  and  (not A298) );
 a39467a <=( a39466a  and  a39463a );
 a39468a <=( a39467a  and  a39460a );
 a39472a <=( A167  and  (not A168) );
 a39473a <=( (not A169)  and  a39472a );
 a39477a <=( (not A200)  and  A199 );
 a39478a <=( A166  and  a39477a );
 a39479a <=( a39478a  and  a39473a );
 a39483a <=( (not A232)  and  A202 );
 a39484a <=( A201  and  a39483a );
 a39487a <=( (not A299)  and  A233 );
 a39490a <=( (not A302)  and  (not A301) );
 a39491a <=( a39490a  and  a39487a );
 a39492a <=( a39491a  and  a39484a );
 a39496a <=( A167  and  (not A168) );
 a39497a <=( (not A169)  and  a39496a );
 a39501a <=( (not A200)  and  A199 );
 a39502a <=( A166  and  a39501a );
 a39503a <=( a39502a  and  a39497a );
 a39507a <=( (not A232)  and  A203 );
 a39508a <=( A201  and  a39507a );
 a39511a <=( (not A299)  and  A233 );
 a39514a <=( (not A302)  and  (not A301) );
 a39515a <=( a39514a  and  a39511a );
 a39516a <=( a39515a  and  a39508a );
 a39520a <=( A167  and  (not A169) );
 a39521a <=( A170  and  a39520a );
 a39525a <=( A200  and  A199 );
 a39526a <=( (not A166)  and  a39525a );
 a39527a <=( a39526a  and  a39521a );
 a39531a <=( A265  and  A233 );
 a39532a <=( A232  and  a39531a );
 a39535a <=( (not A269)  and  (not A268) );
 a39538a <=( A299  and  (not A298) );
 a39539a <=( a39538a  and  a39535a );
 a39540a <=( a39539a  and  a39532a );
 a39544a <=( A167  and  (not A169) );
 a39545a <=( A170  and  a39544a );
 a39549a <=( A200  and  A199 );
 a39550a <=( (not A166)  and  a39549a );
 a39551a <=( a39550a  and  a39545a );
 a39555a <=( (not A236)  and  (not A235) );
 a39556a <=( (not A233)  and  a39555a );
 a39559a <=( A266  and  A265 );
 a39562a <=( A299  and  (not A298) );
 a39563a <=( a39562a  and  a39559a );
 a39564a <=( a39563a  and  a39556a );
 a39568a <=( A167  and  (not A169) );
 a39569a <=( A170  and  a39568a );
 a39573a <=( A200  and  A199 );
 a39574a <=( (not A166)  and  a39573a );
 a39575a <=( a39574a  and  a39569a );
 a39579a <=( (not A236)  and  (not A235) );
 a39580a <=( (not A233)  and  a39579a );
 a39583a <=( (not A267)  and  (not A266) );
 a39586a <=( A299  and  (not A298) );
 a39587a <=( a39586a  and  a39583a );
 a39588a <=( a39587a  and  a39580a );
 a39592a <=( A167  and  (not A169) );
 a39593a <=( A170  and  a39592a );
 a39597a <=( A200  and  A199 );
 a39598a <=( (not A166)  and  a39597a );
 a39599a <=( a39598a  and  a39593a );
 a39603a <=( (not A236)  and  (not A235) );
 a39604a <=( (not A233)  and  a39603a );
 a39607a <=( (not A266)  and  (not A265) );
 a39610a <=( A299  and  (not A298) );
 a39611a <=( a39610a  and  a39607a );
 a39612a <=( a39611a  and  a39604a );
 a39616a <=( A167  and  (not A169) );
 a39617a <=( A170  and  a39616a );
 a39621a <=( A200  and  A199 );
 a39622a <=( (not A166)  and  a39621a );
 a39623a <=( a39622a  and  a39617a );
 a39627a <=( (not A266)  and  (not A234) );
 a39628a <=( (not A233)  and  a39627a );
 a39631a <=( (not A269)  and  (not A268) );
 a39634a <=( A299  and  (not A298) );
 a39635a <=( a39634a  and  a39631a );
 a39636a <=( a39635a  and  a39628a );
 a39640a <=( A167  and  (not A169) );
 a39641a <=( A170  and  a39640a );
 a39645a <=( A200  and  A199 );
 a39646a <=( (not A166)  and  a39645a );
 a39647a <=( a39646a  and  a39641a );
 a39651a <=( A234  and  (not A233) );
 a39652a <=( A232  and  a39651a );
 a39655a <=( A298  and  A235 );
 a39658a <=( (not A302)  and  (not A301) );
 a39659a <=( a39658a  and  a39655a );
 a39660a <=( a39659a  and  a39652a );
 a39664a <=( A167  and  (not A169) );
 a39665a <=( A170  and  a39664a );
 a39669a <=( A200  and  A199 );
 a39670a <=( (not A166)  and  a39669a );
 a39671a <=( a39670a  and  a39665a );
 a39675a <=( A234  and  (not A233) );
 a39676a <=( A232  and  a39675a );
 a39679a <=( A298  and  A236 );
 a39682a <=( (not A302)  and  (not A301) );
 a39683a <=( a39682a  and  a39679a );
 a39684a <=( a39683a  and  a39676a );
 a39688a <=( A167  and  (not A169) );
 a39689a <=( A170  and  a39688a );
 a39693a <=( A200  and  A199 );
 a39694a <=( (not A166)  and  a39693a );
 a39695a <=( a39694a  and  a39689a );
 a39699a <=( (not A266)  and  (not A233) );
 a39700a <=( (not A232)  and  a39699a );
 a39703a <=( (not A269)  and  (not A268) );
 a39706a <=( A299  and  (not A298) );
 a39707a <=( a39706a  and  a39703a );
 a39708a <=( a39707a  and  a39700a );
 a39712a <=( A167  and  (not A169) );
 a39713a <=( A170  and  a39712a );
 a39717a <=( (not A202)  and  (not A200) );
 a39718a <=( (not A166)  and  a39717a );
 a39719a <=( a39718a  and  a39713a );
 a39723a <=( A233  and  A232 );
 a39724a <=( (not A203)  and  a39723a );
 a39727a <=( (not A267)  and  A265 );
 a39730a <=( A299  and  (not A298) );
 a39731a <=( a39730a  and  a39727a );
 a39732a <=( a39731a  and  a39724a );
 a39736a <=( A167  and  (not A169) );
 a39737a <=( A170  and  a39736a );
 a39741a <=( (not A202)  and  (not A200) );
 a39742a <=( (not A166)  and  a39741a );
 a39743a <=( a39742a  and  a39737a );
 a39747a <=( A233  and  A232 );
 a39748a <=( (not A203)  and  a39747a );
 a39751a <=( A266  and  A265 );
 a39754a <=( A299  and  (not A298) );
 a39755a <=( a39754a  and  a39751a );
 a39756a <=( a39755a  and  a39748a );
 a39760a <=( A167  and  (not A169) );
 a39761a <=( A170  and  a39760a );
 a39765a <=( (not A202)  and  (not A200) );
 a39766a <=( (not A166)  and  a39765a );
 a39767a <=( a39766a  and  a39761a );
 a39771a <=( A233  and  A232 );
 a39772a <=( (not A203)  and  a39771a );
 a39775a <=( (not A266)  and  (not A265) );
 a39778a <=( A299  and  (not A298) );
 a39779a <=( a39778a  and  a39775a );
 a39780a <=( a39779a  and  a39772a );
 a39784a <=( A167  and  (not A169) );
 a39785a <=( A170  and  a39784a );
 a39789a <=( (not A202)  and  (not A200) );
 a39790a <=( (not A166)  and  a39789a );
 a39791a <=( a39790a  and  a39785a );
 a39795a <=( A233  and  (not A232) );
 a39796a <=( (not A203)  and  a39795a );
 a39799a <=( (not A266)  and  A265 );
 a39802a <=( A268  and  A267 );
 a39803a <=( a39802a  and  a39799a );
 a39804a <=( a39803a  and  a39796a );
 a39808a <=( A167  and  (not A169) );
 a39809a <=( A170  and  a39808a );
 a39813a <=( (not A202)  and  (not A200) );
 a39814a <=( (not A166)  and  a39813a );
 a39815a <=( a39814a  and  a39809a );
 a39819a <=( A233  and  (not A232) );
 a39820a <=( (not A203)  and  a39819a );
 a39823a <=( (not A266)  and  A265 );
 a39826a <=( A269  and  A267 );
 a39827a <=( a39826a  and  a39823a );
 a39828a <=( a39827a  and  a39820a );
 a39832a <=( A167  and  (not A169) );
 a39833a <=( A170  and  a39832a );
 a39837a <=( (not A202)  and  (not A200) );
 a39838a <=( (not A166)  and  a39837a );
 a39839a <=( a39838a  and  a39833a );
 a39843a <=( (not A234)  and  (not A233) );
 a39844a <=( (not A203)  and  a39843a );
 a39847a <=( A266  and  A265 );
 a39850a <=( A299  and  (not A298) );
 a39851a <=( a39850a  and  a39847a );
 a39852a <=( a39851a  and  a39844a );
 a39856a <=( A167  and  (not A169) );
 a39857a <=( A170  and  a39856a );
 a39861a <=( (not A202)  and  (not A200) );
 a39862a <=( (not A166)  and  a39861a );
 a39863a <=( a39862a  and  a39857a );
 a39867a <=( (not A234)  and  (not A233) );
 a39868a <=( (not A203)  and  a39867a );
 a39871a <=( (not A267)  and  (not A266) );
 a39874a <=( A299  and  (not A298) );
 a39875a <=( a39874a  and  a39871a );
 a39876a <=( a39875a  and  a39868a );
 a39880a <=( A167  and  (not A169) );
 a39881a <=( A170  and  a39880a );
 a39885a <=( (not A202)  and  (not A200) );
 a39886a <=( (not A166)  and  a39885a );
 a39887a <=( a39886a  and  a39881a );
 a39891a <=( (not A234)  and  (not A233) );
 a39892a <=( (not A203)  and  a39891a );
 a39895a <=( (not A266)  and  (not A265) );
 a39898a <=( A299  and  (not A298) );
 a39899a <=( a39898a  and  a39895a );
 a39900a <=( a39899a  and  a39892a );
 a39904a <=( A167  and  (not A169) );
 a39905a <=( A170  and  a39904a );
 a39909a <=( (not A202)  and  (not A200) );
 a39910a <=( (not A166)  and  a39909a );
 a39911a <=( a39910a  and  a39905a );
 a39915a <=( (not A233)  and  A232 );
 a39916a <=( (not A203)  and  a39915a );
 a39919a <=( A235  and  A234 );
 a39922a <=( (not A300)  and  A298 );
 a39923a <=( a39922a  and  a39919a );
 a39924a <=( a39923a  and  a39916a );
 a39928a <=( A167  and  (not A169) );
 a39929a <=( A170  and  a39928a );
 a39933a <=( (not A202)  and  (not A200) );
 a39934a <=( (not A166)  and  a39933a );
 a39935a <=( a39934a  and  a39929a );
 a39939a <=( (not A233)  and  A232 );
 a39940a <=( (not A203)  and  a39939a );
 a39943a <=( A235  and  A234 );
 a39946a <=( A299  and  A298 );
 a39947a <=( a39946a  and  a39943a );
 a39948a <=( a39947a  and  a39940a );
 a39952a <=( A167  and  (not A169) );
 a39953a <=( A170  and  a39952a );
 a39957a <=( (not A202)  and  (not A200) );
 a39958a <=( (not A166)  and  a39957a );
 a39959a <=( a39958a  and  a39953a );
 a39963a <=( (not A233)  and  A232 );
 a39964a <=( (not A203)  and  a39963a );
 a39967a <=( A235  and  A234 );
 a39970a <=( (not A299)  and  (not A298) );
 a39971a <=( a39970a  and  a39967a );
 a39972a <=( a39971a  and  a39964a );
 a39976a <=( A167  and  (not A169) );
 a39977a <=( A170  and  a39976a );
 a39981a <=( (not A202)  and  (not A200) );
 a39982a <=( (not A166)  and  a39981a );
 a39983a <=( a39982a  and  a39977a );
 a39987a <=( (not A233)  and  A232 );
 a39988a <=( (not A203)  and  a39987a );
 a39991a <=( A235  and  A234 );
 a39994a <=( A266  and  (not A265) );
 a39995a <=( a39994a  and  a39991a );
 a39996a <=( a39995a  and  a39988a );
 a40000a <=( A167  and  (not A169) );
 a40001a <=( A170  and  a40000a );
 a40005a <=( (not A202)  and  (not A200) );
 a40006a <=( (not A166)  and  a40005a );
 a40007a <=( a40006a  and  a40001a );
 a40011a <=( (not A233)  and  A232 );
 a40012a <=( (not A203)  and  a40011a );
 a40015a <=( A236  and  A234 );
 a40018a <=( (not A300)  and  A298 );
 a40019a <=( a40018a  and  a40015a );
 a40020a <=( a40019a  and  a40012a );
 a40024a <=( A167  and  (not A169) );
 a40025a <=( A170  and  a40024a );
 a40029a <=( (not A202)  and  (not A200) );
 a40030a <=( (not A166)  and  a40029a );
 a40031a <=( a40030a  and  a40025a );
 a40035a <=( (not A233)  and  A232 );
 a40036a <=( (not A203)  and  a40035a );
 a40039a <=( A236  and  A234 );
 a40042a <=( A299  and  A298 );
 a40043a <=( a40042a  and  a40039a );
 a40044a <=( a40043a  and  a40036a );
 a40048a <=( A167  and  (not A169) );
 a40049a <=( A170  and  a40048a );
 a40053a <=( (not A202)  and  (not A200) );
 a40054a <=( (not A166)  and  a40053a );
 a40055a <=( a40054a  and  a40049a );
 a40059a <=( (not A233)  and  A232 );
 a40060a <=( (not A203)  and  a40059a );
 a40063a <=( A236  and  A234 );
 a40066a <=( (not A299)  and  (not A298) );
 a40067a <=( a40066a  and  a40063a );
 a40068a <=( a40067a  and  a40060a );
 a40072a <=( A167  and  (not A169) );
 a40073a <=( A170  and  a40072a );
 a40077a <=( (not A202)  and  (not A200) );
 a40078a <=( (not A166)  and  a40077a );
 a40079a <=( a40078a  and  a40073a );
 a40083a <=( (not A233)  and  A232 );
 a40084a <=( (not A203)  and  a40083a );
 a40087a <=( A236  and  A234 );
 a40090a <=( A266  and  (not A265) );
 a40091a <=( a40090a  and  a40087a );
 a40092a <=( a40091a  and  a40084a );
 a40096a <=( A167  and  (not A169) );
 a40097a <=( A170  and  a40096a );
 a40101a <=( (not A202)  and  (not A200) );
 a40102a <=( (not A166)  and  a40101a );
 a40103a <=( a40102a  and  a40097a );
 a40107a <=( (not A233)  and  (not A232) );
 a40108a <=( (not A203)  and  a40107a );
 a40111a <=( A266  and  A265 );
 a40114a <=( A299  and  (not A298) );
 a40115a <=( a40114a  and  a40111a );
 a40116a <=( a40115a  and  a40108a );
 a40120a <=( A167  and  (not A169) );
 a40121a <=( A170  and  a40120a );
 a40125a <=( (not A202)  and  (not A200) );
 a40126a <=( (not A166)  and  a40125a );
 a40127a <=( a40126a  and  a40121a );
 a40131a <=( (not A233)  and  (not A232) );
 a40132a <=( (not A203)  and  a40131a );
 a40135a <=( (not A267)  and  (not A266) );
 a40138a <=( A299  and  (not A298) );
 a40139a <=( a40138a  and  a40135a );
 a40140a <=( a40139a  and  a40132a );
 a40144a <=( A167  and  (not A169) );
 a40145a <=( A170  and  a40144a );
 a40149a <=( (not A202)  and  (not A200) );
 a40150a <=( (not A166)  and  a40149a );
 a40151a <=( a40150a  and  a40145a );
 a40155a <=( (not A233)  and  (not A232) );
 a40156a <=( (not A203)  and  a40155a );
 a40159a <=( (not A266)  and  (not A265) );
 a40162a <=( A299  and  (not A298) );
 a40163a <=( a40162a  and  a40159a );
 a40164a <=( a40163a  and  a40156a );
 a40168a <=( A167  and  (not A169) );
 a40169a <=( A170  and  a40168a );
 a40173a <=( (not A201)  and  (not A200) );
 a40174a <=( (not A166)  and  a40173a );
 a40175a <=( a40174a  and  a40169a );
 a40179a <=( A265  and  A233 );
 a40180a <=( A232  and  a40179a );
 a40183a <=( (not A269)  and  (not A268) );
 a40186a <=( A299  and  (not A298) );
 a40187a <=( a40186a  and  a40183a );
 a40188a <=( a40187a  and  a40180a );
 a40192a <=( A167  and  (not A169) );
 a40193a <=( A170  and  a40192a );
 a40197a <=( (not A201)  and  (not A200) );
 a40198a <=( (not A166)  and  a40197a );
 a40199a <=( a40198a  and  a40193a );
 a40203a <=( (not A236)  and  (not A235) );
 a40204a <=( (not A233)  and  a40203a );
 a40207a <=( A266  and  A265 );
 a40210a <=( A299  and  (not A298) );
 a40211a <=( a40210a  and  a40207a );
 a40212a <=( a40211a  and  a40204a );
 a40216a <=( A167  and  (not A169) );
 a40217a <=( A170  and  a40216a );
 a40221a <=( (not A201)  and  (not A200) );
 a40222a <=( (not A166)  and  a40221a );
 a40223a <=( a40222a  and  a40217a );
 a40227a <=( (not A236)  and  (not A235) );
 a40228a <=( (not A233)  and  a40227a );
 a40231a <=( (not A267)  and  (not A266) );
 a40234a <=( A299  and  (not A298) );
 a40235a <=( a40234a  and  a40231a );
 a40236a <=( a40235a  and  a40228a );
 a40240a <=( A167  and  (not A169) );
 a40241a <=( A170  and  a40240a );
 a40245a <=( (not A201)  and  (not A200) );
 a40246a <=( (not A166)  and  a40245a );
 a40247a <=( a40246a  and  a40241a );
 a40251a <=( (not A236)  and  (not A235) );
 a40252a <=( (not A233)  and  a40251a );
 a40255a <=( (not A266)  and  (not A265) );
 a40258a <=( A299  and  (not A298) );
 a40259a <=( a40258a  and  a40255a );
 a40260a <=( a40259a  and  a40252a );
 a40264a <=( A167  and  (not A169) );
 a40265a <=( A170  and  a40264a );
 a40269a <=( (not A201)  and  (not A200) );
 a40270a <=( (not A166)  and  a40269a );
 a40271a <=( a40270a  and  a40265a );
 a40275a <=( (not A266)  and  (not A234) );
 a40276a <=( (not A233)  and  a40275a );
 a40279a <=( (not A269)  and  (not A268) );
 a40282a <=( A299  and  (not A298) );
 a40283a <=( a40282a  and  a40279a );
 a40284a <=( a40283a  and  a40276a );
 a40288a <=( A167  and  (not A169) );
 a40289a <=( A170  and  a40288a );
 a40293a <=( (not A201)  and  (not A200) );
 a40294a <=( (not A166)  and  a40293a );
 a40295a <=( a40294a  and  a40289a );
 a40299a <=( A234  and  (not A233) );
 a40300a <=( A232  and  a40299a );
 a40303a <=( A298  and  A235 );
 a40306a <=( (not A302)  and  (not A301) );
 a40307a <=( a40306a  and  a40303a );
 a40308a <=( a40307a  and  a40300a );
 a40312a <=( A167  and  (not A169) );
 a40313a <=( A170  and  a40312a );
 a40317a <=( (not A201)  and  (not A200) );
 a40318a <=( (not A166)  and  a40317a );
 a40319a <=( a40318a  and  a40313a );
 a40323a <=( A234  and  (not A233) );
 a40324a <=( A232  and  a40323a );
 a40327a <=( A298  and  A236 );
 a40330a <=( (not A302)  and  (not A301) );
 a40331a <=( a40330a  and  a40327a );
 a40332a <=( a40331a  and  a40324a );
 a40336a <=( A167  and  (not A169) );
 a40337a <=( A170  and  a40336a );
 a40341a <=( (not A201)  and  (not A200) );
 a40342a <=( (not A166)  and  a40341a );
 a40343a <=( a40342a  and  a40337a );
 a40347a <=( (not A266)  and  (not A233) );
 a40348a <=( (not A232)  and  a40347a );
 a40351a <=( (not A269)  and  (not A268) );
 a40354a <=( A299  and  (not A298) );
 a40355a <=( a40354a  and  a40351a );
 a40356a <=( a40355a  and  a40348a );
 a40360a <=( A167  and  (not A169) );
 a40361a <=( A170  and  a40360a );
 a40365a <=( (not A200)  and  (not A199) );
 a40366a <=( (not A166)  and  a40365a );
 a40367a <=( a40366a  and  a40361a );
 a40371a <=( A265  and  A233 );
 a40372a <=( A232  and  a40371a );
 a40375a <=( (not A269)  and  (not A268) );
 a40378a <=( A299  and  (not A298) );
 a40379a <=( a40378a  and  a40375a );
 a40380a <=( a40379a  and  a40372a );
 a40384a <=( A167  and  (not A169) );
 a40385a <=( A170  and  a40384a );
 a40389a <=( (not A200)  and  (not A199) );
 a40390a <=( (not A166)  and  a40389a );
 a40391a <=( a40390a  and  a40385a );
 a40395a <=( (not A236)  and  (not A235) );
 a40396a <=( (not A233)  and  a40395a );
 a40399a <=( A266  and  A265 );
 a40402a <=( A299  and  (not A298) );
 a40403a <=( a40402a  and  a40399a );
 a40404a <=( a40403a  and  a40396a );
 a40408a <=( A167  and  (not A169) );
 a40409a <=( A170  and  a40408a );
 a40413a <=( (not A200)  and  (not A199) );
 a40414a <=( (not A166)  and  a40413a );
 a40415a <=( a40414a  and  a40409a );
 a40419a <=( (not A236)  and  (not A235) );
 a40420a <=( (not A233)  and  a40419a );
 a40423a <=( (not A267)  and  (not A266) );
 a40426a <=( A299  and  (not A298) );
 a40427a <=( a40426a  and  a40423a );
 a40428a <=( a40427a  and  a40420a );
 a40432a <=( A167  and  (not A169) );
 a40433a <=( A170  and  a40432a );
 a40437a <=( (not A200)  and  (not A199) );
 a40438a <=( (not A166)  and  a40437a );
 a40439a <=( a40438a  and  a40433a );
 a40443a <=( (not A236)  and  (not A235) );
 a40444a <=( (not A233)  and  a40443a );
 a40447a <=( (not A266)  and  (not A265) );
 a40450a <=( A299  and  (not A298) );
 a40451a <=( a40450a  and  a40447a );
 a40452a <=( a40451a  and  a40444a );
 a40456a <=( A167  and  (not A169) );
 a40457a <=( A170  and  a40456a );
 a40461a <=( (not A200)  and  (not A199) );
 a40462a <=( (not A166)  and  a40461a );
 a40463a <=( a40462a  and  a40457a );
 a40467a <=( (not A266)  and  (not A234) );
 a40468a <=( (not A233)  and  a40467a );
 a40471a <=( (not A269)  and  (not A268) );
 a40474a <=( A299  and  (not A298) );
 a40475a <=( a40474a  and  a40471a );
 a40476a <=( a40475a  and  a40468a );
 a40480a <=( A167  and  (not A169) );
 a40481a <=( A170  and  a40480a );
 a40485a <=( (not A200)  and  (not A199) );
 a40486a <=( (not A166)  and  a40485a );
 a40487a <=( a40486a  and  a40481a );
 a40491a <=( A234  and  (not A233) );
 a40492a <=( A232  and  a40491a );
 a40495a <=( A298  and  A235 );
 a40498a <=( (not A302)  and  (not A301) );
 a40499a <=( a40498a  and  a40495a );
 a40500a <=( a40499a  and  a40492a );
 a40504a <=( A167  and  (not A169) );
 a40505a <=( A170  and  a40504a );
 a40509a <=( (not A200)  and  (not A199) );
 a40510a <=( (not A166)  and  a40509a );
 a40511a <=( a40510a  and  a40505a );
 a40515a <=( A234  and  (not A233) );
 a40516a <=( A232  and  a40515a );
 a40519a <=( A298  and  A236 );
 a40522a <=( (not A302)  and  (not A301) );
 a40523a <=( a40522a  and  a40519a );
 a40524a <=( a40523a  and  a40516a );
 a40528a <=( A167  and  (not A169) );
 a40529a <=( A170  and  a40528a );
 a40533a <=( (not A200)  and  (not A199) );
 a40534a <=( (not A166)  and  a40533a );
 a40535a <=( a40534a  and  a40529a );
 a40539a <=( (not A266)  and  (not A233) );
 a40540a <=( (not A232)  and  a40539a );
 a40543a <=( (not A269)  and  (not A268) );
 a40546a <=( A299  and  (not A298) );
 a40547a <=( a40546a  and  a40543a );
 a40548a <=( a40547a  and  a40540a );
 a40552a <=( (not A167)  and  (not A169) );
 a40553a <=( A170  and  a40552a );
 a40557a <=( A200  and  A199 );
 a40558a <=( A166  and  a40557a );
 a40559a <=( a40558a  and  a40553a );
 a40563a <=( A265  and  A233 );
 a40564a <=( A232  and  a40563a );
 a40567a <=( (not A269)  and  (not A268) );
 a40570a <=( A299  and  (not A298) );
 a40571a <=( a40570a  and  a40567a );
 a40572a <=( a40571a  and  a40564a );
 a40576a <=( (not A167)  and  (not A169) );
 a40577a <=( A170  and  a40576a );
 a40581a <=( A200  and  A199 );
 a40582a <=( A166  and  a40581a );
 a40583a <=( a40582a  and  a40577a );
 a40587a <=( (not A236)  and  (not A235) );
 a40588a <=( (not A233)  and  a40587a );
 a40591a <=( A266  and  A265 );
 a40594a <=( A299  and  (not A298) );
 a40595a <=( a40594a  and  a40591a );
 a40596a <=( a40595a  and  a40588a );
 a40600a <=( (not A167)  and  (not A169) );
 a40601a <=( A170  and  a40600a );
 a40605a <=( A200  and  A199 );
 a40606a <=( A166  and  a40605a );
 a40607a <=( a40606a  and  a40601a );
 a40611a <=( (not A236)  and  (not A235) );
 a40612a <=( (not A233)  and  a40611a );
 a40615a <=( (not A267)  and  (not A266) );
 a40618a <=( A299  and  (not A298) );
 a40619a <=( a40618a  and  a40615a );
 a40620a <=( a40619a  and  a40612a );
 a40624a <=( (not A167)  and  (not A169) );
 a40625a <=( A170  and  a40624a );
 a40629a <=( A200  and  A199 );
 a40630a <=( A166  and  a40629a );
 a40631a <=( a40630a  and  a40625a );
 a40635a <=( (not A236)  and  (not A235) );
 a40636a <=( (not A233)  and  a40635a );
 a40639a <=( (not A266)  and  (not A265) );
 a40642a <=( A299  and  (not A298) );
 a40643a <=( a40642a  and  a40639a );
 a40644a <=( a40643a  and  a40636a );
 a40648a <=( (not A167)  and  (not A169) );
 a40649a <=( A170  and  a40648a );
 a40653a <=( A200  and  A199 );
 a40654a <=( A166  and  a40653a );
 a40655a <=( a40654a  and  a40649a );
 a40659a <=( (not A266)  and  (not A234) );
 a40660a <=( (not A233)  and  a40659a );
 a40663a <=( (not A269)  and  (not A268) );
 a40666a <=( A299  and  (not A298) );
 a40667a <=( a40666a  and  a40663a );
 a40668a <=( a40667a  and  a40660a );
 a40672a <=( (not A167)  and  (not A169) );
 a40673a <=( A170  and  a40672a );
 a40677a <=( A200  and  A199 );
 a40678a <=( A166  and  a40677a );
 a40679a <=( a40678a  and  a40673a );
 a40683a <=( A234  and  (not A233) );
 a40684a <=( A232  and  a40683a );
 a40687a <=( A298  and  A235 );
 a40690a <=( (not A302)  and  (not A301) );
 a40691a <=( a40690a  and  a40687a );
 a40692a <=( a40691a  and  a40684a );
 a40696a <=( (not A167)  and  (not A169) );
 a40697a <=( A170  and  a40696a );
 a40701a <=( A200  and  A199 );
 a40702a <=( A166  and  a40701a );
 a40703a <=( a40702a  and  a40697a );
 a40707a <=( A234  and  (not A233) );
 a40708a <=( A232  and  a40707a );
 a40711a <=( A298  and  A236 );
 a40714a <=( (not A302)  and  (not A301) );
 a40715a <=( a40714a  and  a40711a );
 a40716a <=( a40715a  and  a40708a );
 a40720a <=( (not A167)  and  (not A169) );
 a40721a <=( A170  and  a40720a );
 a40725a <=( A200  and  A199 );
 a40726a <=( A166  and  a40725a );
 a40727a <=( a40726a  and  a40721a );
 a40731a <=( (not A266)  and  (not A233) );
 a40732a <=( (not A232)  and  a40731a );
 a40735a <=( (not A269)  and  (not A268) );
 a40738a <=( A299  and  (not A298) );
 a40739a <=( a40738a  and  a40735a );
 a40740a <=( a40739a  and  a40732a );
 a40744a <=( (not A167)  and  (not A169) );
 a40745a <=( A170  and  a40744a );
 a40749a <=( (not A202)  and  (not A200) );
 a40750a <=( A166  and  a40749a );
 a40751a <=( a40750a  and  a40745a );
 a40755a <=( A233  and  A232 );
 a40756a <=( (not A203)  and  a40755a );
 a40759a <=( (not A267)  and  A265 );
 a40762a <=( A299  and  (not A298) );
 a40763a <=( a40762a  and  a40759a );
 a40764a <=( a40763a  and  a40756a );
 a40768a <=( (not A167)  and  (not A169) );
 a40769a <=( A170  and  a40768a );
 a40773a <=( (not A202)  and  (not A200) );
 a40774a <=( A166  and  a40773a );
 a40775a <=( a40774a  and  a40769a );
 a40779a <=( A233  and  A232 );
 a40780a <=( (not A203)  and  a40779a );
 a40783a <=( A266  and  A265 );
 a40786a <=( A299  and  (not A298) );
 a40787a <=( a40786a  and  a40783a );
 a40788a <=( a40787a  and  a40780a );
 a40792a <=( (not A167)  and  (not A169) );
 a40793a <=( A170  and  a40792a );
 a40797a <=( (not A202)  and  (not A200) );
 a40798a <=( A166  and  a40797a );
 a40799a <=( a40798a  and  a40793a );
 a40803a <=( A233  and  A232 );
 a40804a <=( (not A203)  and  a40803a );
 a40807a <=( (not A266)  and  (not A265) );
 a40810a <=( A299  and  (not A298) );
 a40811a <=( a40810a  and  a40807a );
 a40812a <=( a40811a  and  a40804a );
 a40816a <=( (not A167)  and  (not A169) );
 a40817a <=( A170  and  a40816a );
 a40821a <=( (not A202)  and  (not A200) );
 a40822a <=( A166  and  a40821a );
 a40823a <=( a40822a  and  a40817a );
 a40827a <=( A233  and  (not A232) );
 a40828a <=( (not A203)  and  a40827a );
 a40831a <=( (not A266)  and  A265 );
 a40834a <=( A268  and  A267 );
 a40835a <=( a40834a  and  a40831a );
 a40836a <=( a40835a  and  a40828a );
 a40840a <=( (not A167)  and  (not A169) );
 a40841a <=( A170  and  a40840a );
 a40845a <=( (not A202)  and  (not A200) );
 a40846a <=( A166  and  a40845a );
 a40847a <=( a40846a  and  a40841a );
 a40851a <=( A233  and  (not A232) );
 a40852a <=( (not A203)  and  a40851a );
 a40855a <=( (not A266)  and  A265 );
 a40858a <=( A269  and  A267 );
 a40859a <=( a40858a  and  a40855a );
 a40860a <=( a40859a  and  a40852a );
 a40864a <=( (not A167)  and  (not A169) );
 a40865a <=( A170  and  a40864a );
 a40869a <=( (not A202)  and  (not A200) );
 a40870a <=( A166  and  a40869a );
 a40871a <=( a40870a  and  a40865a );
 a40875a <=( (not A234)  and  (not A233) );
 a40876a <=( (not A203)  and  a40875a );
 a40879a <=( A266  and  A265 );
 a40882a <=( A299  and  (not A298) );
 a40883a <=( a40882a  and  a40879a );
 a40884a <=( a40883a  and  a40876a );
 a40888a <=( (not A167)  and  (not A169) );
 a40889a <=( A170  and  a40888a );
 a40893a <=( (not A202)  and  (not A200) );
 a40894a <=( A166  and  a40893a );
 a40895a <=( a40894a  and  a40889a );
 a40899a <=( (not A234)  and  (not A233) );
 a40900a <=( (not A203)  and  a40899a );
 a40903a <=( (not A267)  and  (not A266) );
 a40906a <=( A299  and  (not A298) );
 a40907a <=( a40906a  and  a40903a );
 a40908a <=( a40907a  and  a40900a );
 a40912a <=( (not A167)  and  (not A169) );
 a40913a <=( A170  and  a40912a );
 a40917a <=( (not A202)  and  (not A200) );
 a40918a <=( A166  and  a40917a );
 a40919a <=( a40918a  and  a40913a );
 a40923a <=( (not A234)  and  (not A233) );
 a40924a <=( (not A203)  and  a40923a );
 a40927a <=( (not A266)  and  (not A265) );
 a40930a <=( A299  and  (not A298) );
 a40931a <=( a40930a  and  a40927a );
 a40932a <=( a40931a  and  a40924a );
 a40936a <=( (not A167)  and  (not A169) );
 a40937a <=( A170  and  a40936a );
 a40941a <=( (not A202)  and  (not A200) );
 a40942a <=( A166  and  a40941a );
 a40943a <=( a40942a  and  a40937a );
 a40947a <=( (not A233)  and  A232 );
 a40948a <=( (not A203)  and  a40947a );
 a40951a <=( A235  and  A234 );
 a40954a <=( (not A300)  and  A298 );
 a40955a <=( a40954a  and  a40951a );
 a40956a <=( a40955a  and  a40948a );
 a40960a <=( (not A167)  and  (not A169) );
 a40961a <=( A170  and  a40960a );
 a40965a <=( (not A202)  and  (not A200) );
 a40966a <=( A166  and  a40965a );
 a40967a <=( a40966a  and  a40961a );
 a40971a <=( (not A233)  and  A232 );
 a40972a <=( (not A203)  and  a40971a );
 a40975a <=( A235  and  A234 );
 a40978a <=( A299  and  A298 );
 a40979a <=( a40978a  and  a40975a );
 a40980a <=( a40979a  and  a40972a );
 a40984a <=( (not A167)  and  (not A169) );
 a40985a <=( A170  and  a40984a );
 a40989a <=( (not A202)  and  (not A200) );
 a40990a <=( A166  and  a40989a );
 a40991a <=( a40990a  and  a40985a );
 a40995a <=( (not A233)  and  A232 );
 a40996a <=( (not A203)  and  a40995a );
 a40999a <=( A235  and  A234 );
 a41002a <=( (not A299)  and  (not A298) );
 a41003a <=( a41002a  and  a40999a );
 a41004a <=( a41003a  and  a40996a );
 a41008a <=( (not A167)  and  (not A169) );
 a41009a <=( A170  and  a41008a );
 a41013a <=( (not A202)  and  (not A200) );
 a41014a <=( A166  and  a41013a );
 a41015a <=( a41014a  and  a41009a );
 a41019a <=( (not A233)  and  A232 );
 a41020a <=( (not A203)  and  a41019a );
 a41023a <=( A235  and  A234 );
 a41026a <=( A266  and  (not A265) );
 a41027a <=( a41026a  and  a41023a );
 a41028a <=( a41027a  and  a41020a );
 a41032a <=( (not A167)  and  (not A169) );
 a41033a <=( A170  and  a41032a );
 a41037a <=( (not A202)  and  (not A200) );
 a41038a <=( A166  and  a41037a );
 a41039a <=( a41038a  and  a41033a );
 a41043a <=( (not A233)  and  A232 );
 a41044a <=( (not A203)  and  a41043a );
 a41047a <=( A236  and  A234 );
 a41050a <=( (not A300)  and  A298 );
 a41051a <=( a41050a  and  a41047a );
 a41052a <=( a41051a  and  a41044a );
 a41056a <=( (not A167)  and  (not A169) );
 a41057a <=( A170  and  a41056a );
 a41061a <=( (not A202)  and  (not A200) );
 a41062a <=( A166  and  a41061a );
 a41063a <=( a41062a  and  a41057a );
 a41067a <=( (not A233)  and  A232 );
 a41068a <=( (not A203)  and  a41067a );
 a41071a <=( A236  and  A234 );
 a41074a <=( A299  and  A298 );
 a41075a <=( a41074a  and  a41071a );
 a41076a <=( a41075a  and  a41068a );
 a41080a <=( (not A167)  and  (not A169) );
 a41081a <=( A170  and  a41080a );
 a41085a <=( (not A202)  and  (not A200) );
 a41086a <=( A166  and  a41085a );
 a41087a <=( a41086a  and  a41081a );
 a41091a <=( (not A233)  and  A232 );
 a41092a <=( (not A203)  and  a41091a );
 a41095a <=( A236  and  A234 );
 a41098a <=( (not A299)  and  (not A298) );
 a41099a <=( a41098a  and  a41095a );
 a41100a <=( a41099a  and  a41092a );
 a41104a <=( (not A167)  and  (not A169) );
 a41105a <=( A170  and  a41104a );
 a41109a <=( (not A202)  and  (not A200) );
 a41110a <=( A166  and  a41109a );
 a41111a <=( a41110a  and  a41105a );
 a41115a <=( (not A233)  and  A232 );
 a41116a <=( (not A203)  and  a41115a );
 a41119a <=( A236  and  A234 );
 a41122a <=( A266  and  (not A265) );
 a41123a <=( a41122a  and  a41119a );
 a41124a <=( a41123a  and  a41116a );
 a41128a <=( (not A167)  and  (not A169) );
 a41129a <=( A170  and  a41128a );
 a41133a <=( (not A202)  and  (not A200) );
 a41134a <=( A166  and  a41133a );
 a41135a <=( a41134a  and  a41129a );
 a41139a <=( (not A233)  and  (not A232) );
 a41140a <=( (not A203)  and  a41139a );
 a41143a <=( A266  and  A265 );
 a41146a <=( A299  and  (not A298) );
 a41147a <=( a41146a  and  a41143a );
 a41148a <=( a41147a  and  a41140a );
 a41152a <=( (not A167)  and  (not A169) );
 a41153a <=( A170  and  a41152a );
 a41157a <=( (not A202)  and  (not A200) );
 a41158a <=( A166  and  a41157a );
 a41159a <=( a41158a  and  a41153a );
 a41163a <=( (not A233)  and  (not A232) );
 a41164a <=( (not A203)  and  a41163a );
 a41167a <=( (not A267)  and  (not A266) );
 a41170a <=( A299  and  (not A298) );
 a41171a <=( a41170a  and  a41167a );
 a41172a <=( a41171a  and  a41164a );
 a41176a <=( (not A167)  and  (not A169) );
 a41177a <=( A170  and  a41176a );
 a41181a <=( (not A202)  and  (not A200) );
 a41182a <=( A166  and  a41181a );
 a41183a <=( a41182a  and  a41177a );
 a41187a <=( (not A233)  and  (not A232) );
 a41188a <=( (not A203)  and  a41187a );
 a41191a <=( (not A266)  and  (not A265) );
 a41194a <=( A299  and  (not A298) );
 a41195a <=( a41194a  and  a41191a );
 a41196a <=( a41195a  and  a41188a );
 a41200a <=( (not A167)  and  (not A169) );
 a41201a <=( A170  and  a41200a );
 a41205a <=( (not A201)  and  (not A200) );
 a41206a <=( A166  and  a41205a );
 a41207a <=( a41206a  and  a41201a );
 a41211a <=( A265  and  A233 );
 a41212a <=( A232  and  a41211a );
 a41215a <=( (not A269)  and  (not A268) );
 a41218a <=( A299  and  (not A298) );
 a41219a <=( a41218a  and  a41215a );
 a41220a <=( a41219a  and  a41212a );
 a41224a <=( (not A167)  and  (not A169) );
 a41225a <=( A170  and  a41224a );
 a41229a <=( (not A201)  and  (not A200) );
 a41230a <=( A166  and  a41229a );
 a41231a <=( a41230a  and  a41225a );
 a41235a <=( (not A236)  and  (not A235) );
 a41236a <=( (not A233)  and  a41235a );
 a41239a <=( A266  and  A265 );
 a41242a <=( A299  and  (not A298) );
 a41243a <=( a41242a  and  a41239a );
 a41244a <=( a41243a  and  a41236a );
 a41248a <=( (not A167)  and  (not A169) );
 a41249a <=( A170  and  a41248a );
 a41253a <=( (not A201)  and  (not A200) );
 a41254a <=( A166  and  a41253a );
 a41255a <=( a41254a  and  a41249a );
 a41259a <=( (not A236)  and  (not A235) );
 a41260a <=( (not A233)  and  a41259a );
 a41263a <=( (not A267)  and  (not A266) );
 a41266a <=( A299  and  (not A298) );
 a41267a <=( a41266a  and  a41263a );
 a41268a <=( a41267a  and  a41260a );
 a41272a <=( (not A167)  and  (not A169) );
 a41273a <=( A170  and  a41272a );
 a41277a <=( (not A201)  and  (not A200) );
 a41278a <=( A166  and  a41277a );
 a41279a <=( a41278a  and  a41273a );
 a41283a <=( (not A236)  and  (not A235) );
 a41284a <=( (not A233)  and  a41283a );
 a41287a <=( (not A266)  and  (not A265) );
 a41290a <=( A299  and  (not A298) );
 a41291a <=( a41290a  and  a41287a );
 a41292a <=( a41291a  and  a41284a );
 a41296a <=( (not A167)  and  (not A169) );
 a41297a <=( A170  and  a41296a );
 a41301a <=( (not A201)  and  (not A200) );
 a41302a <=( A166  and  a41301a );
 a41303a <=( a41302a  and  a41297a );
 a41307a <=( (not A266)  and  (not A234) );
 a41308a <=( (not A233)  and  a41307a );
 a41311a <=( (not A269)  and  (not A268) );
 a41314a <=( A299  and  (not A298) );
 a41315a <=( a41314a  and  a41311a );
 a41316a <=( a41315a  and  a41308a );
 a41320a <=( (not A167)  and  (not A169) );
 a41321a <=( A170  and  a41320a );
 a41325a <=( (not A201)  and  (not A200) );
 a41326a <=( A166  and  a41325a );
 a41327a <=( a41326a  and  a41321a );
 a41331a <=( A234  and  (not A233) );
 a41332a <=( A232  and  a41331a );
 a41335a <=( A298  and  A235 );
 a41338a <=( (not A302)  and  (not A301) );
 a41339a <=( a41338a  and  a41335a );
 a41340a <=( a41339a  and  a41332a );
 a41344a <=( (not A167)  and  (not A169) );
 a41345a <=( A170  and  a41344a );
 a41349a <=( (not A201)  and  (not A200) );
 a41350a <=( A166  and  a41349a );
 a41351a <=( a41350a  and  a41345a );
 a41355a <=( A234  and  (not A233) );
 a41356a <=( A232  and  a41355a );
 a41359a <=( A298  and  A236 );
 a41362a <=( (not A302)  and  (not A301) );
 a41363a <=( a41362a  and  a41359a );
 a41364a <=( a41363a  and  a41356a );
 a41368a <=( (not A167)  and  (not A169) );
 a41369a <=( A170  and  a41368a );
 a41373a <=( (not A201)  and  (not A200) );
 a41374a <=( A166  and  a41373a );
 a41375a <=( a41374a  and  a41369a );
 a41379a <=( (not A266)  and  (not A233) );
 a41380a <=( (not A232)  and  a41379a );
 a41383a <=( (not A269)  and  (not A268) );
 a41386a <=( A299  and  (not A298) );
 a41387a <=( a41386a  and  a41383a );
 a41388a <=( a41387a  and  a41380a );
 a41392a <=( (not A167)  and  (not A169) );
 a41393a <=( A170  and  a41392a );
 a41397a <=( (not A200)  and  (not A199) );
 a41398a <=( A166  and  a41397a );
 a41399a <=( a41398a  and  a41393a );
 a41403a <=( A265  and  A233 );
 a41404a <=( A232  and  a41403a );
 a41407a <=( (not A269)  and  (not A268) );
 a41410a <=( A299  and  (not A298) );
 a41411a <=( a41410a  and  a41407a );
 a41412a <=( a41411a  and  a41404a );
 a41416a <=( (not A167)  and  (not A169) );
 a41417a <=( A170  and  a41416a );
 a41421a <=( (not A200)  and  (not A199) );
 a41422a <=( A166  and  a41421a );
 a41423a <=( a41422a  and  a41417a );
 a41427a <=( (not A236)  and  (not A235) );
 a41428a <=( (not A233)  and  a41427a );
 a41431a <=( A266  and  A265 );
 a41434a <=( A299  and  (not A298) );
 a41435a <=( a41434a  and  a41431a );
 a41436a <=( a41435a  and  a41428a );
 a41440a <=( (not A167)  and  (not A169) );
 a41441a <=( A170  and  a41440a );
 a41445a <=( (not A200)  and  (not A199) );
 a41446a <=( A166  and  a41445a );
 a41447a <=( a41446a  and  a41441a );
 a41451a <=( (not A236)  and  (not A235) );
 a41452a <=( (not A233)  and  a41451a );
 a41455a <=( (not A267)  and  (not A266) );
 a41458a <=( A299  and  (not A298) );
 a41459a <=( a41458a  and  a41455a );
 a41460a <=( a41459a  and  a41452a );
 a41464a <=( (not A167)  and  (not A169) );
 a41465a <=( A170  and  a41464a );
 a41469a <=( (not A200)  and  (not A199) );
 a41470a <=( A166  and  a41469a );
 a41471a <=( a41470a  and  a41465a );
 a41475a <=( (not A236)  and  (not A235) );
 a41476a <=( (not A233)  and  a41475a );
 a41479a <=( (not A266)  and  (not A265) );
 a41482a <=( A299  and  (not A298) );
 a41483a <=( a41482a  and  a41479a );
 a41484a <=( a41483a  and  a41476a );
 a41488a <=( (not A167)  and  (not A169) );
 a41489a <=( A170  and  a41488a );
 a41493a <=( (not A200)  and  (not A199) );
 a41494a <=( A166  and  a41493a );
 a41495a <=( a41494a  and  a41489a );
 a41499a <=( (not A266)  and  (not A234) );
 a41500a <=( (not A233)  and  a41499a );
 a41503a <=( (not A269)  and  (not A268) );
 a41506a <=( A299  and  (not A298) );
 a41507a <=( a41506a  and  a41503a );
 a41508a <=( a41507a  and  a41500a );
 a41512a <=( (not A167)  and  (not A169) );
 a41513a <=( A170  and  a41512a );
 a41517a <=( (not A200)  and  (not A199) );
 a41518a <=( A166  and  a41517a );
 a41519a <=( a41518a  and  a41513a );
 a41523a <=( A234  and  (not A233) );
 a41524a <=( A232  and  a41523a );
 a41527a <=( A298  and  A235 );
 a41530a <=( (not A302)  and  (not A301) );
 a41531a <=( a41530a  and  a41527a );
 a41532a <=( a41531a  and  a41524a );
 a41536a <=( (not A167)  and  (not A169) );
 a41537a <=( A170  and  a41536a );
 a41541a <=( (not A200)  and  (not A199) );
 a41542a <=( A166  and  a41541a );
 a41543a <=( a41542a  and  a41537a );
 a41547a <=( A234  and  (not A233) );
 a41548a <=( A232  and  a41547a );
 a41551a <=( A298  and  A236 );
 a41554a <=( (not A302)  and  (not A301) );
 a41555a <=( a41554a  and  a41551a );
 a41556a <=( a41555a  and  a41548a );
 a41560a <=( (not A167)  and  (not A169) );
 a41561a <=( A170  and  a41560a );
 a41565a <=( (not A200)  and  (not A199) );
 a41566a <=( A166  and  a41565a );
 a41567a <=( a41566a  and  a41561a );
 a41571a <=( (not A266)  and  (not A233) );
 a41572a <=( (not A232)  and  a41571a );
 a41575a <=( (not A269)  and  (not A268) );
 a41578a <=( A299  and  (not A298) );
 a41579a <=( a41578a  and  a41575a );
 a41580a <=( a41579a  and  a41572a );
 a41584a <=( (not A168)  and  (not A169) );
 a41585a <=( (not A170)  and  a41584a );
 a41589a <=( A201  and  (not A200) );
 a41590a <=( A199  and  a41589a );
 a41591a <=( a41590a  and  a41585a );
 a41595a <=( A233  and  A232 );
 a41596a <=( A202  and  a41595a );
 a41599a <=( (not A267)  and  A265 );
 a41602a <=( A299  and  (not A298) );
 a41603a <=( a41602a  and  a41599a );
 a41604a <=( a41603a  and  a41596a );
 a41608a <=( (not A168)  and  (not A169) );
 a41609a <=( (not A170)  and  a41608a );
 a41613a <=( A201  and  (not A200) );
 a41614a <=( A199  and  a41613a );
 a41615a <=( a41614a  and  a41609a );
 a41619a <=( A233  and  A232 );
 a41620a <=( A202  and  a41619a );
 a41623a <=( A266  and  A265 );
 a41626a <=( A299  and  (not A298) );
 a41627a <=( a41626a  and  a41623a );
 a41628a <=( a41627a  and  a41620a );
 a41632a <=( (not A168)  and  (not A169) );
 a41633a <=( (not A170)  and  a41632a );
 a41637a <=( A201  and  (not A200) );
 a41638a <=( A199  and  a41637a );
 a41639a <=( a41638a  and  a41633a );
 a41643a <=( A233  and  A232 );
 a41644a <=( A202  and  a41643a );
 a41647a <=( (not A266)  and  (not A265) );
 a41650a <=( A299  and  (not A298) );
 a41651a <=( a41650a  and  a41647a );
 a41652a <=( a41651a  and  a41644a );
 a41656a <=( (not A168)  and  (not A169) );
 a41657a <=( (not A170)  and  a41656a );
 a41661a <=( A201  and  (not A200) );
 a41662a <=( A199  and  a41661a );
 a41663a <=( a41662a  and  a41657a );
 a41667a <=( A233  and  (not A232) );
 a41668a <=( A202  and  a41667a );
 a41671a <=( (not A266)  and  A265 );
 a41674a <=( A268  and  A267 );
 a41675a <=( a41674a  and  a41671a );
 a41676a <=( a41675a  and  a41668a );
 a41680a <=( (not A168)  and  (not A169) );
 a41681a <=( (not A170)  and  a41680a );
 a41685a <=( A201  and  (not A200) );
 a41686a <=( A199  and  a41685a );
 a41687a <=( a41686a  and  a41681a );
 a41691a <=( A233  and  (not A232) );
 a41692a <=( A202  and  a41691a );
 a41695a <=( (not A266)  and  A265 );
 a41698a <=( A269  and  A267 );
 a41699a <=( a41698a  and  a41695a );
 a41700a <=( a41699a  and  a41692a );
 a41704a <=( (not A168)  and  (not A169) );
 a41705a <=( (not A170)  and  a41704a );
 a41709a <=( A201  and  (not A200) );
 a41710a <=( A199  and  a41709a );
 a41711a <=( a41710a  and  a41705a );
 a41715a <=( (not A234)  and  (not A233) );
 a41716a <=( A202  and  a41715a );
 a41719a <=( A266  and  A265 );
 a41722a <=( A299  and  (not A298) );
 a41723a <=( a41722a  and  a41719a );
 a41724a <=( a41723a  and  a41716a );
 a41728a <=( (not A168)  and  (not A169) );
 a41729a <=( (not A170)  and  a41728a );
 a41733a <=( A201  and  (not A200) );
 a41734a <=( A199  and  a41733a );
 a41735a <=( a41734a  and  a41729a );
 a41739a <=( (not A234)  and  (not A233) );
 a41740a <=( A202  and  a41739a );
 a41743a <=( (not A267)  and  (not A266) );
 a41746a <=( A299  and  (not A298) );
 a41747a <=( a41746a  and  a41743a );
 a41748a <=( a41747a  and  a41740a );
 a41752a <=( (not A168)  and  (not A169) );
 a41753a <=( (not A170)  and  a41752a );
 a41757a <=( A201  and  (not A200) );
 a41758a <=( A199  and  a41757a );
 a41759a <=( a41758a  and  a41753a );
 a41763a <=( (not A234)  and  (not A233) );
 a41764a <=( A202  and  a41763a );
 a41767a <=( (not A266)  and  (not A265) );
 a41770a <=( A299  and  (not A298) );
 a41771a <=( a41770a  and  a41767a );
 a41772a <=( a41771a  and  a41764a );
 a41776a <=( (not A168)  and  (not A169) );
 a41777a <=( (not A170)  and  a41776a );
 a41781a <=( A201  and  (not A200) );
 a41782a <=( A199  and  a41781a );
 a41783a <=( a41782a  and  a41777a );
 a41787a <=( (not A233)  and  A232 );
 a41788a <=( A202  and  a41787a );
 a41791a <=( A235  and  A234 );
 a41794a <=( (not A300)  and  A298 );
 a41795a <=( a41794a  and  a41791a );
 a41796a <=( a41795a  and  a41788a );
 a41800a <=( (not A168)  and  (not A169) );
 a41801a <=( (not A170)  and  a41800a );
 a41805a <=( A201  and  (not A200) );
 a41806a <=( A199  and  a41805a );
 a41807a <=( a41806a  and  a41801a );
 a41811a <=( (not A233)  and  A232 );
 a41812a <=( A202  and  a41811a );
 a41815a <=( A235  and  A234 );
 a41818a <=( A299  and  A298 );
 a41819a <=( a41818a  and  a41815a );
 a41820a <=( a41819a  and  a41812a );
 a41824a <=( (not A168)  and  (not A169) );
 a41825a <=( (not A170)  and  a41824a );
 a41829a <=( A201  and  (not A200) );
 a41830a <=( A199  and  a41829a );
 a41831a <=( a41830a  and  a41825a );
 a41835a <=( (not A233)  and  A232 );
 a41836a <=( A202  and  a41835a );
 a41839a <=( A235  and  A234 );
 a41842a <=( (not A299)  and  (not A298) );
 a41843a <=( a41842a  and  a41839a );
 a41844a <=( a41843a  and  a41836a );
 a41848a <=( (not A168)  and  (not A169) );
 a41849a <=( (not A170)  and  a41848a );
 a41853a <=( A201  and  (not A200) );
 a41854a <=( A199  and  a41853a );
 a41855a <=( a41854a  and  a41849a );
 a41859a <=( (not A233)  and  A232 );
 a41860a <=( A202  and  a41859a );
 a41863a <=( A235  and  A234 );
 a41866a <=( A266  and  (not A265) );
 a41867a <=( a41866a  and  a41863a );
 a41868a <=( a41867a  and  a41860a );
 a41872a <=( (not A168)  and  (not A169) );
 a41873a <=( (not A170)  and  a41872a );
 a41877a <=( A201  and  (not A200) );
 a41878a <=( A199  and  a41877a );
 a41879a <=( a41878a  and  a41873a );
 a41883a <=( (not A233)  and  A232 );
 a41884a <=( A202  and  a41883a );
 a41887a <=( A236  and  A234 );
 a41890a <=( (not A300)  and  A298 );
 a41891a <=( a41890a  and  a41887a );
 a41892a <=( a41891a  and  a41884a );
 a41896a <=( (not A168)  and  (not A169) );
 a41897a <=( (not A170)  and  a41896a );
 a41901a <=( A201  and  (not A200) );
 a41902a <=( A199  and  a41901a );
 a41903a <=( a41902a  and  a41897a );
 a41907a <=( (not A233)  and  A232 );
 a41908a <=( A202  and  a41907a );
 a41911a <=( A236  and  A234 );
 a41914a <=( A299  and  A298 );
 a41915a <=( a41914a  and  a41911a );
 a41916a <=( a41915a  and  a41908a );
 a41920a <=( (not A168)  and  (not A169) );
 a41921a <=( (not A170)  and  a41920a );
 a41925a <=( A201  and  (not A200) );
 a41926a <=( A199  and  a41925a );
 a41927a <=( a41926a  and  a41921a );
 a41931a <=( (not A233)  and  A232 );
 a41932a <=( A202  and  a41931a );
 a41935a <=( A236  and  A234 );
 a41938a <=( (not A299)  and  (not A298) );
 a41939a <=( a41938a  and  a41935a );
 a41940a <=( a41939a  and  a41932a );
 a41944a <=( (not A168)  and  (not A169) );
 a41945a <=( (not A170)  and  a41944a );
 a41949a <=( A201  and  (not A200) );
 a41950a <=( A199  and  a41949a );
 a41951a <=( a41950a  and  a41945a );
 a41955a <=( (not A233)  and  A232 );
 a41956a <=( A202  and  a41955a );
 a41959a <=( A236  and  A234 );
 a41962a <=( A266  and  (not A265) );
 a41963a <=( a41962a  and  a41959a );
 a41964a <=( a41963a  and  a41956a );
 a41968a <=( (not A168)  and  (not A169) );
 a41969a <=( (not A170)  and  a41968a );
 a41973a <=( A201  and  (not A200) );
 a41974a <=( A199  and  a41973a );
 a41975a <=( a41974a  and  a41969a );
 a41979a <=( (not A233)  and  (not A232) );
 a41980a <=( A202  and  a41979a );
 a41983a <=( A266  and  A265 );
 a41986a <=( A299  and  (not A298) );
 a41987a <=( a41986a  and  a41983a );
 a41988a <=( a41987a  and  a41980a );
 a41992a <=( (not A168)  and  (not A169) );
 a41993a <=( (not A170)  and  a41992a );
 a41997a <=( A201  and  (not A200) );
 a41998a <=( A199  and  a41997a );
 a41999a <=( a41998a  and  a41993a );
 a42003a <=( (not A233)  and  (not A232) );
 a42004a <=( A202  and  a42003a );
 a42007a <=( (not A267)  and  (not A266) );
 a42010a <=( A299  and  (not A298) );
 a42011a <=( a42010a  and  a42007a );
 a42012a <=( a42011a  and  a42004a );
 a42016a <=( (not A168)  and  (not A169) );
 a42017a <=( (not A170)  and  a42016a );
 a42021a <=( A201  and  (not A200) );
 a42022a <=( A199  and  a42021a );
 a42023a <=( a42022a  and  a42017a );
 a42027a <=( (not A233)  and  (not A232) );
 a42028a <=( A202  and  a42027a );
 a42031a <=( (not A266)  and  (not A265) );
 a42034a <=( A299  and  (not A298) );
 a42035a <=( a42034a  and  a42031a );
 a42036a <=( a42035a  and  a42028a );
 a42040a <=( (not A168)  and  (not A169) );
 a42041a <=( (not A170)  and  a42040a );
 a42045a <=( A201  and  (not A200) );
 a42046a <=( A199  and  a42045a );
 a42047a <=( a42046a  and  a42041a );
 a42051a <=( A233  and  A232 );
 a42052a <=( A203  and  a42051a );
 a42055a <=( (not A267)  and  A265 );
 a42058a <=( A299  and  (not A298) );
 a42059a <=( a42058a  and  a42055a );
 a42060a <=( a42059a  and  a42052a );
 a42064a <=( (not A168)  and  (not A169) );
 a42065a <=( (not A170)  and  a42064a );
 a42069a <=( A201  and  (not A200) );
 a42070a <=( A199  and  a42069a );
 a42071a <=( a42070a  and  a42065a );
 a42075a <=( A233  and  A232 );
 a42076a <=( A203  and  a42075a );
 a42079a <=( A266  and  A265 );
 a42082a <=( A299  and  (not A298) );
 a42083a <=( a42082a  and  a42079a );
 a42084a <=( a42083a  and  a42076a );
 a42088a <=( (not A168)  and  (not A169) );
 a42089a <=( (not A170)  and  a42088a );
 a42093a <=( A201  and  (not A200) );
 a42094a <=( A199  and  a42093a );
 a42095a <=( a42094a  and  a42089a );
 a42099a <=( A233  and  A232 );
 a42100a <=( A203  and  a42099a );
 a42103a <=( (not A266)  and  (not A265) );
 a42106a <=( A299  and  (not A298) );
 a42107a <=( a42106a  and  a42103a );
 a42108a <=( a42107a  and  a42100a );
 a42112a <=( (not A168)  and  (not A169) );
 a42113a <=( (not A170)  and  a42112a );
 a42117a <=( A201  and  (not A200) );
 a42118a <=( A199  and  a42117a );
 a42119a <=( a42118a  and  a42113a );
 a42123a <=( A233  and  (not A232) );
 a42124a <=( A203  and  a42123a );
 a42127a <=( (not A266)  and  A265 );
 a42130a <=( A268  and  A267 );
 a42131a <=( a42130a  and  a42127a );
 a42132a <=( a42131a  and  a42124a );
 a42136a <=( (not A168)  and  (not A169) );
 a42137a <=( (not A170)  and  a42136a );
 a42141a <=( A201  and  (not A200) );
 a42142a <=( A199  and  a42141a );
 a42143a <=( a42142a  and  a42137a );
 a42147a <=( A233  and  (not A232) );
 a42148a <=( A203  and  a42147a );
 a42151a <=( (not A266)  and  A265 );
 a42154a <=( A269  and  A267 );
 a42155a <=( a42154a  and  a42151a );
 a42156a <=( a42155a  and  a42148a );
 a42160a <=( (not A168)  and  (not A169) );
 a42161a <=( (not A170)  and  a42160a );
 a42165a <=( A201  and  (not A200) );
 a42166a <=( A199  and  a42165a );
 a42167a <=( a42166a  and  a42161a );
 a42171a <=( (not A234)  and  (not A233) );
 a42172a <=( A203  and  a42171a );
 a42175a <=( A266  and  A265 );
 a42178a <=( A299  and  (not A298) );
 a42179a <=( a42178a  and  a42175a );
 a42180a <=( a42179a  and  a42172a );
 a42184a <=( (not A168)  and  (not A169) );
 a42185a <=( (not A170)  and  a42184a );
 a42189a <=( A201  and  (not A200) );
 a42190a <=( A199  and  a42189a );
 a42191a <=( a42190a  and  a42185a );
 a42195a <=( (not A234)  and  (not A233) );
 a42196a <=( A203  and  a42195a );
 a42199a <=( (not A267)  and  (not A266) );
 a42202a <=( A299  and  (not A298) );
 a42203a <=( a42202a  and  a42199a );
 a42204a <=( a42203a  and  a42196a );
 a42208a <=( (not A168)  and  (not A169) );
 a42209a <=( (not A170)  and  a42208a );
 a42213a <=( A201  and  (not A200) );
 a42214a <=( A199  and  a42213a );
 a42215a <=( a42214a  and  a42209a );
 a42219a <=( (not A234)  and  (not A233) );
 a42220a <=( A203  and  a42219a );
 a42223a <=( (not A266)  and  (not A265) );
 a42226a <=( A299  and  (not A298) );
 a42227a <=( a42226a  and  a42223a );
 a42228a <=( a42227a  and  a42220a );
 a42232a <=( (not A168)  and  (not A169) );
 a42233a <=( (not A170)  and  a42232a );
 a42237a <=( A201  and  (not A200) );
 a42238a <=( A199  and  a42237a );
 a42239a <=( a42238a  and  a42233a );
 a42243a <=( (not A233)  and  A232 );
 a42244a <=( A203  and  a42243a );
 a42247a <=( A235  and  A234 );
 a42250a <=( (not A300)  and  A298 );
 a42251a <=( a42250a  and  a42247a );
 a42252a <=( a42251a  and  a42244a );
 a42256a <=( (not A168)  and  (not A169) );
 a42257a <=( (not A170)  and  a42256a );
 a42261a <=( A201  and  (not A200) );
 a42262a <=( A199  and  a42261a );
 a42263a <=( a42262a  and  a42257a );
 a42267a <=( (not A233)  and  A232 );
 a42268a <=( A203  and  a42267a );
 a42271a <=( A235  and  A234 );
 a42274a <=( A299  and  A298 );
 a42275a <=( a42274a  and  a42271a );
 a42276a <=( a42275a  and  a42268a );
 a42280a <=( (not A168)  and  (not A169) );
 a42281a <=( (not A170)  and  a42280a );
 a42285a <=( A201  and  (not A200) );
 a42286a <=( A199  and  a42285a );
 a42287a <=( a42286a  and  a42281a );
 a42291a <=( (not A233)  and  A232 );
 a42292a <=( A203  and  a42291a );
 a42295a <=( A235  and  A234 );
 a42298a <=( (not A299)  and  (not A298) );
 a42299a <=( a42298a  and  a42295a );
 a42300a <=( a42299a  and  a42292a );
 a42304a <=( (not A168)  and  (not A169) );
 a42305a <=( (not A170)  and  a42304a );
 a42309a <=( A201  and  (not A200) );
 a42310a <=( A199  and  a42309a );
 a42311a <=( a42310a  and  a42305a );
 a42315a <=( (not A233)  and  A232 );
 a42316a <=( A203  and  a42315a );
 a42319a <=( A235  and  A234 );
 a42322a <=( A266  and  (not A265) );
 a42323a <=( a42322a  and  a42319a );
 a42324a <=( a42323a  and  a42316a );
 a42328a <=( (not A168)  and  (not A169) );
 a42329a <=( (not A170)  and  a42328a );
 a42333a <=( A201  and  (not A200) );
 a42334a <=( A199  and  a42333a );
 a42335a <=( a42334a  and  a42329a );
 a42339a <=( (not A233)  and  A232 );
 a42340a <=( A203  and  a42339a );
 a42343a <=( A236  and  A234 );
 a42346a <=( (not A300)  and  A298 );
 a42347a <=( a42346a  and  a42343a );
 a42348a <=( a42347a  and  a42340a );
 a42352a <=( (not A168)  and  (not A169) );
 a42353a <=( (not A170)  and  a42352a );
 a42357a <=( A201  and  (not A200) );
 a42358a <=( A199  and  a42357a );
 a42359a <=( a42358a  and  a42353a );
 a42363a <=( (not A233)  and  A232 );
 a42364a <=( A203  and  a42363a );
 a42367a <=( A236  and  A234 );
 a42370a <=( A299  and  A298 );
 a42371a <=( a42370a  and  a42367a );
 a42372a <=( a42371a  and  a42364a );
 a42376a <=( (not A168)  and  (not A169) );
 a42377a <=( (not A170)  and  a42376a );
 a42381a <=( A201  and  (not A200) );
 a42382a <=( A199  and  a42381a );
 a42383a <=( a42382a  and  a42377a );
 a42387a <=( (not A233)  and  A232 );
 a42388a <=( A203  and  a42387a );
 a42391a <=( A236  and  A234 );
 a42394a <=( (not A299)  and  (not A298) );
 a42395a <=( a42394a  and  a42391a );
 a42396a <=( a42395a  and  a42388a );
 a42400a <=( (not A168)  and  (not A169) );
 a42401a <=( (not A170)  and  a42400a );
 a42405a <=( A201  and  (not A200) );
 a42406a <=( A199  and  a42405a );
 a42407a <=( a42406a  and  a42401a );
 a42411a <=( (not A233)  and  A232 );
 a42412a <=( A203  and  a42411a );
 a42415a <=( A236  and  A234 );
 a42418a <=( A266  and  (not A265) );
 a42419a <=( a42418a  and  a42415a );
 a42420a <=( a42419a  and  a42412a );
 a42424a <=( (not A168)  and  (not A169) );
 a42425a <=( (not A170)  and  a42424a );
 a42429a <=( A201  and  (not A200) );
 a42430a <=( A199  and  a42429a );
 a42431a <=( a42430a  and  a42425a );
 a42435a <=( (not A233)  and  (not A232) );
 a42436a <=( A203  and  a42435a );
 a42439a <=( A266  and  A265 );
 a42442a <=( A299  and  (not A298) );
 a42443a <=( a42442a  and  a42439a );
 a42444a <=( a42443a  and  a42436a );
 a42448a <=( (not A168)  and  (not A169) );
 a42449a <=( (not A170)  and  a42448a );
 a42453a <=( A201  and  (not A200) );
 a42454a <=( A199  and  a42453a );
 a42455a <=( a42454a  and  a42449a );
 a42459a <=( (not A233)  and  (not A232) );
 a42460a <=( A203  and  a42459a );
 a42463a <=( (not A267)  and  (not A266) );
 a42466a <=( A299  and  (not A298) );
 a42467a <=( a42466a  and  a42463a );
 a42468a <=( a42467a  and  a42460a );
 a42472a <=( (not A168)  and  (not A169) );
 a42473a <=( (not A170)  and  a42472a );
 a42477a <=( A201  and  (not A200) );
 a42478a <=( A199  and  a42477a );
 a42479a <=( a42478a  and  a42473a );
 a42483a <=( (not A233)  and  (not A232) );
 a42484a <=( A203  and  a42483a );
 a42487a <=( (not A266)  and  (not A265) );
 a42490a <=( A299  and  (not A298) );
 a42491a <=( a42490a  and  a42487a );
 a42492a <=( a42491a  and  a42484a );
 a42496a <=( A199  and  A166 );
 a42497a <=( A168  and  a42496a );
 a42500a <=( (not A233)  and  A200 );
 a42503a <=( (not A236)  and  (not A235) );
 a42504a <=( a42503a  and  a42500a );
 a42505a <=( a42504a  and  a42497a );
 a42509a <=( (not A269)  and  (not A268) );
 a42510a <=( (not A266)  and  a42509a );
 a42513a <=( (not A299)  and  A298 );
 a42516a <=( A301  and  A300 );
 a42517a <=( a42516a  and  a42513a );
 a42518a <=( a42517a  and  a42510a );
 a42522a <=( A199  and  A166 );
 a42523a <=( A168  and  a42522a );
 a42526a <=( (not A233)  and  A200 );
 a42529a <=( (not A236)  and  (not A235) );
 a42530a <=( a42529a  and  a42526a );
 a42531a <=( a42530a  and  a42523a );
 a42535a <=( (not A269)  and  (not A268) );
 a42536a <=( (not A266)  and  a42535a );
 a42539a <=( (not A299)  and  A298 );
 a42542a <=( A302  and  A300 );
 a42543a <=( a42542a  and  a42539a );
 a42544a <=( a42543a  and  a42536a );
 a42548a <=( (not A200)  and  A166 );
 a42549a <=( A168  and  a42548a );
 a42552a <=( (not A203)  and  (not A202) );
 a42555a <=( A233  and  A232 );
 a42556a <=( a42555a  and  a42552a );
 a42557a <=( a42556a  and  a42549a );
 a42561a <=( (not A269)  and  (not A268) );
 a42562a <=( A265  and  a42561a );
 a42565a <=( (not A299)  and  A298 );
 a42568a <=( A301  and  A300 );
 a42569a <=( a42568a  and  a42565a );
 a42570a <=( a42569a  and  a42562a );
 a42574a <=( (not A200)  and  A166 );
 a42575a <=( A168  and  a42574a );
 a42578a <=( (not A203)  and  (not A202) );
 a42581a <=( A233  and  A232 );
 a42582a <=( a42581a  and  a42578a );
 a42583a <=( a42582a  and  a42575a );
 a42587a <=( (not A269)  and  (not A268) );
 a42588a <=( A265  and  a42587a );
 a42591a <=( (not A299)  and  A298 );
 a42594a <=( A302  and  A300 );
 a42595a <=( a42594a  and  a42591a );
 a42596a <=( a42595a  and  a42588a );
 a42600a <=( (not A200)  and  A166 );
 a42601a <=( A168  and  a42600a );
 a42604a <=( (not A203)  and  (not A202) );
 a42607a <=( (not A235)  and  (not A233) );
 a42608a <=( a42607a  and  a42604a );
 a42609a <=( a42608a  and  a42601a );
 a42613a <=( A266  and  A265 );
 a42614a <=( (not A236)  and  a42613a );
 a42617a <=( (not A299)  and  A298 );
 a42620a <=( A301  and  A300 );
 a42621a <=( a42620a  and  a42617a );
 a42622a <=( a42621a  and  a42614a );
 a42626a <=( (not A200)  and  A166 );
 a42627a <=( A168  and  a42626a );
 a42630a <=( (not A203)  and  (not A202) );
 a42633a <=( (not A235)  and  (not A233) );
 a42634a <=( a42633a  and  a42630a );
 a42635a <=( a42634a  and  a42627a );
 a42639a <=( A266  and  A265 );
 a42640a <=( (not A236)  and  a42639a );
 a42643a <=( (not A299)  and  A298 );
 a42646a <=( A302  and  A300 );
 a42647a <=( a42646a  and  a42643a );
 a42648a <=( a42647a  and  a42640a );
 a42652a <=( (not A200)  and  A166 );
 a42653a <=( A168  and  a42652a );
 a42656a <=( (not A203)  and  (not A202) );
 a42659a <=( (not A235)  and  (not A233) );
 a42660a <=( a42659a  and  a42656a );
 a42661a <=( a42660a  and  a42653a );
 a42665a <=( (not A267)  and  (not A266) );
 a42666a <=( (not A236)  and  a42665a );
 a42669a <=( (not A299)  and  A298 );
 a42672a <=( A301  and  A300 );
 a42673a <=( a42672a  and  a42669a );
 a42674a <=( a42673a  and  a42666a );
 a42678a <=( (not A200)  and  A166 );
 a42679a <=( A168  and  a42678a );
 a42682a <=( (not A203)  and  (not A202) );
 a42685a <=( (not A235)  and  (not A233) );
 a42686a <=( a42685a  and  a42682a );
 a42687a <=( a42686a  and  a42679a );
 a42691a <=( (not A267)  and  (not A266) );
 a42692a <=( (not A236)  and  a42691a );
 a42695a <=( (not A299)  and  A298 );
 a42698a <=( A302  and  A300 );
 a42699a <=( a42698a  and  a42695a );
 a42700a <=( a42699a  and  a42692a );
 a42704a <=( (not A200)  and  A166 );
 a42705a <=( A168  and  a42704a );
 a42708a <=( (not A203)  and  (not A202) );
 a42711a <=( (not A235)  and  (not A233) );
 a42712a <=( a42711a  and  a42708a );
 a42713a <=( a42712a  and  a42705a );
 a42717a <=( (not A266)  and  (not A265) );
 a42718a <=( (not A236)  and  a42717a );
 a42721a <=( (not A299)  and  A298 );
 a42724a <=( A301  and  A300 );
 a42725a <=( a42724a  and  a42721a );
 a42726a <=( a42725a  and  a42718a );
 a42730a <=( (not A200)  and  A166 );
 a42731a <=( A168  and  a42730a );
 a42734a <=( (not A203)  and  (not A202) );
 a42737a <=( (not A235)  and  (not A233) );
 a42738a <=( a42737a  and  a42734a );
 a42739a <=( a42738a  and  a42731a );
 a42743a <=( (not A266)  and  (not A265) );
 a42744a <=( (not A236)  and  a42743a );
 a42747a <=( (not A299)  and  A298 );
 a42750a <=( A302  and  A300 );
 a42751a <=( a42750a  and  a42747a );
 a42752a <=( a42751a  and  a42744a );
 a42756a <=( (not A200)  and  A166 );
 a42757a <=( A168  and  a42756a );
 a42760a <=( (not A203)  and  (not A202) );
 a42763a <=( (not A234)  and  (not A233) );
 a42764a <=( a42763a  and  a42760a );
 a42765a <=( a42764a  and  a42757a );
 a42769a <=( (not A269)  and  (not A268) );
 a42770a <=( (not A266)  and  a42769a );
 a42773a <=( (not A299)  and  A298 );
 a42776a <=( A301  and  A300 );
 a42777a <=( a42776a  and  a42773a );
 a42778a <=( a42777a  and  a42770a );
 a42782a <=( (not A200)  and  A166 );
 a42783a <=( A168  and  a42782a );
 a42786a <=( (not A203)  and  (not A202) );
 a42789a <=( (not A234)  and  (not A233) );
 a42790a <=( a42789a  and  a42786a );
 a42791a <=( a42790a  and  a42783a );
 a42795a <=( (not A269)  and  (not A268) );
 a42796a <=( (not A266)  and  a42795a );
 a42799a <=( (not A299)  and  A298 );
 a42802a <=( A302  and  A300 );
 a42803a <=( a42802a  and  a42799a );
 a42804a <=( a42803a  and  a42796a );
 a42808a <=( (not A200)  and  A166 );
 a42809a <=( A168  and  a42808a );
 a42812a <=( (not A203)  and  (not A202) );
 a42815a <=( (not A233)  and  (not A232) );
 a42816a <=( a42815a  and  a42812a );
 a42817a <=( a42816a  and  a42809a );
 a42821a <=( (not A269)  and  (not A268) );
 a42822a <=( (not A266)  and  a42821a );
 a42825a <=( (not A299)  and  A298 );
 a42828a <=( A301  and  A300 );
 a42829a <=( a42828a  and  a42825a );
 a42830a <=( a42829a  and  a42822a );
 a42834a <=( (not A200)  and  A166 );
 a42835a <=( A168  and  a42834a );
 a42838a <=( (not A203)  and  (not A202) );
 a42841a <=( (not A233)  and  (not A232) );
 a42842a <=( a42841a  and  a42838a );
 a42843a <=( a42842a  and  a42835a );
 a42847a <=( (not A269)  and  (not A268) );
 a42848a <=( (not A266)  and  a42847a );
 a42851a <=( (not A299)  and  A298 );
 a42854a <=( A302  and  A300 );
 a42855a <=( a42854a  and  a42851a );
 a42856a <=( a42855a  and  a42848a );
 a42860a <=( (not A200)  and  A166 );
 a42861a <=( A168  and  a42860a );
 a42864a <=( (not A233)  and  (not A201) );
 a42867a <=( (not A236)  and  (not A235) );
 a42868a <=( a42867a  and  a42864a );
 a42869a <=( a42868a  and  a42861a );
 a42873a <=( (not A269)  and  (not A268) );
 a42874a <=( (not A266)  and  a42873a );
 a42877a <=( (not A299)  and  A298 );
 a42880a <=( A301  and  A300 );
 a42881a <=( a42880a  and  a42877a );
 a42882a <=( a42881a  and  a42874a );
 a42886a <=( (not A200)  and  A166 );
 a42887a <=( A168  and  a42886a );
 a42890a <=( (not A233)  and  (not A201) );
 a42893a <=( (not A236)  and  (not A235) );
 a42894a <=( a42893a  and  a42890a );
 a42895a <=( a42894a  and  a42887a );
 a42899a <=( (not A269)  and  (not A268) );
 a42900a <=( (not A266)  and  a42899a );
 a42903a <=( (not A299)  and  A298 );
 a42906a <=( A302  and  A300 );
 a42907a <=( a42906a  and  a42903a );
 a42908a <=( a42907a  and  a42900a );
 a42912a <=( (not A199)  and  A166 );
 a42913a <=( A168  and  a42912a );
 a42916a <=( (not A233)  and  (not A200) );
 a42919a <=( (not A236)  and  (not A235) );
 a42920a <=( a42919a  and  a42916a );
 a42921a <=( a42920a  and  a42913a );
 a42925a <=( (not A269)  and  (not A268) );
 a42926a <=( (not A266)  and  a42925a );
 a42929a <=( (not A299)  and  A298 );
 a42932a <=( A301  and  A300 );
 a42933a <=( a42932a  and  a42929a );
 a42934a <=( a42933a  and  a42926a );
 a42938a <=( (not A199)  and  A166 );
 a42939a <=( A168  and  a42938a );
 a42942a <=( (not A233)  and  (not A200) );
 a42945a <=( (not A236)  and  (not A235) );
 a42946a <=( a42945a  and  a42942a );
 a42947a <=( a42946a  and  a42939a );
 a42951a <=( (not A269)  and  (not A268) );
 a42952a <=( (not A266)  and  a42951a );
 a42955a <=( (not A299)  and  A298 );
 a42958a <=( A302  and  A300 );
 a42959a <=( a42958a  and  a42955a );
 a42960a <=( a42959a  and  a42952a );
 a42964a <=( A199  and  A167 );
 a42965a <=( A168  and  a42964a );
 a42968a <=( (not A233)  and  A200 );
 a42971a <=( (not A236)  and  (not A235) );
 a42972a <=( a42971a  and  a42968a );
 a42973a <=( a42972a  and  a42965a );
 a42977a <=( (not A269)  and  (not A268) );
 a42978a <=( (not A266)  and  a42977a );
 a42981a <=( (not A299)  and  A298 );
 a42984a <=( A301  and  A300 );
 a42985a <=( a42984a  and  a42981a );
 a42986a <=( a42985a  and  a42978a );
 a42990a <=( A199  and  A167 );
 a42991a <=( A168  and  a42990a );
 a42994a <=( (not A233)  and  A200 );
 a42997a <=( (not A236)  and  (not A235) );
 a42998a <=( a42997a  and  a42994a );
 a42999a <=( a42998a  and  a42991a );
 a43003a <=( (not A269)  and  (not A268) );
 a43004a <=( (not A266)  and  a43003a );
 a43007a <=( (not A299)  and  A298 );
 a43010a <=( A302  and  A300 );
 a43011a <=( a43010a  and  a43007a );
 a43012a <=( a43011a  and  a43004a );
 a43016a <=( (not A200)  and  A167 );
 a43017a <=( A168  and  a43016a );
 a43020a <=( (not A203)  and  (not A202) );
 a43023a <=( A233  and  A232 );
 a43024a <=( a43023a  and  a43020a );
 a43025a <=( a43024a  and  a43017a );
 a43029a <=( (not A269)  and  (not A268) );
 a43030a <=( A265  and  a43029a );
 a43033a <=( (not A299)  and  A298 );
 a43036a <=( A301  and  A300 );
 a43037a <=( a43036a  and  a43033a );
 a43038a <=( a43037a  and  a43030a );
 a43042a <=( (not A200)  and  A167 );
 a43043a <=( A168  and  a43042a );
 a43046a <=( (not A203)  and  (not A202) );
 a43049a <=( A233  and  A232 );
 a43050a <=( a43049a  and  a43046a );
 a43051a <=( a43050a  and  a43043a );
 a43055a <=( (not A269)  and  (not A268) );
 a43056a <=( A265  and  a43055a );
 a43059a <=( (not A299)  and  A298 );
 a43062a <=( A302  and  A300 );
 a43063a <=( a43062a  and  a43059a );
 a43064a <=( a43063a  and  a43056a );
 a43068a <=( (not A200)  and  A167 );
 a43069a <=( A168  and  a43068a );
 a43072a <=( (not A203)  and  (not A202) );
 a43075a <=( (not A235)  and  (not A233) );
 a43076a <=( a43075a  and  a43072a );
 a43077a <=( a43076a  and  a43069a );
 a43081a <=( A266  and  A265 );
 a43082a <=( (not A236)  and  a43081a );
 a43085a <=( (not A299)  and  A298 );
 a43088a <=( A301  and  A300 );
 a43089a <=( a43088a  and  a43085a );
 a43090a <=( a43089a  and  a43082a );
 a43094a <=( (not A200)  and  A167 );
 a43095a <=( A168  and  a43094a );
 a43098a <=( (not A203)  and  (not A202) );
 a43101a <=( (not A235)  and  (not A233) );
 a43102a <=( a43101a  and  a43098a );
 a43103a <=( a43102a  and  a43095a );
 a43107a <=( A266  and  A265 );
 a43108a <=( (not A236)  and  a43107a );
 a43111a <=( (not A299)  and  A298 );
 a43114a <=( A302  and  A300 );
 a43115a <=( a43114a  and  a43111a );
 a43116a <=( a43115a  and  a43108a );
 a43120a <=( (not A200)  and  A167 );
 a43121a <=( A168  and  a43120a );
 a43124a <=( (not A203)  and  (not A202) );
 a43127a <=( (not A235)  and  (not A233) );
 a43128a <=( a43127a  and  a43124a );
 a43129a <=( a43128a  and  a43121a );
 a43133a <=( (not A267)  and  (not A266) );
 a43134a <=( (not A236)  and  a43133a );
 a43137a <=( (not A299)  and  A298 );
 a43140a <=( A301  and  A300 );
 a43141a <=( a43140a  and  a43137a );
 a43142a <=( a43141a  and  a43134a );
 a43146a <=( (not A200)  and  A167 );
 a43147a <=( A168  and  a43146a );
 a43150a <=( (not A203)  and  (not A202) );
 a43153a <=( (not A235)  and  (not A233) );
 a43154a <=( a43153a  and  a43150a );
 a43155a <=( a43154a  and  a43147a );
 a43159a <=( (not A267)  and  (not A266) );
 a43160a <=( (not A236)  and  a43159a );
 a43163a <=( (not A299)  and  A298 );
 a43166a <=( A302  and  A300 );
 a43167a <=( a43166a  and  a43163a );
 a43168a <=( a43167a  and  a43160a );
 a43172a <=( (not A200)  and  A167 );
 a43173a <=( A168  and  a43172a );
 a43176a <=( (not A203)  and  (not A202) );
 a43179a <=( (not A235)  and  (not A233) );
 a43180a <=( a43179a  and  a43176a );
 a43181a <=( a43180a  and  a43173a );
 a43185a <=( (not A266)  and  (not A265) );
 a43186a <=( (not A236)  and  a43185a );
 a43189a <=( (not A299)  and  A298 );
 a43192a <=( A301  and  A300 );
 a43193a <=( a43192a  and  a43189a );
 a43194a <=( a43193a  and  a43186a );
 a43198a <=( (not A200)  and  A167 );
 a43199a <=( A168  and  a43198a );
 a43202a <=( (not A203)  and  (not A202) );
 a43205a <=( (not A235)  and  (not A233) );
 a43206a <=( a43205a  and  a43202a );
 a43207a <=( a43206a  and  a43199a );
 a43211a <=( (not A266)  and  (not A265) );
 a43212a <=( (not A236)  and  a43211a );
 a43215a <=( (not A299)  and  A298 );
 a43218a <=( A302  and  A300 );
 a43219a <=( a43218a  and  a43215a );
 a43220a <=( a43219a  and  a43212a );
 a43224a <=( (not A200)  and  A167 );
 a43225a <=( A168  and  a43224a );
 a43228a <=( (not A203)  and  (not A202) );
 a43231a <=( (not A234)  and  (not A233) );
 a43232a <=( a43231a  and  a43228a );
 a43233a <=( a43232a  and  a43225a );
 a43237a <=( (not A269)  and  (not A268) );
 a43238a <=( (not A266)  and  a43237a );
 a43241a <=( (not A299)  and  A298 );
 a43244a <=( A301  and  A300 );
 a43245a <=( a43244a  and  a43241a );
 a43246a <=( a43245a  and  a43238a );
 a43250a <=( (not A200)  and  A167 );
 a43251a <=( A168  and  a43250a );
 a43254a <=( (not A203)  and  (not A202) );
 a43257a <=( (not A234)  and  (not A233) );
 a43258a <=( a43257a  and  a43254a );
 a43259a <=( a43258a  and  a43251a );
 a43263a <=( (not A269)  and  (not A268) );
 a43264a <=( (not A266)  and  a43263a );
 a43267a <=( (not A299)  and  A298 );
 a43270a <=( A302  and  A300 );
 a43271a <=( a43270a  and  a43267a );
 a43272a <=( a43271a  and  a43264a );
 a43276a <=( (not A200)  and  A167 );
 a43277a <=( A168  and  a43276a );
 a43280a <=( (not A203)  and  (not A202) );
 a43283a <=( (not A233)  and  (not A232) );
 a43284a <=( a43283a  and  a43280a );
 a43285a <=( a43284a  and  a43277a );
 a43289a <=( (not A269)  and  (not A268) );
 a43290a <=( (not A266)  and  a43289a );
 a43293a <=( (not A299)  and  A298 );
 a43296a <=( A301  and  A300 );
 a43297a <=( a43296a  and  a43293a );
 a43298a <=( a43297a  and  a43290a );
 a43302a <=( (not A200)  and  A167 );
 a43303a <=( A168  and  a43302a );
 a43306a <=( (not A203)  and  (not A202) );
 a43309a <=( (not A233)  and  (not A232) );
 a43310a <=( a43309a  and  a43306a );
 a43311a <=( a43310a  and  a43303a );
 a43315a <=( (not A269)  and  (not A268) );
 a43316a <=( (not A266)  and  a43315a );
 a43319a <=( (not A299)  and  A298 );
 a43322a <=( A302  and  A300 );
 a43323a <=( a43322a  and  a43319a );
 a43324a <=( a43323a  and  a43316a );
 a43328a <=( (not A200)  and  A167 );
 a43329a <=( A168  and  a43328a );
 a43332a <=( (not A233)  and  (not A201) );
 a43335a <=( (not A236)  and  (not A235) );
 a43336a <=( a43335a  and  a43332a );
 a43337a <=( a43336a  and  a43329a );
 a43341a <=( (not A269)  and  (not A268) );
 a43342a <=( (not A266)  and  a43341a );
 a43345a <=( (not A299)  and  A298 );
 a43348a <=( A301  and  A300 );
 a43349a <=( a43348a  and  a43345a );
 a43350a <=( a43349a  and  a43342a );
 a43354a <=( (not A200)  and  A167 );
 a43355a <=( A168  and  a43354a );
 a43358a <=( (not A233)  and  (not A201) );
 a43361a <=( (not A236)  and  (not A235) );
 a43362a <=( a43361a  and  a43358a );
 a43363a <=( a43362a  and  a43355a );
 a43367a <=( (not A269)  and  (not A268) );
 a43368a <=( (not A266)  and  a43367a );
 a43371a <=( (not A299)  and  A298 );
 a43374a <=( A302  and  A300 );
 a43375a <=( a43374a  and  a43371a );
 a43376a <=( a43375a  and  a43368a );
 a43380a <=( (not A199)  and  A167 );
 a43381a <=( A168  and  a43380a );
 a43384a <=( (not A233)  and  (not A200) );
 a43387a <=( (not A236)  and  (not A235) );
 a43388a <=( a43387a  and  a43384a );
 a43389a <=( a43388a  and  a43381a );
 a43393a <=( (not A269)  and  (not A268) );
 a43394a <=( (not A266)  and  a43393a );
 a43397a <=( (not A299)  and  A298 );
 a43400a <=( A301  and  A300 );
 a43401a <=( a43400a  and  a43397a );
 a43402a <=( a43401a  and  a43394a );
 a43406a <=( (not A199)  and  A167 );
 a43407a <=( A168  and  a43406a );
 a43410a <=( (not A233)  and  (not A200) );
 a43413a <=( (not A236)  and  (not A235) );
 a43414a <=( a43413a  and  a43410a );
 a43415a <=( a43414a  and  a43407a );
 a43419a <=( (not A269)  and  (not A268) );
 a43420a <=( (not A266)  and  a43419a );
 a43423a <=( (not A299)  and  A298 );
 a43426a <=( A302  and  A300 );
 a43427a <=( a43426a  and  a43423a );
 a43428a <=( a43427a  and  a43420a );
 a43432a <=( (not A166)  and  (not A167) );
 a43433a <=( A170  and  a43432a );
 a43436a <=( A200  and  (not A199) );
 a43439a <=( A233  and  A232 );
 a43440a <=( a43439a  and  a43436a );
 a43441a <=( a43440a  and  a43433a );
 a43445a <=( (not A269)  and  (not A268) );
 a43446a <=( A265  and  a43445a );
 a43449a <=( (not A299)  and  A298 );
 a43452a <=( A301  and  A300 );
 a43453a <=( a43452a  and  a43449a );
 a43454a <=( a43453a  and  a43446a );
 a43458a <=( (not A166)  and  (not A167) );
 a43459a <=( A170  and  a43458a );
 a43462a <=( A200  and  (not A199) );
 a43465a <=( A233  and  A232 );
 a43466a <=( a43465a  and  a43462a );
 a43467a <=( a43466a  and  a43459a );
 a43471a <=( (not A269)  and  (not A268) );
 a43472a <=( A265  and  a43471a );
 a43475a <=( (not A299)  and  A298 );
 a43478a <=( A302  and  A300 );
 a43479a <=( a43478a  and  a43475a );
 a43480a <=( a43479a  and  a43472a );
 a43484a <=( (not A166)  and  (not A167) );
 a43485a <=( A170  and  a43484a );
 a43488a <=( A200  and  (not A199) );
 a43491a <=( (not A235)  and  (not A233) );
 a43492a <=( a43491a  and  a43488a );
 a43493a <=( a43492a  and  a43485a );
 a43497a <=( A266  and  A265 );
 a43498a <=( (not A236)  and  a43497a );
 a43501a <=( (not A299)  and  A298 );
 a43504a <=( A301  and  A300 );
 a43505a <=( a43504a  and  a43501a );
 a43506a <=( a43505a  and  a43498a );
 a43510a <=( (not A166)  and  (not A167) );
 a43511a <=( A170  and  a43510a );
 a43514a <=( A200  and  (not A199) );
 a43517a <=( (not A235)  and  (not A233) );
 a43518a <=( a43517a  and  a43514a );
 a43519a <=( a43518a  and  a43511a );
 a43523a <=( A266  and  A265 );
 a43524a <=( (not A236)  and  a43523a );
 a43527a <=( (not A299)  and  A298 );
 a43530a <=( A302  and  A300 );
 a43531a <=( a43530a  and  a43527a );
 a43532a <=( a43531a  and  a43524a );
 a43536a <=( (not A166)  and  (not A167) );
 a43537a <=( A170  and  a43536a );
 a43540a <=( A200  and  (not A199) );
 a43543a <=( (not A235)  and  (not A233) );
 a43544a <=( a43543a  and  a43540a );
 a43545a <=( a43544a  and  a43537a );
 a43549a <=( (not A267)  and  (not A266) );
 a43550a <=( (not A236)  and  a43549a );
 a43553a <=( (not A299)  and  A298 );
 a43556a <=( A301  and  A300 );
 a43557a <=( a43556a  and  a43553a );
 a43558a <=( a43557a  and  a43550a );
 a43562a <=( (not A166)  and  (not A167) );
 a43563a <=( A170  and  a43562a );
 a43566a <=( A200  and  (not A199) );
 a43569a <=( (not A235)  and  (not A233) );
 a43570a <=( a43569a  and  a43566a );
 a43571a <=( a43570a  and  a43563a );
 a43575a <=( (not A267)  and  (not A266) );
 a43576a <=( (not A236)  and  a43575a );
 a43579a <=( (not A299)  and  A298 );
 a43582a <=( A302  and  A300 );
 a43583a <=( a43582a  and  a43579a );
 a43584a <=( a43583a  and  a43576a );
 a43588a <=( (not A166)  and  (not A167) );
 a43589a <=( A170  and  a43588a );
 a43592a <=( A200  and  (not A199) );
 a43595a <=( (not A235)  and  (not A233) );
 a43596a <=( a43595a  and  a43592a );
 a43597a <=( a43596a  and  a43589a );
 a43601a <=( (not A266)  and  (not A265) );
 a43602a <=( (not A236)  and  a43601a );
 a43605a <=( (not A299)  and  A298 );
 a43608a <=( A301  and  A300 );
 a43609a <=( a43608a  and  a43605a );
 a43610a <=( a43609a  and  a43602a );
 a43614a <=( (not A166)  and  (not A167) );
 a43615a <=( A170  and  a43614a );
 a43618a <=( A200  and  (not A199) );
 a43621a <=( (not A235)  and  (not A233) );
 a43622a <=( a43621a  and  a43618a );
 a43623a <=( a43622a  and  a43615a );
 a43627a <=( (not A266)  and  (not A265) );
 a43628a <=( (not A236)  and  a43627a );
 a43631a <=( (not A299)  and  A298 );
 a43634a <=( A302  and  A300 );
 a43635a <=( a43634a  and  a43631a );
 a43636a <=( a43635a  and  a43628a );
 a43640a <=( (not A166)  and  (not A167) );
 a43641a <=( A170  and  a43640a );
 a43644a <=( A200  and  (not A199) );
 a43647a <=( (not A234)  and  (not A233) );
 a43648a <=( a43647a  and  a43644a );
 a43649a <=( a43648a  and  a43641a );
 a43653a <=( (not A269)  and  (not A268) );
 a43654a <=( (not A266)  and  a43653a );
 a43657a <=( (not A299)  and  A298 );
 a43660a <=( A301  and  A300 );
 a43661a <=( a43660a  and  a43657a );
 a43662a <=( a43661a  and  a43654a );
 a43666a <=( (not A166)  and  (not A167) );
 a43667a <=( A170  and  a43666a );
 a43670a <=( A200  and  (not A199) );
 a43673a <=( (not A234)  and  (not A233) );
 a43674a <=( a43673a  and  a43670a );
 a43675a <=( a43674a  and  a43667a );
 a43679a <=( (not A269)  and  (not A268) );
 a43680a <=( (not A266)  and  a43679a );
 a43683a <=( (not A299)  and  A298 );
 a43686a <=( A302  and  A300 );
 a43687a <=( a43686a  and  a43683a );
 a43688a <=( a43687a  and  a43680a );
 a43692a <=( (not A166)  and  (not A167) );
 a43693a <=( A170  and  a43692a );
 a43696a <=( A200  and  (not A199) );
 a43699a <=( (not A233)  and  (not A232) );
 a43700a <=( a43699a  and  a43696a );
 a43701a <=( a43700a  and  a43693a );
 a43705a <=( (not A269)  and  (not A268) );
 a43706a <=( (not A266)  and  a43705a );
 a43709a <=( (not A299)  and  A298 );
 a43712a <=( A301  and  A300 );
 a43713a <=( a43712a  and  a43709a );
 a43714a <=( a43713a  and  a43706a );
 a43718a <=( (not A166)  and  (not A167) );
 a43719a <=( A170  and  a43718a );
 a43722a <=( A200  and  (not A199) );
 a43725a <=( (not A233)  and  (not A232) );
 a43726a <=( a43725a  and  a43722a );
 a43727a <=( a43726a  and  a43719a );
 a43731a <=( (not A269)  and  (not A268) );
 a43732a <=( (not A266)  and  a43731a );
 a43735a <=( (not A299)  and  A298 );
 a43738a <=( A302  and  A300 );
 a43739a <=( a43738a  and  a43735a );
 a43740a <=( a43739a  and  a43732a );
 a43744a <=( (not A166)  and  (not A167) );
 a43745a <=( A170  and  a43744a );
 a43748a <=( (not A200)  and  A199 );
 a43751a <=( A202  and  A201 );
 a43752a <=( a43751a  and  a43748a );
 a43753a <=( a43752a  and  a43745a );
 a43757a <=( A265  and  A233 );
 a43758a <=( A232  and  a43757a );
 a43761a <=( (not A269)  and  (not A268) );
 a43764a <=( A299  and  (not A298) );
 a43765a <=( a43764a  and  a43761a );
 a43766a <=( a43765a  and  a43758a );
 a43770a <=( (not A166)  and  (not A167) );
 a43771a <=( A170  and  a43770a );
 a43774a <=( (not A200)  and  A199 );
 a43777a <=( A202  and  A201 );
 a43778a <=( a43777a  and  a43774a );
 a43779a <=( a43778a  and  a43771a );
 a43783a <=( (not A236)  and  (not A235) );
 a43784a <=( (not A233)  and  a43783a );
 a43787a <=( A266  and  A265 );
 a43790a <=( A299  and  (not A298) );
 a43791a <=( a43790a  and  a43787a );
 a43792a <=( a43791a  and  a43784a );
 a43796a <=( (not A166)  and  (not A167) );
 a43797a <=( A170  and  a43796a );
 a43800a <=( (not A200)  and  A199 );
 a43803a <=( A202  and  A201 );
 a43804a <=( a43803a  and  a43800a );
 a43805a <=( a43804a  and  a43797a );
 a43809a <=( (not A236)  and  (not A235) );
 a43810a <=( (not A233)  and  a43809a );
 a43813a <=( (not A267)  and  (not A266) );
 a43816a <=( A299  and  (not A298) );
 a43817a <=( a43816a  and  a43813a );
 a43818a <=( a43817a  and  a43810a );
 a43822a <=( (not A166)  and  (not A167) );
 a43823a <=( A170  and  a43822a );
 a43826a <=( (not A200)  and  A199 );
 a43829a <=( A202  and  A201 );
 a43830a <=( a43829a  and  a43826a );
 a43831a <=( a43830a  and  a43823a );
 a43835a <=( (not A236)  and  (not A235) );
 a43836a <=( (not A233)  and  a43835a );
 a43839a <=( (not A266)  and  (not A265) );
 a43842a <=( A299  and  (not A298) );
 a43843a <=( a43842a  and  a43839a );
 a43844a <=( a43843a  and  a43836a );
 a43848a <=( (not A166)  and  (not A167) );
 a43849a <=( A170  and  a43848a );
 a43852a <=( (not A200)  and  A199 );
 a43855a <=( A202  and  A201 );
 a43856a <=( a43855a  and  a43852a );
 a43857a <=( a43856a  and  a43849a );
 a43861a <=( (not A266)  and  (not A234) );
 a43862a <=( (not A233)  and  a43861a );
 a43865a <=( (not A269)  and  (not A268) );
 a43868a <=( A299  and  (not A298) );
 a43869a <=( a43868a  and  a43865a );
 a43870a <=( a43869a  and  a43862a );
 a43874a <=( (not A166)  and  (not A167) );
 a43875a <=( A170  and  a43874a );
 a43878a <=( (not A200)  and  A199 );
 a43881a <=( A202  and  A201 );
 a43882a <=( a43881a  and  a43878a );
 a43883a <=( a43882a  and  a43875a );
 a43887a <=( A234  and  (not A233) );
 a43888a <=( A232  and  a43887a );
 a43891a <=( A298  and  A235 );
 a43894a <=( (not A302)  and  (not A301) );
 a43895a <=( a43894a  and  a43891a );
 a43896a <=( a43895a  and  a43888a );
 a43900a <=( (not A166)  and  (not A167) );
 a43901a <=( A170  and  a43900a );
 a43904a <=( (not A200)  and  A199 );
 a43907a <=( A202  and  A201 );
 a43908a <=( a43907a  and  a43904a );
 a43909a <=( a43908a  and  a43901a );
 a43913a <=( A234  and  (not A233) );
 a43914a <=( A232  and  a43913a );
 a43917a <=( A298  and  A236 );
 a43920a <=( (not A302)  and  (not A301) );
 a43921a <=( a43920a  and  a43917a );
 a43922a <=( a43921a  and  a43914a );
 a43926a <=( (not A166)  and  (not A167) );
 a43927a <=( A170  and  a43926a );
 a43930a <=( (not A200)  and  A199 );
 a43933a <=( A202  and  A201 );
 a43934a <=( a43933a  and  a43930a );
 a43935a <=( a43934a  and  a43927a );
 a43939a <=( (not A266)  and  (not A233) );
 a43940a <=( (not A232)  and  a43939a );
 a43943a <=( (not A269)  and  (not A268) );
 a43946a <=( A299  and  (not A298) );
 a43947a <=( a43946a  and  a43943a );
 a43948a <=( a43947a  and  a43940a );
 a43952a <=( (not A166)  and  (not A167) );
 a43953a <=( A170  and  a43952a );
 a43956a <=( (not A200)  and  A199 );
 a43959a <=( A203  and  A201 );
 a43960a <=( a43959a  and  a43956a );
 a43961a <=( a43960a  and  a43953a );
 a43965a <=( A265  and  A233 );
 a43966a <=( A232  and  a43965a );
 a43969a <=( (not A269)  and  (not A268) );
 a43972a <=( A299  and  (not A298) );
 a43973a <=( a43972a  and  a43969a );
 a43974a <=( a43973a  and  a43966a );
 a43978a <=( (not A166)  and  (not A167) );
 a43979a <=( A170  and  a43978a );
 a43982a <=( (not A200)  and  A199 );
 a43985a <=( A203  and  A201 );
 a43986a <=( a43985a  and  a43982a );
 a43987a <=( a43986a  and  a43979a );
 a43991a <=( (not A236)  and  (not A235) );
 a43992a <=( (not A233)  and  a43991a );
 a43995a <=( A266  and  A265 );
 a43998a <=( A299  and  (not A298) );
 a43999a <=( a43998a  and  a43995a );
 a44000a <=( a43999a  and  a43992a );
 a44004a <=( (not A166)  and  (not A167) );
 a44005a <=( A170  and  a44004a );
 a44008a <=( (not A200)  and  A199 );
 a44011a <=( A203  and  A201 );
 a44012a <=( a44011a  and  a44008a );
 a44013a <=( a44012a  and  a44005a );
 a44017a <=( (not A236)  and  (not A235) );
 a44018a <=( (not A233)  and  a44017a );
 a44021a <=( (not A267)  and  (not A266) );
 a44024a <=( A299  and  (not A298) );
 a44025a <=( a44024a  and  a44021a );
 a44026a <=( a44025a  and  a44018a );
 a44030a <=( (not A166)  and  (not A167) );
 a44031a <=( A170  and  a44030a );
 a44034a <=( (not A200)  and  A199 );
 a44037a <=( A203  and  A201 );
 a44038a <=( a44037a  and  a44034a );
 a44039a <=( a44038a  and  a44031a );
 a44043a <=( (not A236)  and  (not A235) );
 a44044a <=( (not A233)  and  a44043a );
 a44047a <=( (not A266)  and  (not A265) );
 a44050a <=( A299  and  (not A298) );
 a44051a <=( a44050a  and  a44047a );
 a44052a <=( a44051a  and  a44044a );
 a44056a <=( (not A166)  and  (not A167) );
 a44057a <=( A170  and  a44056a );
 a44060a <=( (not A200)  and  A199 );
 a44063a <=( A203  and  A201 );
 a44064a <=( a44063a  and  a44060a );
 a44065a <=( a44064a  and  a44057a );
 a44069a <=( (not A266)  and  (not A234) );
 a44070a <=( (not A233)  and  a44069a );
 a44073a <=( (not A269)  and  (not A268) );
 a44076a <=( A299  and  (not A298) );
 a44077a <=( a44076a  and  a44073a );
 a44078a <=( a44077a  and  a44070a );
 a44082a <=( (not A166)  and  (not A167) );
 a44083a <=( A170  and  a44082a );
 a44086a <=( (not A200)  and  A199 );
 a44089a <=( A203  and  A201 );
 a44090a <=( a44089a  and  a44086a );
 a44091a <=( a44090a  and  a44083a );
 a44095a <=( A234  and  (not A233) );
 a44096a <=( A232  and  a44095a );
 a44099a <=( A298  and  A235 );
 a44102a <=( (not A302)  and  (not A301) );
 a44103a <=( a44102a  and  a44099a );
 a44104a <=( a44103a  and  a44096a );
 a44108a <=( (not A166)  and  (not A167) );
 a44109a <=( A170  and  a44108a );
 a44112a <=( (not A200)  and  A199 );
 a44115a <=( A203  and  A201 );
 a44116a <=( a44115a  and  a44112a );
 a44117a <=( a44116a  and  a44109a );
 a44121a <=( A234  and  (not A233) );
 a44122a <=( A232  and  a44121a );
 a44125a <=( A298  and  A236 );
 a44128a <=( (not A302)  and  (not A301) );
 a44129a <=( a44128a  and  a44125a );
 a44130a <=( a44129a  and  a44122a );
 a44134a <=( (not A166)  and  (not A167) );
 a44135a <=( A170  and  a44134a );
 a44138a <=( (not A200)  and  A199 );
 a44141a <=( A203  and  A201 );
 a44142a <=( a44141a  and  a44138a );
 a44143a <=( a44142a  and  a44135a );
 a44147a <=( (not A266)  and  (not A233) );
 a44148a <=( (not A232)  and  a44147a );
 a44151a <=( (not A269)  and  (not A268) );
 a44154a <=( A299  and  (not A298) );
 a44155a <=( a44154a  and  a44151a );
 a44156a <=( a44155a  and  a44148a );
 a44160a <=( A167  and  (not A168) );
 a44161a <=( A170  and  a44160a );
 a44164a <=( (not A199)  and  A166 );
 a44167a <=( A232  and  A200 );
 a44168a <=( a44167a  and  a44164a );
 a44169a <=( a44168a  and  a44161a );
 a44173a <=( (not A267)  and  A265 );
 a44174a <=( A233  and  a44173a );
 a44177a <=( (not A299)  and  A298 );
 a44180a <=( A301  and  A300 );
 a44181a <=( a44180a  and  a44177a );
 a44182a <=( a44181a  and  a44174a );
 a44186a <=( A167  and  (not A168) );
 a44187a <=( A170  and  a44186a );
 a44190a <=( (not A199)  and  A166 );
 a44193a <=( A232  and  A200 );
 a44194a <=( a44193a  and  a44190a );
 a44195a <=( a44194a  and  a44187a );
 a44199a <=( (not A267)  and  A265 );
 a44200a <=( A233  and  a44199a );
 a44203a <=( (not A299)  and  A298 );
 a44206a <=( A302  and  A300 );
 a44207a <=( a44206a  and  a44203a );
 a44208a <=( a44207a  and  a44200a );
 a44212a <=( A167  and  (not A168) );
 a44213a <=( A170  and  a44212a );
 a44216a <=( (not A199)  and  A166 );
 a44219a <=( A232  and  A200 );
 a44220a <=( a44219a  and  a44216a );
 a44221a <=( a44220a  and  a44213a );
 a44225a <=( A266  and  A265 );
 a44226a <=( A233  and  a44225a );
 a44229a <=( (not A299)  and  A298 );
 a44232a <=( A301  and  A300 );
 a44233a <=( a44232a  and  a44229a );
 a44234a <=( a44233a  and  a44226a );
 a44238a <=( A167  and  (not A168) );
 a44239a <=( A170  and  a44238a );
 a44242a <=( (not A199)  and  A166 );
 a44245a <=( A232  and  A200 );
 a44246a <=( a44245a  and  a44242a );
 a44247a <=( a44246a  and  a44239a );
 a44251a <=( A266  and  A265 );
 a44252a <=( A233  and  a44251a );
 a44255a <=( (not A299)  and  A298 );
 a44258a <=( A302  and  A300 );
 a44259a <=( a44258a  and  a44255a );
 a44260a <=( a44259a  and  a44252a );
 a44264a <=( A167  and  (not A168) );
 a44265a <=( A170  and  a44264a );
 a44268a <=( (not A199)  and  A166 );
 a44271a <=( A232  and  A200 );
 a44272a <=( a44271a  and  a44268a );
 a44273a <=( a44272a  and  a44265a );
 a44277a <=( (not A266)  and  (not A265) );
 a44278a <=( A233  and  a44277a );
 a44281a <=( (not A299)  and  A298 );
 a44284a <=( A301  and  A300 );
 a44285a <=( a44284a  and  a44281a );
 a44286a <=( a44285a  and  a44278a );
 a44290a <=( A167  and  (not A168) );
 a44291a <=( A170  and  a44290a );
 a44294a <=( (not A199)  and  A166 );
 a44297a <=( A232  and  A200 );
 a44298a <=( a44297a  and  a44294a );
 a44299a <=( a44298a  and  a44291a );
 a44303a <=( (not A266)  and  (not A265) );
 a44304a <=( A233  and  a44303a );
 a44307a <=( (not A299)  and  A298 );
 a44310a <=( A302  and  A300 );
 a44311a <=( a44310a  and  a44307a );
 a44312a <=( a44311a  and  a44304a );
 a44316a <=( A167  and  (not A168) );
 a44317a <=( A170  and  a44316a );
 a44320a <=( (not A199)  and  A166 );
 a44323a <=( (not A233)  and  A200 );
 a44324a <=( a44323a  and  a44320a );
 a44325a <=( a44324a  and  a44317a );
 a44329a <=( (not A266)  and  (not A236) );
 a44330a <=( (not A235)  and  a44329a );
 a44333a <=( (not A269)  and  (not A268) );
 a44336a <=( A299  and  (not A298) );
 a44337a <=( a44336a  and  a44333a );
 a44338a <=( a44337a  and  a44330a );
 a44342a <=( A167  and  (not A168) );
 a44343a <=( A170  and  a44342a );
 a44346a <=( (not A199)  and  A166 );
 a44349a <=( (not A233)  and  A200 );
 a44350a <=( a44349a  and  a44346a );
 a44351a <=( a44350a  and  a44343a );
 a44355a <=( A266  and  A265 );
 a44356a <=( (not A234)  and  a44355a );
 a44359a <=( (not A299)  and  A298 );
 a44362a <=( A301  and  A300 );
 a44363a <=( a44362a  and  a44359a );
 a44364a <=( a44363a  and  a44356a );
 a44368a <=( A167  and  (not A168) );
 a44369a <=( A170  and  a44368a );
 a44372a <=( (not A199)  and  A166 );
 a44375a <=( (not A233)  and  A200 );
 a44376a <=( a44375a  and  a44372a );
 a44377a <=( a44376a  and  a44369a );
 a44381a <=( A266  and  A265 );
 a44382a <=( (not A234)  and  a44381a );
 a44385a <=( (not A299)  and  A298 );
 a44388a <=( A302  and  A300 );
 a44389a <=( a44388a  and  a44385a );
 a44390a <=( a44389a  and  a44382a );
 a44394a <=( A167  and  (not A168) );
 a44395a <=( A170  and  a44394a );
 a44398a <=( (not A199)  and  A166 );
 a44401a <=( (not A233)  and  A200 );
 a44402a <=( a44401a  and  a44398a );
 a44403a <=( a44402a  and  a44395a );
 a44407a <=( (not A267)  and  (not A266) );
 a44408a <=( (not A234)  and  a44407a );
 a44411a <=( (not A299)  and  A298 );
 a44414a <=( A301  and  A300 );
 a44415a <=( a44414a  and  a44411a );
 a44416a <=( a44415a  and  a44408a );
 a44420a <=( A167  and  (not A168) );
 a44421a <=( A170  and  a44420a );
 a44424a <=( (not A199)  and  A166 );
 a44427a <=( (not A233)  and  A200 );
 a44428a <=( a44427a  and  a44424a );
 a44429a <=( a44428a  and  a44421a );
 a44433a <=( (not A267)  and  (not A266) );
 a44434a <=( (not A234)  and  a44433a );
 a44437a <=( (not A299)  and  A298 );
 a44440a <=( A302  and  A300 );
 a44441a <=( a44440a  and  a44437a );
 a44442a <=( a44441a  and  a44434a );
 a44446a <=( A167  and  (not A168) );
 a44447a <=( A170  and  a44446a );
 a44450a <=( (not A199)  and  A166 );
 a44453a <=( (not A233)  and  A200 );
 a44454a <=( a44453a  and  a44450a );
 a44455a <=( a44454a  and  a44447a );
 a44459a <=( (not A266)  and  (not A265) );
 a44460a <=( (not A234)  and  a44459a );
 a44463a <=( (not A299)  and  A298 );
 a44466a <=( A301  and  A300 );
 a44467a <=( a44466a  and  a44463a );
 a44468a <=( a44467a  and  a44460a );
 a44472a <=( A167  and  (not A168) );
 a44473a <=( A170  and  a44472a );
 a44476a <=( (not A199)  and  A166 );
 a44479a <=( (not A233)  and  A200 );
 a44480a <=( a44479a  and  a44476a );
 a44481a <=( a44480a  and  a44473a );
 a44485a <=( (not A266)  and  (not A265) );
 a44486a <=( (not A234)  and  a44485a );
 a44489a <=( (not A299)  and  A298 );
 a44492a <=( A302  and  A300 );
 a44493a <=( a44492a  and  a44489a );
 a44494a <=( a44493a  and  a44486a );
 a44498a <=( A167  and  (not A168) );
 a44499a <=( A170  and  a44498a );
 a44502a <=( (not A199)  and  A166 );
 a44505a <=( A232  and  A200 );
 a44506a <=( a44505a  and  a44502a );
 a44507a <=( a44506a  and  a44499a );
 a44511a <=( A235  and  A234 );
 a44512a <=( (not A233)  and  a44511a );
 a44515a <=( (not A266)  and  A265 );
 a44518a <=( A268  and  A267 );
 a44519a <=( a44518a  and  a44515a );
 a44520a <=( a44519a  and  a44512a );
 a44524a <=( A167  and  (not A168) );
 a44525a <=( A170  and  a44524a );
 a44528a <=( (not A199)  and  A166 );
 a44531a <=( A232  and  A200 );
 a44532a <=( a44531a  and  a44528a );
 a44533a <=( a44532a  and  a44525a );
 a44537a <=( A235  and  A234 );
 a44538a <=( (not A233)  and  a44537a );
 a44541a <=( (not A266)  and  A265 );
 a44544a <=( A269  and  A267 );
 a44545a <=( a44544a  and  a44541a );
 a44546a <=( a44545a  and  a44538a );
 a44550a <=( A167  and  (not A168) );
 a44551a <=( A170  and  a44550a );
 a44554a <=( (not A199)  and  A166 );
 a44557a <=( A232  and  A200 );
 a44558a <=( a44557a  and  a44554a );
 a44559a <=( a44558a  and  a44551a );
 a44563a <=( A236  and  A234 );
 a44564a <=( (not A233)  and  a44563a );
 a44567a <=( (not A266)  and  A265 );
 a44570a <=( A268  and  A267 );
 a44571a <=( a44570a  and  a44567a );
 a44572a <=( a44571a  and  a44564a );
 a44576a <=( A167  and  (not A168) );
 a44577a <=( A170  and  a44576a );
 a44580a <=( (not A199)  and  A166 );
 a44583a <=( A232  and  A200 );
 a44584a <=( a44583a  and  a44580a );
 a44585a <=( a44584a  and  a44577a );
 a44589a <=( A236  and  A234 );
 a44590a <=( (not A233)  and  a44589a );
 a44593a <=( (not A266)  and  A265 );
 a44596a <=( A269  and  A267 );
 a44597a <=( a44596a  and  a44593a );
 a44598a <=( a44597a  and  a44590a );
 a44602a <=( A167  and  (not A168) );
 a44603a <=( A170  and  a44602a );
 a44606a <=( (not A199)  and  A166 );
 a44609a <=( (not A232)  and  A200 );
 a44610a <=( a44609a  and  a44606a );
 a44611a <=( a44610a  and  a44603a );
 a44615a <=( A266  and  A265 );
 a44616a <=( (not A233)  and  a44615a );
 a44619a <=( (not A299)  and  A298 );
 a44622a <=( A301  and  A300 );
 a44623a <=( a44622a  and  a44619a );
 a44624a <=( a44623a  and  a44616a );
 a44628a <=( A167  and  (not A168) );
 a44629a <=( A170  and  a44628a );
 a44632a <=( (not A199)  and  A166 );
 a44635a <=( (not A232)  and  A200 );
 a44636a <=( a44635a  and  a44632a );
 a44637a <=( a44636a  and  a44629a );
 a44641a <=( A266  and  A265 );
 a44642a <=( (not A233)  and  a44641a );
 a44645a <=( (not A299)  and  A298 );
 a44648a <=( A302  and  A300 );
 a44649a <=( a44648a  and  a44645a );
 a44650a <=( a44649a  and  a44642a );
 a44654a <=( A167  and  (not A168) );
 a44655a <=( A170  and  a44654a );
 a44658a <=( (not A199)  and  A166 );
 a44661a <=( (not A232)  and  A200 );
 a44662a <=( a44661a  and  a44658a );
 a44663a <=( a44662a  and  a44655a );
 a44667a <=( (not A267)  and  (not A266) );
 a44668a <=( (not A233)  and  a44667a );
 a44671a <=( (not A299)  and  A298 );
 a44674a <=( A301  and  A300 );
 a44675a <=( a44674a  and  a44671a );
 a44676a <=( a44675a  and  a44668a );
 a44680a <=( A167  and  (not A168) );
 a44681a <=( A170  and  a44680a );
 a44684a <=( (not A199)  and  A166 );
 a44687a <=( (not A232)  and  A200 );
 a44688a <=( a44687a  and  a44684a );
 a44689a <=( a44688a  and  a44681a );
 a44693a <=( (not A267)  and  (not A266) );
 a44694a <=( (not A233)  and  a44693a );
 a44697a <=( (not A299)  and  A298 );
 a44700a <=( A302  and  A300 );
 a44701a <=( a44700a  and  a44697a );
 a44702a <=( a44701a  and  a44694a );
 a44706a <=( A167  and  (not A168) );
 a44707a <=( A170  and  a44706a );
 a44710a <=( (not A199)  and  A166 );
 a44713a <=( (not A232)  and  A200 );
 a44714a <=( a44713a  and  a44710a );
 a44715a <=( a44714a  and  a44707a );
 a44719a <=( (not A266)  and  (not A265) );
 a44720a <=( (not A233)  and  a44719a );
 a44723a <=( (not A299)  and  A298 );
 a44726a <=( A301  and  A300 );
 a44727a <=( a44726a  and  a44723a );
 a44728a <=( a44727a  and  a44720a );
 a44732a <=( A167  and  (not A168) );
 a44733a <=( A170  and  a44732a );
 a44736a <=( (not A199)  and  A166 );
 a44739a <=( (not A232)  and  A200 );
 a44740a <=( a44739a  and  a44736a );
 a44741a <=( a44740a  and  a44733a );
 a44745a <=( (not A266)  and  (not A265) );
 a44746a <=( (not A233)  and  a44745a );
 a44749a <=( (not A299)  and  A298 );
 a44752a <=( A302  and  A300 );
 a44753a <=( a44752a  and  a44749a );
 a44754a <=( a44753a  and  a44746a );
 a44758a <=( A167  and  (not A168) );
 a44759a <=( (not A170)  and  a44758a );
 a44762a <=( (not A199)  and  (not A166) );
 a44765a <=( A232  and  A200 );
 a44766a <=( a44765a  and  a44762a );
 a44767a <=( a44766a  and  a44759a );
 a44771a <=( (not A267)  and  A265 );
 a44772a <=( A233  and  a44771a );
 a44775a <=( (not A299)  and  A298 );
 a44778a <=( A301  and  A300 );
 a44779a <=( a44778a  and  a44775a );
 a44780a <=( a44779a  and  a44772a );
 a44784a <=( A167  and  (not A168) );
 a44785a <=( (not A170)  and  a44784a );
 a44788a <=( (not A199)  and  (not A166) );
 a44791a <=( A232  and  A200 );
 a44792a <=( a44791a  and  a44788a );
 a44793a <=( a44792a  and  a44785a );
 a44797a <=( (not A267)  and  A265 );
 a44798a <=( A233  and  a44797a );
 a44801a <=( (not A299)  and  A298 );
 a44804a <=( A302  and  A300 );
 a44805a <=( a44804a  and  a44801a );
 a44806a <=( a44805a  and  a44798a );
 a44810a <=( A167  and  (not A168) );
 a44811a <=( (not A170)  and  a44810a );
 a44814a <=( (not A199)  and  (not A166) );
 a44817a <=( A232  and  A200 );
 a44818a <=( a44817a  and  a44814a );
 a44819a <=( a44818a  and  a44811a );
 a44823a <=( A266  and  A265 );
 a44824a <=( A233  and  a44823a );
 a44827a <=( (not A299)  and  A298 );
 a44830a <=( A301  and  A300 );
 a44831a <=( a44830a  and  a44827a );
 a44832a <=( a44831a  and  a44824a );
 a44836a <=( A167  and  (not A168) );
 a44837a <=( (not A170)  and  a44836a );
 a44840a <=( (not A199)  and  (not A166) );
 a44843a <=( A232  and  A200 );
 a44844a <=( a44843a  and  a44840a );
 a44845a <=( a44844a  and  a44837a );
 a44849a <=( A266  and  A265 );
 a44850a <=( A233  and  a44849a );
 a44853a <=( (not A299)  and  A298 );
 a44856a <=( A302  and  A300 );
 a44857a <=( a44856a  and  a44853a );
 a44858a <=( a44857a  and  a44850a );
 a44862a <=( A167  and  (not A168) );
 a44863a <=( (not A170)  and  a44862a );
 a44866a <=( (not A199)  and  (not A166) );
 a44869a <=( A232  and  A200 );
 a44870a <=( a44869a  and  a44866a );
 a44871a <=( a44870a  and  a44863a );
 a44875a <=( (not A266)  and  (not A265) );
 a44876a <=( A233  and  a44875a );
 a44879a <=( (not A299)  and  A298 );
 a44882a <=( A301  and  A300 );
 a44883a <=( a44882a  and  a44879a );
 a44884a <=( a44883a  and  a44876a );
 a44888a <=( A167  and  (not A168) );
 a44889a <=( (not A170)  and  a44888a );
 a44892a <=( (not A199)  and  (not A166) );
 a44895a <=( A232  and  A200 );
 a44896a <=( a44895a  and  a44892a );
 a44897a <=( a44896a  and  a44889a );
 a44901a <=( (not A266)  and  (not A265) );
 a44902a <=( A233  and  a44901a );
 a44905a <=( (not A299)  and  A298 );
 a44908a <=( A302  and  A300 );
 a44909a <=( a44908a  and  a44905a );
 a44910a <=( a44909a  and  a44902a );
 a44914a <=( A167  and  (not A168) );
 a44915a <=( (not A170)  and  a44914a );
 a44918a <=( (not A199)  and  (not A166) );
 a44921a <=( (not A233)  and  A200 );
 a44922a <=( a44921a  and  a44918a );
 a44923a <=( a44922a  and  a44915a );
 a44927a <=( (not A266)  and  (not A236) );
 a44928a <=( (not A235)  and  a44927a );
 a44931a <=( (not A269)  and  (not A268) );
 a44934a <=( A299  and  (not A298) );
 a44935a <=( a44934a  and  a44931a );
 a44936a <=( a44935a  and  a44928a );
 a44940a <=( A167  and  (not A168) );
 a44941a <=( (not A170)  and  a44940a );
 a44944a <=( (not A199)  and  (not A166) );
 a44947a <=( (not A233)  and  A200 );
 a44948a <=( a44947a  and  a44944a );
 a44949a <=( a44948a  and  a44941a );
 a44953a <=( A266  and  A265 );
 a44954a <=( (not A234)  and  a44953a );
 a44957a <=( (not A299)  and  A298 );
 a44960a <=( A301  and  A300 );
 a44961a <=( a44960a  and  a44957a );
 a44962a <=( a44961a  and  a44954a );
 a44966a <=( A167  and  (not A168) );
 a44967a <=( (not A170)  and  a44966a );
 a44970a <=( (not A199)  and  (not A166) );
 a44973a <=( (not A233)  and  A200 );
 a44974a <=( a44973a  and  a44970a );
 a44975a <=( a44974a  and  a44967a );
 a44979a <=( A266  and  A265 );
 a44980a <=( (not A234)  and  a44979a );
 a44983a <=( (not A299)  and  A298 );
 a44986a <=( A302  and  A300 );
 a44987a <=( a44986a  and  a44983a );
 a44988a <=( a44987a  and  a44980a );
 a44992a <=( A167  and  (not A168) );
 a44993a <=( (not A170)  and  a44992a );
 a44996a <=( (not A199)  and  (not A166) );
 a44999a <=( (not A233)  and  A200 );
 a45000a <=( a44999a  and  a44996a );
 a45001a <=( a45000a  and  a44993a );
 a45005a <=( (not A267)  and  (not A266) );
 a45006a <=( (not A234)  and  a45005a );
 a45009a <=( (not A299)  and  A298 );
 a45012a <=( A301  and  A300 );
 a45013a <=( a45012a  and  a45009a );
 a45014a <=( a45013a  and  a45006a );
 a45018a <=( A167  and  (not A168) );
 a45019a <=( (not A170)  and  a45018a );
 a45022a <=( (not A199)  and  (not A166) );
 a45025a <=( (not A233)  and  A200 );
 a45026a <=( a45025a  and  a45022a );
 a45027a <=( a45026a  and  a45019a );
 a45031a <=( (not A267)  and  (not A266) );
 a45032a <=( (not A234)  and  a45031a );
 a45035a <=( (not A299)  and  A298 );
 a45038a <=( A302  and  A300 );
 a45039a <=( a45038a  and  a45035a );
 a45040a <=( a45039a  and  a45032a );
 a45044a <=( A167  and  (not A168) );
 a45045a <=( (not A170)  and  a45044a );
 a45048a <=( (not A199)  and  (not A166) );
 a45051a <=( (not A233)  and  A200 );
 a45052a <=( a45051a  and  a45048a );
 a45053a <=( a45052a  and  a45045a );
 a45057a <=( (not A266)  and  (not A265) );
 a45058a <=( (not A234)  and  a45057a );
 a45061a <=( (not A299)  and  A298 );
 a45064a <=( A301  and  A300 );
 a45065a <=( a45064a  and  a45061a );
 a45066a <=( a45065a  and  a45058a );
 a45070a <=( A167  and  (not A168) );
 a45071a <=( (not A170)  and  a45070a );
 a45074a <=( (not A199)  and  (not A166) );
 a45077a <=( (not A233)  and  A200 );
 a45078a <=( a45077a  and  a45074a );
 a45079a <=( a45078a  and  a45071a );
 a45083a <=( (not A266)  and  (not A265) );
 a45084a <=( (not A234)  and  a45083a );
 a45087a <=( (not A299)  and  A298 );
 a45090a <=( A302  and  A300 );
 a45091a <=( a45090a  and  a45087a );
 a45092a <=( a45091a  and  a45084a );
 a45096a <=( A167  and  (not A168) );
 a45097a <=( (not A170)  and  a45096a );
 a45100a <=( (not A199)  and  (not A166) );
 a45103a <=( A232  and  A200 );
 a45104a <=( a45103a  and  a45100a );
 a45105a <=( a45104a  and  a45097a );
 a45109a <=( A235  and  A234 );
 a45110a <=( (not A233)  and  a45109a );
 a45113a <=( (not A266)  and  A265 );
 a45116a <=( A268  and  A267 );
 a45117a <=( a45116a  and  a45113a );
 a45118a <=( a45117a  and  a45110a );
 a45122a <=( A167  and  (not A168) );
 a45123a <=( (not A170)  and  a45122a );
 a45126a <=( (not A199)  and  (not A166) );
 a45129a <=( A232  and  A200 );
 a45130a <=( a45129a  and  a45126a );
 a45131a <=( a45130a  and  a45123a );
 a45135a <=( A235  and  A234 );
 a45136a <=( (not A233)  and  a45135a );
 a45139a <=( (not A266)  and  A265 );
 a45142a <=( A269  and  A267 );
 a45143a <=( a45142a  and  a45139a );
 a45144a <=( a45143a  and  a45136a );
 a45148a <=( A167  and  (not A168) );
 a45149a <=( (not A170)  and  a45148a );
 a45152a <=( (not A199)  and  (not A166) );
 a45155a <=( A232  and  A200 );
 a45156a <=( a45155a  and  a45152a );
 a45157a <=( a45156a  and  a45149a );
 a45161a <=( A236  and  A234 );
 a45162a <=( (not A233)  and  a45161a );
 a45165a <=( (not A266)  and  A265 );
 a45168a <=( A268  and  A267 );
 a45169a <=( a45168a  and  a45165a );
 a45170a <=( a45169a  and  a45162a );
 a45174a <=( A167  and  (not A168) );
 a45175a <=( (not A170)  and  a45174a );
 a45178a <=( (not A199)  and  (not A166) );
 a45181a <=( A232  and  A200 );
 a45182a <=( a45181a  and  a45178a );
 a45183a <=( a45182a  and  a45175a );
 a45187a <=( A236  and  A234 );
 a45188a <=( (not A233)  and  a45187a );
 a45191a <=( (not A266)  and  A265 );
 a45194a <=( A269  and  A267 );
 a45195a <=( a45194a  and  a45191a );
 a45196a <=( a45195a  and  a45188a );
 a45200a <=( A167  and  (not A168) );
 a45201a <=( (not A170)  and  a45200a );
 a45204a <=( (not A199)  and  (not A166) );
 a45207a <=( (not A232)  and  A200 );
 a45208a <=( a45207a  and  a45204a );
 a45209a <=( a45208a  and  a45201a );
 a45213a <=( A266  and  A265 );
 a45214a <=( (not A233)  and  a45213a );
 a45217a <=( (not A299)  and  A298 );
 a45220a <=( A301  and  A300 );
 a45221a <=( a45220a  and  a45217a );
 a45222a <=( a45221a  and  a45214a );
 a45226a <=( A167  and  (not A168) );
 a45227a <=( (not A170)  and  a45226a );
 a45230a <=( (not A199)  and  (not A166) );
 a45233a <=( (not A232)  and  A200 );
 a45234a <=( a45233a  and  a45230a );
 a45235a <=( a45234a  and  a45227a );
 a45239a <=( A266  and  A265 );
 a45240a <=( (not A233)  and  a45239a );
 a45243a <=( (not A299)  and  A298 );
 a45246a <=( A302  and  A300 );
 a45247a <=( a45246a  and  a45243a );
 a45248a <=( a45247a  and  a45240a );
 a45252a <=( A167  and  (not A168) );
 a45253a <=( (not A170)  and  a45252a );
 a45256a <=( (not A199)  and  (not A166) );
 a45259a <=( (not A232)  and  A200 );
 a45260a <=( a45259a  and  a45256a );
 a45261a <=( a45260a  and  a45253a );
 a45265a <=( (not A267)  and  (not A266) );
 a45266a <=( (not A233)  and  a45265a );
 a45269a <=( (not A299)  and  A298 );
 a45272a <=( A301  and  A300 );
 a45273a <=( a45272a  and  a45269a );
 a45274a <=( a45273a  and  a45266a );
 a45278a <=( A167  and  (not A168) );
 a45279a <=( (not A170)  and  a45278a );
 a45282a <=( (not A199)  and  (not A166) );
 a45285a <=( (not A232)  and  A200 );
 a45286a <=( a45285a  and  a45282a );
 a45287a <=( a45286a  and  a45279a );
 a45291a <=( (not A267)  and  (not A266) );
 a45292a <=( (not A233)  and  a45291a );
 a45295a <=( (not A299)  and  A298 );
 a45298a <=( A302  and  A300 );
 a45299a <=( a45298a  and  a45295a );
 a45300a <=( a45299a  and  a45292a );
 a45304a <=( A167  and  (not A168) );
 a45305a <=( (not A170)  and  a45304a );
 a45308a <=( (not A199)  and  (not A166) );
 a45311a <=( (not A232)  and  A200 );
 a45312a <=( a45311a  and  a45308a );
 a45313a <=( a45312a  and  a45305a );
 a45317a <=( (not A266)  and  (not A265) );
 a45318a <=( (not A233)  and  a45317a );
 a45321a <=( (not A299)  and  A298 );
 a45324a <=( A301  and  A300 );
 a45325a <=( a45324a  and  a45321a );
 a45326a <=( a45325a  and  a45318a );
 a45330a <=( A167  and  (not A168) );
 a45331a <=( (not A170)  and  a45330a );
 a45334a <=( (not A199)  and  (not A166) );
 a45337a <=( (not A232)  and  A200 );
 a45338a <=( a45337a  and  a45334a );
 a45339a <=( a45338a  and  a45331a );
 a45343a <=( (not A266)  and  (not A265) );
 a45344a <=( (not A233)  and  a45343a );
 a45347a <=( (not A299)  and  A298 );
 a45350a <=( A302  and  A300 );
 a45351a <=( a45350a  and  a45347a );
 a45352a <=( a45351a  and  a45344a );
 a45356a <=( (not A167)  and  (not A168) );
 a45357a <=( (not A170)  and  a45356a );
 a45360a <=( (not A199)  and  A166 );
 a45363a <=( A232  and  A200 );
 a45364a <=( a45363a  and  a45360a );
 a45365a <=( a45364a  and  a45357a );
 a45369a <=( (not A267)  and  A265 );
 a45370a <=( A233  and  a45369a );
 a45373a <=( (not A299)  and  A298 );
 a45376a <=( A301  and  A300 );
 a45377a <=( a45376a  and  a45373a );
 a45378a <=( a45377a  and  a45370a );
 a45382a <=( (not A167)  and  (not A168) );
 a45383a <=( (not A170)  and  a45382a );
 a45386a <=( (not A199)  and  A166 );
 a45389a <=( A232  and  A200 );
 a45390a <=( a45389a  and  a45386a );
 a45391a <=( a45390a  and  a45383a );
 a45395a <=( (not A267)  and  A265 );
 a45396a <=( A233  and  a45395a );
 a45399a <=( (not A299)  and  A298 );
 a45402a <=( A302  and  A300 );
 a45403a <=( a45402a  and  a45399a );
 a45404a <=( a45403a  and  a45396a );
 a45408a <=( (not A167)  and  (not A168) );
 a45409a <=( (not A170)  and  a45408a );
 a45412a <=( (not A199)  and  A166 );
 a45415a <=( A232  and  A200 );
 a45416a <=( a45415a  and  a45412a );
 a45417a <=( a45416a  and  a45409a );
 a45421a <=( A266  and  A265 );
 a45422a <=( A233  and  a45421a );
 a45425a <=( (not A299)  and  A298 );
 a45428a <=( A301  and  A300 );
 a45429a <=( a45428a  and  a45425a );
 a45430a <=( a45429a  and  a45422a );
 a45434a <=( (not A167)  and  (not A168) );
 a45435a <=( (not A170)  and  a45434a );
 a45438a <=( (not A199)  and  A166 );
 a45441a <=( A232  and  A200 );
 a45442a <=( a45441a  and  a45438a );
 a45443a <=( a45442a  and  a45435a );
 a45447a <=( A266  and  A265 );
 a45448a <=( A233  and  a45447a );
 a45451a <=( (not A299)  and  A298 );
 a45454a <=( A302  and  A300 );
 a45455a <=( a45454a  and  a45451a );
 a45456a <=( a45455a  and  a45448a );
 a45460a <=( (not A167)  and  (not A168) );
 a45461a <=( (not A170)  and  a45460a );
 a45464a <=( (not A199)  and  A166 );
 a45467a <=( A232  and  A200 );
 a45468a <=( a45467a  and  a45464a );
 a45469a <=( a45468a  and  a45461a );
 a45473a <=( (not A266)  and  (not A265) );
 a45474a <=( A233  and  a45473a );
 a45477a <=( (not A299)  and  A298 );
 a45480a <=( A301  and  A300 );
 a45481a <=( a45480a  and  a45477a );
 a45482a <=( a45481a  and  a45474a );
 a45486a <=( (not A167)  and  (not A168) );
 a45487a <=( (not A170)  and  a45486a );
 a45490a <=( (not A199)  and  A166 );
 a45493a <=( A232  and  A200 );
 a45494a <=( a45493a  and  a45490a );
 a45495a <=( a45494a  and  a45487a );
 a45499a <=( (not A266)  and  (not A265) );
 a45500a <=( A233  and  a45499a );
 a45503a <=( (not A299)  and  A298 );
 a45506a <=( A302  and  A300 );
 a45507a <=( a45506a  and  a45503a );
 a45508a <=( a45507a  and  a45500a );
 a45512a <=( (not A167)  and  (not A168) );
 a45513a <=( (not A170)  and  a45512a );
 a45516a <=( (not A199)  and  A166 );
 a45519a <=( (not A233)  and  A200 );
 a45520a <=( a45519a  and  a45516a );
 a45521a <=( a45520a  and  a45513a );
 a45525a <=( (not A266)  and  (not A236) );
 a45526a <=( (not A235)  and  a45525a );
 a45529a <=( (not A269)  and  (not A268) );
 a45532a <=( A299  and  (not A298) );
 a45533a <=( a45532a  and  a45529a );
 a45534a <=( a45533a  and  a45526a );
 a45538a <=( (not A167)  and  (not A168) );
 a45539a <=( (not A170)  and  a45538a );
 a45542a <=( (not A199)  and  A166 );
 a45545a <=( (not A233)  and  A200 );
 a45546a <=( a45545a  and  a45542a );
 a45547a <=( a45546a  and  a45539a );
 a45551a <=( A266  and  A265 );
 a45552a <=( (not A234)  and  a45551a );
 a45555a <=( (not A299)  and  A298 );
 a45558a <=( A301  and  A300 );
 a45559a <=( a45558a  and  a45555a );
 a45560a <=( a45559a  and  a45552a );
 a45564a <=( (not A167)  and  (not A168) );
 a45565a <=( (not A170)  and  a45564a );
 a45568a <=( (not A199)  and  A166 );
 a45571a <=( (not A233)  and  A200 );
 a45572a <=( a45571a  and  a45568a );
 a45573a <=( a45572a  and  a45565a );
 a45577a <=( A266  and  A265 );
 a45578a <=( (not A234)  and  a45577a );
 a45581a <=( (not A299)  and  A298 );
 a45584a <=( A302  and  A300 );
 a45585a <=( a45584a  and  a45581a );
 a45586a <=( a45585a  and  a45578a );
 a45590a <=( (not A167)  and  (not A168) );
 a45591a <=( (not A170)  and  a45590a );
 a45594a <=( (not A199)  and  A166 );
 a45597a <=( (not A233)  and  A200 );
 a45598a <=( a45597a  and  a45594a );
 a45599a <=( a45598a  and  a45591a );
 a45603a <=( (not A267)  and  (not A266) );
 a45604a <=( (not A234)  and  a45603a );
 a45607a <=( (not A299)  and  A298 );
 a45610a <=( A301  and  A300 );
 a45611a <=( a45610a  and  a45607a );
 a45612a <=( a45611a  and  a45604a );
 a45616a <=( (not A167)  and  (not A168) );
 a45617a <=( (not A170)  and  a45616a );
 a45620a <=( (not A199)  and  A166 );
 a45623a <=( (not A233)  and  A200 );
 a45624a <=( a45623a  and  a45620a );
 a45625a <=( a45624a  and  a45617a );
 a45629a <=( (not A267)  and  (not A266) );
 a45630a <=( (not A234)  and  a45629a );
 a45633a <=( (not A299)  and  A298 );
 a45636a <=( A302  and  A300 );
 a45637a <=( a45636a  and  a45633a );
 a45638a <=( a45637a  and  a45630a );
 a45642a <=( (not A167)  and  (not A168) );
 a45643a <=( (not A170)  and  a45642a );
 a45646a <=( (not A199)  and  A166 );
 a45649a <=( (not A233)  and  A200 );
 a45650a <=( a45649a  and  a45646a );
 a45651a <=( a45650a  and  a45643a );
 a45655a <=( (not A266)  and  (not A265) );
 a45656a <=( (not A234)  and  a45655a );
 a45659a <=( (not A299)  and  A298 );
 a45662a <=( A301  and  A300 );
 a45663a <=( a45662a  and  a45659a );
 a45664a <=( a45663a  and  a45656a );
 a45668a <=( (not A167)  and  (not A168) );
 a45669a <=( (not A170)  and  a45668a );
 a45672a <=( (not A199)  and  A166 );
 a45675a <=( (not A233)  and  A200 );
 a45676a <=( a45675a  and  a45672a );
 a45677a <=( a45676a  and  a45669a );
 a45681a <=( (not A266)  and  (not A265) );
 a45682a <=( (not A234)  and  a45681a );
 a45685a <=( (not A299)  and  A298 );
 a45688a <=( A302  and  A300 );
 a45689a <=( a45688a  and  a45685a );
 a45690a <=( a45689a  and  a45682a );
 a45694a <=( (not A167)  and  (not A168) );
 a45695a <=( (not A170)  and  a45694a );
 a45698a <=( (not A199)  and  A166 );
 a45701a <=( A232  and  A200 );
 a45702a <=( a45701a  and  a45698a );
 a45703a <=( a45702a  and  a45695a );
 a45707a <=( A235  and  A234 );
 a45708a <=( (not A233)  and  a45707a );
 a45711a <=( (not A266)  and  A265 );
 a45714a <=( A268  and  A267 );
 a45715a <=( a45714a  and  a45711a );
 a45716a <=( a45715a  and  a45708a );
 a45720a <=( (not A167)  and  (not A168) );
 a45721a <=( (not A170)  and  a45720a );
 a45724a <=( (not A199)  and  A166 );
 a45727a <=( A232  and  A200 );
 a45728a <=( a45727a  and  a45724a );
 a45729a <=( a45728a  and  a45721a );
 a45733a <=( A235  and  A234 );
 a45734a <=( (not A233)  and  a45733a );
 a45737a <=( (not A266)  and  A265 );
 a45740a <=( A269  and  A267 );
 a45741a <=( a45740a  and  a45737a );
 a45742a <=( a45741a  and  a45734a );
 a45746a <=( (not A167)  and  (not A168) );
 a45747a <=( (not A170)  and  a45746a );
 a45750a <=( (not A199)  and  A166 );
 a45753a <=( A232  and  A200 );
 a45754a <=( a45753a  and  a45750a );
 a45755a <=( a45754a  and  a45747a );
 a45759a <=( A236  and  A234 );
 a45760a <=( (not A233)  and  a45759a );
 a45763a <=( (not A266)  and  A265 );
 a45766a <=( A268  and  A267 );
 a45767a <=( a45766a  and  a45763a );
 a45768a <=( a45767a  and  a45760a );
 a45772a <=( (not A167)  and  (not A168) );
 a45773a <=( (not A170)  and  a45772a );
 a45776a <=( (not A199)  and  A166 );
 a45779a <=( A232  and  A200 );
 a45780a <=( a45779a  and  a45776a );
 a45781a <=( a45780a  and  a45773a );
 a45785a <=( A236  and  A234 );
 a45786a <=( (not A233)  and  a45785a );
 a45789a <=( (not A266)  and  A265 );
 a45792a <=( A269  and  A267 );
 a45793a <=( a45792a  and  a45789a );
 a45794a <=( a45793a  and  a45786a );
 a45798a <=( (not A167)  and  (not A168) );
 a45799a <=( (not A170)  and  a45798a );
 a45802a <=( (not A199)  and  A166 );
 a45805a <=( (not A232)  and  A200 );
 a45806a <=( a45805a  and  a45802a );
 a45807a <=( a45806a  and  a45799a );
 a45811a <=( A266  and  A265 );
 a45812a <=( (not A233)  and  a45811a );
 a45815a <=( (not A299)  and  A298 );
 a45818a <=( A301  and  A300 );
 a45819a <=( a45818a  and  a45815a );
 a45820a <=( a45819a  and  a45812a );
 a45824a <=( (not A167)  and  (not A168) );
 a45825a <=( (not A170)  and  a45824a );
 a45828a <=( (not A199)  and  A166 );
 a45831a <=( (not A232)  and  A200 );
 a45832a <=( a45831a  and  a45828a );
 a45833a <=( a45832a  and  a45825a );
 a45837a <=( A266  and  A265 );
 a45838a <=( (not A233)  and  a45837a );
 a45841a <=( (not A299)  and  A298 );
 a45844a <=( A302  and  A300 );
 a45845a <=( a45844a  and  a45841a );
 a45846a <=( a45845a  and  a45838a );
 a45850a <=( (not A167)  and  (not A168) );
 a45851a <=( (not A170)  and  a45850a );
 a45854a <=( (not A199)  and  A166 );
 a45857a <=( (not A232)  and  A200 );
 a45858a <=( a45857a  and  a45854a );
 a45859a <=( a45858a  and  a45851a );
 a45863a <=( (not A267)  and  (not A266) );
 a45864a <=( (not A233)  and  a45863a );
 a45867a <=( (not A299)  and  A298 );
 a45870a <=( A301  and  A300 );
 a45871a <=( a45870a  and  a45867a );
 a45872a <=( a45871a  and  a45864a );
 a45876a <=( (not A167)  and  (not A168) );
 a45877a <=( (not A170)  and  a45876a );
 a45880a <=( (not A199)  and  A166 );
 a45883a <=( (not A232)  and  A200 );
 a45884a <=( a45883a  and  a45880a );
 a45885a <=( a45884a  and  a45877a );
 a45889a <=( (not A267)  and  (not A266) );
 a45890a <=( (not A233)  and  a45889a );
 a45893a <=( (not A299)  and  A298 );
 a45896a <=( A302  and  A300 );
 a45897a <=( a45896a  and  a45893a );
 a45898a <=( a45897a  and  a45890a );
 a45902a <=( (not A167)  and  (not A168) );
 a45903a <=( (not A170)  and  a45902a );
 a45906a <=( (not A199)  and  A166 );
 a45909a <=( (not A232)  and  A200 );
 a45910a <=( a45909a  and  a45906a );
 a45911a <=( a45910a  and  a45903a );
 a45915a <=( (not A266)  and  (not A265) );
 a45916a <=( (not A233)  and  a45915a );
 a45919a <=( (not A299)  and  A298 );
 a45922a <=( A301  and  A300 );
 a45923a <=( a45922a  and  a45919a );
 a45924a <=( a45923a  and  a45916a );
 a45928a <=( (not A167)  and  (not A168) );
 a45929a <=( (not A170)  and  a45928a );
 a45932a <=( (not A199)  and  A166 );
 a45935a <=( (not A232)  and  A200 );
 a45936a <=( a45935a  and  a45932a );
 a45937a <=( a45936a  and  a45929a );
 a45941a <=( (not A266)  and  (not A265) );
 a45942a <=( (not A233)  and  a45941a );
 a45945a <=( (not A299)  and  A298 );
 a45948a <=( A302  and  A300 );
 a45949a <=( a45948a  and  a45945a );
 a45950a <=( a45949a  and  a45942a );
 a45954a <=( A167  and  (not A168) );
 a45955a <=( A169  and  a45954a );
 a45958a <=( (not A199)  and  (not A166) );
 a45961a <=( A232  and  A200 );
 a45962a <=( a45961a  and  a45958a );
 a45963a <=( a45962a  and  a45955a );
 a45967a <=( (not A267)  and  A265 );
 a45968a <=( A233  and  a45967a );
 a45971a <=( (not A299)  and  A298 );
 a45974a <=( A301  and  A300 );
 a45975a <=( a45974a  and  a45971a );
 a45976a <=( a45975a  and  a45968a );
 a45980a <=( A167  and  (not A168) );
 a45981a <=( A169  and  a45980a );
 a45984a <=( (not A199)  and  (not A166) );
 a45987a <=( A232  and  A200 );
 a45988a <=( a45987a  and  a45984a );
 a45989a <=( a45988a  and  a45981a );
 a45993a <=( (not A267)  and  A265 );
 a45994a <=( A233  and  a45993a );
 a45997a <=( (not A299)  and  A298 );
 a46000a <=( A302  and  A300 );
 a46001a <=( a46000a  and  a45997a );
 a46002a <=( a46001a  and  a45994a );
 a46006a <=( A167  and  (not A168) );
 a46007a <=( A169  and  a46006a );
 a46010a <=( (not A199)  and  (not A166) );
 a46013a <=( A232  and  A200 );
 a46014a <=( a46013a  and  a46010a );
 a46015a <=( a46014a  and  a46007a );
 a46019a <=( A266  and  A265 );
 a46020a <=( A233  and  a46019a );
 a46023a <=( (not A299)  and  A298 );
 a46026a <=( A301  and  A300 );
 a46027a <=( a46026a  and  a46023a );
 a46028a <=( a46027a  and  a46020a );
 a46032a <=( A167  and  (not A168) );
 a46033a <=( A169  and  a46032a );
 a46036a <=( (not A199)  and  (not A166) );
 a46039a <=( A232  and  A200 );
 a46040a <=( a46039a  and  a46036a );
 a46041a <=( a46040a  and  a46033a );
 a46045a <=( A266  and  A265 );
 a46046a <=( A233  and  a46045a );
 a46049a <=( (not A299)  and  A298 );
 a46052a <=( A302  and  A300 );
 a46053a <=( a46052a  and  a46049a );
 a46054a <=( a46053a  and  a46046a );
 a46058a <=( A167  and  (not A168) );
 a46059a <=( A169  and  a46058a );
 a46062a <=( (not A199)  and  (not A166) );
 a46065a <=( A232  and  A200 );
 a46066a <=( a46065a  and  a46062a );
 a46067a <=( a46066a  and  a46059a );
 a46071a <=( (not A266)  and  (not A265) );
 a46072a <=( A233  and  a46071a );
 a46075a <=( (not A299)  and  A298 );
 a46078a <=( A301  and  A300 );
 a46079a <=( a46078a  and  a46075a );
 a46080a <=( a46079a  and  a46072a );
 a46084a <=( A167  and  (not A168) );
 a46085a <=( A169  and  a46084a );
 a46088a <=( (not A199)  and  (not A166) );
 a46091a <=( A232  and  A200 );
 a46092a <=( a46091a  and  a46088a );
 a46093a <=( a46092a  and  a46085a );
 a46097a <=( (not A266)  and  (not A265) );
 a46098a <=( A233  and  a46097a );
 a46101a <=( (not A299)  and  A298 );
 a46104a <=( A302  and  A300 );
 a46105a <=( a46104a  and  a46101a );
 a46106a <=( a46105a  and  a46098a );
 a46110a <=( A167  and  (not A168) );
 a46111a <=( A169  and  a46110a );
 a46114a <=( (not A199)  and  (not A166) );
 a46117a <=( (not A233)  and  A200 );
 a46118a <=( a46117a  and  a46114a );
 a46119a <=( a46118a  and  a46111a );
 a46123a <=( (not A266)  and  (not A236) );
 a46124a <=( (not A235)  and  a46123a );
 a46127a <=( (not A269)  and  (not A268) );
 a46130a <=( A299  and  (not A298) );
 a46131a <=( a46130a  and  a46127a );
 a46132a <=( a46131a  and  a46124a );
 a46136a <=( A167  and  (not A168) );
 a46137a <=( A169  and  a46136a );
 a46140a <=( (not A199)  and  (not A166) );
 a46143a <=( (not A233)  and  A200 );
 a46144a <=( a46143a  and  a46140a );
 a46145a <=( a46144a  and  a46137a );
 a46149a <=( A266  and  A265 );
 a46150a <=( (not A234)  and  a46149a );
 a46153a <=( (not A299)  and  A298 );
 a46156a <=( A301  and  A300 );
 a46157a <=( a46156a  and  a46153a );
 a46158a <=( a46157a  and  a46150a );
 a46162a <=( A167  and  (not A168) );
 a46163a <=( A169  and  a46162a );
 a46166a <=( (not A199)  and  (not A166) );
 a46169a <=( (not A233)  and  A200 );
 a46170a <=( a46169a  and  a46166a );
 a46171a <=( a46170a  and  a46163a );
 a46175a <=( A266  and  A265 );
 a46176a <=( (not A234)  and  a46175a );
 a46179a <=( (not A299)  and  A298 );
 a46182a <=( A302  and  A300 );
 a46183a <=( a46182a  and  a46179a );
 a46184a <=( a46183a  and  a46176a );
 a46188a <=( A167  and  (not A168) );
 a46189a <=( A169  and  a46188a );
 a46192a <=( (not A199)  and  (not A166) );
 a46195a <=( (not A233)  and  A200 );
 a46196a <=( a46195a  and  a46192a );
 a46197a <=( a46196a  and  a46189a );
 a46201a <=( (not A267)  and  (not A266) );
 a46202a <=( (not A234)  and  a46201a );
 a46205a <=( (not A299)  and  A298 );
 a46208a <=( A301  and  A300 );
 a46209a <=( a46208a  and  a46205a );
 a46210a <=( a46209a  and  a46202a );
 a46214a <=( A167  and  (not A168) );
 a46215a <=( A169  and  a46214a );
 a46218a <=( (not A199)  and  (not A166) );
 a46221a <=( (not A233)  and  A200 );
 a46222a <=( a46221a  and  a46218a );
 a46223a <=( a46222a  and  a46215a );
 a46227a <=( (not A267)  and  (not A266) );
 a46228a <=( (not A234)  and  a46227a );
 a46231a <=( (not A299)  and  A298 );
 a46234a <=( A302  and  A300 );
 a46235a <=( a46234a  and  a46231a );
 a46236a <=( a46235a  and  a46228a );
 a46240a <=( A167  and  (not A168) );
 a46241a <=( A169  and  a46240a );
 a46244a <=( (not A199)  and  (not A166) );
 a46247a <=( (not A233)  and  A200 );
 a46248a <=( a46247a  and  a46244a );
 a46249a <=( a46248a  and  a46241a );
 a46253a <=( (not A266)  and  (not A265) );
 a46254a <=( (not A234)  and  a46253a );
 a46257a <=( (not A299)  and  A298 );
 a46260a <=( A301  and  A300 );
 a46261a <=( a46260a  and  a46257a );
 a46262a <=( a46261a  and  a46254a );
 a46266a <=( A167  and  (not A168) );
 a46267a <=( A169  and  a46266a );
 a46270a <=( (not A199)  and  (not A166) );
 a46273a <=( (not A233)  and  A200 );
 a46274a <=( a46273a  and  a46270a );
 a46275a <=( a46274a  and  a46267a );
 a46279a <=( (not A266)  and  (not A265) );
 a46280a <=( (not A234)  and  a46279a );
 a46283a <=( (not A299)  and  A298 );
 a46286a <=( A302  and  A300 );
 a46287a <=( a46286a  and  a46283a );
 a46288a <=( a46287a  and  a46280a );
 a46292a <=( A167  and  (not A168) );
 a46293a <=( A169  and  a46292a );
 a46296a <=( (not A199)  and  (not A166) );
 a46299a <=( A232  and  A200 );
 a46300a <=( a46299a  and  a46296a );
 a46301a <=( a46300a  and  a46293a );
 a46305a <=( A235  and  A234 );
 a46306a <=( (not A233)  and  a46305a );
 a46309a <=( (not A266)  and  A265 );
 a46312a <=( A268  and  A267 );
 a46313a <=( a46312a  and  a46309a );
 a46314a <=( a46313a  and  a46306a );
 a46318a <=( A167  and  (not A168) );
 a46319a <=( A169  and  a46318a );
 a46322a <=( (not A199)  and  (not A166) );
 a46325a <=( A232  and  A200 );
 a46326a <=( a46325a  and  a46322a );
 a46327a <=( a46326a  and  a46319a );
 a46331a <=( A235  and  A234 );
 a46332a <=( (not A233)  and  a46331a );
 a46335a <=( (not A266)  and  A265 );
 a46338a <=( A269  and  A267 );
 a46339a <=( a46338a  and  a46335a );
 a46340a <=( a46339a  and  a46332a );
 a46344a <=( A167  and  (not A168) );
 a46345a <=( A169  and  a46344a );
 a46348a <=( (not A199)  and  (not A166) );
 a46351a <=( A232  and  A200 );
 a46352a <=( a46351a  and  a46348a );
 a46353a <=( a46352a  and  a46345a );
 a46357a <=( A236  and  A234 );
 a46358a <=( (not A233)  and  a46357a );
 a46361a <=( (not A266)  and  A265 );
 a46364a <=( A268  and  A267 );
 a46365a <=( a46364a  and  a46361a );
 a46366a <=( a46365a  and  a46358a );
 a46370a <=( A167  and  (not A168) );
 a46371a <=( A169  and  a46370a );
 a46374a <=( (not A199)  and  (not A166) );
 a46377a <=( A232  and  A200 );
 a46378a <=( a46377a  and  a46374a );
 a46379a <=( a46378a  and  a46371a );
 a46383a <=( A236  and  A234 );
 a46384a <=( (not A233)  and  a46383a );
 a46387a <=( (not A266)  and  A265 );
 a46390a <=( A269  and  A267 );
 a46391a <=( a46390a  and  a46387a );
 a46392a <=( a46391a  and  a46384a );
 a46396a <=( A167  and  (not A168) );
 a46397a <=( A169  and  a46396a );
 a46400a <=( (not A199)  and  (not A166) );
 a46403a <=( (not A232)  and  A200 );
 a46404a <=( a46403a  and  a46400a );
 a46405a <=( a46404a  and  a46397a );
 a46409a <=( A266  and  A265 );
 a46410a <=( (not A233)  and  a46409a );
 a46413a <=( (not A299)  and  A298 );
 a46416a <=( A301  and  A300 );
 a46417a <=( a46416a  and  a46413a );
 a46418a <=( a46417a  and  a46410a );
 a46422a <=( A167  and  (not A168) );
 a46423a <=( A169  and  a46422a );
 a46426a <=( (not A199)  and  (not A166) );
 a46429a <=( (not A232)  and  A200 );
 a46430a <=( a46429a  and  a46426a );
 a46431a <=( a46430a  and  a46423a );
 a46435a <=( A266  and  A265 );
 a46436a <=( (not A233)  and  a46435a );
 a46439a <=( (not A299)  and  A298 );
 a46442a <=( A302  and  A300 );
 a46443a <=( a46442a  and  a46439a );
 a46444a <=( a46443a  and  a46436a );
 a46448a <=( A167  and  (not A168) );
 a46449a <=( A169  and  a46448a );
 a46452a <=( (not A199)  and  (not A166) );
 a46455a <=( (not A232)  and  A200 );
 a46456a <=( a46455a  and  a46452a );
 a46457a <=( a46456a  and  a46449a );
 a46461a <=( (not A267)  and  (not A266) );
 a46462a <=( (not A233)  and  a46461a );
 a46465a <=( (not A299)  and  A298 );
 a46468a <=( A301  and  A300 );
 a46469a <=( a46468a  and  a46465a );
 a46470a <=( a46469a  and  a46462a );
 a46474a <=( A167  and  (not A168) );
 a46475a <=( A169  and  a46474a );
 a46478a <=( (not A199)  and  (not A166) );
 a46481a <=( (not A232)  and  A200 );
 a46482a <=( a46481a  and  a46478a );
 a46483a <=( a46482a  and  a46475a );
 a46487a <=( (not A267)  and  (not A266) );
 a46488a <=( (not A233)  and  a46487a );
 a46491a <=( (not A299)  and  A298 );
 a46494a <=( A302  and  A300 );
 a46495a <=( a46494a  and  a46491a );
 a46496a <=( a46495a  and  a46488a );
 a46500a <=( A167  and  (not A168) );
 a46501a <=( A169  and  a46500a );
 a46504a <=( (not A199)  and  (not A166) );
 a46507a <=( (not A232)  and  A200 );
 a46508a <=( a46507a  and  a46504a );
 a46509a <=( a46508a  and  a46501a );
 a46513a <=( (not A266)  and  (not A265) );
 a46514a <=( (not A233)  and  a46513a );
 a46517a <=( (not A299)  and  A298 );
 a46520a <=( A301  and  A300 );
 a46521a <=( a46520a  and  a46517a );
 a46522a <=( a46521a  and  a46514a );
 a46526a <=( A167  and  (not A168) );
 a46527a <=( A169  and  a46526a );
 a46530a <=( (not A199)  and  (not A166) );
 a46533a <=( (not A232)  and  A200 );
 a46534a <=( a46533a  and  a46530a );
 a46535a <=( a46534a  and  a46527a );
 a46539a <=( (not A266)  and  (not A265) );
 a46540a <=( (not A233)  and  a46539a );
 a46543a <=( (not A299)  and  A298 );
 a46546a <=( A302  and  A300 );
 a46547a <=( a46546a  and  a46543a );
 a46548a <=( a46547a  and  a46540a );
 a46552a <=( A167  and  (not A168) );
 a46553a <=( A169  and  a46552a );
 a46556a <=( A199  and  (not A166) );
 a46559a <=( A201  and  (not A200) );
 a46560a <=( a46559a  and  a46556a );
 a46561a <=( a46560a  and  a46553a );
 a46565a <=( A233  and  A232 );
 a46566a <=( A202  and  a46565a );
 a46569a <=( (not A267)  and  A265 );
 a46572a <=( A299  and  (not A298) );
 a46573a <=( a46572a  and  a46569a );
 a46574a <=( a46573a  and  a46566a );
 a46578a <=( A167  and  (not A168) );
 a46579a <=( A169  and  a46578a );
 a46582a <=( A199  and  (not A166) );
 a46585a <=( A201  and  (not A200) );
 a46586a <=( a46585a  and  a46582a );
 a46587a <=( a46586a  and  a46579a );
 a46591a <=( A233  and  A232 );
 a46592a <=( A202  and  a46591a );
 a46595a <=( A266  and  A265 );
 a46598a <=( A299  and  (not A298) );
 a46599a <=( a46598a  and  a46595a );
 a46600a <=( a46599a  and  a46592a );
 a46604a <=( A167  and  (not A168) );
 a46605a <=( A169  and  a46604a );
 a46608a <=( A199  and  (not A166) );
 a46611a <=( A201  and  (not A200) );
 a46612a <=( a46611a  and  a46608a );
 a46613a <=( a46612a  and  a46605a );
 a46617a <=( A233  and  A232 );
 a46618a <=( A202  and  a46617a );
 a46621a <=( (not A266)  and  (not A265) );
 a46624a <=( A299  and  (not A298) );
 a46625a <=( a46624a  and  a46621a );
 a46626a <=( a46625a  and  a46618a );
 a46630a <=( A167  and  (not A168) );
 a46631a <=( A169  and  a46630a );
 a46634a <=( A199  and  (not A166) );
 a46637a <=( A201  and  (not A200) );
 a46638a <=( a46637a  and  a46634a );
 a46639a <=( a46638a  and  a46631a );
 a46643a <=( A233  and  (not A232) );
 a46644a <=( A202  and  a46643a );
 a46647a <=( (not A266)  and  A265 );
 a46650a <=( A268  and  A267 );
 a46651a <=( a46650a  and  a46647a );
 a46652a <=( a46651a  and  a46644a );
 a46656a <=( A167  and  (not A168) );
 a46657a <=( A169  and  a46656a );
 a46660a <=( A199  and  (not A166) );
 a46663a <=( A201  and  (not A200) );
 a46664a <=( a46663a  and  a46660a );
 a46665a <=( a46664a  and  a46657a );
 a46669a <=( A233  and  (not A232) );
 a46670a <=( A202  and  a46669a );
 a46673a <=( (not A266)  and  A265 );
 a46676a <=( A269  and  A267 );
 a46677a <=( a46676a  and  a46673a );
 a46678a <=( a46677a  and  a46670a );
 a46682a <=( A167  and  (not A168) );
 a46683a <=( A169  and  a46682a );
 a46686a <=( A199  and  (not A166) );
 a46689a <=( A201  and  (not A200) );
 a46690a <=( a46689a  and  a46686a );
 a46691a <=( a46690a  and  a46683a );
 a46695a <=( (not A234)  and  (not A233) );
 a46696a <=( A202  and  a46695a );
 a46699a <=( A266  and  A265 );
 a46702a <=( A299  and  (not A298) );
 a46703a <=( a46702a  and  a46699a );
 a46704a <=( a46703a  and  a46696a );
 a46708a <=( A167  and  (not A168) );
 a46709a <=( A169  and  a46708a );
 a46712a <=( A199  and  (not A166) );
 a46715a <=( A201  and  (not A200) );
 a46716a <=( a46715a  and  a46712a );
 a46717a <=( a46716a  and  a46709a );
 a46721a <=( (not A234)  and  (not A233) );
 a46722a <=( A202  and  a46721a );
 a46725a <=( (not A267)  and  (not A266) );
 a46728a <=( A299  and  (not A298) );
 a46729a <=( a46728a  and  a46725a );
 a46730a <=( a46729a  and  a46722a );
 a46734a <=( A167  and  (not A168) );
 a46735a <=( A169  and  a46734a );
 a46738a <=( A199  and  (not A166) );
 a46741a <=( A201  and  (not A200) );
 a46742a <=( a46741a  and  a46738a );
 a46743a <=( a46742a  and  a46735a );
 a46747a <=( (not A234)  and  (not A233) );
 a46748a <=( A202  and  a46747a );
 a46751a <=( (not A266)  and  (not A265) );
 a46754a <=( A299  and  (not A298) );
 a46755a <=( a46754a  and  a46751a );
 a46756a <=( a46755a  and  a46748a );
 a46760a <=( A167  and  (not A168) );
 a46761a <=( A169  and  a46760a );
 a46764a <=( A199  and  (not A166) );
 a46767a <=( A201  and  (not A200) );
 a46768a <=( a46767a  and  a46764a );
 a46769a <=( a46768a  and  a46761a );
 a46773a <=( (not A233)  and  A232 );
 a46774a <=( A202  and  a46773a );
 a46777a <=( A235  and  A234 );
 a46780a <=( (not A300)  and  A298 );
 a46781a <=( a46780a  and  a46777a );
 a46782a <=( a46781a  and  a46774a );
 a46786a <=( A167  and  (not A168) );
 a46787a <=( A169  and  a46786a );
 a46790a <=( A199  and  (not A166) );
 a46793a <=( A201  and  (not A200) );
 a46794a <=( a46793a  and  a46790a );
 a46795a <=( a46794a  and  a46787a );
 a46799a <=( (not A233)  and  A232 );
 a46800a <=( A202  and  a46799a );
 a46803a <=( A235  and  A234 );
 a46806a <=( A299  and  A298 );
 a46807a <=( a46806a  and  a46803a );
 a46808a <=( a46807a  and  a46800a );
 a46812a <=( A167  and  (not A168) );
 a46813a <=( A169  and  a46812a );
 a46816a <=( A199  and  (not A166) );
 a46819a <=( A201  and  (not A200) );
 a46820a <=( a46819a  and  a46816a );
 a46821a <=( a46820a  and  a46813a );
 a46825a <=( (not A233)  and  A232 );
 a46826a <=( A202  and  a46825a );
 a46829a <=( A235  and  A234 );
 a46832a <=( (not A299)  and  (not A298) );
 a46833a <=( a46832a  and  a46829a );
 a46834a <=( a46833a  and  a46826a );
 a46838a <=( A167  and  (not A168) );
 a46839a <=( A169  and  a46838a );
 a46842a <=( A199  and  (not A166) );
 a46845a <=( A201  and  (not A200) );
 a46846a <=( a46845a  and  a46842a );
 a46847a <=( a46846a  and  a46839a );
 a46851a <=( (not A233)  and  A232 );
 a46852a <=( A202  and  a46851a );
 a46855a <=( A235  and  A234 );
 a46858a <=( A266  and  (not A265) );
 a46859a <=( a46858a  and  a46855a );
 a46860a <=( a46859a  and  a46852a );
 a46864a <=( A167  and  (not A168) );
 a46865a <=( A169  and  a46864a );
 a46868a <=( A199  and  (not A166) );
 a46871a <=( A201  and  (not A200) );
 a46872a <=( a46871a  and  a46868a );
 a46873a <=( a46872a  and  a46865a );
 a46877a <=( (not A233)  and  A232 );
 a46878a <=( A202  and  a46877a );
 a46881a <=( A236  and  A234 );
 a46884a <=( (not A300)  and  A298 );
 a46885a <=( a46884a  and  a46881a );
 a46886a <=( a46885a  and  a46878a );
 a46890a <=( A167  and  (not A168) );
 a46891a <=( A169  and  a46890a );
 a46894a <=( A199  and  (not A166) );
 a46897a <=( A201  and  (not A200) );
 a46898a <=( a46897a  and  a46894a );
 a46899a <=( a46898a  and  a46891a );
 a46903a <=( (not A233)  and  A232 );
 a46904a <=( A202  and  a46903a );
 a46907a <=( A236  and  A234 );
 a46910a <=( A299  and  A298 );
 a46911a <=( a46910a  and  a46907a );
 a46912a <=( a46911a  and  a46904a );
 a46916a <=( A167  and  (not A168) );
 a46917a <=( A169  and  a46916a );
 a46920a <=( A199  and  (not A166) );
 a46923a <=( A201  and  (not A200) );
 a46924a <=( a46923a  and  a46920a );
 a46925a <=( a46924a  and  a46917a );
 a46929a <=( (not A233)  and  A232 );
 a46930a <=( A202  and  a46929a );
 a46933a <=( A236  and  A234 );
 a46936a <=( (not A299)  and  (not A298) );
 a46937a <=( a46936a  and  a46933a );
 a46938a <=( a46937a  and  a46930a );
 a46942a <=( A167  and  (not A168) );
 a46943a <=( A169  and  a46942a );
 a46946a <=( A199  and  (not A166) );
 a46949a <=( A201  and  (not A200) );
 a46950a <=( a46949a  and  a46946a );
 a46951a <=( a46950a  and  a46943a );
 a46955a <=( (not A233)  and  A232 );
 a46956a <=( A202  and  a46955a );
 a46959a <=( A236  and  A234 );
 a46962a <=( A266  and  (not A265) );
 a46963a <=( a46962a  and  a46959a );
 a46964a <=( a46963a  and  a46956a );
 a46968a <=( A167  and  (not A168) );
 a46969a <=( A169  and  a46968a );
 a46972a <=( A199  and  (not A166) );
 a46975a <=( A201  and  (not A200) );
 a46976a <=( a46975a  and  a46972a );
 a46977a <=( a46976a  and  a46969a );
 a46981a <=( (not A233)  and  (not A232) );
 a46982a <=( A202  and  a46981a );
 a46985a <=( A266  and  A265 );
 a46988a <=( A299  and  (not A298) );
 a46989a <=( a46988a  and  a46985a );
 a46990a <=( a46989a  and  a46982a );
 a46994a <=( A167  and  (not A168) );
 a46995a <=( A169  and  a46994a );
 a46998a <=( A199  and  (not A166) );
 a47001a <=( A201  and  (not A200) );
 a47002a <=( a47001a  and  a46998a );
 a47003a <=( a47002a  and  a46995a );
 a47007a <=( (not A233)  and  (not A232) );
 a47008a <=( A202  and  a47007a );
 a47011a <=( (not A267)  and  (not A266) );
 a47014a <=( A299  and  (not A298) );
 a47015a <=( a47014a  and  a47011a );
 a47016a <=( a47015a  and  a47008a );
 a47020a <=( A167  and  (not A168) );
 a47021a <=( A169  and  a47020a );
 a47024a <=( A199  and  (not A166) );
 a47027a <=( A201  and  (not A200) );
 a47028a <=( a47027a  and  a47024a );
 a47029a <=( a47028a  and  a47021a );
 a47033a <=( (not A233)  and  (not A232) );
 a47034a <=( A202  and  a47033a );
 a47037a <=( (not A266)  and  (not A265) );
 a47040a <=( A299  and  (not A298) );
 a47041a <=( a47040a  and  a47037a );
 a47042a <=( a47041a  and  a47034a );
 a47046a <=( A167  and  (not A168) );
 a47047a <=( A169  and  a47046a );
 a47050a <=( A199  and  (not A166) );
 a47053a <=( A201  and  (not A200) );
 a47054a <=( a47053a  and  a47050a );
 a47055a <=( a47054a  and  a47047a );
 a47059a <=( A233  and  A232 );
 a47060a <=( A203  and  a47059a );
 a47063a <=( (not A267)  and  A265 );
 a47066a <=( A299  and  (not A298) );
 a47067a <=( a47066a  and  a47063a );
 a47068a <=( a47067a  and  a47060a );
 a47072a <=( A167  and  (not A168) );
 a47073a <=( A169  and  a47072a );
 a47076a <=( A199  and  (not A166) );
 a47079a <=( A201  and  (not A200) );
 a47080a <=( a47079a  and  a47076a );
 a47081a <=( a47080a  and  a47073a );
 a47085a <=( A233  and  A232 );
 a47086a <=( A203  and  a47085a );
 a47089a <=( A266  and  A265 );
 a47092a <=( A299  and  (not A298) );
 a47093a <=( a47092a  and  a47089a );
 a47094a <=( a47093a  and  a47086a );
 a47098a <=( A167  and  (not A168) );
 a47099a <=( A169  and  a47098a );
 a47102a <=( A199  and  (not A166) );
 a47105a <=( A201  and  (not A200) );
 a47106a <=( a47105a  and  a47102a );
 a47107a <=( a47106a  and  a47099a );
 a47111a <=( A233  and  A232 );
 a47112a <=( A203  and  a47111a );
 a47115a <=( (not A266)  and  (not A265) );
 a47118a <=( A299  and  (not A298) );
 a47119a <=( a47118a  and  a47115a );
 a47120a <=( a47119a  and  a47112a );
 a47124a <=( A167  and  (not A168) );
 a47125a <=( A169  and  a47124a );
 a47128a <=( A199  and  (not A166) );
 a47131a <=( A201  and  (not A200) );
 a47132a <=( a47131a  and  a47128a );
 a47133a <=( a47132a  and  a47125a );
 a47137a <=( A233  and  (not A232) );
 a47138a <=( A203  and  a47137a );
 a47141a <=( (not A266)  and  A265 );
 a47144a <=( A268  and  A267 );
 a47145a <=( a47144a  and  a47141a );
 a47146a <=( a47145a  and  a47138a );
 a47150a <=( A167  and  (not A168) );
 a47151a <=( A169  and  a47150a );
 a47154a <=( A199  and  (not A166) );
 a47157a <=( A201  and  (not A200) );
 a47158a <=( a47157a  and  a47154a );
 a47159a <=( a47158a  and  a47151a );
 a47163a <=( A233  and  (not A232) );
 a47164a <=( A203  and  a47163a );
 a47167a <=( (not A266)  and  A265 );
 a47170a <=( A269  and  A267 );
 a47171a <=( a47170a  and  a47167a );
 a47172a <=( a47171a  and  a47164a );
 a47176a <=( A167  and  (not A168) );
 a47177a <=( A169  and  a47176a );
 a47180a <=( A199  and  (not A166) );
 a47183a <=( A201  and  (not A200) );
 a47184a <=( a47183a  and  a47180a );
 a47185a <=( a47184a  and  a47177a );
 a47189a <=( (not A234)  and  (not A233) );
 a47190a <=( A203  and  a47189a );
 a47193a <=( A266  and  A265 );
 a47196a <=( A299  and  (not A298) );
 a47197a <=( a47196a  and  a47193a );
 a47198a <=( a47197a  and  a47190a );
 a47202a <=( A167  and  (not A168) );
 a47203a <=( A169  and  a47202a );
 a47206a <=( A199  and  (not A166) );
 a47209a <=( A201  and  (not A200) );
 a47210a <=( a47209a  and  a47206a );
 a47211a <=( a47210a  and  a47203a );
 a47215a <=( (not A234)  and  (not A233) );
 a47216a <=( A203  and  a47215a );
 a47219a <=( (not A267)  and  (not A266) );
 a47222a <=( A299  and  (not A298) );
 a47223a <=( a47222a  and  a47219a );
 a47224a <=( a47223a  and  a47216a );
 a47228a <=( A167  and  (not A168) );
 a47229a <=( A169  and  a47228a );
 a47232a <=( A199  and  (not A166) );
 a47235a <=( A201  and  (not A200) );
 a47236a <=( a47235a  and  a47232a );
 a47237a <=( a47236a  and  a47229a );
 a47241a <=( (not A234)  and  (not A233) );
 a47242a <=( A203  and  a47241a );
 a47245a <=( (not A266)  and  (not A265) );
 a47248a <=( A299  and  (not A298) );
 a47249a <=( a47248a  and  a47245a );
 a47250a <=( a47249a  and  a47242a );
 a47254a <=( A167  and  (not A168) );
 a47255a <=( A169  and  a47254a );
 a47258a <=( A199  and  (not A166) );
 a47261a <=( A201  and  (not A200) );
 a47262a <=( a47261a  and  a47258a );
 a47263a <=( a47262a  and  a47255a );
 a47267a <=( (not A233)  and  A232 );
 a47268a <=( A203  and  a47267a );
 a47271a <=( A235  and  A234 );
 a47274a <=( (not A300)  and  A298 );
 a47275a <=( a47274a  and  a47271a );
 a47276a <=( a47275a  and  a47268a );
 a47280a <=( A167  and  (not A168) );
 a47281a <=( A169  and  a47280a );
 a47284a <=( A199  and  (not A166) );
 a47287a <=( A201  and  (not A200) );
 a47288a <=( a47287a  and  a47284a );
 a47289a <=( a47288a  and  a47281a );
 a47293a <=( (not A233)  and  A232 );
 a47294a <=( A203  and  a47293a );
 a47297a <=( A235  and  A234 );
 a47300a <=( A299  and  A298 );
 a47301a <=( a47300a  and  a47297a );
 a47302a <=( a47301a  and  a47294a );
 a47306a <=( A167  and  (not A168) );
 a47307a <=( A169  and  a47306a );
 a47310a <=( A199  and  (not A166) );
 a47313a <=( A201  and  (not A200) );
 a47314a <=( a47313a  and  a47310a );
 a47315a <=( a47314a  and  a47307a );
 a47319a <=( (not A233)  and  A232 );
 a47320a <=( A203  and  a47319a );
 a47323a <=( A235  and  A234 );
 a47326a <=( (not A299)  and  (not A298) );
 a47327a <=( a47326a  and  a47323a );
 a47328a <=( a47327a  and  a47320a );
 a47332a <=( A167  and  (not A168) );
 a47333a <=( A169  and  a47332a );
 a47336a <=( A199  and  (not A166) );
 a47339a <=( A201  and  (not A200) );
 a47340a <=( a47339a  and  a47336a );
 a47341a <=( a47340a  and  a47333a );
 a47345a <=( (not A233)  and  A232 );
 a47346a <=( A203  and  a47345a );
 a47349a <=( A235  and  A234 );
 a47352a <=( A266  and  (not A265) );
 a47353a <=( a47352a  and  a47349a );
 a47354a <=( a47353a  and  a47346a );
 a47358a <=( A167  and  (not A168) );
 a47359a <=( A169  and  a47358a );
 a47362a <=( A199  and  (not A166) );
 a47365a <=( A201  and  (not A200) );
 a47366a <=( a47365a  and  a47362a );
 a47367a <=( a47366a  and  a47359a );
 a47371a <=( (not A233)  and  A232 );
 a47372a <=( A203  and  a47371a );
 a47375a <=( A236  and  A234 );
 a47378a <=( (not A300)  and  A298 );
 a47379a <=( a47378a  and  a47375a );
 a47380a <=( a47379a  and  a47372a );
 a47384a <=( A167  and  (not A168) );
 a47385a <=( A169  and  a47384a );
 a47388a <=( A199  and  (not A166) );
 a47391a <=( A201  and  (not A200) );
 a47392a <=( a47391a  and  a47388a );
 a47393a <=( a47392a  and  a47385a );
 a47397a <=( (not A233)  and  A232 );
 a47398a <=( A203  and  a47397a );
 a47401a <=( A236  and  A234 );
 a47404a <=( A299  and  A298 );
 a47405a <=( a47404a  and  a47401a );
 a47406a <=( a47405a  and  a47398a );
 a47410a <=( A167  and  (not A168) );
 a47411a <=( A169  and  a47410a );
 a47414a <=( A199  and  (not A166) );
 a47417a <=( A201  and  (not A200) );
 a47418a <=( a47417a  and  a47414a );
 a47419a <=( a47418a  and  a47411a );
 a47423a <=( (not A233)  and  A232 );
 a47424a <=( A203  and  a47423a );
 a47427a <=( A236  and  A234 );
 a47430a <=( (not A299)  and  (not A298) );
 a47431a <=( a47430a  and  a47427a );
 a47432a <=( a47431a  and  a47424a );
 a47436a <=( A167  and  (not A168) );
 a47437a <=( A169  and  a47436a );
 a47440a <=( A199  and  (not A166) );
 a47443a <=( A201  and  (not A200) );
 a47444a <=( a47443a  and  a47440a );
 a47445a <=( a47444a  and  a47437a );
 a47449a <=( (not A233)  and  A232 );
 a47450a <=( A203  and  a47449a );
 a47453a <=( A236  and  A234 );
 a47456a <=( A266  and  (not A265) );
 a47457a <=( a47456a  and  a47453a );
 a47458a <=( a47457a  and  a47450a );
 a47462a <=( A167  and  (not A168) );
 a47463a <=( A169  and  a47462a );
 a47466a <=( A199  and  (not A166) );
 a47469a <=( A201  and  (not A200) );
 a47470a <=( a47469a  and  a47466a );
 a47471a <=( a47470a  and  a47463a );
 a47475a <=( (not A233)  and  (not A232) );
 a47476a <=( A203  and  a47475a );
 a47479a <=( A266  and  A265 );
 a47482a <=( A299  and  (not A298) );
 a47483a <=( a47482a  and  a47479a );
 a47484a <=( a47483a  and  a47476a );
 a47488a <=( A167  and  (not A168) );
 a47489a <=( A169  and  a47488a );
 a47492a <=( A199  and  (not A166) );
 a47495a <=( A201  and  (not A200) );
 a47496a <=( a47495a  and  a47492a );
 a47497a <=( a47496a  and  a47489a );
 a47501a <=( (not A233)  and  (not A232) );
 a47502a <=( A203  and  a47501a );
 a47505a <=( (not A267)  and  (not A266) );
 a47508a <=( A299  and  (not A298) );
 a47509a <=( a47508a  and  a47505a );
 a47510a <=( a47509a  and  a47502a );
 a47514a <=( A167  and  (not A168) );
 a47515a <=( A169  and  a47514a );
 a47518a <=( A199  and  (not A166) );
 a47521a <=( A201  and  (not A200) );
 a47522a <=( a47521a  and  a47518a );
 a47523a <=( a47522a  and  a47515a );
 a47527a <=( (not A233)  and  (not A232) );
 a47528a <=( A203  and  a47527a );
 a47531a <=( (not A266)  and  (not A265) );
 a47534a <=( A299  and  (not A298) );
 a47535a <=( a47534a  and  a47531a );
 a47536a <=( a47535a  and  a47528a );
 a47540a <=( (not A167)  and  (not A168) );
 a47541a <=( A169  and  a47540a );
 a47544a <=( (not A199)  and  A166 );
 a47547a <=( A232  and  A200 );
 a47548a <=( a47547a  and  a47544a );
 a47549a <=( a47548a  and  a47541a );
 a47553a <=( (not A267)  and  A265 );
 a47554a <=( A233  and  a47553a );
 a47557a <=( (not A299)  and  A298 );
 a47560a <=( A301  and  A300 );
 a47561a <=( a47560a  and  a47557a );
 a47562a <=( a47561a  and  a47554a );
 a47566a <=( (not A167)  and  (not A168) );
 a47567a <=( A169  and  a47566a );
 a47570a <=( (not A199)  and  A166 );
 a47573a <=( A232  and  A200 );
 a47574a <=( a47573a  and  a47570a );
 a47575a <=( a47574a  and  a47567a );
 a47579a <=( (not A267)  and  A265 );
 a47580a <=( A233  and  a47579a );
 a47583a <=( (not A299)  and  A298 );
 a47586a <=( A302  and  A300 );
 a47587a <=( a47586a  and  a47583a );
 a47588a <=( a47587a  and  a47580a );
 a47592a <=( (not A167)  and  (not A168) );
 a47593a <=( A169  and  a47592a );
 a47596a <=( (not A199)  and  A166 );
 a47599a <=( A232  and  A200 );
 a47600a <=( a47599a  and  a47596a );
 a47601a <=( a47600a  and  a47593a );
 a47605a <=( A266  and  A265 );
 a47606a <=( A233  and  a47605a );
 a47609a <=( (not A299)  and  A298 );
 a47612a <=( A301  and  A300 );
 a47613a <=( a47612a  and  a47609a );
 a47614a <=( a47613a  and  a47606a );
 a47618a <=( (not A167)  and  (not A168) );
 a47619a <=( A169  and  a47618a );
 a47622a <=( (not A199)  and  A166 );
 a47625a <=( A232  and  A200 );
 a47626a <=( a47625a  and  a47622a );
 a47627a <=( a47626a  and  a47619a );
 a47631a <=( A266  and  A265 );
 a47632a <=( A233  and  a47631a );
 a47635a <=( (not A299)  and  A298 );
 a47638a <=( A302  and  A300 );
 a47639a <=( a47638a  and  a47635a );
 a47640a <=( a47639a  and  a47632a );
 a47644a <=( (not A167)  and  (not A168) );
 a47645a <=( A169  and  a47644a );
 a47648a <=( (not A199)  and  A166 );
 a47651a <=( A232  and  A200 );
 a47652a <=( a47651a  and  a47648a );
 a47653a <=( a47652a  and  a47645a );
 a47657a <=( (not A266)  and  (not A265) );
 a47658a <=( A233  and  a47657a );
 a47661a <=( (not A299)  and  A298 );
 a47664a <=( A301  and  A300 );
 a47665a <=( a47664a  and  a47661a );
 a47666a <=( a47665a  and  a47658a );
 a47670a <=( (not A167)  and  (not A168) );
 a47671a <=( A169  and  a47670a );
 a47674a <=( (not A199)  and  A166 );
 a47677a <=( A232  and  A200 );
 a47678a <=( a47677a  and  a47674a );
 a47679a <=( a47678a  and  a47671a );
 a47683a <=( (not A266)  and  (not A265) );
 a47684a <=( A233  and  a47683a );
 a47687a <=( (not A299)  and  A298 );
 a47690a <=( A302  and  A300 );
 a47691a <=( a47690a  and  a47687a );
 a47692a <=( a47691a  and  a47684a );
 a47696a <=( (not A167)  and  (not A168) );
 a47697a <=( A169  and  a47696a );
 a47700a <=( (not A199)  and  A166 );
 a47703a <=( (not A233)  and  A200 );
 a47704a <=( a47703a  and  a47700a );
 a47705a <=( a47704a  and  a47697a );
 a47709a <=( (not A266)  and  (not A236) );
 a47710a <=( (not A235)  and  a47709a );
 a47713a <=( (not A269)  and  (not A268) );
 a47716a <=( A299  and  (not A298) );
 a47717a <=( a47716a  and  a47713a );
 a47718a <=( a47717a  and  a47710a );
 a47722a <=( (not A167)  and  (not A168) );
 a47723a <=( A169  and  a47722a );
 a47726a <=( (not A199)  and  A166 );
 a47729a <=( (not A233)  and  A200 );
 a47730a <=( a47729a  and  a47726a );
 a47731a <=( a47730a  and  a47723a );
 a47735a <=( A266  and  A265 );
 a47736a <=( (not A234)  and  a47735a );
 a47739a <=( (not A299)  and  A298 );
 a47742a <=( A301  and  A300 );
 a47743a <=( a47742a  and  a47739a );
 a47744a <=( a47743a  and  a47736a );
 a47748a <=( (not A167)  and  (not A168) );
 a47749a <=( A169  and  a47748a );
 a47752a <=( (not A199)  and  A166 );
 a47755a <=( (not A233)  and  A200 );
 a47756a <=( a47755a  and  a47752a );
 a47757a <=( a47756a  and  a47749a );
 a47761a <=( A266  and  A265 );
 a47762a <=( (not A234)  and  a47761a );
 a47765a <=( (not A299)  and  A298 );
 a47768a <=( A302  and  A300 );
 a47769a <=( a47768a  and  a47765a );
 a47770a <=( a47769a  and  a47762a );
 a47774a <=( (not A167)  and  (not A168) );
 a47775a <=( A169  and  a47774a );
 a47778a <=( (not A199)  and  A166 );
 a47781a <=( (not A233)  and  A200 );
 a47782a <=( a47781a  and  a47778a );
 a47783a <=( a47782a  and  a47775a );
 a47787a <=( (not A267)  and  (not A266) );
 a47788a <=( (not A234)  and  a47787a );
 a47791a <=( (not A299)  and  A298 );
 a47794a <=( A301  and  A300 );
 a47795a <=( a47794a  and  a47791a );
 a47796a <=( a47795a  and  a47788a );
 a47800a <=( (not A167)  and  (not A168) );
 a47801a <=( A169  and  a47800a );
 a47804a <=( (not A199)  and  A166 );
 a47807a <=( (not A233)  and  A200 );
 a47808a <=( a47807a  and  a47804a );
 a47809a <=( a47808a  and  a47801a );
 a47813a <=( (not A267)  and  (not A266) );
 a47814a <=( (not A234)  and  a47813a );
 a47817a <=( (not A299)  and  A298 );
 a47820a <=( A302  and  A300 );
 a47821a <=( a47820a  and  a47817a );
 a47822a <=( a47821a  and  a47814a );
 a47826a <=( (not A167)  and  (not A168) );
 a47827a <=( A169  and  a47826a );
 a47830a <=( (not A199)  and  A166 );
 a47833a <=( (not A233)  and  A200 );
 a47834a <=( a47833a  and  a47830a );
 a47835a <=( a47834a  and  a47827a );
 a47839a <=( (not A266)  and  (not A265) );
 a47840a <=( (not A234)  and  a47839a );
 a47843a <=( (not A299)  and  A298 );
 a47846a <=( A301  and  A300 );
 a47847a <=( a47846a  and  a47843a );
 a47848a <=( a47847a  and  a47840a );
 a47852a <=( (not A167)  and  (not A168) );
 a47853a <=( A169  and  a47852a );
 a47856a <=( (not A199)  and  A166 );
 a47859a <=( (not A233)  and  A200 );
 a47860a <=( a47859a  and  a47856a );
 a47861a <=( a47860a  and  a47853a );
 a47865a <=( (not A266)  and  (not A265) );
 a47866a <=( (not A234)  and  a47865a );
 a47869a <=( (not A299)  and  A298 );
 a47872a <=( A302  and  A300 );
 a47873a <=( a47872a  and  a47869a );
 a47874a <=( a47873a  and  a47866a );
 a47878a <=( (not A167)  and  (not A168) );
 a47879a <=( A169  and  a47878a );
 a47882a <=( (not A199)  and  A166 );
 a47885a <=( A232  and  A200 );
 a47886a <=( a47885a  and  a47882a );
 a47887a <=( a47886a  and  a47879a );
 a47891a <=( A235  and  A234 );
 a47892a <=( (not A233)  and  a47891a );
 a47895a <=( (not A266)  and  A265 );
 a47898a <=( A268  and  A267 );
 a47899a <=( a47898a  and  a47895a );
 a47900a <=( a47899a  and  a47892a );
 a47904a <=( (not A167)  and  (not A168) );
 a47905a <=( A169  and  a47904a );
 a47908a <=( (not A199)  and  A166 );
 a47911a <=( A232  and  A200 );
 a47912a <=( a47911a  and  a47908a );
 a47913a <=( a47912a  and  a47905a );
 a47917a <=( A235  and  A234 );
 a47918a <=( (not A233)  and  a47917a );
 a47921a <=( (not A266)  and  A265 );
 a47924a <=( A269  and  A267 );
 a47925a <=( a47924a  and  a47921a );
 a47926a <=( a47925a  and  a47918a );
 a47930a <=( (not A167)  and  (not A168) );
 a47931a <=( A169  and  a47930a );
 a47934a <=( (not A199)  and  A166 );
 a47937a <=( A232  and  A200 );
 a47938a <=( a47937a  and  a47934a );
 a47939a <=( a47938a  and  a47931a );
 a47943a <=( A236  and  A234 );
 a47944a <=( (not A233)  and  a47943a );
 a47947a <=( (not A266)  and  A265 );
 a47950a <=( A268  and  A267 );
 a47951a <=( a47950a  and  a47947a );
 a47952a <=( a47951a  and  a47944a );
 a47956a <=( (not A167)  and  (not A168) );
 a47957a <=( A169  and  a47956a );
 a47960a <=( (not A199)  and  A166 );
 a47963a <=( A232  and  A200 );
 a47964a <=( a47963a  and  a47960a );
 a47965a <=( a47964a  and  a47957a );
 a47969a <=( A236  and  A234 );
 a47970a <=( (not A233)  and  a47969a );
 a47973a <=( (not A266)  and  A265 );
 a47976a <=( A269  and  A267 );
 a47977a <=( a47976a  and  a47973a );
 a47978a <=( a47977a  and  a47970a );
 a47982a <=( (not A167)  and  (not A168) );
 a47983a <=( A169  and  a47982a );
 a47986a <=( (not A199)  and  A166 );
 a47989a <=( (not A232)  and  A200 );
 a47990a <=( a47989a  and  a47986a );
 a47991a <=( a47990a  and  a47983a );
 a47995a <=( A266  and  A265 );
 a47996a <=( (not A233)  and  a47995a );
 a47999a <=( (not A299)  and  A298 );
 a48002a <=( A301  and  A300 );
 a48003a <=( a48002a  and  a47999a );
 a48004a <=( a48003a  and  a47996a );
 a48008a <=( (not A167)  and  (not A168) );
 a48009a <=( A169  and  a48008a );
 a48012a <=( (not A199)  and  A166 );
 a48015a <=( (not A232)  and  A200 );
 a48016a <=( a48015a  and  a48012a );
 a48017a <=( a48016a  and  a48009a );
 a48021a <=( A266  and  A265 );
 a48022a <=( (not A233)  and  a48021a );
 a48025a <=( (not A299)  and  A298 );
 a48028a <=( A302  and  A300 );
 a48029a <=( a48028a  and  a48025a );
 a48030a <=( a48029a  and  a48022a );
 a48034a <=( (not A167)  and  (not A168) );
 a48035a <=( A169  and  a48034a );
 a48038a <=( (not A199)  and  A166 );
 a48041a <=( (not A232)  and  A200 );
 a48042a <=( a48041a  and  a48038a );
 a48043a <=( a48042a  and  a48035a );
 a48047a <=( (not A267)  and  (not A266) );
 a48048a <=( (not A233)  and  a48047a );
 a48051a <=( (not A299)  and  A298 );
 a48054a <=( A301  and  A300 );
 a48055a <=( a48054a  and  a48051a );
 a48056a <=( a48055a  and  a48048a );
 a48060a <=( (not A167)  and  (not A168) );
 a48061a <=( A169  and  a48060a );
 a48064a <=( (not A199)  and  A166 );
 a48067a <=( (not A232)  and  A200 );
 a48068a <=( a48067a  and  a48064a );
 a48069a <=( a48068a  and  a48061a );
 a48073a <=( (not A267)  and  (not A266) );
 a48074a <=( (not A233)  and  a48073a );
 a48077a <=( (not A299)  and  A298 );
 a48080a <=( A302  and  A300 );
 a48081a <=( a48080a  and  a48077a );
 a48082a <=( a48081a  and  a48074a );
 a48086a <=( (not A167)  and  (not A168) );
 a48087a <=( A169  and  a48086a );
 a48090a <=( (not A199)  and  A166 );
 a48093a <=( (not A232)  and  A200 );
 a48094a <=( a48093a  and  a48090a );
 a48095a <=( a48094a  and  a48087a );
 a48099a <=( (not A266)  and  (not A265) );
 a48100a <=( (not A233)  and  a48099a );
 a48103a <=( (not A299)  and  A298 );
 a48106a <=( A301  and  A300 );
 a48107a <=( a48106a  and  a48103a );
 a48108a <=( a48107a  and  a48100a );
 a48112a <=( (not A167)  and  (not A168) );
 a48113a <=( A169  and  a48112a );
 a48116a <=( (not A199)  and  A166 );
 a48119a <=( (not A232)  and  A200 );
 a48120a <=( a48119a  and  a48116a );
 a48121a <=( a48120a  and  a48113a );
 a48125a <=( (not A266)  and  (not A265) );
 a48126a <=( (not A233)  and  a48125a );
 a48129a <=( (not A299)  and  A298 );
 a48132a <=( A302  and  A300 );
 a48133a <=( a48132a  and  a48129a );
 a48134a <=( a48133a  and  a48126a );
 a48138a <=( (not A167)  and  (not A168) );
 a48139a <=( A169  and  a48138a );
 a48142a <=( A199  and  A166 );
 a48145a <=( A201  and  (not A200) );
 a48146a <=( a48145a  and  a48142a );
 a48147a <=( a48146a  and  a48139a );
 a48151a <=( A233  and  A232 );
 a48152a <=( A202  and  a48151a );
 a48155a <=( (not A267)  and  A265 );
 a48158a <=( A299  and  (not A298) );
 a48159a <=( a48158a  and  a48155a );
 a48160a <=( a48159a  and  a48152a );
 a48164a <=( (not A167)  and  (not A168) );
 a48165a <=( A169  and  a48164a );
 a48168a <=( A199  and  A166 );
 a48171a <=( A201  and  (not A200) );
 a48172a <=( a48171a  and  a48168a );
 a48173a <=( a48172a  and  a48165a );
 a48177a <=( A233  and  A232 );
 a48178a <=( A202  and  a48177a );
 a48181a <=( A266  and  A265 );
 a48184a <=( A299  and  (not A298) );
 a48185a <=( a48184a  and  a48181a );
 a48186a <=( a48185a  and  a48178a );
 a48190a <=( (not A167)  and  (not A168) );
 a48191a <=( A169  and  a48190a );
 a48194a <=( A199  and  A166 );
 a48197a <=( A201  and  (not A200) );
 a48198a <=( a48197a  and  a48194a );
 a48199a <=( a48198a  and  a48191a );
 a48203a <=( A233  and  A232 );
 a48204a <=( A202  and  a48203a );
 a48207a <=( (not A266)  and  (not A265) );
 a48210a <=( A299  and  (not A298) );
 a48211a <=( a48210a  and  a48207a );
 a48212a <=( a48211a  and  a48204a );
 a48216a <=( (not A167)  and  (not A168) );
 a48217a <=( A169  and  a48216a );
 a48220a <=( A199  and  A166 );
 a48223a <=( A201  and  (not A200) );
 a48224a <=( a48223a  and  a48220a );
 a48225a <=( a48224a  and  a48217a );
 a48229a <=( A233  and  (not A232) );
 a48230a <=( A202  and  a48229a );
 a48233a <=( (not A266)  and  A265 );
 a48236a <=( A268  and  A267 );
 a48237a <=( a48236a  and  a48233a );
 a48238a <=( a48237a  and  a48230a );
 a48242a <=( (not A167)  and  (not A168) );
 a48243a <=( A169  and  a48242a );
 a48246a <=( A199  and  A166 );
 a48249a <=( A201  and  (not A200) );
 a48250a <=( a48249a  and  a48246a );
 a48251a <=( a48250a  and  a48243a );
 a48255a <=( A233  and  (not A232) );
 a48256a <=( A202  and  a48255a );
 a48259a <=( (not A266)  and  A265 );
 a48262a <=( A269  and  A267 );
 a48263a <=( a48262a  and  a48259a );
 a48264a <=( a48263a  and  a48256a );
 a48268a <=( (not A167)  and  (not A168) );
 a48269a <=( A169  and  a48268a );
 a48272a <=( A199  and  A166 );
 a48275a <=( A201  and  (not A200) );
 a48276a <=( a48275a  and  a48272a );
 a48277a <=( a48276a  and  a48269a );
 a48281a <=( (not A234)  and  (not A233) );
 a48282a <=( A202  and  a48281a );
 a48285a <=( A266  and  A265 );
 a48288a <=( A299  and  (not A298) );
 a48289a <=( a48288a  and  a48285a );
 a48290a <=( a48289a  and  a48282a );
 a48294a <=( (not A167)  and  (not A168) );
 a48295a <=( A169  and  a48294a );
 a48298a <=( A199  and  A166 );
 a48301a <=( A201  and  (not A200) );
 a48302a <=( a48301a  and  a48298a );
 a48303a <=( a48302a  and  a48295a );
 a48307a <=( (not A234)  and  (not A233) );
 a48308a <=( A202  and  a48307a );
 a48311a <=( (not A267)  and  (not A266) );
 a48314a <=( A299  and  (not A298) );
 a48315a <=( a48314a  and  a48311a );
 a48316a <=( a48315a  and  a48308a );
 a48320a <=( (not A167)  and  (not A168) );
 a48321a <=( A169  and  a48320a );
 a48324a <=( A199  and  A166 );
 a48327a <=( A201  and  (not A200) );
 a48328a <=( a48327a  and  a48324a );
 a48329a <=( a48328a  and  a48321a );
 a48333a <=( (not A234)  and  (not A233) );
 a48334a <=( A202  and  a48333a );
 a48337a <=( (not A266)  and  (not A265) );
 a48340a <=( A299  and  (not A298) );
 a48341a <=( a48340a  and  a48337a );
 a48342a <=( a48341a  and  a48334a );
 a48346a <=( (not A167)  and  (not A168) );
 a48347a <=( A169  and  a48346a );
 a48350a <=( A199  and  A166 );
 a48353a <=( A201  and  (not A200) );
 a48354a <=( a48353a  and  a48350a );
 a48355a <=( a48354a  and  a48347a );
 a48359a <=( (not A233)  and  A232 );
 a48360a <=( A202  and  a48359a );
 a48363a <=( A235  and  A234 );
 a48366a <=( (not A300)  and  A298 );
 a48367a <=( a48366a  and  a48363a );
 a48368a <=( a48367a  and  a48360a );
 a48372a <=( (not A167)  and  (not A168) );
 a48373a <=( A169  and  a48372a );
 a48376a <=( A199  and  A166 );
 a48379a <=( A201  and  (not A200) );
 a48380a <=( a48379a  and  a48376a );
 a48381a <=( a48380a  and  a48373a );
 a48385a <=( (not A233)  and  A232 );
 a48386a <=( A202  and  a48385a );
 a48389a <=( A235  and  A234 );
 a48392a <=( A299  and  A298 );
 a48393a <=( a48392a  and  a48389a );
 a48394a <=( a48393a  and  a48386a );
 a48398a <=( (not A167)  and  (not A168) );
 a48399a <=( A169  and  a48398a );
 a48402a <=( A199  and  A166 );
 a48405a <=( A201  and  (not A200) );
 a48406a <=( a48405a  and  a48402a );
 a48407a <=( a48406a  and  a48399a );
 a48411a <=( (not A233)  and  A232 );
 a48412a <=( A202  and  a48411a );
 a48415a <=( A235  and  A234 );
 a48418a <=( (not A299)  and  (not A298) );
 a48419a <=( a48418a  and  a48415a );
 a48420a <=( a48419a  and  a48412a );
 a48424a <=( (not A167)  and  (not A168) );
 a48425a <=( A169  and  a48424a );
 a48428a <=( A199  and  A166 );
 a48431a <=( A201  and  (not A200) );
 a48432a <=( a48431a  and  a48428a );
 a48433a <=( a48432a  and  a48425a );
 a48437a <=( (not A233)  and  A232 );
 a48438a <=( A202  and  a48437a );
 a48441a <=( A235  and  A234 );
 a48444a <=( A266  and  (not A265) );
 a48445a <=( a48444a  and  a48441a );
 a48446a <=( a48445a  and  a48438a );
 a48450a <=( (not A167)  and  (not A168) );
 a48451a <=( A169  and  a48450a );
 a48454a <=( A199  and  A166 );
 a48457a <=( A201  and  (not A200) );
 a48458a <=( a48457a  and  a48454a );
 a48459a <=( a48458a  and  a48451a );
 a48463a <=( (not A233)  and  A232 );
 a48464a <=( A202  and  a48463a );
 a48467a <=( A236  and  A234 );
 a48470a <=( (not A300)  and  A298 );
 a48471a <=( a48470a  and  a48467a );
 a48472a <=( a48471a  and  a48464a );
 a48476a <=( (not A167)  and  (not A168) );
 a48477a <=( A169  and  a48476a );
 a48480a <=( A199  and  A166 );
 a48483a <=( A201  and  (not A200) );
 a48484a <=( a48483a  and  a48480a );
 a48485a <=( a48484a  and  a48477a );
 a48489a <=( (not A233)  and  A232 );
 a48490a <=( A202  and  a48489a );
 a48493a <=( A236  and  A234 );
 a48496a <=( A299  and  A298 );
 a48497a <=( a48496a  and  a48493a );
 a48498a <=( a48497a  and  a48490a );
 a48502a <=( (not A167)  and  (not A168) );
 a48503a <=( A169  and  a48502a );
 a48506a <=( A199  and  A166 );
 a48509a <=( A201  and  (not A200) );
 a48510a <=( a48509a  and  a48506a );
 a48511a <=( a48510a  and  a48503a );
 a48515a <=( (not A233)  and  A232 );
 a48516a <=( A202  and  a48515a );
 a48519a <=( A236  and  A234 );
 a48522a <=( (not A299)  and  (not A298) );
 a48523a <=( a48522a  and  a48519a );
 a48524a <=( a48523a  and  a48516a );
 a48528a <=( (not A167)  and  (not A168) );
 a48529a <=( A169  and  a48528a );
 a48532a <=( A199  and  A166 );
 a48535a <=( A201  and  (not A200) );
 a48536a <=( a48535a  and  a48532a );
 a48537a <=( a48536a  and  a48529a );
 a48541a <=( (not A233)  and  A232 );
 a48542a <=( A202  and  a48541a );
 a48545a <=( A236  and  A234 );
 a48548a <=( A266  and  (not A265) );
 a48549a <=( a48548a  and  a48545a );
 a48550a <=( a48549a  and  a48542a );
 a48554a <=( (not A167)  and  (not A168) );
 a48555a <=( A169  and  a48554a );
 a48558a <=( A199  and  A166 );
 a48561a <=( A201  and  (not A200) );
 a48562a <=( a48561a  and  a48558a );
 a48563a <=( a48562a  and  a48555a );
 a48567a <=( (not A233)  and  (not A232) );
 a48568a <=( A202  and  a48567a );
 a48571a <=( A266  and  A265 );
 a48574a <=( A299  and  (not A298) );
 a48575a <=( a48574a  and  a48571a );
 a48576a <=( a48575a  and  a48568a );
 a48580a <=( (not A167)  and  (not A168) );
 a48581a <=( A169  and  a48580a );
 a48584a <=( A199  and  A166 );
 a48587a <=( A201  and  (not A200) );
 a48588a <=( a48587a  and  a48584a );
 a48589a <=( a48588a  and  a48581a );
 a48593a <=( (not A233)  and  (not A232) );
 a48594a <=( A202  and  a48593a );
 a48597a <=( (not A267)  and  (not A266) );
 a48600a <=( A299  and  (not A298) );
 a48601a <=( a48600a  and  a48597a );
 a48602a <=( a48601a  and  a48594a );
 a48606a <=( (not A167)  and  (not A168) );
 a48607a <=( A169  and  a48606a );
 a48610a <=( A199  and  A166 );
 a48613a <=( A201  and  (not A200) );
 a48614a <=( a48613a  and  a48610a );
 a48615a <=( a48614a  and  a48607a );
 a48619a <=( (not A233)  and  (not A232) );
 a48620a <=( A202  and  a48619a );
 a48623a <=( (not A266)  and  (not A265) );
 a48626a <=( A299  and  (not A298) );
 a48627a <=( a48626a  and  a48623a );
 a48628a <=( a48627a  and  a48620a );
 a48632a <=( (not A167)  and  (not A168) );
 a48633a <=( A169  and  a48632a );
 a48636a <=( A199  and  A166 );
 a48639a <=( A201  and  (not A200) );
 a48640a <=( a48639a  and  a48636a );
 a48641a <=( a48640a  and  a48633a );
 a48645a <=( A233  and  A232 );
 a48646a <=( A203  and  a48645a );
 a48649a <=( (not A267)  and  A265 );
 a48652a <=( A299  and  (not A298) );
 a48653a <=( a48652a  and  a48649a );
 a48654a <=( a48653a  and  a48646a );
 a48658a <=( (not A167)  and  (not A168) );
 a48659a <=( A169  and  a48658a );
 a48662a <=( A199  and  A166 );
 a48665a <=( A201  and  (not A200) );
 a48666a <=( a48665a  and  a48662a );
 a48667a <=( a48666a  and  a48659a );
 a48671a <=( A233  and  A232 );
 a48672a <=( A203  and  a48671a );
 a48675a <=( A266  and  A265 );
 a48678a <=( A299  and  (not A298) );
 a48679a <=( a48678a  and  a48675a );
 a48680a <=( a48679a  and  a48672a );
 a48684a <=( (not A167)  and  (not A168) );
 a48685a <=( A169  and  a48684a );
 a48688a <=( A199  and  A166 );
 a48691a <=( A201  and  (not A200) );
 a48692a <=( a48691a  and  a48688a );
 a48693a <=( a48692a  and  a48685a );
 a48697a <=( A233  and  A232 );
 a48698a <=( A203  and  a48697a );
 a48701a <=( (not A266)  and  (not A265) );
 a48704a <=( A299  and  (not A298) );
 a48705a <=( a48704a  and  a48701a );
 a48706a <=( a48705a  and  a48698a );
 a48710a <=( (not A167)  and  (not A168) );
 a48711a <=( A169  and  a48710a );
 a48714a <=( A199  and  A166 );
 a48717a <=( A201  and  (not A200) );
 a48718a <=( a48717a  and  a48714a );
 a48719a <=( a48718a  and  a48711a );
 a48723a <=( A233  and  (not A232) );
 a48724a <=( A203  and  a48723a );
 a48727a <=( (not A266)  and  A265 );
 a48730a <=( A268  and  A267 );
 a48731a <=( a48730a  and  a48727a );
 a48732a <=( a48731a  and  a48724a );
 a48736a <=( (not A167)  and  (not A168) );
 a48737a <=( A169  and  a48736a );
 a48740a <=( A199  and  A166 );
 a48743a <=( A201  and  (not A200) );
 a48744a <=( a48743a  and  a48740a );
 a48745a <=( a48744a  and  a48737a );
 a48749a <=( A233  and  (not A232) );
 a48750a <=( A203  and  a48749a );
 a48753a <=( (not A266)  and  A265 );
 a48756a <=( A269  and  A267 );
 a48757a <=( a48756a  and  a48753a );
 a48758a <=( a48757a  and  a48750a );
 a48762a <=( (not A167)  and  (not A168) );
 a48763a <=( A169  and  a48762a );
 a48766a <=( A199  and  A166 );
 a48769a <=( A201  and  (not A200) );
 a48770a <=( a48769a  and  a48766a );
 a48771a <=( a48770a  and  a48763a );
 a48775a <=( (not A234)  and  (not A233) );
 a48776a <=( A203  and  a48775a );
 a48779a <=( A266  and  A265 );
 a48782a <=( A299  and  (not A298) );
 a48783a <=( a48782a  and  a48779a );
 a48784a <=( a48783a  and  a48776a );
 a48788a <=( (not A167)  and  (not A168) );
 a48789a <=( A169  and  a48788a );
 a48792a <=( A199  and  A166 );
 a48795a <=( A201  and  (not A200) );
 a48796a <=( a48795a  and  a48792a );
 a48797a <=( a48796a  and  a48789a );
 a48801a <=( (not A234)  and  (not A233) );
 a48802a <=( A203  and  a48801a );
 a48805a <=( (not A267)  and  (not A266) );
 a48808a <=( A299  and  (not A298) );
 a48809a <=( a48808a  and  a48805a );
 a48810a <=( a48809a  and  a48802a );
 a48814a <=( (not A167)  and  (not A168) );
 a48815a <=( A169  and  a48814a );
 a48818a <=( A199  and  A166 );
 a48821a <=( A201  and  (not A200) );
 a48822a <=( a48821a  and  a48818a );
 a48823a <=( a48822a  and  a48815a );
 a48827a <=( (not A234)  and  (not A233) );
 a48828a <=( A203  and  a48827a );
 a48831a <=( (not A266)  and  (not A265) );
 a48834a <=( A299  and  (not A298) );
 a48835a <=( a48834a  and  a48831a );
 a48836a <=( a48835a  and  a48828a );
 a48840a <=( (not A167)  and  (not A168) );
 a48841a <=( A169  and  a48840a );
 a48844a <=( A199  and  A166 );
 a48847a <=( A201  and  (not A200) );
 a48848a <=( a48847a  and  a48844a );
 a48849a <=( a48848a  and  a48841a );
 a48853a <=( (not A233)  and  A232 );
 a48854a <=( A203  and  a48853a );
 a48857a <=( A235  and  A234 );
 a48860a <=( (not A300)  and  A298 );
 a48861a <=( a48860a  and  a48857a );
 a48862a <=( a48861a  and  a48854a );
 a48866a <=( (not A167)  and  (not A168) );
 a48867a <=( A169  and  a48866a );
 a48870a <=( A199  and  A166 );
 a48873a <=( A201  and  (not A200) );
 a48874a <=( a48873a  and  a48870a );
 a48875a <=( a48874a  and  a48867a );
 a48879a <=( (not A233)  and  A232 );
 a48880a <=( A203  and  a48879a );
 a48883a <=( A235  and  A234 );
 a48886a <=( A299  and  A298 );
 a48887a <=( a48886a  and  a48883a );
 a48888a <=( a48887a  and  a48880a );
 a48892a <=( (not A167)  and  (not A168) );
 a48893a <=( A169  and  a48892a );
 a48896a <=( A199  and  A166 );
 a48899a <=( A201  and  (not A200) );
 a48900a <=( a48899a  and  a48896a );
 a48901a <=( a48900a  and  a48893a );
 a48905a <=( (not A233)  and  A232 );
 a48906a <=( A203  and  a48905a );
 a48909a <=( A235  and  A234 );
 a48912a <=( (not A299)  and  (not A298) );
 a48913a <=( a48912a  and  a48909a );
 a48914a <=( a48913a  and  a48906a );
 a48918a <=( (not A167)  and  (not A168) );
 a48919a <=( A169  and  a48918a );
 a48922a <=( A199  and  A166 );
 a48925a <=( A201  and  (not A200) );
 a48926a <=( a48925a  and  a48922a );
 a48927a <=( a48926a  and  a48919a );
 a48931a <=( (not A233)  and  A232 );
 a48932a <=( A203  and  a48931a );
 a48935a <=( A235  and  A234 );
 a48938a <=( A266  and  (not A265) );
 a48939a <=( a48938a  and  a48935a );
 a48940a <=( a48939a  and  a48932a );
 a48944a <=( (not A167)  and  (not A168) );
 a48945a <=( A169  and  a48944a );
 a48948a <=( A199  and  A166 );
 a48951a <=( A201  and  (not A200) );
 a48952a <=( a48951a  and  a48948a );
 a48953a <=( a48952a  and  a48945a );
 a48957a <=( (not A233)  and  A232 );
 a48958a <=( A203  and  a48957a );
 a48961a <=( A236  and  A234 );
 a48964a <=( (not A300)  and  A298 );
 a48965a <=( a48964a  and  a48961a );
 a48966a <=( a48965a  and  a48958a );
 a48970a <=( (not A167)  and  (not A168) );
 a48971a <=( A169  and  a48970a );
 a48974a <=( A199  and  A166 );
 a48977a <=( A201  and  (not A200) );
 a48978a <=( a48977a  and  a48974a );
 a48979a <=( a48978a  and  a48971a );
 a48983a <=( (not A233)  and  A232 );
 a48984a <=( A203  and  a48983a );
 a48987a <=( A236  and  A234 );
 a48990a <=( A299  and  A298 );
 a48991a <=( a48990a  and  a48987a );
 a48992a <=( a48991a  and  a48984a );
 a48996a <=( (not A167)  and  (not A168) );
 a48997a <=( A169  and  a48996a );
 a49000a <=( A199  and  A166 );
 a49003a <=( A201  and  (not A200) );
 a49004a <=( a49003a  and  a49000a );
 a49005a <=( a49004a  and  a48997a );
 a49009a <=( (not A233)  and  A232 );
 a49010a <=( A203  and  a49009a );
 a49013a <=( A236  and  A234 );
 a49016a <=( (not A299)  and  (not A298) );
 a49017a <=( a49016a  and  a49013a );
 a49018a <=( a49017a  and  a49010a );
 a49022a <=( (not A167)  and  (not A168) );
 a49023a <=( A169  and  a49022a );
 a49026a <=( A199  and  A166 );
 a49029a <=( A201  and  (not A200) );
 a49030a <=( a49029a  and  a49026a );
 a49031a <=( a49030a  and  a49023a );
 a49035a <=( (not A233)  and  A232 );
 a49036a <=( A203  and  a49035a );
 a49039a <=( A236  and  A234 );
 a49042a <=( A266  and  (not A265) );
 a49043a <=( a49042a  and  a49039a );
 a49044a <=( a49043a  and  a49036a );
 a49048a <=( (not A167)  and  (not A168) );
 a49049a <=( A169  and  a49048a );
 a49052a <=( A199  and  A166 );
 a49055a <=( A201  and  (not A200) );
 a49056a <=( a49055a  and  a49052a );
 a49057a <=( a49056a  and  a49049a );
 a49061a <=( (not A233)  and  (not A232) );
 a49062a <=( A203  and  a49061a );
 a49065a <=( A266  and  A265 );
 a49068a <=( A299  and  (not A298) );
 a49069a <=( a49068a  and  a49065a );
 a49070a <=( a49069a  and  a49062a );
 a49074a <=( (not A167)  and  (not A168) );
 a49075a <=( A169  and  a49074a );
 a49078a <=( A199  and  A166 );
 a49081a <=( A201  and  (not A200) );
 a49082a <=( a49081a  and  a49078a );
 a49083a <=( a49082a  and  a49075a );
 a49087a <=( (not A233)  and  (not A232) );
 a49088a <=( A203  and  a49087a );
 a49091a <=( (not A267)  and  (not A266) );
 a49094a <=( A299  and  (not A298) );
 a49095a <=( a49094a  and  a49091a );
 a49096a <=( a49095a  and  a49088a );
 a49100a <=( (not A167)  and  (not A168) );
 a49101a <=( A169  and  a49100a );
 a49104a <=( A199  and  A166 );
 a49107a <=( A201  and  (not A200) );
 a49108a <=( a49107a  and  a49104a );
 a49109a <=( a49108a  and  a49101a );
 a49113a <=( (not A233)  and  (not A232) );
 a49114a <=( A203  and  a49113a );
 a49117a <=( (not A266)  and  (not A265) );
 a49120a <=( A299  and  (not A298) );
 a49121a <=( a49120a  and  a49117a );
 a49122a <=( a49121a  and  a49114a );
 a49126a <=( (not A168)  and  A169 );
 a49127a <=( A170  and  a49126a );
 a49130a <=( (not A200)  and  A199 );
 a49133a <=( A202  and  A201 );
 a49134a <=( a49133a  and  a49130a );
 a49135a <=( a49134a  and  a49127a );
 a49139a <=( A265  and  A233 );
 a49140a <=( A232  and  a49139a );
 a49143a <=( (not A269)  and  (not A268) );
 a49146a <=( A299  and  (not A298) );
 a49147a <=( a49146a  and  a49143a );
 a49148a <=( a49147a  and  a49140a );
 a49152a <=( (not A168)  and  A169 );
 a49153a <=( A170  and  a49152a );
 a49156a <=( (not A200)  and  A199 );
 a49159a <=( A202  and  A201 );
 a49160a <=( a49159a  and  a49156a );
 a49161a <=( a49160a  and  a49153a );
 a49165a <=( (not A236)  and  (not A235) );
 a49166a <=( (not A233)  and  a49165a );
 a49169a <=( A266  and  A265 );
 a49172a <=( A299  and  (not A298) );
 a49173a <=( a49172a  and  a49169a );
 a49174a <=( a49173a  and  a49166a );
 a49178a <=( (not A168)  and  A169 );
 a49179a <=( A170  and  a49178a );
 a49182a <=( (not A200)  and  A199 );
 a49185a <=( A202  and  A201 );
 a49186a <=( a49185a  and  a49182a );
 a49187a <=( a49186a  and  a49179a );
 a49191a <=( (not A236)  and  (not A235) );
 a49192a <=( (not A233)  and  a49191a );
 a49195a <=( (not A267)  and  (not A266) );
 a49198a <=( A299  and  (not A298) );
 a49199a <=( a49198a  and  a49195a );
 a49200a <=( a49199a  and  a49192a );
 a49204a <=( (not A168)  and  A169 );
 a49205a <=( A170  and  a49204a );
 a49208a <=( (not A200)  and  A199 );
 a49211a <=( A202  and  A201 );
 a49212a <=( a49211a  and  a49208a );
 a49213a <=( a49212a  and  a49205a );
 a49217a <=( (not A236)  and  (not A235) );
 a49218a <=( (not A233)  and  a49217a );
 a49221a <=( (not A266)  and  (not A265) );
 a49224a <=( A299  and  (not A298) );
 a49225a <=( a49224a  and  a49221a );
 a49226a <=( a49225a  and  a49218a );
 a49230a <=( (not A168)  and  A169 );
 a49231a <=( A170  and  a49230a );
 a49234a <=( (not A200)  and  A199 );
 a49237a <=( A202  and  A201 );
 a49238a <=( a49237a  and  a49234a );
 a49239a <=( a49238a  and  a49231a );
 a49243a <=( (not A266)  and  (not A234) );
 a49244a <=( (not A233)  and  a49243a );
 a49247a <=( (not A269)  and  (not A268) );
 a49250a <=( A299  and  (not A298) );
 a49251a <=( a49250a  and  a49247a );
 a49252a <=( a49251a  and  a49244a );
 a49256a <=( (not A168)  and  A169 );
 a49257a <=( A170  and  a49256a );
 a49260a <=( (not A200)  and  A199 );
 a49263a <=( A202  and  A201 );
 a49264a <=( a49263a  and  a49260a );
 a49265a <=( a49264a  and  a49257a );
 a49269a <=( A234  and  (not A233) );
 a49270a <=( A232  and  a49269a );
 a49273a <=( A298  and  A235 );
 a49276a <=( (not A302)  and  (not A301) );
 a49277a <=( a49276a  and  a49273a );
 a49278a <=( a49277a  and  a49270a );
 a49282a <=( (not A168)  and  A169 );
 a49283a <=( A170  and  a49282a );
 a49286a <=( (not A200)  and  A199 );
 a49289a <=( A202  and  A201 );
 a49290a <=( a49289a  and  a49286a );
 a49291a <=( a49290a  and  a49283a );
 a49295a <=( A234  and  (not A233) );
 a49296a <=( A232  and  a49295a );
 a49299a <=( A298  and  A236 );
 a49302a <=( (not A302)  and  (not A301) );
 a49303a <=( a49302a  and  a49299a );
 a49304a <=( a49303a  and  a49296a );
 a49308a <=( (not A168)  and  A169 );
 a49309a <=( A170  and  a49308a );
 a49312a <=( (not A200)  and  A199 );
 a49315a <=( A202  and  A201 );
 a49316a <=( a49315a  and  a49312a );
 a49317a <=( a49316a  and  a49309a );
 a49321a <=( (not A266)  and  (not A233) );
 a49322a <=( (not A232)  and  a49321a );
 a49325a <=( (not A269)  and  (not A268) );
 a49328a <=( A299  and  (not A298) );
 a49329a <=( a49328a  and  a49325a );
 a49330a <=( a49329a  and  a49322a );
 a49334a <=( (not A168)  and  A169 );
 a49335a <=( A170  and  a49334a );
 a49338a <=( (not A200)  and  A199 );
 a49341a <=( A203  and  A201 );
 a49342a <=( a49341a  and  a49338a );
 a49343a <=( a49342a  and  a49335a );
 a49347a <=( A265  and  A233 );
 a49348a <=( A232  and  a49347a );
 a49351a <=( (not A269)  and  (not A268) );
 a49354a <=( A299  and  (not A298) );
 a49355a <=( a49354a  and  a49351a );
 a49356a <=( a49355a  and  a49348a );
 a49360a <=( (not A168)  and  A169 );
 a49361a <=( A170  and  a49360a );
 a49364a <=( (not A200)  and  A199 );
 a49367a <=( A203  and  A201 );
 a49368a <=( a49367a  and  a49364a );
 a49369a <=( a49368a  and  a49361a );
 a49373a <=( (not A236)  and  (not A235) );
 a49374a <=( (not A233)  and  a49373a );
 a49377a <=( A266  and  A265 );
 a49380a <=( A299  and  (not A298) );
 a49381a <=( a49380a  and  a49377a );
 a49382a <=( a49381a  and  a49374a );
 a49386a <=( (not A168)  and  A169 );
 a49387a <=( A170  and  a49386a );
 a49390a <=( (not A200)  and  A199 );
 a49393a <=( A203  and  A201 );
 a49394a <=( a49393a  and  a49390a );
 a49395a <=( a49394a  and  a49387a );
 a49399a <=( (not A236)  and  (not A235) );
 a49400a <=( (not A233)  and  a49399a );
 a49403a <=( (not A267)  and  (not A266) );
 a49406a <=( A299  and  (not A298) );
 a49407a <=( a49406a  and  a49403a );
 a49408a <=( a49407a  and  a49400a );
 a49412a <=( (not A168)  and  A169 );
 a49413a <=( A170  and  a49412a );
 a49416a <=( (not A200)  and  A199 );
 a49419a <=( A203  and  A201 );
 a49420a <=( a49419a  and  a49416a );
 a49421a <=( a49420a  and  a49413a );
 a49425a <=( (not A236)  and  (not A235) );
 a49426a <=( (not A233)  and  a49425a );
 a49429a <=( (not A266)  and  (not A265) );
 a49432a <=( A299  and  (not A298) );
 a49433a <=( a49432a  and  a49429a );
 a49434a <=( a49433a  and  a49426a );
 a49438a <=( (not A168)  and  A169 );
 a49439a <=( A170  and  a49438a );
 a49442a <=( (not A200)  and  A199 );
 a49445a <=( A203  and  A201 );
 a49446a <=( a49445a  and  a49442a );
 a49447a <=( a49446a  and  a49439a );
 a49451a <=( (not A266)  and  (not A234) );
 a49452a <=( (not A233)  and  a49451a );
 a49455a <=( (not A269)  and  (not A268) );
 a49458a <=( A299  and  (not A298) );
 a49459a <=( a49458a  and  a49455a );
 a49460a <=( a49459a  and  a49452a );
 a49464a <=( (not A168)  and  A169 );
 a49465a <=( A170  and  a49464a );
 a49468a <=( (not A200)  and  A199 );
 a49471a <=( A203  and  A201 );
 a49472a <=( a49471a  and  a49468a );
 a49473a <=( a49472a  and  a49465a );
 a49477a <=( A234  and  (not A233) );
 a49478a <=( A232  and  a49477a );
 a49481a <=( A298  and  A235 );
 a49484a <=( (not A302)  and  (not A301) );
 a49485a <=( a49484a  and  a49481a );
 a49486a <=( a49485a  and  a49478a );
 a49490a <=( (not A168)  and  A169 );
 a49491a <=( A170  and  a49490a );
 a49494a <=( (not A200)  and  A199 );
 a49497a <=( A203  and  A201 );
 a49498a <=( a49497a  and  a49494a );
 a49499a <=( a49498a  and  a49491a );
 a49503a <=( A234  and  (not A233) );
 a49504a <=( A232  and  a49503a );
 a49507a <=( A298  and  A236 );
 a49510a <=( (not A302)  and  (not A301) );
 a49511a <=( a49510a  and  a49507a );
 a49512a <=( a49511a  and  a49504a );
 a49516a <=( (not A168)  and  A169 );
 a49517a <=( A170  and  a49516a );
 a49520a <=( (not A200)  and  A199 );
 a49523a <=( A203  and  A201 );
 a49524a <=( a49523a  and  a49520a );
 a49525a <=( a49524a  and  a49517a );
 a49529a <=( (not A266)  and  (not A233) );
 a49530a <=( (not A232)  and  a49529a );
 a49533a <=( (not A269)  and  (not A268) );
 a49536a <=( A299  and  (not A298) );
 a49537a <=( a49536a  and  a49533a );
 a49538a <=( a49537a  and  a49530a );
 a49542a <=( A167  and  A169 );
 a49543a <=( (not A170)  and  a49542a );
 a49546a <=( A199  and  A166 );
 a49549a <=( A232  and  A200 );
 a49550a <=( a49549a  and  a49546a );
 a49551a <=( a49550a  and  a49543a );
 a49555a <=( (not A267)  and  A265 );
 a49556a <=( A233  and  a49555a );
 a49559a <=( (not A299)  and  A298 );
 a49562a <=( A301  and  A300 );
 a49563a <=( a49562a  and  a49559a );
 a49564a <=( a49563a  and  a49556a );
 a49568a <=( A167  and  A169 );
 a49569a <=( (not A170)  and  a49568a );
 a49572a <=( A199  and  A166 );
 a49575a <=( A232  and  A200 );
 a49576a <=( a49575a  and  a49572a );
 a49577a <=( a49576a  and  a49569a );
 a49581a <=( (not A267)  and  A265 );
 a49582a <=( A233  and  a49581a );
 a49585a <=( (not A299)  and  A298 );
 a49588a <=( A302  and  A300 );
 a49589a <=( a49588a  and  a49585a );
 a49590a <=( a49589a  and  a49582a );
 a49594a <=( A167  and  A169 );
 a49595a <=( (not A170)  and  a49594a );
 a49598a <=( A199  and  A166 );
 a49601a <=( A232  and  A200 );
 a49602a <=( a49601a  and  a49598a );
 a49603a <=( a49602a  and  a49595a );
 a49607a <=( A266  and  A265 );
 a49608a <=( A233  and  a49607a );
 a49611a <=( (not A299)  and  A298 );
 a49614a <=( A301  and  A300 );
 a49615a <=( a49614a  and  a49611a );
 a49616a <=( a49615a  and  a49608a );
 a49620a <=( A167  and  A169 );
 a49621a <=( (not A170)  and  a49620a );
 a49624a <=( A199  and  A166 );
 a49627a <=( A232  and  A200 );
 a49628a <=( a49627a  and  a49624a );
 a49629a <=( a49628a  and  a49621a );
 a49633a <=( A266  and  A265 );
 a49634a <=( A233  and  a49633a );
 a49637a <=( (not A299)  and  A298 );
 a49640a <=( A302  and  A300 );
 a49641a <=( a49640a  and  a49637a );
 a49642a <=( a49641a  and  a49634a );
 a49646a <=( A167  and  A169 );
 a49647a <=( (not A170)  and  a49646a );
 a49650a <=( A199  and  A166 );
 a49653a <=( A232  and  A200 );
 a49654a <=( a49653a  and  a49650a );
 a49655a <=( a49654a  and  a49647a );
 a49659a <=( (not A266)  and  (not A265) );
 a49660a <=( A233  and  a49659a );
 a49663a <=( (not A299)  and  A298 );
 a49666a <=( A301  and  A300 );
 a49667a <=( a49666a  and  a49663a );
 a49668a <=( a49667a  and  a49660a );
 a49672a <=( A167  and  A169 );
 a49673a <=( (not A170)  and  a49672a );
 a49676a <=( A199  and  A166 );
 a49679a <=( A232  and  A200 );
 a49680a <=( a49679a  and  a49676a );
 a49681a <=( a49680a  and  a49673a );
 a49685a <=( (not A266)  and  (not A265) );
 a49686a <=( A233  and  a49685a );
 a49689a <=( (not A299)  and  A298 );
 a49692a <=( A302  and  A300 );
 a49693a <=( a49692a  and  a49689a );
 a49694a <=( a49693a  and  a49686a );
 a49698a <=( A167  and  A169 );
 a49699a <=( (not A170)  and  a49698a );
 a49702a <=( A199  and  A166 );
 a49705a <=( (not A233)  and  A200 );
 a49706a <=( a49705a  and  a49702a );
 a49707a <=( a49706a  and  a49699a );
 a49711a <=( (not A266)  and  (not A236) );
 a49712a <=( (not A235)  and  a49711a );
 a49715a <=( (not A269)  and  (not A268) );
 a49718a <=( A299  and  (not A298) );
 a49719a <=( a49718a  and  a49715a );
 a49720a <=( a49719a  and  a49712a );
 a49724a <=( A167  and  A169 );
 a49725a <=( (not A170)  and  a49724a );
 a49728a <=( A199  and  A166 );
 a49731a <=( (not A233)  and  A200 );
 a49732a <=( a49731a  and  a49728a );
 a49733a <=( a49732a  and  a49725a );
 a49737a <=( A266  and  A265 );
 a49738a <=( (not A234)  and  a49737a );
 a49741a <=( (not A299)  and  A298 );
 a49744a <=( A301  and  A300 );
 a49745a <=( a49744a  and  a49741a );
 a49746a <=( a49745a  and  a49738a );
 a49750a <=( A167  and  A169 );
 a49751a <=( (not A170)  and  a49750a );
 a49754a <=( A199  and  A166 );
 a49757a <=( (not A233)  and  A200 );
 a49758a <=( a49757a  and  a49754a );
 a49759a <=( a49758a  and  a49751a );
 a49763a <=( A266  and  A265 );
 a49764a <=( (not A234)  and  a49763a );
 a49767a <=( (not A299)  and  A298 );
 a49770a <=( A302  and  A300 );
 a49771a <=( a49770a  and  a49767a );
 a49772a <=( a49771a  and  a49764a );
 a49776a <=( A167  and  A169 );
 a49777a <=( (not A170)  and  a49776a );
 a49780a <=( A199  and  A166 );
 a49783a <=( (not A233)  and  A200 );
 a49784a <=( a49783a  and  a49780a );
 a49785a <=( a49784a  and  a49777a );
 a49789a <=( (not A267)  and  (not A266) );
 a49790a <=( (not A234)  and  a49789a );
 a49793a <=( (not A299)  and  A298 );
 a49796a <=( A301  and  A300 );
 a49797a <=( a49796a  and  a49793a );
 a49798a <=( a49797a  and  a49790a );
 a49802a <=( A167  and  A169 );
 a49803a <=( (not A170)  and  a49802a );
 a49806a <=( A199  and  A166 );
 a49809a <=( (not A233)  and  A200 );
 a49810a <=( a49809a  and  a49806a );
 a49811a <=( a49810a  and  a49803a );
 a49815a <=( (not A267)  and  (not A266) );
 a49816a <=( (not A234)  and  a49815a );
 a49819a <=( (not A299)  and  A298 );
 a49822a <=( A302  and  A300 );
 a49823a <=( a49822a  and  a49819a );
 a49824a <=( a49823a  and  a49816a );
 a49828a <=( A167  and  A169 );
 a49829a <=( (not A170)  and  a49828a );
 a49832a <=( A199  and  A166 );
 a49835a <=( (not A233)  and  A200 );
 a49836a <=( a49835a  and  a49832a );
 a49837a <=( a49836a  and  a49829a );
 a49841a <=( (not A266)  and  (not A265) );
 a49842a <=( (not A234)  and  a49841a );
 a49845a <=( (not A299)  and  A298 );
 a49848a <=( A301  and  A300 );
 a49849a <=( a49848a  and  a49845a );
 a49850a <=( a49849a  and  a49842a );
 a49854a <=( A167  and  A169 );
 a49855a <=( (not A170)  and  a49854a );
 a49858a <=( A199  and  A166 );
 a49861a <=( (not A233)  and  A200 );
 a49862a <=( a49861a  and  a49858a );
 a49863a <=( a49862a  and  a49855a );
 a49867a <=( (not A266)  and  (not A265) );
 a49868a <=( (not A234)  and  a49867a );
 a49871a <=( (not A299)  and  A298 );
 a49874a <=( A302  and  A300 );
 a49875a <=( a49874a  and  a49871a );
 a49876a <=( a49875a  and  a49868a );
 a49880a <=( A167  and  A169 );
 a49881a <=( (not A170)  and  a49880a );
 a49884a <=( A199  and  A166 );
 a49887a <=( A232  and  A200 );
 a49888a <=( a49887a  and  a49884a );
 a49889a <=( a49888a  and  a49881a );
 a49893a <=( A235  and  A234 );
 a49894a <=( (not A233)  and  a49893a );
 a49897a <=( (not A266)  and  A265 );
 a49900a <=( A268  and  A267 );
 a49901a <=( a49900a  and  a49897a );
 a49902a <=( a49901a  and  a49894a );
 a49906a <=( A167  and  A169 );
 a49907a <=( (not A170)  and  a49906a );
 a49910a <=( A199  and  A166 );
 a49913a <=( A232  and  A200 );
 a49914a <=( a49913a  and  a49910a );
 a49915a <=( a49914a  and  a49907a );
 a49919a <=( A235  and  A234 );
 a49920a <=( (not A233)  and  a49919a );
 a49923a <=( (not A266)  and  A265 );
 a49926a <=( A269  and  A267 );
 a49927a <=( a49926a  and  a49923a );
 a49928a <=( a49927a  and  a49920a );
 a49932a <=( A167  and  A169 );
 a49933a <=( (not A170)  and  a49932a );
 a49936a <=( A199  and  A166 );
 a49939a <=( A232  and  A200 );
 a49940a <=( a49939a  and  a49936a );
 a49941a <=( a49940a  and  a49933a );
 a49945a <=( A236  and  A234 );
 a49946a <=( (not A233)  and  a49945a );
 a49949a <=( (not A266)  and  A265 );
 a49952a <=( A268  and  A267 );
 a49953a <=( a49952a  and  a49949a );
 a49954a <=( a49953a  and  a49946a );
 a49958a <=( A167  and  A169 );
 a49959a <=( (not A170)  and  a49958a );
 a49962a <=( A199  and  A166 );
 a49965a <=( A232  and  A200 );
 a49966a <=( a49965a  and  a49962a );
 a49967a <=( a49966a  and  a49959a );
 a49971a <=( A236  and  A234 );
 a49972a <=( (not A233)  and  a49971a );
 a49975a <=( (not A266)  and  A265 );
 a49978a <=( A269  and  A267 );
 a49979a <=( a49978a  and  a49975a );
 a49980a <=( a49979a  and  a49972a );
 a49984a <=( A167  and  A169 );
 a49985a <=( (not A170)  and  a49984a );
 a49988a <=( A199  and  A166 );
 a49991a <=( (not A232)  and  A200 );
 a49992a <=( a49991a  and  a49988a );
 a49993a <=( a49992a  and  a49985a );
 a49997a <=( A266  and  A265 );
 a49998a <=( (not A233)  and  a49997a );
 a50001a <=( (not A299)  and  A298 );
 a50004a <=( A301  and  A300 );
 a50005a <=( a50004a  and  a50001a );
 a50006a <=( a50005a  and  a49998a );
 a50010a <=( A167  and  A169 );
 a50011a <=( (not A170)  and  a50010a );
 a50014a <=( A199  and  A166 );
 a50017a <=( (not A232)  and  A200 );
 a50018a <=( a50017a  and  a50014a );
 a50019a <=( a50018a  and  a50011a );
 a50023a <=( A266  and  A265 );
 a50024a <=( (not A233)  and  a50023a );
 a50027a <=( (not A299)  and  A298 );
 a50030a <=( A302  and  A300 );
 a50031a <=( a50030a  and  a50027a );
 a50032a <=( a50031a  and  a50024a );
 a50036a <=( A167  and  A169 );
 a50037a <=( (not A170)  and  a50036a );
 a50040a <=( A199  and  A166 );
 a50043a <=( (not A232)  and  A200 );
 a50044a <=( a50043a  and  a50040a );
 a50045a <=( a50044a  and  a50037a );
 a50049a <=( (not A267)  and  (not A266) );
 a50050a <=( (not A233)  and  a50049a );
 a50053a <=( (not A299)  and  A298 );
 a50056a <=( A301  and  A300 );
 a50057a <=( a50056a  and  a50053a );
 a50058a <=( a50057a  and  a50050a );
 a50062a <=( A167  and  A169 );
 a50063a <=( (not A170)  and  a50062a );
 a50066a <=( A199  and  A166 );
 a50069a <=( (not A232)  and  A200 );
 a50070a <=( a50069a  and  a50066a );
 a50071a <=( a50070a  and  a50063a );
 a50075a <=( (not A267)  and  (not A266) );
 a50076a <=( (not A233)  and  a50075a );
 a50079a <=( (not A299)  and  A298 );
 a50082a <=( A302  and  A300 );
 a50083a <=( a50082a  and  a50079a );
 a50084a <=( a50083a  and  a50076a );
 a50088a <=( A167  and  A169 );
 a50089a <=( (not A170)  and  a50088a );
 a50092a <=( A199  and  A166 );
 a50095a <=( (not A232)  and  A200 );
 a50096a <=( a50095a  and  a50092a );
 a50097a <=( a50096a  and  a50089a );
 a50101a <=( (not A266)  and  (not A265) );
 a50102a <=( (not A233)  and  a50101a );
 a50105a <=( (not A299)  and  A298 );
 a50108a <=( A301  and  A300 );
 a50109a <=( a50108a  and  a50105a );
 a50110a <=( a50109a  and  a50102a );
 a50114a <=( A167  and  A169 );
 a50115a <=( (not A170)  and  a50114a );
 a50118a <=( A199  and  A166 );
 a50121a <=( (not A232)  and  A200 );
 a50122a <=( a50121a  and  a50118a );
 a50123a <=( a50122a  and  a50115a );
 a50127a <=( (not A266)  and  (not A265) );
 a50128a <=( (not A233)  and  a50127a );
 a50131a <=( (not A299)  and  A298 );
 a50134a <=( A302  and  A300 );
 a50135a <=( a50134a  and  a50131a );
 a50136a <=( a50135a  and  a50128a );
 a50140a <=( A167  and  A169 );
 a50141a <=( (not A170)  and  a50140a );
 a50144a <=( (not A200)  and  A166 );
 a50147a <=( (not A203)  and  (not A202) );
 a50148a <=( a50147a  and  a50144a );
 a50149a <=( a50148a  and  a50141a );
 a50153a <=( A265  and  A233 );
 a50154a <=( A232  and  a50153a );
 a50157a <=( (not A269)  and  (not A268) );
 a50160a <=( A299  and  (not A298) );
 a50161a <=( a50160a  and  a50157a );
 a50162a <=( a50161a  and  a50154a );
 a50166a <=( A167  and  A169 );
 a50167a <=( (not A170)  and  a50166a );
 a50170a <=( (not A200)  and  A166 );
 a50173a <=( (not A203)  and  (not A202) );
 a50174a <=( a50173a  and  a50170a );
 a50175a <=( a50174a  and  a50167a );
 a50179a <=( (not A236)  and  (not A235) );
 a50180a <=( (not A233)  and  a50179a );
 a50183a <=( A266  and  A265 );
 a50186a <=( A299  and  (not A298) );
 a50187a <=( a50186a  and  a50183a );
 a50188a <=( a50187a  and  a50180a );
 a50192a <=( A167  and  A169 );
 a50193a <=( (not A170)  and  a50192a );
 a50196a <=( (not A200)  and  A166 );
 a50199a <=( (not A203)  and  (not A202) );
 a50200a <=( a50199a  and  a50196a );
 a50201a <=( a50200a  and  a50193a );
 a50205a <=( (not A236)  and  (not A235) );
 a50206a <=( (not A233)  and  a50205a );
 a50209a <=( (not A267)  and  (not A266) );
 a50212a <=( A299  and  (not A298) );
 a50213a <=( a50212a  and  a50209a );
 a50214a <=( a50213a  and  a50206a );
 a50218a <=( A167  and  A169 );
 a50219a <=( (not A170)  and  a50218a );
 a50222a <=( (not A200)  and  A166 );
 a50225a <=( (not A203)  and  (not A202) );
 a50226a <=( a50225a  and  a50222a );
 a50227a <=( a50226a  and  a50219a );
 a50231a <=( (not A236)  and  (not A235) );
 a50232a <=( (not A233)  and  a50231a );
 a50235a <=( (not A266)  and  (not A265) );
 a50238a <=( A299  and  (not A298) );
 a50239a <=( a50238a  and  a50235a );
 a50240a <=( a50239a  and  a50232a );
 a50244a <=( A167  and  A169 );
 a50245a <=( (not A170)  and  a50244a );
 a50248a <=( (not A200)  and  A166 );
 a50251a <=( (not A203)  and  (not A202) );
 a50252a <=( a50251a  and  a50248a );
 a50253a <=( a50252a  and  a50245a );
 a50257a <=( (not A266)  and  (not A234) );
 a50258a <=( (not A233)  and  a50257a );
 a50261a <=( (not A269)  and  (not A268) );
 a50264a <=( A299  and  (not A298) );
 a50265a <=( a50264a  and  a50261a );
 a50266a <=( a50265a  and  a50258a );
 a50270a <=( A167  and  A169 );
 a50271a <=( (not A170)  and  a50270a );
 a50274a <=( (not A200)  and  A166 );
 a50277a <=( (not A203)  and  (not A202) );
 a50278a <=( a50277a  and  a50274a );
 a50279a <=( a50278a  and  a50271a );
 a50283a <=( A234  and  (not A233) );
 a50284a <=( A232  and  a50283a );
 a50287a <=( A298  and  A235 );
 a50290a <=( (not A302)  and  (not A301) );
 a50291a <=( a50290a  and  a50287a );
 a50292a <=( a50291a  and  a50284a );
 a50296a <=( A167  and  A169 );
 a50297a <=( (not A170)  and  a50296a );
 a50300a <=( (not A200)  and  A166 );
 a50303a <=( (not A203)  and  (not A202) );
 a50304a <=( a50303a  and  a50300a );
 a50305a <=( a50304a  and  a50297a );
 a50309a <=( A234  and  (not A233) );
 a50310a <=( A232  and  a50309a );
 a50313a <=( A298  and  A236 );
 a50316a <=( (not A302)  and  (not A301) );
 a50317a <=( a50316a  and  a50313a );
 a50318a <=( a50317a  and  a50310a );
 a50322a <=( A167  and  A169 );
 a50323a <=( (not A170)  and  a50322a );
 a50326a <=( (not A200)  and  A166 );
 a50329a <=( (not A203)  and  (not A202) );
 a50330a <=( a50329a  and  a50326a );
 a50331a <=( a50330a  and  a50323a );
 a50335a <=( (not A266)  and  (not A233) );
 a50336a <=( (not A232)  and  a50335a );
 a50339a <=( (not A269)  and  (not A268) );
 a50342a <=( A299  and  (not A298) );
 a50343a <=( a50342a  and  a50339a );
 a50344a <=( a50343a  and  a50336a );
 a50348a <=( A167  and  A169 );
 a50349a <=( (not A170)  and  a50348a );
 a50352a <=( (not A200)  and  A166 );
 a50355a <=( A232  and  (not A201) );
 a50356a <=( a50355a  and  a50352a );
 a50357a <=( a50356a  and  a50349a );
 a50361a <=( (not A267)  and  A265 );
 a50362a <=( A233  and  a50361a );
 a50365a <=( (not A299)  and  A298 );
 a50368a <=( A301  and  A300 );
 a50369a <=( a50368a  and  a50365a );
 a50370a <=( a50369a  and  a50362a );
 a50374a <=( A167  and  A169 );
 a50375a <=( (not A170)  and  a50374a );
 a50378a <=( (not A200)  and  A166 );
 a50381a <=( A232  and  (not A201) );
 a50382a <=( a50381a  and  a50378a );
 a50383a <=( a50382a  and  a50375a );
 a50387a <=( (not A267)  and  A265 );
 a50388a <=( A233  and  a50387a );
 a50391a <=( (not A299)  and  A298 );
 a50394a <=( A302  and  A300 );
 a50395a <=( a50394a  and  a50391a );
 a50396a <=( a50395a  and  a50388a );
 a50400a <=( A167  and  A169 );
 a50401a <=( (not A170)  and  a50400a );
 a50404a <=( (not A200)  and  A166 );
 a50407a <=( A232  and  (not A201) );
 a50408a <=( a50407a  and  a50404a );
 a50409a <=( a50408a  and  a50401a );
 a50413a <=( A266  and  A265 );
 a50414a <=( A233  and  a50413a );
 a50417a <=( (not A299)  and  A298 );
 a50420a <=( A301  and  A300 );
 a50421a <=( a50420a  and  a50417a );
 a50422a <=( a50421a  and  a50414a );
 a50426a <=( A167  and  A169 );
 a50427a <=( (not A170)  and  a50426a );
 a50430a <=( (not A200)  and  A166 );
 a50433a <=( A232  and  (not A201) );
 a50434a <=( a50433a  and  a50430a );
 a50435a <=( a50434a  and  a50427a );
 a50439a <=( A266  and  A265 );
 a50440a <=( A233  and  a50439a );
 a50443a <=( (not A299)  and  A298 );
 a50446a <=( A302  and  A300 );
 a50447a <=( a50446a  and  a50443a );
 a50448a <=( a50447a  and  a50440a );
 a50452a <=( A167  and  A169 );
 a50453a <=( (not A170)  and  a50452a );
 a50456a <=( (not A200)  and  A166 );
 a50459a <=( A232  and  (not A201) );
 a50460a <=( a50459a  and  a50456a );
 a50461a <=( a50460a  and  a50453a );
 a50465a <=( (not A266)  and  (not A265) );
 a50466a <=( A233  and  a50465a );
 a50469a <=( (not A299)  and  A298 );
 a50472a <=( A301  and  A300 );
 a50473a <=( a50472a  and  a50469a );
 a50474a <=( a50473a  and  a50466a );
 a50478a <=( A167  and  A169 );
 a50479a <=( (not A170)  and  a50478a );
 a50482a <=( (not A200)  and  A166 );
 a50485a <=( A232  and  (not A201) );
 a50486a <=( a50485a  and  a50482a );
 a50487a <=( a50486a  and  a50479a );
 a50491a <=( (not A266)  and  (not A265) );
 a50492a <=( A233  and  a50491a );
 a50495a <=( (not A299)  and  A298 );
 a50498a <=( A302  and  A300 );
 a50499a <=( a50498a  and  a50495a );
 a50500a <=( a50499a  and  a50492a );
 a50504a <=( A167  and  A169 );
 a50505a <=( (not A170)  and  a50504a );
 a50508a <=( (not A200)  and  A166 );
 a50511a <=( (not A233)  and  (not A201) );
 a50512a <=( a50511a  and  a50508a );
 a50513a <=( a50512a  and  a50505a );
 a50517a <=( (not A266)  and  (not A236) );
 a50518a <=( (not A235)  and  a50517a );
 a50521a <=( (not A269)  and  (not A268) );
 a50524a <=( A299  and  (not A298) );
 a50525a <=( a50524a  and  a50521a );
 a50526a <=( a50525a  and  a50518a );
 a50530a <=( A167  and  A169 );
 a50531a <=( (not A170)  and  a50530a );
 a50534a <=( (not A200)  and  A166 );
 a50537a <=( (not A233)  and  (not A201) );
 a50538a <=( a50537a  and  a50534a );
 a50539a <=( a50538a  and  a50531a );
 a50543a <=( A266  and  A265 );
 a50544a <=( (not A234)  and  a50543a );
 a50547a <=( (not A299)  and  A298 );
 a50550a <=( A301  and  A300 );
 a50551a <=( a50550a  and  a50547a );
 a50552a <=( a50551a  and  a50544a );
 a50556a <=( A167  and  A169 );
 a50557a <=( (not A170)  and  a50556a );
 a50560a <=( (not A200)  and  A166 );
 a50563a <=( (not A233)  and  (not A201) );
 a50564a <=( a50563a  and  a50560a );
 a50565a <=( a50564a  and  a50557a );
 a50569a <=( A266  and  A265 );
 a50570a <=( (not A234)  and  a50569a );
 a50573a <=( (not A299)  and  A298 );
 a50576a <=( A302  and  A300 );
 a50577a <=( a50576a  and  a50573a );
 a50578a <=( a50577a  and  a50570a );
 a50582a <=( A167  and  A169 );
 a50583a <=( (not A170)  and  a50582a );
 a50586a <=( (not A200)  and  A166 );
 a50589a <=( (not A233)  and  (not A201) );
 a50590a <=( a50589a  and  a50586a );
 a50591a <=( a50590a  and  a50583a );
 a50595a <=( (not A267)  and  (not A266) );
 a50596a <=( (not A234)  and  a50595a );
 a50599a <=( (not A299)  and  A298 );
 a50602a <=( A301  and  A300 );
 a50603a <=( a50602a  and  a50599a );
 a50604a <=( a50603a  and  a50596a );
 a50608a <=( A167  and  A169 );
 a50609a <=( (not A170)  and  a50608a );
 a50612a <=( (not A200)  and  A166 );
 a50615a <=( (not A233)  and  (not A201) );
 a50616a <=( a50615a  and  a50612a );
 a50617a <=( a50616a  and  a50609a );
 a50621a <=( (not A267)  and  (not A266) );
 a50622a <=( (not A234)  and  a50621a );
 a50625a <=( (not A299)  and  A298 );
 a50628a <=( A302  and  A300 );
 a50629a <=( a50628a  and  a50625a );
 a50630a <=( a50629a  and  a50622a );
 a50634a <=( A167  and  A169 );
 a50635a <=( (not A170)  and  a50634a );
 a50638a <=( (not A200)  and  A166 );
 a50641a <=( (not A233)  and  (not A201) );
 a50642a <=( a50641a  and  a50638a );
 a50643a <=( a50642a  and  a50635a );
 a50647a <=( (not A266)  and  (not A265) );
 a50648a <=( (not A234)  and  a50647a );
 a50651a <=( (not A299)  and  A298 );
 a50654a <=( A301  and  A300 );
 a50655a <=( a50654a  and  a50651a );
 a50656a <=( a50655a  and  a50648a );
 a50660a <=( A167  and  A169 );
 a50661a <=( (not A170)  and  a50660a );
 a50664a <=( (not A200)  and  A166 );
 a50667a <=( (not A233)  and  (not A201) );
 a50668a <=( a50667a  and  a50664a );
 a50669a <=( a50668a  and  a50661a );
 a50673a <=( (not A266)  and  (not A265) );
 a50674a <=( (not A234)  and  a50673a );
 a50677a <=( (not A299)  and  A298 );
 a50680a <=( A302  and  A300 );
 a50681a <=( a50680a  and  a50677a );
 a50682a <=( a50681a  and  a50674a );
 a50686a <=( A167  and  A169 );
 a50687a <=( (not A170)  and  a50686a );
 a50690a <=( (not A200)  and  A166 );
 a50693a <=( A232  and  (not A201) );
 a50694a <=( a50693a  and  a50690a );
 a50695a <=( a50694a  and  a50687a );
 a50699a <=( A235  and  A234 );
 a50700a <=( (not A233)  and  a50699a );
 a50703a <=( (not A266)  and  A265 );
 a50706a <=( A268  and  A267 );
 a50707a <=( a50706a  and  a50703a );
 a50708a <=( a50707a  and  a50700a );
 a50712a <=( A167  and  A169 );
 a50713a <=( (not A170)  and  a50712a );
 a50716a <=( (not A200)  and  A166 );
 a50719a <=( A232  and  (not A201) );
 a50720a <=( a50719a  and  a50716a );
 a50721a <=( a50720a  and  a50713a );
 a50725a <=( A235  and  A234 );
 a50726a <=( (not A233)  and  a50725a );
 a50729a <=( (not A266)  and  A265 );
 a50732a <=( A269  and  A267 );
 a50733a <=( a50732a  and  a50729a );
 a50734a <=( a50733a  and  a50726a );
 a50738a <=( A167  and  A169 );
 a50739a <=( (not A170)  and  a50738a );
 a50742a <=( (not A200)  and  A166 );
 a50745a <=( A232  and  (not A201) );
 a50746a <=( a50745a  and  a50742a );
 a50747a <=( a50746a  and  a50739a );
 a50751a <=( A236  and  A234 );
 a50752a <=( (not A233)  and  a50751a );
 a50755a <=( (not A266)  and  A265 );
 a50758a <=( A268  and  A267 );
 a50759a <=( a50758a  and  a50755a );
 a50760a <=( a50759a  and  a50752a );
 a50764a <=( A167  and  A169 );
 a50765a <=( (not A170)  and  a50764a );
 a50768a <=( (not A200)  and  A166 );
 a50771a <=( A232  and  (not A201) );
 a50772a <=( a50771a  and  a50768a );
 a50773a <=( a50772a  and  a50765a );
 a50777a <=( A236  and  A234 );
 a50778a <=( (not A233)  and  a50777a );
 a50781a <=( (not A266)  and  A265 );
 a50784a <=( A269  and  A267 );
 a50785a <=( a50784a  and  a50781a );
 a50786a <=( a50785a  and  a50778a );
 a50790a <=( A167  and  A169 );
 a50791a <=( (not A170)  and  a50790a );
 a50794a <=( (not A200)  and  A166 );
 a50797a <=( (not A232)  and  (not A201) );
 a50798a <=( a50797a  and  a50794a );
 a50799a <=( a50798a  and  a50791a );
 a50803a <=( A266  and  A265 );
 a50804a <=( (not A233)  and  a50803a );
 a50807a <=( (not A299)  and  A298 );
 a50810a <=( A301  and  A300 );
 a50811a <=( a50810a  and  a50807a );
 a50812a <=( a50811a  and  a50804a );
 a50816a <=( A167  and  A169 );
 a50817a <=( (not A170)  and  a50816a );
 a50820a <=( (not A200)  and  A166 );
 a50823a <=( (not A232)  and  (not A201) );
 a50824a <=( a50823a  and  a50820a );
 a50825a <=( a50824a  and  a50817a );
 a50829a <=( A266  and  A265 );
 a50830a <=( (not A233)  and  a50829a );
 a50833a <=( (not A299)  and  A298 );
 a50836a <=( A302  and  A300 );
 a50837a <=( a50836a  and  a50833a );
 a50838a <=( a50837a  and  a50830a );
 a50842a <=( A167  and  A169 );
 a50843a <=( (not A170)  and  a50842a );
 a50846a <=( (not A200)  and  A166 );
 a50849a <=( (not A232)  and  (not A201) );
 a50850a <=( a50849a  and  a50846a );
 a50851a <=( a50850a  and  a50843a );
 a50855a <=( (not A267)  and  (not A266) );
 a50856a <=( (not A233)  and  a50855a );
 a50859a <=( (not A299)  and  A298 );
 a50862a <=( A301  and  A300 );
 a50863a <=( a50862a  and  a50859a );
 a50864a <=( a50863a  and  a50856a );
 a50868a <=( A167  and  A169 );
 a50869a <=( (not A170)  and  a50868a );
 a50872a <=( (not A200)  and  A166 );
 a50875a <=( (not A232)  and  (not A201) );
 a50876a <=( a50875a  and  a50872a );
 a50877a <=( a50876a  and  a50869a );
 a50881a <=( (not A267)  and  (not A266) );
 a50882a <=( (not A233)  and  a50881a );
 a50885a <=( (not A299)  and  A298 );
 a50888a <=( A302  and  A300 );
 a50889a <=( a50888a  and  a50885a );
 a50890a <=( a50889a  and  a50882a );
 a50894a <=( A167  and  A169 );
 a50895a <=( (not A170)  and  a50894a );
 a50898a <=( (not A200)  and  A166 );
 a50901a <=( (not A232)  and  (not A201) );
 a50902a <=( a50901a  and  a50898a );
 a50903a <=( a50902a  and  a50895a );
 a50907a <=( (not A266)  and  (not A265) );
 a50908a <=( (not A233)  and  a50907a );
 a50911a <=( (not A299)  and  A298 );
 a50914a <=( A301  and  A300 );
 a50915a <=( a50914a  and  a50911a );
 a50916a <=( a50915a  and  a50908a );
 a50920a <=( A167  and  A169 );
 a50921a <=( (not A170)  and  a50920a );
 a50924a <=( (not A200)  and  A166 );
 a50927a <=( (not A232)  and  (not A201) );
 a50928a <=( a50927a  and  a50924a );
 a50929a <=( a50928a  and  a50921a );
 a50933a <=( (not A266)  and  (not A265) );
 a50934a <=( (not A233)  and  a50933a );
 a50937a <=( (not A299)  and  A298 );
 a50940a <=( A302  and  A300 );
 a50941a <=( a50940a  and  a50937a );
 a50942a <=( a50941a  and  a50934a );
 a50946a <=( A167  and  A169 );
 a50947a <=( (not A170)  and  a50946a );
 a50950a <=( (not A199)  and  A166 );
 a50953a <=( A232  and  (not A200) );
 a50954a <=( a50953a  and  a50950a );
 a50955a <=( a50954a  and  a50947a );
 a50959a <=( (not A267)  and  A265 );
 a50960a <=( A233  and  a50959a );
 a50963a <=( (not A299)  and  A298 );
 a50966a <=( A301  and  A300 );
 a50967a <=( a50966a  and  a50963a );
 a50968a <=( a50967a  and  a50960a );
 a50972a <=( A167  and  A169 );
 a50973a <=( (not A170)  and  a50972a );
 a50976a <=( (not A199)  and  A166 );
 a50979a <=( A232  and  (not A200) );
 a50980a <=( a50979a  and  a50976a );
 a50981a <=( a50980a  and  a50973a );
 a50985a <=( (not A267)  and  A265 );
 a50986a <=( A233  and  a50985a );
 a50989a <=( (not A299)  and  A298 );
 a50992a <=( A302  and  A300 );
 a50993a <=( a50992a  and  a50989a );
 a50994a <=( a50993a  and  a50986a );
 a50998a <=( A167  and  A169 );
 a50999a <=( (not A170)  and  a50998a );
 a51002a <=( (not A199)  and  A166 );
 a51005a <=( A232  and  (not A200) );
 a51006a <=( a51005a  and  a51002a );
 a51007a <=( a51006a  and  a50999a );
 a51011a <=( A266  and  A265 );
 a51012a <=( A233  and  a51011a );
 a51015a <=( (not A299)  and  A298 );
 a51018a <=( A301  and  A300 );
 a51019a <=( a51018a  and  a51015a );
 a51020a <=( a51019a  and  a51012a );
 a51024a <=( A167  and  A169 );
 a51025a <=( (not A170)  and  a51024a );
 a51028a <=( (not A199)  and  A166 );
 a51031a <=( A232  and  (not A200) );
 a51032a <=( a51031a  and  a51028a );
 a51033a <=( a51032a  and  a51025a );
 a51037a <=( A266  and  A265 );
 a51038a <=( A233  and  a51037a );
 a51041a <=( (not A299)  and  A298 );
 a51044a <=( A302  and  A300 );
 a51045a <=( a51044a  and  a51041a );
 a51046a <=( a51045a  and  a51038a );
 a51050a <=( A167  and  A169 );
 a51051a <=( (not A170)  and  a51050a );
 a51054a <=( (not A199)  and  A166 );
 a51057a <=( A232  and  (not A200) );
 a51058a <=( a51057a  and  a51054a );
 a51059a <=( a51058a  and  a51051a );
 a51063a <=( (not A266)  and  (not A265) );
 a51064a <=( A233  and  a51063a );
 a51067a <=( (not A299)  and  A298 );
 a51070a <=( A301  and  A300 );
 a51071a <=( a51070a  and  a51067a );
 a51072a <=( a51071a  and  a51064a );
 a51076a <=( A167  and  A169 );
 a51077a <=( (not A170)  and  a51076a );
 a51080a <=( (not A199)  and  A166 );
 a51083a <=( A232  and  (not A200) );
 a51084a <=( a51083a  and  a51080a );
 a51085a <=( a51084a  and  a51077a );
 a51089a <=( (not A266)  and  (not A265) );
 a51090a <=( A233  and  a51089a );
 a51093a <=( (not A299)  and  A298 );
 a51096a <=( A302  and  A300 );
 a51097a <=( a51096a  and  a51093a );
 a51098a <=( a51097a  and  a51090a );
 a51102a <=( A167  and  A169 );
 a51103a <=( (not A170)  and  a51102a );
 a51106a <=( (not A199)  and  A166 );
 a51109a <=( (not A233)  and  (not A200) );
 a51110a <=( a51109a  and  a51106a );
 a51111a <=( a51110a  and  a51103a );
 a51115a <=( (not A266)  and  (not A236) );
 a51116a <=( (not A235)  and  a51115a );
 a51119a <=( (not A269)  and  (not A268) );
 a51122a <=( A299  and  (not A298) );
 a51123a <=( a51122a  and  a51119a );
 a51124a <=( a51123a  and  a51116a );
 a51128a <=( A167  and  A169 );
 a51129a <=( (not A170)  and  a51128a );
 a51132a <=( (not A199)  and  A166 );
 a51135a <=( (not A233)  and  (not A200) );
 a51136a <=( a51135a  and  a51132a );
 a51137a <=( a51136a  and  a51129a );
 a51141a <=( A266  and  A265 );
 a51142a <=( (not A234)  and  a51141a );
 a51145a <=( (not A299)  and  A298 );
 a51148a <=( A301  and  A300 );
 a51149a <=( a51148a  and  a51145a );
 a51150a <=( a51149a  and  a51142a );
 a51154a <=( A167  and  A169 );
 a51155a <=( (not A170)  and  a51154a );
 a51158a <=( (not A199)  and  A166 );
 a51161a <=( (not A233)  and  (not A200) );
 a51162a <=( a51161a  and  a51158a );
 a51163a <=( a51162a  and  a51155a );
 a51167a <=( A266  and  A265 );
 a51168a <=( (not A234)  and  a51167a );
 a51171a <=( (not A299)  and  A298 );
 a51174a <=( A302  and  A300 );
 a51175a <=( a51174a  and  a51171a );
 a51176a <=( a51175a  and  a51168a );
 a51180a <=( A167  and  A169 );
 a51181a <=( (not A170)  and  a51180a );
 a51184a <=( (not A199)  and  A166 );
 a51187a <=( (not A233)  and  (not A200) );
 a51188a <=( a51187a  and  a51184a );
 a51189a <=( a51188a  and  a51181a );
 a51193a <=( (not A267)  and  (not A266) );
 a51194a <=( (not A234)  and  a51193a );
 a51197a <=( (not A299)  and  A298 );
 a51200a <=( A301  and  A300 );
 a51201a <=( a51200a  and  a51197a );
 a51202a <=( a51201a  and  a51194a );
 a51206a <=( A167  and  A169 );
 a51207a <=( (not A170)  and  a51206a );
 a51210a <=( (not A199)  and  A166 );
 a51213a <=( (not A233)  and  (not A200) );
 a51214a <=( a51213a  and  a51210a );
 a51215a <=( a51214a  and  a51207a );
 a51219a <=( (not A267)  and  (not A266) );
 a51220a <=( (not A234)  and  a51219a );
 a51223a <=( (not A299)  and  A298 );
 a51226a <=( A302  and  A300 );
 a51227a <=( a51226a  and  a51223a );
 a51228a <=( a51227a  and  a51220a );
 a51232a <=( A167  and  A169 );
 a51233a <=( (not A170)  and  a51232a );
 a51236a <=( (not A199)  and  A166 );
 a51239a <=( (not A233)  and  (not A200) );
 a51240a <=( a51239a  and  a51236a );
 a51241a <=( a51240a  and  a51233a );
 a51245a <=( (not A266)  and  (not A265) );
 a51246a <=( (not A234)  and  a51245a );
 a51249a <=( (not A299)  and  A298 );
 a51252a <=( A301  and  A300 );
 a51253a <=( a51252a  and  a51249a );
 a51254a <=( a51253a  and  a51246a );
 a51258a <=( A167  and  A169 );
 a51259a <=( (not A170)  and  a51258a );
 a51262a <=( (not A199)  and  A166 );
 a51265a <=( (not A233)  and  (not A200) );
 a51266a <=( a51265a  and  a51262a );
 a51267a <=( a51266a  and  a51259a );
 a51271a <=( (not A266)  and  (not A265) );
 a51272a <=( (not A234)  and  a51271a );
 a51275a <=( (not A299)  and  A298 );
 a51278a <=( A302  and  A300 );
 a51279a <=( a51278a  and  a51275a );
 a51280a <=( a51279a  and  a51272a );
 a51284a <=( A167  and  A169 );
 a51285a <=( (not A170)  and  a51284a );
 a51288a <=( (not A199)  and  A166 );
 a51291a <=( A232  and  (not A200) );
 a51292a <=( a51291a  and  a51288a );
 a51293a <=( a51292a  and  a51285a );
 a51297a <=( A235  and  A234 );
 a51298a <=( (not A233)  and  a51297a );
 a51301a <=( (not A266)  and  A265 );
 a51304a <=( A268  and  A267 );
 a51305a <=( a51304a  and  a51301a );
 a51306a <=( a51305a  and  a51298a );
 a51310a <=( A167  and  A169 );
 a51311a <=( (not A170)  and  a51310a );
 a51314a <=( (not A199)  and  A166 );
 a51317a <=( A232  and  (not A200) );
 a51318a <=( a51317a  and  a51314a );
 a51319a <=( a51318a  and  a51311a );
 a51323a <=( A235  and  A234 );
 a51324a <=( (not A233)  and  a51323a );
 a51327a <=( (not A266)  and  A265 );
 a51330a <=( A269  and  A267 );
 a51331a <=( a51330a  and  a51327a );
 a51332a <=( a51331a  and  a51324a );
 a51336a <=( A167  and  A169 );
 a51337a <=( (not A170)  and  a51336a );
 a51340a <=( (not A199)  and  A166 );
 a51343a <=( A232  and  (not A200) );
 a51344a <=( a51343a  and  a51340a );
 a51345a <=( a51344a  and  a51337a );
 a51349a <=( A236  and  A234 );
 a51350a <=( (not A233)  and  a51349a );
 a51353a <=( (not A266)  and  A265 );
 a51356a <=( A268  and  A267 );
 a51357a <=( a51356a  and  a51353a );
 a51358a <=( a51357a  and  a51350a );
 a51362a <=( A167  and  A169 );
 a51363a <=( (not A170)  and  a51362a );
 a51366a <=( (not A199)  and  A166 );
 a51369a <=( A232  and  (not A200) );
 a51370a <=( a51369a  and  a51366a );
 a51371a <=( a51370a  and  a51363a );
 a51375a <=( A236  and  A234 );
 a51376a <=( (not A233)  and  a51375a );
 a51379a <=( (not A266)  and  A265 );
 a51382a <=( A269  and  A267 );
 a51383a <=( a51382a  and  a51379a );
 a51384a <=( a51383a  and  a51376a );
 a51388a <=( A167  and  A169 );
 a51389a <=( (not A170)  and  a51388a );
 a51392a <=( (not A199)  and  A166 );
 a51395a <=( (not A232)  and  (not A200) );
 a51396a <=( a51395a  and  a51392a );
 a51397a <=( a51396a  and  a51389a );
 a51401a <=( A266  and  A265 );
 a51402a <=( (not A233)  and  a51401a );
 a51405a <=( (not A299)  and  A298 );
 a51408a <=( A301  and  A300 );
 a51409a <=( a51408a  and  a51405a );
 a51410a <=( a51409a  and  a51402a );
 a51414a <=( A167  and  A169 );
 a51415a <=( (not A170)  and  a51414a );
 a51418a <=( (not A199)  and  A166 );
 a51421a <=( (not A232)  and  (not A200) );
 a51422a <=( a51421a  and  a51418a );
 a51423a <=( a51422a  and  a51415a );
 a51427a <=( A266  and  A265 );
 a51428a <=( (not A233)  and  a51427a );
 a51431a <=( (not A299)  and  A298 );
 a51434a <=( A302  and  A300 );
 a51435a <=( a51434a  and  a51431a );
 a51436a <=( a51435a  and  a51428a );
 a51440a <=( A167  and  A169 );
 a51441a <=( (not A170)  and  a51440a );
 a51444a <=( (not A199)  and  A166 );
 a51447a <=( (not A232)  and  (not A200) );
 a51448a <=( a51447a  and  a51444a );
 a51449a <=( a51448a  and  a51441a );
 a51453a <=( (not A267)  and  (not A266) );
 a51454a <=( (not A233)  and  a51453a );
 a51457a <=( (not A299)  and  A298 );
 a51460a <=( A301  and  A300 );
 a51461a <=( a51460a  and  a51457a );
 a51462a <=( a51461a  and  a51454a );
 a51466a <=( A167  and  A169 );
 a51467a <=( (not A170)  and  a51466a );
 a51470a <=( (not A199)  and  A166 );
 a51473a <=( (not A232)  and  (not A200) );
 a51474a <=( a51473a  and  a51470a );
 a51475a <=( a51474a  and  a51467a );
 a51479a <=( (not A267)  and  (not A266) );
 a51480a <=( (not A233)  and  a51479a );
 a51483a <=( (not A299)  and  A298 );
 a51486a <=( A302  and  A300 );
 a51487a <=( a51486a  and  a51483a );
 a51488a <=( a51487a  and  a51480a );
 a51492a <=( A167  and  A169 );
 a51493a <=( (not A170)  and  a51492a );
 a51496a <=( (not A199)  and  A166 );
 a51499a <=( (not A232)  and  (not A200) );
 a51500a <=( a51499a  and  a51496a );
 a51501a <=( a51500a  and  a51493a );
 a51505a <=( (not A266)  and  (not A265) );
 a51506a <=( (not A233)  and  a51505a );
 a51509a <=( (not A299)  and  A298 );
 a51512a <=( A301  and  A300 );
 a51513a <=( a51512a  and  a51509a );
 a51514a <=( a51513a  and  a51506a );
 a51518a <=( A167  and  A169 );
 a51519a <=( (not A170)  and  a51518a );
 a51522a <=( (not A199)  and  A166 );
 a51525a <=( (not A232)  and  (not A200) );
 a51526a <=( a51525a  and  a51522a );
 a51527a <=( a51526a  and  a51519a );
 a51531a <=( (not A266)  and  (not A265) );
 a51532a <=( (not A233)  and  a51531a );
 a51535a <=( (not A299)  and  A298 );
 a51538a <=( A302  and  A300 );
 a51539a <=( a51538a  and  a51535a );
 a51540a <=( a51539a  and  a51532a );
 a51544a <=( (not A167)  and  A169 );
 a51545a <=( (not A170)  and  a51544a );
 a51548a <=( A199  and  (not A166) );
 a51551a <=( A232  and  A200 );
 a51552a <=( a51551a  and  a51548a );
 a51553a <=( a51552a  and  a51545a );
 a51557a <=( (not A267)  and  A265 );
 a51558a <=( A233  and  a51557a );
 a51561a <=( (not A299)  and  A298 );
 a51564a <=( A301  and  A300 );
 a51565a <=( a51564a  and  a51561a );
 a51566a <=( a51565a  and  a51558a );
 a51570a <=( (not A167)  and  A169 );
 a51571a <=( (not A170)  and  a51570a );
 a51574a <=( A199  and  (not A166) );
 a51577a <=( A232  and  A200 );
 a51578a <=( a51577a  and  a51574a );
 a51579a <=( a51578a  and  a51571a );
 a51583a <=( (not A267)  and  A265 );
 a51584a <=( A233  and  a51583a );
 a51587a <=( (not A299)  and  A298 );
 a51590a <=( A302  and  A300 );
 a51591a <=( a51590a  and  a51587a );
 a51592a <=( a51591a  and  a51584a );
 a51596a <=( (not A167)  and  A169 );
 a51597a <=( (not A170)  and  a51596a );
 a51600a <=( A199  and  (not A166) );
 a51603a <=( A232  and  A200 );
 a51604a <=( a51603a  and  a51600a );
 a51605a <=( a51604a  and  a51597a );
 a51609a <=( A266  and  A265 );
 a51610a <=( A233  and  a51609a );
 a51613a <=( (not A299)  and  A298 );
 a51616a <=( A301  and  A300 );
 a51617a <=( a51616a  and  a51613a );
 a51618a <=( a51617a  and  a51610a );
 a51622a <=( (not A167)  and  A169 );
 a51623a <=( (not A170)  and  a51622a );
 a51626a <=( A199  and  (not A166) );
 a51629a <=( A232  and  A200 );
 a51630a <=( a51629a  and  a51626a );
 a51631a <=( a51630a  and  a51623a );
 a51635a <=( A266  and  A265 );
 a51636a <=( A233  and  a51635a );
 a51639a <=( (not A299)  and  A298 );
 a51642a <=( A302  and  A300 );
 a51643a <=( a51642a  and  a51639a );
 a51644a <=( a51643a  and  a51636a );
 a51648a <=( (not A167)  and  A169 );
 a51649a <=( (not A170)  and  a51648a );
 a51652a <=( A199  and  (not A166) );
 a51655a <=( A232  and  A200 );
 a51656a <=( a51655a  and  a51652a );
 a51657a <=( a51656a  and  a51649a );
 a51661a <=( (not A266)  and  (not A265) );
 a51662a <=( A233  and  a51661a );
 a51665a <=( (not A299)  and  A298 );
 a51668a <=( A301  and  A300 );
 a51669a <=( a51668a  and  a51665a );
 a51670a <=( a51669a  and  a51662a );
 a51674a <=( (not A167)  and  A169 );
 a51675a <=( (not A170)  and  a51674a );
 a51678a <=( A199  and  (not A166) );
 a51681a <=( A232  and  A200 );
 a51682a <=( a51681a  and  a51678a );
 a51683a <=( a51682a  and  a51675a );
 a51687a <=( (not A266)  and  (not A265) );
 a51688a <=( A233  and  a51687a );
 a51691a <=( (not A299)  and  A298 );
 a51694a <=( A302  and  A300 );
 a51695a <=( a51694a  and  a51691a );
 a51696a <=( a51695a  and  a51688a );
 a51700a <=( (not A167)  and  A169 );
 a51701a <=( (not A170)  and  a51700a );
 a51704a <=( A199  and  (not A166) );
 a51707a <=( (not A233)  and  A200 );
 a51708a <=( a51707a  and  a51704a );
 a51709a <=( a51708a  and  a51701a );
 a51713a <=( (not A266)  and  (not A236) );
 a51714a <=( (not A235)  and  a51713a );
 a51717a <=( (not A269)  and  (not A268) );
 a51720a <=( A299  and  (not A298) );
 a51721a <=( a51720a  and  a51717a );
 a51722a <=( a51721a  and  a51714a );
 a51726a <=( (not A167)  and  A169 );
 a51727a <=( (not A170)  and  a51726a );
 a51730a <=( A199  and  (not A166) );
 a51733a <=( (not A233)  and  A200 );
 a51734a <=( a51733a  and  a51730a );
 a51735a <=( a51734a  and  a51727a );
 a51739a <=( A266  and  A265 );
 a51740a <=( (not A234)  and  a51739a );
 a51743a <=( (not A299)  and  A298 );
 a51746a <=( A301  and  A300 );
 a51747a <=( a51746a  and  a51743a );
 a51748a <=( a51747a  and  a51740a );
 a51752a <=( (not A167)  and  A169 );
 a51753a <=( (not A170)  and  a51752a );
 a51756a <=( A199  and  (not A166) );
 a51759a <=( (not A233)  and  A200 );
 a51760a <=( a51759a  and  a51756a );
 a51761a <=( a51760a  and  a51753a );
 a51765a <=( A266  and  A265 );
 a51766a <=( (not A234)  and  a51765a );
 a51769a <=( (not A299)  and  A298 );
 a51772a <=( A302  and  A300 );
 a51773a <=( a51772a  and  a51769a );
 a51774a <=( a51773a  and  a51766a );
 a51778a <=( (not A167)  and  A169 );
 a51779a <=( (not A170)  and  a51778a );
 a51782a <=( A199  and  (not A166) );
 a51785a <=( (not A233)  and  A200 );
 a51786a <=( a51785a  and  a51782a );
 a51787a <=( a51786a  and  a51779a );
 a51791a <=( (not A267)  and  (not A266) );
 a51792a <=( (not A234)  and  a51791a );
 a51795a <=( (not A299)  and  A298 );
 a51798a <=( A301  and  A300 );
 a51799a <=( a51798a  and  a51795a );
 a51800a <=( a51799a  and  a51792a );
 a51804a <=( (not A167)  and  A169 );
 a51805a <=( (not A170)  and  a51804a );
 a51808a <=( A199  and  (not A166) );
 a51811a <=( (not A233)  and  A200 );
 a51812a <=( a51811a  and  a51808a );
 a51813a <=( a51812a  and  a51805a );
 a51817a <=( (not A267)  and  (not A266) );
 a51818a <=( (not A234)  and  a51817a );
 a51821a <=( (not A299)  and  A298 );
 a51824a <=( A302  and  A300 );
 a51825a <=( a51824a  and  a51821a );
 a51826a <=( a51825a  and  a51818a );
 a51830a <=( (not A167)  and  A169 );
 a51831a <=( (not A170)  and  a51830a );
 a51834a <=( A199  and  (not A166) );
 a51837a <=( (not A233)  and  A200 );
 a51838a <=( a51837a  and  a51834a );
 a51839a <=( a51838a  and  a51831a );
 a51843a <=( (not A266)  and  (not A265) );
 a51844a <=( (not A234)  and  a51843a );
 a51847a <=( (not A299)  and  A298 );
 a51850a <=( A301  and  A300 );
 a51851a <=( a51850a  and  a51847a );
 a51852a <=( a51851a  and  a51844a );
 a51856a <=( (not A167)  and  A169 );
 a51857a <=( (not A170)  and  a51856a );
 a51860a <=( A199  and  (not A166) );
 a51863a <=( (not A233)  and  A200 );
 a51864a <=( a51863a  and  a51860a );
 a51865a <=( a51864a  and  a51857a );
 a51869a <=( (not A266)  and  (not A265) );
 a51870a <=( (not A234)  and  a51869a );
 a51873a <=( (not A299)  and  A298 );
 a51876a <=( A302  and  A300 );
 a51877a <=( a51876a  and  a51873a );
 a51878a <=( a51877a  and  a51870a );
 a51882a <=( (not A167)  and  A169 );
 a51883a <=( (not A170)  and  a51882a );
 a51886a <=( A199  and  (not A166) );
 a51889a <=( A232  and  A200 );
 a51890a <=( a51889a  and  a51886a );
 a51891a <=( a51890a  and  a51883a );
 a51895a <=( A235  and  A234 );
 a51896a <=( (not A233)  and  a51895a );
 a51899a <=( (not A266)  and  A265 );
 a51902a <=( A268  and  A267 );
 a51903a <=( a51902a  and  a51899a );
 a51904a <=( a51903a  and  a51896a );
 a51908a <=( (not A167)  and  A169 );
 a51909a <=( (not A170)  and  a51908a );
 a51912a <=( A199  and  (not A166) );
 a51915a <=( A232  and  A200 );
 a51916a <=( a51915a  and  a51912a );
 a51917a <=( a51916a  and  a51909a );
 a51921a <=( A235  and  A234 );
 a51922a <=( (not A233)  and  a51921a );
 a51925a <=( (not A266)  and  A265 );
 a51928a <=( A269  and  A267 );
 a51929a <=( a51928a  and  a51925a );
 a51930a <=( a51929a  and  a51922a );
 a51934a <=( (not A167)  and  A169 );
 a51935a <=( (not A170)  and  a51934a );
 a51938a <=( A199  and  (not A166) );
 a51941a <=( A232  and  A200 );
 a51942a <=( a51941a  and  a51938a );
 a51943a <=( a51942a  and  a51935a );
 a51947a <=( A236  and  A234 );
 a51948a <=( (not A233)  and  a51947a );
 a51951a <=( (not A266)  and  A265 );
 a51954a <=( A268  and  A267 );
 a51955a <=( a51954a  and  a51951a );
 a51956a <=( a51955a  and  a51948a );
 a51960a <=( (not A167)  and  A169 );
 a51961a <=( (not A170)  and  a51960a );
 a51964a <=( A199  and  (not A166) );
 a51967a <=( A232  and  A200 );
 a51968a <=( a51967a  and  a51964a );
 a51969a <=( a51968a  and  a51961a );
 a51973a <=( A236  and  A234 );
 a51974a <=( (not A233)  and  a51973a );
 a51977a <=( (not A266)  and  A265 );
 a51980a <=( A269  and  A267 );
 a51981a <=( a51980a  and  a51977a );
 a51982a <=( a51981a  and  a51974a );
 a51986a <=( (not A167)  and  A169 );
 a51987a <=( (not A170)  and  a51986a );
 a51990a <=( A199  and  (not A166) );
 a51993a <=( (not A232)  and  A200 );
 a51994a <=( a51993a  and  a51990a );
 a51995a <=( a51994a  and  a51987a );
 a51999a <=( A266  and  A265 );
 a52000a <=( (not A233)  and  a51999a );
 a52003a <=( (not A299)  and  A298 );
 a52006a <=( A301  and  A300 );
 a52007a <=( a52006a  and  a52003a );
 a52008a <=( a52007a  and  a52000a );
 a52012a <=( (not A167)  and  A169 );
 a52013a <=( (not A170)  and  a52012a );
 a52016a <=( A199  and  (not A166) );
 a52019a <=( (not A232)  and  A200 );
 a52020a <=( a52019a  and  a52016a );
 a52021a <=( a52020a  and  a52013a );
 a52025a <=( A266  and  A265 );
 a52026a <=( (not A233)  and  a52025a );
 a52029a <=( (not A299)  and  A298 );
 a52032a <=( A302  and  A300 );
 a52033a <=( a52032a  and  a52029a );
 a52034a <=( a52033a  and  a52026a );
 a52038a <=( (not A167)  and  A169 );
 a52039a <=( (not A170)  and  a52038a );
 a52042a <=( A199  and  (not A166) );
 a52045a <=( (not A232)  and  A200 );
 a52046a <=( a52045a  and  a52042a );
 a52047a <=( a52046a  and  a52039a );
 a52051a <=( (not A267)  and  (not A266) );
 a52052a <=( (not A233)  and  a52051a );
 a52055a <=( (not A299)  and  A298 );
 a52058a <=( A301  and  A300 );
 a52059a <=( a52058a  and  a52055a );
 a52060a <=( a52059a  and  a52052a );
 a52064a <=( (not A167)  and  A169 );
 a52065a <=( (not A170)  and  a52064a );
 a52068a <=( A199  and  (not A166) );
 a52071a <=( (not A232)  and  A200 );
 a52072a <=( a52071a  and  a52068a );
 a52073a <=( a52072a  and  a52065a );
 a52077a <=( (not A267)  and  (not A266) );
 a52078a <=( (not A233)  and  a52077a );
 a52081a <=( (not A299)  and  A298 );
 a52084a <=( A302  and  A300 );
 a52085a <=( a52084a  and  a52081a );
 a52086a <=( a52085a  and  a52078a );
 a52090a <=( (not A167)  and  A169 );
 a52091a <=( (not A170)  and  a52090a );
 a52094a <=( A199  and  (not A166) );
 a52097a <=( (not A232)  and  A200 );
 a52098a <=( a52097a  and  a52094a );
 a52099a <=( a52098a  and  a52091a );
 a52103a <=( (not A266)  and  (not A265) );
 a52104a <=( (not A233)  and  a52103a );
 a52107a <=( (not A299)  and  A298 );
 a52110a <=( A301  and  A300 );
 a52111a <=( a52110a  and  a52107a );
 a52112a <=( a52111a  and  a52104a );
 a52116a <=( (not A167)  and  A169 );
 a52117a <=( (not A170)  and  a52116a );
 a52120a <=( A199  and  (not A166) );
 a52123a <=( (not A232)  and  A200 );
 a52124a <=( a52123a  and  a52120a );
 a52125a <=( a52124a  and  a52117a );
 a52129a <=( (not A266)  and  (not A265) );
 a52130a <=( (not A233)  and  a52129a );
 a52133a <=( (not A299)  and  A298 );
 a52136a <=( A302  and  A300 );
 a52137a <=( a52136a  and  a52133a );
 a52138a <=( a52137a  and  a52130a );
 a52142a <=( (not A167)  and  A169 );
 a52143a <=( (not A170)  and  a52142a );
 a52146a <=( (not A200)  and  (not A166) );
 a52149a <=( (not A203)  and  (not A202) );
 a52150a <=( a52149a  and  a52146a );
 a52151a <=( a52150a  and  a52143a );
 a52155a <=( A265  and  A233 );
 a52156a <=( A232  and  a52155a );
 a52159a <=( (not A269)  and  (not A268) );
 a52162a <=( A299  and  (not A298) );
 a52163a <=( a52162a  and  a52159a );
 a52164a <=( a52163a  and  a52156a );
 a52168a <=( (not A167)  and  A169 );
 a52169a <=( (not A170)  and  a52168a );
 a52172a <=( (not A200)  and  (not A166) );
 a52175a <=( (not A203)  and  (not A202) );
 a52176a <=( a52175a  and  a52172a );
 a52177a <=( a52176a  and  a52169a );
 a52181a <=( (not A236)  and  (not A235) );
 a52182a <=( (not A233)  and  a52181a );
 a52185a <=( A266  and  A265 );
 a52188a <=( A299  and  (not A298) );
 a52189a <=( a52188a  and  a52185a );
 a52190a <=( a52189a  and  a52182a );
 a52194a <=( (not A167)  and  A169 );
 a52195a <=( (not A170)  and  a52194a );
 a52198a <=( (not A200)  and  (not A166) );
 a52201a <=( (not A203)  and  (not A202) );
 a52202a <=( a52201a  and  a52198a );
 a52203a <=( a52202a  and  a52195a );
 a52207a <=( (not A236)  and  (not A235) );
 a52208a <=( (not A233)  and  a52207a );
 a52211a <=( (not A267)  and  (not A266) );
 a52214a <=( A299  and  (not A298) );
 a52215a <=( a52214a  and  a52211a );
 a52216a <=( a52215a  and  a52208a );
 a52220a <=( (not A167)  and  A169 );
 a52221a <=( (not A170)  and  a52220a );
 a52224a <=( (not A200)  and  (not A166) );
 a52227a <=( (not A203)  and  (not A202) );
 a52228a <=( a52227a  and  a52224a );
 a52229a <=( a52228a  and  a52221a );
 a52233a <=( (not A236)  and  (not A235) );
 a52234a <=( (not A233)  and  a52233a );
 a52237a <=( (not A266)  and  (not A265) );
 a52240a <=( A299  and  (not A298) );
 a52241a <=( a52240a  and  a52237a );
 a52242a <=( a52241a  and  a52234a );
 a52246a <=( (not A167)  and  A169 );
 a52247a <=( (not A170)  and  a52246a );
 a52250a <=( (not A200)  and  (not A166) );
 a52253a <=( (not A203)  and  (not A202) );
 a52254a <=( a52253a  and  a52250a );
 a52255a <=( a52254a  and  a52247a );
 a52259a <=( (not A266)  and  (not A234) );
 a52260a <=( (not A233)  and  a52259a );
 a52263a <=( (not A269)  and  (not A268) );
 a52266a <=( A299  and  (not A298) );
 a52267a <=( a52266a  and  a52263a );
 a52268a <=( a52267a  and  a52260a );
 a52272a <=( (not A167)  and  A169 );
 a52273a <=( (not A170)  and  a52272a );
 a52276a <=( (not A200)  and  (not A166) );
 a52279a <=( (not A203)  and  (not A202) );
 a52280a <=( a52279a  and  a52276a );
 a52281a <=( a52280a  and  a52273a );
 a52285a <=( A234  and  (not A233) );
 a52286a <=( A232  and  a52285a );
 a52289a <=( A298  and  A235 );
 a52292a <=( (not A302)  and  (not A301) );
 a52293a <=( a52292a  and  a52289a );
 a52294a <=( a52293a  and  a52286a );
 a52298a <=( (not A167)  and  A169 );
 a52299a <=( (not A170)  and  a52298a );
 a52302a <=( (not A200)  and  (not A166) );
 a52305a <=( (not A203)  and  (not A202) );
 a52306a <=( a52305a  and  a52302a );
 a52307a <=( a52306a  and  a52299a );
 a52311a <=( A234  and  (not A233) );
 a52312a <=( A232  and  a52311a );
 a52315a <=( A298  and  A236 );
 a52318a <=( (not A302)  and  (not A301) );
 a52319a <=( a52318a  and  a52315a );
 a52320a <=( a52319a  and  a52312a );
 a52324a <=( (not A167)  and  A169 );
 a52325a <=( (not A170)  and  a52324a );
 a52328a <=( (not A200)  and  (not A166) );
 a52331a <=( (not A203)  and  (not A202) );
 a52332a <=( a52331a  and  a52328a );
 a52333a <=( a52332a  and  a52325a );
 a52337a <=( (not A266)  and  (not A233) );
 a52338a <=( (not A232)  and  a52337a );
 a52341a <=( (not A269)  and  (not A268) );
 a52344a <=( A299  and  (not A298) );
 a52345a <=( a52344a  and  a52341a );
 a52346a <=( a52345a  and  a52338a );
 a52350a <=( (not A167)  and  A169 );
 a52351a <=( (not A170)  and  a52350a );
 a52354a <=( (not A200)  and  (not A166) );
 a52357a <=( A232  and  (not A201) );
 a52358a <=( a52357a  and  a52354a );
 a52359a <=( a52358a  and  a52351a );
 a52363a <=( (not A267)  and  A265 );
 a52364a <=( A233  and  a52363a );
 a52367a <=( (not A299)  and  A298 );
 a52370a <=( A301  and  A300 );
 a52371a <=( a52370a  and  a52367a );
 a52372a <=( a52371a  and  a52364a );
 a52376a <=( (not A167)  and  A169 );
 a52377a <=( (not A170)  and  a52376a );
 a52380a <=( (not A200)  and  (not A166) );
 a52383a <=( A232  and  (not A201) );
 a52384a <=( a52383a  and  a52380a );
 a52385a <=( a52384a  and  a52377a );
 a52389a <=( (not A267)  and  A265 );
 a52390a <=( A233  and  a52389a );
 a52393a <=( (not A299)  and  A298 );
 a52396a <=( A302  and  A300 );
 a52397a <=( a52396a  and  a52393a );
 a52398a <=( a52397a  and  a52390a );
 a52402a <=( (not A167)  and  A169 );
 a52403a <=( (not A170)  and  a52402a );
 a52406a <=( (not A200)  and  (not A166) );
 a52409a <=( A232  and  (not A201) );
 a52410a <=( a52409a  and  a52406a );
 a52411a <=( a52410a  and  a52403a );
 a52415a <=( A266  and  A265 );
 a52416a <=( A233  and  a52415a );
 a52419a <=( (not A299)  and  A298 );
 a52422a <=( A301  and  A300 );
 a52423a <=( a52422a  and  a52419a );
 a52424a <=( a52423a  and  a52416a );
 a52428a <=( (not A167)  and  A169 );
 a52429a <=( (not A170)  and  a52428a );
 a52432a <=( (not A200)  and  (not A166) );
 a52435a <=( A232  and  (not A201) );
 a52436a <=( a52435a  and  a52432a );
 a52437a <=( a52436a  and  a52429a );
 a52441a <=( A266  and  A265 );
 a52442a <=( A233  and  a52441a );
 a52445a <=( (not A299)  and  A298 );
 a52448a <=( A302  and  A300 );
 a52449a <=( a52448a  and  a52445a );
 a52450a <=( a52449a  and  a52442a );
 a52454a <=( (not A167)  and  A169 );
 a52455a <=( (not A170)  and  a52454a );
 a52458a <=( (not A200)  and  (not A166) );
 a52461a <=( A232  and  (not A201) );
 a52462a <=( a52461a  and  a52458a );
 a52463a <=( a52462a  and  a52455a );
 a52467a <=( (not A266)  and  (not A265) );
 a52468a <=( A233  and  a52467a );
 a52471a <=( (not A299)  and  A298 );
 a52474a <=( A301  and  A300 );
 a52475a <=( a52474a  and  a52471a );
 a52476a <=( a52475a  and  a52468a );
 a52480a <=( (not A167)  and  A169 );
 a52481a <=( (not A170)  and  a52480a );
 a52484a <=( (not A200)  and  (not A166) );
 a52487a <=( A232  and  (not A201) );
 a52488a <=( a52487a  and  a52484a );
 a52489a <=( a52488a  and  a52481a );
 a52493a <=( (not A266)  and  (not A265) );
 a52494a <=( A233  and  a52493a );
 a52497a <=( (not A299)  and  A298 );
 a52500a <=( A302  and  A300 );
 a52501a <=( a52500a  and  a52497a );
 a52502a <=( a52501a  and  a52494a );
 a52506a <=( (not A167)  and  A169 );
 a52507a <=( (not A170)  and  a52506a );
 a52510a <=( (not A200)  and  (not A166) );
 a52513a <=( (not A233)  and  (not A201) );
 a52514a <=( a52513a  and  a52510a );
 a52515a <=( a52514a  and  a52507a );
 a52519a <=( (not A266)  and  (not A236) );
 a52520a <=( (not A235)  and  a52519a );
 a52523a <=( (not A269)  and  (not A268) );
 a52526a <=( A299  and  (not A298) );
 a52527a <=( a52526a  and  a52523a );
 a52528a <=( a52527a  and  a52520a );
 a52532a <=( (not A167)  and  A169 );
 a52533a <=( (not A170)  and  a52532a );
 a52536a <=( (not A200)  and  (not A166) );
 a52539a <=( (not A233)  and  (not A201) );
 a52540a <=( a52539a  and  a52536a );
 a52541a <=( a52540a  and  a52533a );
 a52545a <=( A266  and  A265 );
 a52546a <=( (not A234)  and  a52545a );
 a52549a <=( (not A299)  and  A298 );
 a52552a <=( A301  and  A300 );
 a52553a <=( a52552a  and  a52549a );
 a52554a <=( a52553a  and  a52546a );
 a52558a <=( (not A167)  and  A169 );
 a52559a <=( (not A170)  and  a52558a );
 a52562a <=( (not A200)  and  (not A166) );
 a52565a <=( (not A233)  and  (not A201) );
 a52566a <=( a52565a  and  a52562a );
 a52567a <=( a52566a  and  a52559a );
 a52571a <=( A266  and  A265 );
 a52572a <=( (not A234)  and  a52571a );
 a52575a <=( (not A299)  and  A298 );
 a52578a <=( A302  and  A300 );
 a52579a <=( a52578a  and  a52575a );
 a52580a <=( a52579a  and  a52572a );
 a52584a <=( (not A167)  and  A169 );
 a52585a <=( (not A170)  and  a52584a );
 a52588a <=( (not A200)  and  (not A166) );
 a52591a <=( (not A233)  and  (not A201) );
 a52592a <=( a52591a  and  a52588a );
 a52593a <=( a52592a  and  a52585a );
 a52597a <=( (not A267)  and  (not A266) );
 a52598a <=( (not A234)  and  a52597a );
 a52601a <=( (not A299)  and  A298 );
 a52604a <=( A301  and  A300 );
 a52605a <=( a52604a  and  a52601a );
 a52606a <=( a52605a  and  a52598a );
 a52610a <=( (not A167)  and  A169 );
 a52611a <=( (not A170)  and  a52610a );
 a52614a <=( (not A200)  and  (not A166) );
 a52617a <=( (not A233)  and  (not A201) );
 a52618a <=( a52617a  and  a52614a );
 a52619a <=( a52618a  and  a52611a );
 a52623a <=( (not A267)  and  (not A266) );
 a52624a <=( (not A234)  and  a52623a );
 a52627a <=( (not A299)  and  A298 );
 a52630a <=( A302  and  A300 );
 a52631a <=( a52630a  and  a52627a );
 a52632a <=( a52631a  and  a52624a );
 a52636a <=( (not A167)  and  A169 );
 a52637a <=( (not A170)  and  a52636a );
 a52640a <=( (not A200)  and  (not A166) );
 a52643a <=( (not A233)  and  (not A201) );
 a52644a <=( a52643a  and  a52640a );
 a52645a <=( a52644a  and  a52637a );
 a52649a <=( (not A266)  and  (not A265) );
 a52650a <=( (not A234)  and  a52649a );
 a52653a <=( (not A299)  and  A298 );
 a52656a <=( A301  and  A300 );
 a52657a <=( a52656a  and  a52653a );
 a52658a <=( a52657a  and  a52650a );
 a52662a <=( (not A167)  and  A169 );
 a52663a <=( (not A170)  and  a52662a );
 a52666a <=( (not A200)  and  (not A166) );
 a52669a <=( (not A233)  and  (not A201) );
 a52670a <=( a52669a  and  a52666a );
 a52671a <=( a52670a  and  a52663a );
 a52675a <=( (not A266)  and  (not A265) );
 a52676a <=( (not A234)  and  a52675a );
 a52679a <=( (not A299)  and  A298 );
 a52682a <=( A302  and  A300 );
 a52683a <=( a52682a  and  a52679a );
 a52684a <=( a52683a  and  a52676a );
 a52688a <=( (not A167)  and  A169 );
 a52689a <=( (not A170)  and  a52688a );
 a52692a <=( (not A200)  and  (not A166) );
 a52695a <=( A232  and  (not A201) );
 a52696a <=( a52695a  and  a52692a );
 a52697a <=( a52696a  and  a52689a );
 a52701a <=( A235  and  A234 );
 a52702a <=( (not A233)  and  a52701a );
 a52705a <=( (not A266)  and  A265 );
 a52708a <=( A268  and  A267 );
 a52709a <=( a52708a  and  a52705a );
 a52710a <=( a52709a  and  a52702a );
 a52714a <=( (not A167)  and  A169 );
 a52715a <=( (not A170)  and  a52714a );
 a52718a <=( (not A200)  and  (not A166) );
 a52721a <=( A232  and  (not A201) );
 a52722a <=( a52721a  and  a52718a );
 a52723a <=( a52722a  and  a52715a );
 a52727a <=( A235  and  A234 );
 a52728a <=( (not A233)  and  a52727a );
 a52731a <=( (not A266)  and  A265 );
 a52734a <=( A269  and  A267 );
 a52735a <=( a52734a  and  a52731a );
 a52736a <=( a52735a  and  a52728a );
 a52740a <=( (not A167)  and  A169 );
 a52741a <=( (not A170)  and  a52740a );
 a52744a <=( (not A200)  and  (not A166) );
 a52747a <=( A232  and  (not A201) );
 a52748a <=( a52747a  and  a52744a );
 a52749a <=( a52748a  and  a52741a );
 a52753a <=( A236  and  A234 );
 a52754a <=( (not A233)  and  a52753a );
 a52757a <=( (not A266)  and  A265 );
 a52760a <=( A268  and  A267 );
 a52761a <=( a52760a  and  a52757a );
 a52762a <=( a52761a  and  a52754a );
 a52766a <=( (not A167)  and  A169 );
 a52767a <=( (not A170)  and  a52766a );
 a52770a <=( (not A200)  and  (not A166) );
 a52773a <=( A232  and  (not A201) );
 a52774a <=( a52773a  and  a52770a );
 a52775a <=( a52774a  and  a52767a );
 a52779a <=( A236  and  A234 );
 a52780a <=( (not A233)  and  a52779a );
 a52783a <=( (not A266)  and  A265 );
 a52786a <=( A269  and  A267 );
 a52787a <=( a52786a  and  a52783a );
 a52788a <=( a52787a  and  a52780a );
 a52792a <=( (not A167)  and  A169 );
 a52793a <=( (not A170)  and  a52792a );
 a52796a <=( (not A200)  and  (not A166) );
 a52799a <=( (not A232)  and  (not A201) );
 a52800a <=( a52799a  and  a52796a );
 a52801a <=( a52800a  and  a52793a );
 a52805a <=( A266  and  A265 );
 a52806a <=( (not A233)  and  a52805a );
 a52809a <=( (not A299)  and  A298 );
 a52812a <=( A301  and  A300 );
 a52813a <=( a52812a  and  a52809a );
 a52814a <=( a52813a  and  a52806a );
 a52818a <=( (not A167)  and  A169 );
 a52819a <=( (not A170)  and  a52818a );
 a52822a <=( (not A200)  and  (not A166) );
 a52825a <=( (not A232)  and  (not A201) );
 a52826a <=( a52825a  and  a52822a );
 a52827a <=( a52826a  and  a52819a );
 a52831a <=( A266  and  A265 );
 a52832a <=( (not A233)  and  a52831a );
 a52835a <=( (not A299)  and  A298 );
 a52838a <=( A302  and  A300 );
 a52839a <=( a52838a  and  a52835a );
 a52840a <=( a52839a  and  a52832a );
 a52844a <=( (not A167)  and  A169 );
 a52845a <=( (not A170)  and  a52844a );
 a52848a <=( (not A200)  and  (not A166) );
 a52851a <=( (not A232)  and  (not A201) );
 a52852a <=( a52851a  and  a52848a );
 a52853a <=( a52852a  and  a52845a );
 a52857a <=( (not A267)  and  (not A266) );
 a52858a <=( (not A233)  and  a52857a );
 a52861a <=( (not A299)  and  A298 );
 a52864a <=( A301  and  A300 );
 a52865a <=( a52864a  and  a52861a );
 a52866a <=( a52865a  and  a52858a );
 a52870a <=( (not A167)  and  A169 );
 a52871a <=( (not A170)  and  a52870a );
 a52874a <=( (not A200)  and  (not A166) );
 a52877a <=( (not A232)  and  (not A201) );
 a52878a <=( a52877a  and  a52874a );
 a52879a <=( a52878a  and  a52871a );
 a52883a <=( (not A267)  and  (not A266) );
 a52884a <=( (not A233)  and  a52883a );
 a52887a <=( (not A299)  and  A298 );
 a52890a <=( A302  and  A300 );
 a52891a <=( a52890a  and  a52887a );
 a52892a <=( a52891a  and  a52884a );
 a52896a <=( (not A167)  and  A169 );
 a52897a <=( (not A170)  and  a52896a );
 a52900a <=( (not A200)  and  (not A166) );
 a52903a <=( (not A232)  and  (not A201) );
 a52904a <=( a52903a  and  a52900a );
 a52905a <=( a52904a  and  a52897a );
 a52909a <=( (not A266)  and  (not A265) );
 a52910a <=( (not A233)  and  a52909a );
 a52913a <=( (not A299)  and  A298 );
 a52916a <=( A301  and  A300 );
 a52917a <=( a52916a  and  a52913a );
 a52918a <=( a52917a  and  a52910a );
 a52922a <=( (not A167)  and  A169 );
 a52923a <=( (not A170)  and  a52922a );
 a52926a <=( (not A200)  and  (not A166) );
 a52929a <=( (not A232)  and  (not A201) );
 a52930a <=( a52929a  and  a52926a );
 a52931a <=( a52930a  and  a52923a );
 a52935a <=( (not A266)  and  (not A265) );
 a52936a <=( (not A233)  and  a52935a );
 a52939a <=( (not A299)  and  A298 );
 a52942a <=( A302  and  A300 );
 a52943a <=( a52942a  and  a52939a );
 a52944a <=( a52943a  and  a52936a );
 a52948a <=( (not A167)  and  A169 );
 a52949a <=( (not A170)  and  a52948a );
 a52952a <=( (not A199)  and  (not A166) );
 a52955a <=( A232  and  (not A200) );
 a52956a <=( a52955a  and  a52952a );
 a52957a <=( a52956a  and  a52949a );
 a52961a <=( (not A267)  and  A265 );
 a52962a <=( A233  and  a52961a );
 a52965a <=( (not A299)  and  A298 );
 a52968a <=( A301  and  A300 );
 a52969a <=( a52968a  and  a52965a );
 a52970a <=( a52969a  and  a52962a );
 a52974a <=( (not A167)  and  A169 );
 a52975a <=( (not A170)  and  a52974a );
 a52978a <=( (not A199)  and  (not A166) );
 a52981a <=( A232  and  (not A200) );
 a52982a <=( a52981a  and  a52978a );
 a52983a <=( a52982a  and  a52975a );
 a52987a <=( (not A267)  and  A265 );
 a52988a <=( A233  and  a52987a );
 a52991a <=( (not A299)  and  A298 );
 a52994a <=( A302  and  A300 );
 a52995a <=( a52994a  and  a52991a );
 a52996a <=( a52995a  and  a52988a );
 a53000a <=( (not A167)  and  A169 );
 a53001a <=( (not A170)  and  a53000a );
 a53004a <=( (not A199)  and  (not A166) );
 a53007a <=( A232  and  (not A200) );
 a53008a <=( a53007a  and  a53004a );
 a53009a <=( a53008a  and  a53001a );
 a53013a <=( A266  and  A265 );
 a53014a <=( A233  and  a53013a );
 a53017a <=( (not A299)  and  A298 );
 a53020a <=( A301  and  A300 );
 a53021a <=( a53020a  and  a53017a );
 a53022a <=( a53021a  and  a53014a );
 a53026a <=( (not A167)  and  A169 );
 a53027a <=( (not A170)  and  a53026a );
 a53030a <=( (not A199)  and  (not A166) );
 a53033a <=( A232  and  (not A200) );
 a53034a <=( a53033a  and  a53030a );
 a53035a <=( a53034a  and  a53027a );
 a53039a <=( A266  and  A265 );
 a53040a <=( A233  and  a53039a );
 a53043a <=( (not A299)  and  A298 );
 a53046a <=( A302  and  A300 );
 a53047a <=( a53046a  and  a53043a );
 a53048a <=( a53047a  and  a53040a );
 a53052a <=( (not A167)  and  A169 );
 a53053a <=( (not A170)  and  a53052a );
 a53056a <=( (not A199)  and  (not A166) );
 a53059a <=( A232  and  (not A200) );
 a53060a <=( a53059a  and  a53056a );
 a53061a <=( a53060a  and  a53053a );
 a53065a <=( (not A266)  and  (not A265) );
 a53066a <=( A233  and  a53065a );
 a53069a <=( (not A299)  and  A298 );
 a53072a <=( A301  and  A300 );
 a53073a <=( a53072a  and  a53069a );
 a53074a <=( a53073a  and  a53066a );
 a53078a <=( (not A167)  and  A169 );
 a53079a <=( (not A170)  and  a53078a );
 a53082a <=( (not A199)  and  (not A166) );
 a53085a <=( A232  and  (not A200) );
 a53086a <=( a53085a  and  a53082a );
 a53087a <=( a53086a  and  a53079a );
 a53091a <=( (not A266)  and  (not A265) );
 a53092a <=( A233  and  a53091a );
 a53095a <=( (not A299)  and  A298 );
 a53098a <=( A302  and  A300 );
 a53099a <=( a53098a  and  a53095a );
 a53100a <=( a53099a  and  a53092a );
 a53104a <=( (not A167)  and  A169 );
 a53105a <=( (not A170)  and  a53104a );
 a53108a <=( (not A199)  and  (not A166) );
 a53111a <=( (not A233)  and  (not A200) );
 a53112a <=( a53111a  and  a53108a );
 a53113a <=( a53112a  and  a53105a );
 a53117a <=( (not A266)  and  (not A236) );
 a53118a <=( (not A235)  and  a53117a );
 a53121a <=( (not A269)  and  (not A268) );
 a53124a <=( A299  and  (not A298) );
 a53125a <=( a53124a  and  a53121a );
 a53126a <=( a53125a  and  a53118a );
 a53130a <=( (not A167)  and  A169 );
 a53131a <=( (not A170)  and  a53130a );
 a53134a <=( (not A199)  and  (not A166) );
 a53137a <=( (not A233)  and  (not A200) );
 a53138a <=( a53137a  and  a53134a );
 a53139a <=( a53138a  and  a53131a );
 a53143a <=( A266  and  A265 );
 a53144a <=( (not A234)  and  a53143a );
 a53147a <=( (not A299)  and  A298 );
 a53150a <=( A301  and  A300 );
 a53151a <=( a53150a  and  a53147a );
 a53152a <=( a53151a  and  a53144a );
 a53156a <=( (not A167)  and  A169 );
 a53157a <=( (not A170)  and  a53156a );
 a53160a <=( (not A199)  and  (not A166) );
 a53163a <=( (not A233)  and  (not A200) );
 a53164a <=( a53163a  and  a53160a );
 a53165a <=( a53164a  and  a53157a );
 a53169a <=( A266  and  A265 );
 a53170a <=( (not A234)  and  a53169a );
 a53173a <=( (not A299)  and  A298 );
 a53176a <=( A302  and  A300 );
 a53177a <=( a53176a  and  a53173a );
 a53178a <=( a53177a  and  a53170a );
 a53182a <=( (not A167)  and  A169 );
 a53183a <=( (not A170)  and  a53182a );
 a53186a <=( (not A199)  and  (not A166) );
 a53189a <=( (not A233)  and  (not A200) );
 a53190a <=( a53189a  and  a53186a );
 a53191a <=( a53190a  and  a53183a );
 a53195a <=( (not A267)  and  (not A266) );
 a53196a <=( (not A234)  and  a53195a );
 a53199a <=( (not A299)  and  A298 );
 a53202a <=( A301  and  A300 );
 a53203a <=( a53202a  and  a53199a );
 a53204a <=( a53203a  and  a53196a );
 a53208a <=( (not A167)  and  A169 );
 a53209a <=( (not A170)  and  a53208a );
 a53212a <=( (not A199)  and  (not A166) );
 a53215a <=( (not A233)  and  (not A200) );
 a53216a <=( a53215a  and  a53212a );
 a53217a <=( a53216a  and  a53209a );
 a53221a <=( (not A267)  and  (not A266) );
 a53222a <=( (not A234)  and  a53221a );
 a53225a <=( (not A299)  and  A298 );
 a53228a <=( A302  and  A300 );
 a53229a <=( a53228a  and  a53225a );
 a53230a <=( a53229a  and  a53222a );
 a53234a <=( (not A167)  and  A169 );
 a53235a <=( (not A170)  and  a53234a );
 a53238a <=( (not A199)  and  (not A166) );
 a53241a <=( (not A233)  and  (not A200) );
 a53242a <=( a53241a  and  a53238a );
 a53243a <=( a53242a  and  a53235a );
 a53247a <=( (not A266)  and  (not A265) );
 a53248a <=( (not A234)  and  a53247a );
 a53251a <=( (not A299)  and  A298 );
 a53254a <=( A301  and  A300 );
 a53255a <=( a53254a  and  a53251a );
 a53256a <=( a53255a  and  a53248a );
 a53260a <=( (not A167)  and  A169 );
 a53261a <=( (not A170)  and  a53260a );
 a53264a <=( (not A199)  and  (not A166) );
 a53267a <=( (not A233)  and  (not A200) );
 a53268a <=( a53267a  and  a53264a );
 a53269a <=( a53268a  and  a53261a );
 a53273a <=( (not A266)  and  (not A265) );
 a53274a <=( (not A234)  and  a53273a );
 a53277a <=( (not A299)  and  A298 );
 a53280a <=( A302  and  A300 );
 a53281a <=( a53280a  and  a53277a );
 a53282a <=( a53281a  and  a53274a );
 a53286a <=( (not A167)  and  A169 );
 a53287a <=( (not A170)  and  a53286a );
 a53290a <=( (not A199)  and  (not A166) );
 a53293a <=( A232  and  (not A200) );
 a53294a <=( a53293a  and  a53290a );
 a53295a <=( a53294a  and  a53287a );
 a53299a <=( A235  and  A234 );
 a53300a <=( (not A233)  and  a53299a );
 a53303a <=( (not A266)  and  A265 );
 a53306a <=( A268  and  A267 );
 a53307a <=( a53306a  and  a53303a );
 a53308a <=( a53307a  and  a53300a );
 a53312a <=( (not A167)  and  A169 );
 a53313a <=( (not A170)  and  a53312a );
 a53316a <=( (not A199)  and  (not A166) );
 a53319a <=( A232  and  (not A200) );
 a53320a <=( a53319a  and  a53316a );
 a53321a <=( a53320a  and  a53313a );
 a53325a <=( A235  and  A234 );
 a53326a <=( (not A233)  and  a53325a );
 a53329a <=( (not A266)  and  A265 );
 a53332a <=( A269  and  A267 );
 a53333a <=( a53332a  and  a53329a );
 a53334a <=( a53333a  and  a53326a );
 a53338a <=( (not A167)  and  A169 );
 a53339a <=( (not A170)  and  a53338a );
 a53342a <=( (not A199)  and  (not A166) );
 a53345a <=( A232  and  (not A200) );
 a53346a <=( a53345a  and  a53342a );
 a53347a <=( a53346a  and  a53339a );
 a53351a <=( A236  and  A234 );
 a53352a <=( (not A233)  and  a53351a );
 a53355a <=( (not A266)  and  A265 );
 a53358a <=( A268  and  A267 );
 a53359a <=( a53358a  and  a53355a );
 a53360a <=( a53359a  and  a53352a );
 a53364a <=( (not A167)  and  A169 );
 a53365a <=( (not A170)  and  a53364a );
 a53368a <=( (not A199)  and  (not A166) );
 a53371a <=( A232  and  (not A200) );
 a53372a <=( a53371a  and  a53368a );
 a53373a <=( a53372a  and  a53365a );
 a53377a <=( A236  and  A234 );
 a53378a <=( (not A233)  and  a53377a );
 a53381a <=( (not A266)  and  A265 );
 a53384a <=( A269  and  A267 );
 a53385a <=( a53384a  and  a53381a );
 a53386a <=( a53385a  and  a53378a );
 a53390a <=( (not A167)  and  A169 );
 a53391a <=( (not A170)  and  a53390a );
 a53394a <=( (not A199)  and  (not A166) );
 a53397a <=( (not A232)  and  (not A200) );
 a53398a <=( a53397a  and  a53394a );
 a53399a <=( a53398a  and  a53391a );
 a53403a <=( A266  and  A265 );
 a53404a <=( (not A233)  and  a53403a );
 a53407a <=( (not A299)  and  A298 );
 a53410a <=( A301  and  A300 );
 a53411a <=( a53410a  and  a53407a );
 a53412a <=( a53411a  and  a53404a );
 a53416a <=( (not A167)  and  A169 );
 a53417a <=( (not A170)  and  a53416a );
 a53420a <=( (not A199)  and  (not A166) );
 a53423a <=( (not A232)  and  (not A200) );
 a53424a <=( a53423a  and  a53420a );
 a53425a <=( a53424a  and  a53417a );
 a53429a <=( A266  and  A265 );
 a53430a <=( (not A233)  and  a53429a );
 a53433a <=( (not A299)  and  A298 );
 a53436a <=( A302  and  A300 );
 a53437a <=( a53436a  and  a53433a );
 a53438a <=( a53437a  and  a53430a );
 a53442a <=( (not A167)  and  A169 );
 a53443a <=( (not A170)  and  a53442a );
 a53446a <=( (not A199)  and  (not A166) );
 a53449a <=( (not A232)  and  (not A200) );
 a53450a <=( a53449a  and  a53446a );
 a53451a <=( a53450a  and  a53443a );
 a53455a <=( (not A267)  and  (not A266) );
 a53456a <=( (not A233)  and  a53455a );
 a53459a <=( (not A299)  and  A298 );
 a53462a <=( A301  and  A300 );
 a53463a <=( a53462a  and  a53459a );
 a53464a <=( a53463a  and  a53456a );
 a53468a <=( (not A167)  and  A169 );
 a53469a <=( (not A170)  and  a53468a );
 a53472a <=( (not A199)  and  (not A166) );
 a53475a <=( (not A232)  and  (not A200) );
 a53476a <=( a53475a  and  a53472a );
 a53477a <=( a53476a  and  a53469a );
 a53481a <=( (not A267)  and  (not A266) );
 a53482a <=( (not A233)  and  a53481a );
 a53485a <=( (not A299)  and  A298 );
 a53488a <=( A302  and  A300 );
 a53489a <=( a53488a  and  a53485a );
 a53490a <=( a53489a  and  a53482a );
 a53494a <=( (not A167)  and  A169 );
 a53495a <=( (not A170)  and  a53494a );
 a53498a <=( (not A199)  and  (not A166) );
 a53501a <=( (not A232)  and  (not A200) );
 a53502a <=( a53501a  and  a53498a );
 a53503a <=( a53502a  and  a53495a );
 a53507a <=( (not A266)  and  (not A265) );
 a53508a <=( (not A233)  and  a53507a );
 a53511a <=( (not A299)  and  A298 );
 a53514a <=( A301  and  A300 );
 a53515a <=( a53514a  and  a53511a );
 a53516a <=( a53515a  and  a53508a );
 a53520a <=( (not A167)  and  A169 );
 a53521a <=( (not A170)  and  a53520a );
 a53524a <=( (not A199)  and  (not A166) );
 a53527a <=( (not A232)  and  (not A200) );
 a53528a <=( a53527a  and  a53524a );
 a53529a <=( a53528a  and  a53521a );
 a53533a <=( (not A266)  and  (not A265) );
 a53534a <=( (not A233)  and  a53533a );
 a53537a <=( (not A299)  and  A298 );
 a53540a <=( A302  and  A300 );
 a53541a <=( a53540a  and  a53537a );
 a53542a <=( a53541a  and  a53534a );
 a53546a <=( (not A166)  and  (not A167) );
 a53547a <=( (not A169)  and  a53546a );
 a53550a <=( A200  and  (not A199) );
 a53553a <=( A233  and  A232 );
 a53554a <=( a53553a  and  a53550a );
 a53555a <=( a53554a  and  a53547a );
 a53559a <=( (not A269)  and  (not A268) );
 a53560a <=( A265  and  a53559a );
 a53563a <=( (not A299)  and  A298 );
 a53566a <=( A301  and  A300 );
 a53567a <=( a53566a  and  a53563a );
 a53568a <=( a53567a  and  a53560a );
 a53572a <=( (not A166)  and  (not A167) );
 a53573a <=( (not A169)  and  a53572a );
 a53576a <=( A200  and  (not A199) );
 a53579a <=( A233  and  A232 );
 a53580a <=( a53579a  and  a53576a );
 a53581a <=( a53580a  and  a53573a );
 a53585a <=( (not A269)  and  (not A268) );
 a53586a <=( A265  and  a53585a );
 a53589a <=( (not A299)  and  A298 );
 a53592a <=( A302  and  A300 );
 a53593a <=( a53592a  and  a53589a );
 a53594a <=( a53593a  and  a53586a );
 a53598a <=( (not A166)  and  (not A167) );
 a53599a <=( (not A169)  and  a53598a );
 a53602a <=( A200  and  (not A199) );
 a53605a <=( (not A235)  and  (not A233) );
 a53606a <=( a53605a  and  a53602a );
 a53607a <=( a53606a  and  a53599a );
 a53611a <=( A266  and  A265 );
 a53612a <=( (not A236)  and  a53611a );
 a53615a <=( (not A299)  and  A298 );
 a53618a <=( A301  and  A300 );
 a53619a <=( a53618a  and  a53615a );
 a53620a <=( a53619a  and  a53612a );
 a53624a <=( (not A166)  and  (not A167) );
 a53625a <=( (not A169)  and  a53624a );
 a53628a <=( A200  and  (not A199) );
 a53631a <=( (not A235)  and  (not A233) );
 a53632a <=( a53631a  and  a53628a );
 a53633a <=( a53632a  and  a53625a );
 a53637a <=( A266  and  A265 );
 a53638a <=( (not A236)  and  a53637a );
 a53641a <=( (not A299)  and  A298 );
 a53644a <=( A302  and  A300 );
 a53645a <=( a53644a  and  a53641a );
 a53646a <=( a53645a  and  a53638a );
 a53650a <=( (not A166)  and  (not A167) );
 a53651a <=( (not A169)  and  a53650a );
 a53654a <=( A200  and  (not A199) );
 a53657a <=( (not A235)  and  (not A233) );
 a53658a <=( a53657a  and  a53654a );
 a53659a <=( a53658a  and  a53651a );
 a53663a <=( (not A267)  and  (not A266) );
 a53664a <=( (not A236)  and  a53663a );
 a53667a <=( (not A299)  and  A298 );
 a53670a <=( A301  and  A300 );
 a53671a <=( a53670a  and  a53667a );
 a53672a <=( a53671a  and  a53664a );
 a53676a <=( (not A166)  and  (not A167) );
 a53677a <=( (not A169)  and  a53676a );
 a53680a <=( A200  and  (not A199) );
 a53683a <=( (not A235)  and  (not A233) );
 a53684a <=( a53683a  and  a53680a );
 a53685a <=( a53684a  and  a53677a );
 a53689a <=( (not A267)  and  (not A266) );
 a53690a <=( (not A236)  and  a53689a );
 a53693a <=( (not A299)  and  A298 );
 a53696a <=( A302  and  A300 );
 a53697a <=( a53696a  and  a53693a );
 a53698a <=( a53697a  and  a53690a );
 a53702a <=( (not A166)  and  (not A167) );
 a53703a <=( (not A169)  and  a53702a );
 a53706a <=( A200  and  (not A199) );
 a53709a <=( (not A235)  and  (not A233) );
 a53710a <=( a53709a  and  a53706a );
 a53711a <=( a53710a  and  a53703a );
 a53715a <=( (not A266)  and  (not A265) );
 a53716a <=( (not A236)  and  a53715a );
 a53719a <=( (not A299)  and  A298 );
 a53722a <=( A301  and  A300 );
 a53723a <=( a53722a  and  a53719a );
 a53724a <=( a53723a  and  a53716a );
 a53728a <=( (not A166)  and  (not A167) );
 a53729a <=( (not A169)  and  a53728a );
 a53732a <=( A200  and  (not A199) );
 a53735a <=( (not A235)  and  (not A233) );
 a53736a <=( a53735a  and  a53732a );
 a53737a <=( a53736a  and  a53729a );
 a53741a <=( (not A266)  and  (not A265) );
 a53742a <=( (not A236)  and  a53741a );
 a53745a <=( (not A299)  and  A298 );
 a53748a <=( A302  and  A300 );
 a53749a <=( a53748a  and  a53745a );
 a53750a <=( a53749a  and  a53742a );
 a53754a <=( (not A166)  and  (not A167) );
 a53755a <=( (not A169)  and  a53754a );
 a53758a <=( A200  and  (not A199) );
 a53761a <=( (not A234)  and  (not A233) );
 a53762a <=( a53761a  and  a53758a );
 a53763a <=( a53762a  and  a53755a );
 a53767a <=( (not A269)  and  (not A268) );
 a53768a <=( (not A266)  and  a53767a );
 a53771a <=( (not A299)  and  A298 );
 a53774a <=( A301  and  A300 );
 a53775a <=( a53774a  and  a53771a );
 a53776a <=( a53775a  and  a53768a );
 a53780a <=( (not A166)  and  (not A167) );
 a53781a <=( (not A169)  and  a53780a );
 a53784a <=( A200  and  (not A199) );
 a53787a <=( (not A234)  and  (not A233) );
 a53788a <=( a53787a  and  a53784a );
 a53789a <=( a53788a  and  a53781a );
 a53793a <=( (not A269)  and  (not A268) );
 a53794a <=( (not A266)  and  a53793a );
 a53797a <=( (not A299)  and  A298 );
 a53800a <=( A302  and  A300 );
 a53801a <=( a53800a  and  a53797a );
 a53802a <=( a53801a  and  a53794a );
 a53806a <=( (not A166)  and  (not A167) );
 a53807a <=( (not A169)  and  a53806a );
 a53810a <=( A200  and  (not A199) );
 a53813a <=( (not A233)  and  (not A232) );
 a53814a <=( a53813a  and  a53810a );
 a53815a <=( a53814a  and  a53807a );
 a53819a <=( (not A269)  and  (not A268) );
 a53820a <=( (not A266)  and  a53819a );
 a53823a <=( (not A299)  and  A298 );
 a53826a <=( A301  and  A300 );
 a53827a <=( a53826a  and  a53823a );
 a53828a <=( a53827a  and  a53820a );
 a53832a <=( (not A166)  and  (not A167) );
 a53833a <=( (not A169)  and  a53832a );
 a53836a <=( A200  and  (not A199) );
 a53839a <=( (not A233)  and  (not A232) );
 a53840a <=( a53839a  and  a53836a );
 a53841a <=( a53840a  and  a53833a );
 a53845a <=( (not A269)  and  (not A268) );
 a53846a <=( (not A266)  and  a53845a );
 a53849a <=( (not A299)  and  A298 );
 a53852a <=( A302  and  A300 );
 a53853a <=( a53852a  and  a53849a );
 a53854a <=( a53853a  and  a53846a );
 a53858a <=( (not A166)  and  (not A167) );
 a53859a <=( (not A169)  and  a53858a );
 a53862a <=( (not A200)  and  A199 );
 a53865a <=( A202  and  A201 );
 a53866a <=( a53865a  and  a53862a );
 a53867a <=( a53866a  and  a53859a );
 a53871a <=( A265  and  A233 );
 a53872a <=( A232  and  a53871a );
 a53875a <=( (not A269)  and  (not A268) );
 a53878a <=( A299  and  (not A298) );
 a53879a <=( a53878a  and  a53875a );
 a53880a <=( a53879a  and  a53872a );
 a53884a <=( (not A166)  and  (not A167) );
 a53885a <=( (not A169)  and  a53884a );
 a53888a <=( (not A200)  and  A199 );
 a53891a <=( A202  and  A201 );
 a53892a <=( a53891a  and  a53888a );
 a53893a <=( a53892a  and  a53885a );
 a53897a <=( (not A236)  and  (not A235) );
 a53898a <=( (not A233)  and  a53897a );
 a53901a <=( A266  and  A265 );
 a53904a <=( A299  and  (not A298) );
 a53905a <=( a53904a  and  a53901a );
 a53906a <=( a53905a  and  a53898a );
 a53910a <=( (not A166)  and  (not A167) );
 a53911a <=( (not A169)  and  a53910a );
 a53914a <=( (not A200)  and  A199 );
 a53917a <=( A202  and  A201 );
 a53918a <=( a53917a  and  a53914a );
 a53919a <=( a53918a  and  a53911a );
 a53923a <=( (not A236)  and  (not A235) );
 a53924a <=( (not A233)  and  a53923a );
 a53927a <=( (not A267)  and  (not A266) );
 a53930a <=( A299  and  (not A298) );
 a53931a <=( a53930a  and  a53927a );
 a53932a <=( a53931a  and  a53924a );
 a53936a <=( (not A166)  and  (not A167) );
 a53937a <=( (not A169)  and  a53936a );
 a53940a <=( (not A200)  and  A199 );
 a53943a <=( A202  and  A201 );
 a53944a <=( a53943a  and  a53940a );
 a53945a <=( a53944a  and  a53937a );
 a53949a <=( (not A236)  and  (not A235) );
 a53950a <=( (not A233)  and  a53949a );
 a53953a <=( (not A266)  and  (not A265) );
 a53956a <=( A299  and  (not A298) );
 a53957a <=( a53956a  and  a53953a );
 a53958a <=( a53957a  and  a53950a );
 a53962a <=( (not A166)  and  (not A167) );
 a53963a <=( (not A169)  and  a53962a );
 a53966a <=( (not A200)  and  A199 );
 a53969a <=( A202  and  A201 );
 a53970a <=( a53969a  and  a53966a );
 a53971a <=( a53970a  and  a53963a );
 a53975a <=( (not A266)  and  (not A234) );
 a53976a <=( (not A233)  and  a53975a );
 a53979a <=( (not A269)  and  (not A268) );
 a53982a <=( A299  and  (not A298) );
 a53983a <=( a53982a  and  a53979a );
 a53984a <=( a53983a  and  a53976a );
 a53988a <=( (not A166)  and  (not A167) );
 a53989a <=( (not A169)  and  a53988a );
 a53992a <=( (not A200)  and  A199 );
 a53995a <=( A202  and  A201 );
 a53996a <=( a53995a  and  a53992a );
 a53997a <=( a53996a  and  a53989a );
 a54001a <=( A234  and  (not A233) );
 a54002a <=( A232  and  a54001a );
 a54005a <=( A298  and  A235 );
 a54008a <=( (not A302)  and  (not A301) );
 a54009a <=( a54008a  and  a54005a );
 a54010a <=( a54009a  and  a54002a );
 a54014a <=( (not A166)  and  (not A167) );
 a54015a <=( (not A169)  and  a54014a );
 a54018a <=( (not A200)  and  A199 );
 a54021a <=( A202  and  A201 );
 a54022a <=( a54021a  and  a54018a );
 a54023a <=( a54022a  and  a54015a );
 a54027a <=( A234  and  (not A233) );
 a54028a <=( A232  and  a54027a );
 a54031a <=( A298  and  A236 );
 a54034a <=( (not A302)  and  (not A301) );
 a54035a <=( a54034a  and  a54031a );
 a54036a <=( a54035a  and  a54028a );
 a54040a <=( (not A166)  and  (not A167) );
 a54041a <=( (not A169)  and  a54040a );
 a54044a <=( (not A200)  and  A199 );
 a54047a <=( A202  and  A201 );
 a54048a <=( a54047a  and  a54044a );
 a54049a <=( a54048a  and  a54041a );
 a54053a <=( (not A266)  and  (not A233) );
 a54054a <=( (not A232)  and  a54053a );
 a54057a <=( (not A269)  and  (not A268) );
 a54060a <=( A299  and  (not A298) );
 a54061a <=( a54060a  and  a54057a );
 a54062a <=( a54061a  and  a54054a );
 a54066a <=( (not A166)  and  (not A167) );
 a54067a <=( (not A169)  and  a54066a );
 a54070a <=( (not A200)  and  A199 );
 a54073a <=( A203  and  A201 );
 a54074a <=( a54073a  and  a54070a );
 a54075a <=( a54074a  and  a54067a );
 a54079a <=( A265  and  A233 );
 a54080a <=( A232  and  a54079a );
 a54083a <=( (not A269)  and  (not A268) );
 a54086a <=( A299  and  (not A298) );
 a54087a <=( a54086a  and  a54083a );
 a54088a <=( a54087a  and  a54080a );
 a54092a <=( (not A166)  and  (not A167) );
 a54093a <=( (not A169)  and  a54092a );
 a54096a <=( (not A200)  and  A199 );
 a54099a <=( A203  and  A201 );
 a54100a <=( a54099a  and  a54096a );
 a54101a <=( a54100a  and  a54093a );
 a54105a <=( (not A236)  and  (not A235) );
 a54106a <=( (not A233)  and  a54105a );
 a54109a <=( A266  and  A265 );
 a54112a <=( A299  and  (not A298) );
 a54113a <=( a54112a  and  a54109a );
 a54114a <=( a54113a  and  a54106a );
 a54118a <=( (not A166)  and  (not A167) );
 a54119a <=( (not A169)  and  a54118a );
 a54122a <=( (not A200)  and  A199 );
 a54125a <=( A203  and  A201 );
 a54126a <=( a54125a  and  a54122a );
 a54127a <=( a54126a  and  a54119a );
 a54131a <=( (not A236)  and  (not A235) );
 a54132a <=( (not A233)  and  a54131a );
 a54135a <=( (not A267)  and  (not A266) );
 a54138a <=( A299  and  (not A298) );
 a54139a <=( a54138a  and  a54135a );
 a54140a <=( a54139a  and  a54132a );
 a54144a <=( (not A166)  and  (not A167) );
 a54145a <=( (not A169)  and  a54144a );
 a54148a <=( (not A200)  and  A199 );
 a54151a <=( A203  and  A201 );
 a54152a <=( a54151a  and  a54148a );
 a54153a <=( a54152a  and  a54145a );
 a54157a <=( (not A236)  and  (not A235) );
 a54158a <=( (not A233)  and  a54157a );
 a54161a <=( (not A266)  and  (not A265) );
 a54164a <=( A299  and  (not A298) );
 a54165a <=( a54164a  and  a54161a );
 a54166a <=( a54165a  and  a54158a );
 a54170a <=( (not A166)  and  (not A167) );
 a54171a <=( (not A169)  and  a54170a );
 a54174a <=( (not A200)  and  A199 );
 a54177a <=( A203  and  A201 );
 a54178a <=( a54177a  and  a54174a );
 a54179a <=( a54178a  and  a54171a );
 a54183a <=( (not A266)  and  (not A234) );
 a54184a <=( (not A233)  and  a54183a );
 a54187a <=( (not A269)  and  (not A268) );
 a54190a <=( A299  and  (not A298) );
 a54191a <=( a54190a  and  a54187a );
 a54192a <=( a54191a  and  a54184a );
 a54196a <=( (not A166)  and  (not A167) );
 a54197a <=( (not A169)  and  a54196a );
 a54200a <=( (not A200)  and  A199 );
 a54203a <=( A203  and  A201 );
 a54204a <=( a54203a  and  a54200a );
 a54205a <=( a54204a  and  a54197a );
 a54209a <=( A234  and  (not A233) );
 a54210a <=( A232  and  a54209a );
 a54213a <=( A298  and  A235 );
 a54216a <=( (not A302)  and  (not A301) );
 a54217a <=( a54216a  and  a54213a );
 a54218a <=( a54217a  and  a54210a );
 a54222a <=( (not A166)  and  (not A167) );
 a54223a <=( (not A169)  and  a54222a );
 a54226a <=( (not A200)  and  A199 );
 a54229a <=( A203  and  A201 );
 a54230a <=( a54229a  and  a54226a );
 a54231a <=( a54230a  and  a54223a );
 a54235a <=( A234  and  (not A233) );
 a54236a <=( A232  and  a54235a );
 a54239a <=( A298  and  A236 );
 a54242a <=( (not A302)  and  (not A301) );
 a54243a <=( a54242a  and  a54239a );
 a54244a <=( a54243a  and  a54236a );
 a54248a <=( (not A166)  and  (not A167) );
 a54249a <=( (not A169)  and  a54248a );
 a54252a <=( (not A200)  and  A199 );
 a54255a <=( A203  and  A201 );
 a54256a <=( a54255a  and  a54252a );
 a54257a <=( a54256a  and  a54249a );
 a54261a <=( (not A266)  and  (not A233) );
 a54262a <=( (not A232)  and  a54261a );
 a54265a <=( (not A269)  and  (not A268) );
 a54268a <=( A299  and  (not A298) );
 a54269a <=( a54268a  and  a54265a );
 a54270a <=( a54269a  and  a54262a );
 a54274a <=( A167  and  (not A168) );
 a54275a <=( (not A169)  and  a54274a );
 a54278a <=( (not A199)  and  A166 );
 a54281a <=( A232  and  A200 );
 a54282a <=( a54281a  and  a54278a );
 a54283a <=( a54282a  and  a54275a );
 a54287a <=( (not A267)  and  A265 );
 a54288a <=( A233  and  a54287a );
 a54291a <=( (not A299)  and  A298 );
 a54294a <=( A301  and  A300 );
 a54295a <=( a54294a  and  a54291a );
 a54296a <=( a54295a  and  a54288a );
 a54300a <=( A167  and  (not A168) );
 a54301a <=( (not A169)  and  a54300a );
 a54304a <=( (not A199)  and  A166 );
 a54307a <=( A232  and  A200 );
 a54308a <=( a54307a  and  a54304a );
 a54309a <=( a54308a  and  a54301a );
 a54313a <=( (not A267)  and  A265 );
 a54314a <=( A233  and  a54313a );
 a54317a <=( (not A299)  and  A298 );
 a54320a <=( A302  and  A300 );
 a54321a <=( a54320a  and  a54317a );
 a54322a <=( a54321a  and  a54314a );
 a54326a <=( A167  and  (not A168) );
 a54327a <=( (not A169)  and  a54326a );
 a54330a <=( (not A199)  and  A166 );
 a54333a <=( A232  and  A200 );
 a54334a <=( a54333a  and  a54330a );
 a54335a <=( a54334a  and  a54327a );
 a54339a <=( A266  and  A265 );
 a54340a <=( A233  and  a54339a );
 a54343a <=( (not A299)  and  A298 );
 a54346a <=( A301  and  A300 );
 a54347a <=( a54346a  and  a54343a );
 a54348a <=( a54347a  and  a54340a );
 a54352a <=( A167  and  (not A168) );
 a54353a <=( (not A169)  and  a54352a );
 a54356a <=( (not A199)  and  A166 );
 a54359a <=( A232  and  A200 );
 a54360a <=( a54359a  and  a54356a );
 a54361a <=( a54360a  and  a54353a );
 a54365a <=( A266  and  A265 );
 a54366a <=( A233  and  a54365a );
 a54369a <=( (not A299)  and  A298 );
 a54372a <=( A302  and  A300 );
 a54373a <=( a54372a  and  a54369a );
 a54374a <=( a54373a  and  a54366a );
 a54378a <=( A167  and  (not A168) );
 a54379a <=( (not A169)  and  a54378a );
 a54382a <=( (not A199)  and  A166 );
 a54385a <=( A232  and  A200 );
 a54386a <=( a54385a  and  a54382a );
 a54387a <=( a54386a  and  a54379a );
 a54391a <=( (not A266)  and  (not A265) );
 a54392a <=( A233  and  a54391a );
 a54395a <=( (not A299)  and  A298 );
 a54398a <=( A301  and  A300 );
 a54399a <=( a54398a  and  a54395a );
 a54400a <=( a54399a  and  a54392a );
 a54404a <=( A167  and  (not A168) );
 a54405a <=( (not A169)  and  a54404a );
 a54408a <=( (not A199)  and  A166 );
 a54411a <=( A232  and  A200 );
 a54412a <=( a54411a  and  a54408a );
 a54413a <=( a54412a  and  a54405a );
 a54417a <=( (not A266)  and  (not A265) );
 a54418a <=( A233  and  a54417a );
 a54421a <=( (not A299)  and  A298 );
 a54424a <=( A302  and  A300 );
 a54425a <=( a54424a  and  a54421a );
 a54426a <=( a54425a  and  a54418a );
 a54430a <=( A167  and  (not A168) );
 a54431a <=( (not A169)  and  a54430a );
 a54434a <=( (not A199)  and  A166 );
 a54437a <=( (not A233)  and  A200 );
 a54438a <=( a54437a  and  a54434a );
 a54439a <=( a54438a  and  a54431a );
 a54443a <=( (not A266)  and  (not A236) );
 a54444a <=( (not A235)  and  a54443a );
 a54447a <=( (not A269)  and  (not A268) );
 a54450a <=( A299  and  (not A298) );
 a54451a <=( a54450a  and  a54447a );
 a54452a <=( a54451a  and  a54444a );
 a54456a <=( A167  and  (not A168) );
 a54457a <=( (not A169)  and  a54456a );
 a54460a <=( (not A199)  and  A166 );
 a54463a <=( (not A233)  and  A200 );
 a54464a <=( a54463a  and  a54460a );
 a54465a <=( a54464a  and  a54457a );
 a54469a <=( A266  and  A265 );
 a54470a <=( (not A234)  and  a54469a );
 a54473a <=( (not A299)  and  A298 );
 a54476a <=( A301  and  A300 );
 a54477a <=( a54476a  and  a54473a );
 a54478a <=( a54477a  and  a54470a );
 a54482a <=( A167  and  (not A168) );
 a54483a <=( (not A169)  and  a54482a );
 a54486a <=( (not A199)  and  A166 );
 a54489a <=( (not A233)  and  A200 );
 a54490a <=( a54489a  and  a54486a );
 a54491a <=( a54490a  and  a54483a );
 a54495a <=( A266  and  A265 );
 a54496a <=( (not A234)  and  a54495a );
 a54499a <=( (not A299)  and  A298 );
 a54502a <=( A302  and  A300 );
 a54503a <=( a54502a  and  a54499a );
 a54504a <=( a54503a  and  a54496a );
 a54508a <=( A167  and  (not A168) );
 a54509a <=( (not A169)  and  a54508a );
 a54512a <=( (not A199)  and  A166 );
 a54515a <=( (not A233)  and  A200 );
 a54516a <=( a54515a  and  a54512a );
 a54517a <=( a54516a  and  a54509a );
 a54521a <=( (not A267)  and  (not A266) );
 a54522a <=( (not A234)  and  a54521a );
 a54525a <=( (not A299)  and  A298 );
 a54528a <=( A301  and  A300 );
 a54529a <=( a54528a  and  a54525a );
 a54530a <=( a54529a  and  a54522a );
 a54534a <=( A167  and  (not A168) );
 a54535a <=( (not A169)  and  a54534a );
 a54538a <=( (not A199)  and  A166 );
 a54541a <=( (not A233)  and  A200 );
 a54542a <=( a54541a  and  a54538a );
 a54543a <=( a54542a  and  a54535a );
 a54547a <=( (not A267)  and  (not A266) );
 a54548a <=( (not A234)  and  a54547a );
 a54551a <=( (not A299)  and  A298 );
 a54554a <=( A302  and  A300 );
 a54555a <=( a54554a  and  a54551a );
 a54556a <=( a54555a  and  a54548a );
 a54560a <=( A167  and  (not A168) );
 a54561a <=( (not A169)  and  a54560a );
 a54564a <=( (not A199)  and  A166 );
 a54567a <=( (not A233)  and  A200 );
 a54568a <=( a54567a  and  a54564a );
 a54569a <=( a54568a  and  a54561a );
 a54573a <=( (not A266)  and  (not A265) );
 a54574a <=( (not A234)  and  a54573a );
 a54577a <=( (not A299)  and  A298 );
 a54580a <=( A301  and  A300 );
 a54581a <=( a54580a  and  a54577a );
 a54582a <=( a54581a  and  a54574a );
 a54586a <=( A167  and  (not A168) );
 a54587a <=( (not A169)  and  a54586a );
 a54590a <=( (not A199)  and  A166 );
 a54593a <=( (not A233)  and  A200 );
 a54594a <=( a54593a  and  a54590a );
 a54595a <=( a54594a  and  a54587a );
 a54599a <=( (not A266)  and  (not A265) );
 a54600a <=( (not A234)  and  a54599a );
 a54603a <=( (not A299)  and  A298 );
 a54606a <=( A302  and  A300 );
 a54607a <=( a54606a  and  a54603a );
 a54608a <=( a54607a  and  a54600a );
 a54612a <=( A167  and  (not A168) );
 a54613a <=( (not A169)  and  a54612a );
 a54616a <=( (not A199)  and  A166 );
 a54619a <=( A232  and  A200 );
 a54620a <=( a54619a  and  a54616a );
 a54621a <=( a54620a  and  a54613a );
 a54625a <=( A235  and  A234 );
 a54626a <=( (not A233)  and  a54625a );
 a54629a <=( (not A266)  and  A265 );
 a54632a <=( A268  and  A267 );
 a54633a <=( a54632a  and  a54629a );
 a54634a <=( a54633a  and  a54626a );
 a54638a <=( A167  and  (not A168) );
 a54639a <=( (not A169)  and  a54638a );
 a54642a <=( (not A199)  and  A166 );
 a54645a <=( A232  and  A200 );
 a54646a <=( a54645a  and  a54642a );
 a54647a <=( a54646a  and  a54639a );
 a54651a <=( A235  and  A234 );
 a54652a <=( (not A233)  and  a54651a );
 a54655a <=( (not A266)  and  A265 );
 a54658a <=( A269  and  A267 );
 a54659a <=( a54658a  and  a54655a );
 a54660a <=( a54659a  and  a54652a );
 a54664a <=( A167  and  (not A168) );
 a54665a <=( (not A169)  and  a54664a );
 a54668a <=( (not A199)  and  A166 );
 a54671a <=( A232  and  A200 );
 a54672a <=( a54671a  and  a54668a );
 a54673a <=( a54672a  and  a54665a );
 a54677a <=( A236  and  A234 );
 a54678a <=( (not A233)  and  a54677a );
 a54681a <=( (not A266)  and  A265 );
 a54684a <=( A268  and  A267 );
 a54685a <=( a54684a  and  a54681a );
 a54686a <=( a54685a  and  a54678a );
 a54690a <=( A167  and  (not A168) );
 a54691a <=( (not A169)  and  a54690a );
 a54694a <=( (not A199)  and  A166 );
 a54697a <=( A232  and  A200 );
 a54698a <=( a54697a  and  a54694a );
 a54699a <=( a54698a  and  a54691a );
 a54703a <=( A236  and  A234 );
 a54704a <=( (not A233)  and  a54703a );
 a54707a <=( (not A266)  and  A265 );
 a54710a <=( A269  and  A267 );
 a54711a <=( a54710a  and  a54707a );
 a54712a <=( a54711a  and  a54704a );
 a54716a <=( A167  and  (not A168) );
 a54717a <=( (not A169)  and  a54716a );
 a54720a <=( (not A199)  and  A166 );
 a54723a <=( (not A232)  and  A200 );
 a54724a <=( a54723a  and  a54720a );
 a54725a <=( a54724a  and  a54717a );
 a54729a <=( A266  and  A265 );
 a54730a <=( (not A233)  and  a54729a );
 a54733a <=( (not A299)  and  A298 );
 a54736a <=( A301  and  A300 );
 a54737a <=( a54736a  and  a54733a );
 a54738a <=( a54737a  and  a54730a );
 a54742a <=( A167  and  (not A168) );
 a54743a <=( (not A169)  and  a54742a );
 a54746a <=( (not A199)  and  A166 );
 a54749a <=( (not A232)  and  A200 );
 a54750a <=( a54749a  and  a54746a );
 a54751a <=( a54750a  and  a54743a );
 a54755a <=( A266  and  A265 );
 a54756a <=( (not A233)  and  a54755a );
 a54759a <=( (not A299)  and  A298 );
 a54762a <=( A302  and  A300 );
 a54763a <=( a54762a  and  a54759a );
 a54764a <=( a54763a  and  a54756a );
 a54768a <=( A167  and  (not A168) );
 a54769a <=( (not A169)  and  a54768a );
 a54772a <=( (not A199)  and  A166 );
 a54775a <=( (not A232)  and  A200 );
 a54776a <=( a54775a  and  a54772a );
 a54777a <=( a54776a  and  a54769a );
 a54781a <=( (not A267)  and  (not A266) );
 a54782a <=( (not A233)  and  a54781a );
 a54785a <=( (not A299)  and  A298 );
 a54788a <=( A301  and  A300 );
 a54789a <=( a54788a  and  a54785a );
 a54790a <=( a54789a  and  a54782a );
 a54794a <=( A167  and  (not A168) );
 a54795a <=( (not A169)  and  a54794a );
 a54798a <=( (not A199)  and  A166 );
 a54801a <=( (not A232)  and  A200 );
 a54802a <=( a54801a  and  a54798a );
 a54803a <=( a54802a  and  a54795a );
 a54807a <=( (not A267)  and  (not A266) );
 a54808a <=( (not A233)  and  a54807a );
 a54811a <=( (not A299)  and  A298 );
 a54814a <=( A302  and  A300 );
 a54815a <=( a54814a  and  a54811a );
 a54816a <=( a54815a  and  a54808a );
 a54820a <=( A167  and  (not A168) );
 a54821a <=( (not A169)  and  a54820a );
 a54824a <=( (not A199)  and  A166 );
 a54827a <=( (not A232)  and  A200 );
 a54828a <=( a54827a  and  a54824a );
 a54829a <=( a54828a  and  a54821a );
 a54833a <=( (not A266)  and  (not A265) );
 a54834a <=( (not A233)  and  a54833a );
 a54837a <=( (not A299)  and  A298 );
 a54840a <=( A301  and  A300 );
 a54841a <=( a54840a  and  a54837a );
 a54842a <=( a54841a  and  a54834a );
 a54846a <=( A167  and  (not A168) );
 a54847a <=( (not A169)  and  a54846a );
 a54850a <=( (not A199)  and  A166 );
 a54853a <=( (not A232)  and  A200 );
 a54854a <=( a54853a  and  a54850a );
 a54855a <=( a54854a  and  a54847a );
 a54859a <=( (not A266)  and  (not A265) );
 a54860a <=( (not A233)  and  a54859a );
 a54863a <=( (not A299)  and  A298 );
 a54866a <=( A302  and  A300 );
 a54867a <=( a54866a  and  a54863a );
 a54868a <=( a54867a  and  a54860a );
 a54872a <=( A167  and  (not A168) );
 a54873a <=( (not A169)  and  a54872a );
 a54876a <=( A199  and  A166 );
 a54879a <=( A201  and  (not A200) );
 a54880a <=( a54879a  and  a54876a );
 a54881a <=( a54880a  and  a54873a );
 a54885a <=( A233  and  A232 );
 a54886a <=( A202  and  a54885a );
 a54889a <=( (not A267)  and  A265 );
 a54892a <=( A299  and  (not A298) );
 a54893a <=( a54892a  and  a54889a );
 a54894a <=( a54893a  and  a54886a );
 a54898a <=( A167  and  (not A168) );
 a54899a <=( (not A169)  and  a54898a );
 a54902a <=( A199  and  A166 );
 a54905a <=( A201  and  (not A200) );
 a54906a <=( a54905a  and  a54902a );
 a54907a <=( a54906a  and  a54899a );
 a54911a <=( A233  and  A232 );
 a54912a <=( A202  and  a54911a );
 a54915a <=( A266  and  A265 );
 a54918a <=( A299  and  (not A298) );
 a54919a <=( a54918a  and  a54915a );
 a54920a <=( a54919a  and  a54912a );
 a54924a <=( A167  and  (not A168) );
 a54925a <=( (not A169)  and  a54924a );
 a54928a <=( A199  and  A166 );
 a54931a <=( A201  and  (not A200) );
 a54932a <=( a54931a  and  a54928a );
 a54933a <=( a54932a  and  a54925a );
 a54937a <=( A233  and  A232 );
 a54938a <=( A202  and  a54937a );
 a54941a <=( (not A266)  and  (not A265) );
 a54944a <=( A299  and  (not A298) );
 a54945a <=( a54944a  and  a54941a );
 a54946a <=( a54945a  and  a54938a );
 a54950a <=( A167  and  (not A168) );
 a54951a <=( (not A169)  and  a54950a );
 a54954a <=( A199  and  A166 );
 a54957a <=( A201  and  (not A200) );
 a54958a <=( a54957a  and  a54954a );
 a54959a <=( a54958a  and  a54951a );
 a54963a <=( A233  and  (not A232) );
 a54964a <=( A202  and  a54963a );
 a54967a <=( (not A266)  and  A265 );
 a54970a <=( A268  and  A267 );
 a54971a <=( a54970a  and  a54967a );
 a54972a <=( a54971a  and  a54964a );
 a54976a <=( A167  and  (not A168) );
 a54977a <=( (not A169)  and  a54976a );
 a54980a <=( A199  and  A166 );
 a54983a <=( A201  and  (not A200) );
 a54984a <=( a54983a  and  a54980a );
 a54985a <=( a54984a  and  a54977a );
 a54989a <=( A233  and  (not A232) );
 a54990a <=( A202  and  a54989a );
 a54993a <=( (not A266)  and  A265 );
 a54996a <=( A269  and  A267 );
 a54997a <=( a54996a  and  a54993a );
 a54998a <=( a54997a  and  a54990a );
 a55002a <=( A167  and  (not A168) );
 a55003a <=( (not A169)  and  a55002a );
 a55006a <=( A199  and  A166 );
 a55009a <=( A201  and  (not A200) );
 a55010a <=( a55009a  and  a55006a );
 a55011a <=( a55010a  and  a55003a );
 a55015a <=( (not A234)  and  (not A233) );
 a55016a <=( A202  and  a55015a );
 a55019a <=( A266  and  A265 );
 a55022a <=( A299  and  (not A298) );
 a55023a <=( a55022a  and  a55019a );
 a55024a <=( a55023a  and  a55016a );
 a55028a <=( A167  and  (not A168) );
 a55029a <=( (not A169)  and  a55028a );
 a55032a <=( A199  and  A166 );
 a55035a <=( A201  and  (not A200) );
 a55036a <=( a55035a  and  a55032a );
 a55037a <=( a55036a  and  a55029a );
 a55041a <=( (not A234)  and  (not A233) );
 a55042a <=( A202  and  a55041a );
 a55045a <=( (not A267)  and  (not A266) );
 a55048a <=( A299  and  (not A298) );
 a55049a <=( a55048a  and  a55045a );
 a55050a <=( a55049a  and  a55042a );
 a55054a <=( A167  and  (not A168) );
 a55055a <=( (not A169)  and  a55054a );
 a55058a <=( A199  and  A166 );
 a55061a <=( A201  and  (not A200) );
 a55062a <=( a55061a  and  a55058a );
 a55063a <=( a55062a  and  a55055a );
 a55067a <=( (not A234)  and  (not A233) );
 a55068a <=( A202  and  a55067a );
 a55071a <=( (not A266)  and  (not A265) );
 a55074a <=( A299  and  (not A298) );
 a55075a <=( a55074a  and  a55071a );
 a55076a <=( a55075a  and  a55068a );
 a55080a <=( A167  and  (not A168) );
 a55081a <=( (not A169)  and  a55080a );
 a55084a <=( A199  and  A166 );
 a55087a <=( A201  and  (not A200) );
 a55088a <=( a55087a  and  a55084a );
 a55089a <=( a55088a  and  a55081a );
 a55093a <=( (not A233)  and  A232 );
 a55094a <=( A202  and  a55093a );
 a55097a <=( A235  and  A234 );
 a55100a <=( (not A300)  and  A298 );
 a55101a <=( a55100a  and  a55097a );
 a55102a <=( a55101a  and  a55094a );
 a55106a <=( A167  and  (not A168) );
 a55107a <=( (not A169)  and  a55106a );
 a55110a <=( A199  and  A166 );
 a55113a <=( A201  and  (not A200) );
 a55114a <=( a55113a  and  a55110a );
 a55115a <=( a55114a  and  a55107a );
 a55119a <=( (not A233)  and  A232 );
 a55120a <=( A202  and  a55119a );
 a55123a <=( A235  and  A234 );
 a55126a <=( A299  and  A298 );
 a55127a <=( a55126a  and  a55123a );
 a55128a <=( a55127a  and  a55120a );
 a55132a <=( A167  and  (not A168) );
 a55133a <=( (not A169)  and  a55132a );
 a55136a <=( A199  and  A166 );
 a55139a <=( A201  and  (not A200) );
 a55140a <=( a55139a  and  a55136a );
 a55141a <=( a55140a  and  a55133a );
 a55145a <=( (not A233)  and  A232 );
 a55146a <=( A202  and  a55145a );
 a55149a <=( A235  and  A234 );
 a55152a <=( (not A299)  and  (not A298) );
 a55153a <=( a55152a  and  a55149a );
 a55154a <=( a55153a  and  a55146a );
 a55158a <=( A167  and  (not A168) );
 a55159a <=( (not A169)  and  a55158a );
 a55162a <=( A199  and  A166 );
 a55165a <=( A201  and  (not A200) );
 a55166a <=( a55165a  and  a55162a );
 a55167a <=( a55166a  and  a55159a );
 a55171a <=( (not A233)  and  A232 );
 a55172a <=( A202  and  a55171a );
 a55175a <=( A235  and  A234 );
 a55178a <=( A266  and  (not A265) );
 a55179a <=( a55178a  and  a55175a );
 a55180a <=( a55179a  and  a55172a );
 a55184a <=( A167  and  (not A168) );
 a55185a <=( (not A169)  and  a55184a );
 a55188a <=( A199  and  A166 );
 a55191a <=( A201  and  (not A200) );
 a55192a <=( a55191a  and  a55188a );
 a55193a <=( a55192a  and  a55185a );
 a55197a <=( (not A233)  and  A232 );
 a55198a <=( A202  and  a55197a );
 a55201a <=( A236  and  A234 );
 a55204a <=( (not A300)  and  A298 );
 a55205a <=( a55204a  and  a55201a );
 a55206a <=( a55205a  and  a55198a );
 a55210a <=( A167  and  (not A168) );
 a55211a <=( (not A169)  and  a55210a );
 a55214a <=( A199  and  A166 );
 a55217a <=( A201  and  (not A200) );
 a55218a <=( a55217a  and  a55214a );
 a55219a <=( a55218a  and  a55211a );
 a55223a <=( (not A233)  and  A232 );
 a55224a <=( A202  and  a55223a );
 a55227a <=( A236  and  A234 );
 a55230a <=( A299  and  A298 );
 a55231a <=( a55230a  and  a55227a );
 a55232a <=( a55231a  and  a55224a );
 a55236a <=( A167  and  (not A168) );
 a55237a <=( (not A169)  and  a55236a );
 a55240a <=( A199  and  A166 );
 a55243a <=( A201  and  (not A200) );
 a55244a <=( a55243a  and  a55240a );
 a55245a <=( a55244a  and  a55237a );
 a55249a <=( (not A233)  and  A232 );
 a55250a <=( A202  and  a55249a );
 a55253a <=( A236  and  A234 );
 a55256a <=( (not A299)  and  (not A298) );
 a55257a <=( a55256a  and  a55253a );
 a55258a <=( a55257a  and  a55250a );
 a55262a <=( A167  and  (not A168) );
 a55263a <=( (not A169)  and  a55262a );
 a55266a <=( A199  and  A166 );
 a55269a <=( A201  and  (not A200) );
 a55270a <=( a55269a  and  a55266a );
 a55271a <=( a55270a  and  a55263a );
 a55275a <=( (not A233)  and  A232 );
 a55276a <=( A202  and  a55275a );
 a55279a <=( A236  and  A234 );
 a55282a <=( A266  and  (not A265) );
 a55283a <=( a55282a  and  a55279a );
 a55284a <=( a55283a  and  a55276a );
 a55288a <=( A167  and  (not A168) );
 a55289a <=( (not A169)  and  a55288a );
 a55292a <=( A199  and  A166 );
 a55295a <=( A201  and  (not A200) );
 a55296a <=( a55295a  and  a55292a );
 a55297a <=( a55296a  and  a55289a );
 a55301a <=( (not A233)  and  (not A232) );
 a55302a <=( A202  and  a55301a );
 a55305a <=( A266  and  A265 );
 a55308a <=( A299  and  (not A298) );
 a55309a <=( a55308a  and  a55305a );
 a55310a <=( a55309a  and  a55302a );
 a55314a <=( A167  and  (not A168) );
 a55315a <=( (not A169)  and  a55314a );
 a55318a <=( A199  and  A166 );
 a55321a <=( A201  and  (not A200) );
 a55322a <=( a55321a  and  a55318a );
 a55323a <=( a55322a  and  a55315a );
 a55327a <=( (not A233)  and  (not A232) );
 a55328a <=( A202  and  a55327a );
 a55331a <=( (not A267)  and  (not A266) );
 a55334a <=( A299  and  (not A298) );
 a55335a <=( a55334a  and  a55331a );
 a55336a <=( a55335a  and  a55328a );
 a55340a <=( A167  and  (not A168) );
 a55341a <=( (not A169)  and  a55340a );
 a55344a <=( A199  and  A166 );
 a55347a <=( A201  and  (not A200) );
 a55348a <=( a55347a  and  a55344a );
 a55349a <=( a55348a  and  a55341a );
 a55353a <=( (not A233)  and  (not A232) );
 a55354a <=( A202  and  a55353a );
 a55357a <=( (not A266)  and  (not A265) );
 a55360a <=( A299  and  (not A298) );
 a55361a <=( a55360a  and  a55357a );
 a55362a <=( a55361a  and  a55354a );
 a55366a <=( A167  and  (not A168) );
 a55367a <=( (not A169)  and  a55366a );
 a55370a <=( A199  and  A166 );
 a55373a <=( A201  and  (not A200) );
 a55374a <=( a55373a  and  a55370a );
 a55375a <=( a55374a  and  a55367a );
 a55379a <=( A233  and  A232 );
 a55380a <=( A203  and  a55379a );
 a55383a <=( (not A267)  and  A265 );
 a55386a <=( A299  and  (not A298) );
 a55387a <=( a55386a  and  a55383a );
 a55388a <=( a55387a  and  a55380a );
 a55392a <=( A167  and  (not A168) );
 a55393a <=( (not A169)  and  a55392a );
 a55396a <=( A199  and  A166 );
 a55399a <=( A201  and  (not A200) );
 a55400a <=( a55399a  and  a55396a );
 a55401a <=( a55400a  and  a55393a );
 a55405a <=( A233  and  A232 );
 a55406a <=( A203  and  a55405a );
 a55409a <=( A266  and  A265 );
 a55412a <=( A299  and  (not A298) );
 a55413a <=( a55412a  and  a55409a );
 a55414a <=( a55413a  and  a55406a );
 a55418a <=( A167  and  (not A168) );
 a55419a <=( (not A169)  and  a55418a );
 a55422a <=( A199  and  A166 );
 a55425a <=( A201  and  (not A200) );
 a55426a <=( a55425a  and  a55422a );
 a55427a <=( a55426a  and  a55419a );
 a55431a <=( A233  and  A232 );
 a55432a <=( A203  and  a55431a );
 a55435a <=( (not A266)  and  (not A265) );
 a55438a <=( A299  and  (not A298) );
 a55439a <=( a55438a  and  a55435a );
 a55440a <=( a55439a  and  a55432a );
 a55444a <=( A167  and  (not A168) );
 a55445a <=( (not A169)  and  a55444a );
 a55448a <=( A199  and  A166 );
 a55451a <=( A201  and  (not A200) );
 a55452a <=( a55451a  and  a55448a );
 a55453a <=( a55452a  and  a55445a );
 a55457a <=( A233  and  (not A232) );
 a55458a <=( A203  and  a55457a );
 a55461a <=( (not A266)  and  A265 );
 a55464a <=( A268  and  A267 );
 a55465a <=( a55464a  and  a55461a );
 a55466a <=( a55465a  and  a55458a );
 a55470a <=( A167  and  (not A168) );
 a55471a <=( (not A169)  and  a55470a );
 a55474a <=( A199  and  A166 );
 a55477a <=( A201  and  (not A200) );
 a55478a <=( a55477a  and  a55474a );
 a55479a <=( a55478a  and  a55471a );
 a55483a <=( A233  and  (not A232) );
 a55484a <=( A203  and  a55483a );
 a55487a <=( (not A266)  and  A265 );
 a55490a <=( A269  and  A267 );
 a55491a <=( a55490a  and  a55487a );
 a55492a <=( a55491a  and  a55484a );
 a55496a <=( A167  and  (not A168) );
 a55497a <=( (not A169)  and  a55496a );
 a55500a <=( A199  and  A166 );
 a55503a <=( A201  and  (not A200) );
 a55504a <=( a55503a  and  a55500a );
 a55505a <=( a55504a  and  a55497a );
 a55509a <=( (not A234)  and  (not A233) );
 a55510a <=( A203  and  a55509a );
 a55513a <=( A266  and  A265 );
 a55516a <=( A299  and  (not A298) );
 a55517a <=( a55516a  and  a55513a );
 a55518a <=( a55517a  and  a55510a );
 a55522a <=( A167  and  (not A168) );
 a55523a <=( (not A169)  and  a55522a );
 a55526a <=( A199  and  A166 );
 a55529a <=( A201  and  (not A200) );
 a55530a <=( a55529a  and  a55526a );
 a55531a <=( a55530a  and  a55523a );
 a55535a <=( (not A234)  and  (not A233) );
 a55536a <=( A203  and  a55535a );
 a55539a <=( (not A267)  and  (not A266) );
 a55542a <=( A299  and  (not A298) );
 a55543a <=( a55542a  and  a55539a );
 a55544a <=( a55543a  and  a55536a );
 a55548a <=( A167  and  (not A168) );
 a55549a <=( (not A169)  and  a55548a );
 a55552a <=( A199  and  A166 );
 a55555a <=( A201  and  (not A200) );
 a55556a <=( a55555a  and  a55552a );
 a55557a <=( a55556a  and  a55549a );
 a55561a <=( (not A234)  and  (not A233) );
 a55562a <=( A203  and  a55561a );
 a55565a <=( (not A266)  and  (not A265) );
 a55568a <=( A299  and  (not A298) );
 a55569a <=( a55568a  and  a55565a );
 a55570a <=( a55569a  and  a55562a );
 a55574a <=( A167  and  (not A168) );
 a55575a <=( (not A169)  and  a55574a );
 a55578a <=( A199  and  A166 );
 a55581a <=( A201  and  (not A200) );
 a55582a <=( a55581a  and  a55578a );
 a55583a <=( a55582a  and  a55575a );
 a55587a <=( (not A233)  and  A232 );
 a55588a <=( A203  and  a55587a );
 a55591a <=( A235  and  A234 );
 a55594a <=( (not A300)  and  A298 );
 a55595a <=( a55594a  and  a55591a );
 a55596a <=( a55595a  and  a55588a );
 a55600a <=( A167  and  (not A168) );
 a55601a <=( (not A169)  and  a55600a );
 a55604a <=( A199  and  A166 );
 a55607a <=( A201  and  (not A200) );
 a55608a <=( a55607a  and  a55604a );
 a55609a <=( a55608a  and  a55601a );
 a55613a <=( (not A233)  and  A232 );
 a55614a <=( A203  and  a55613a );
 a55617a <=( A235  and  A234 );
 a55620a <=( A299  and  A298 );
 a55621a <=( a55620a  and  a55617a );
 a55622a <=( a55621a  and  a55614a );
 a55626a <=( A167  and  (not A168) );
 a55627a <=( (not A169)  and  a55626a );
 a55630a <=( A199  and  A166 );
 a55633a <=( A201  and  (not A200) );
 a55634a <=( a55633a  and  a55630a );
 a55635a <=( a55634a  and  a55627a );
 a55639a <=( (not A233)  and  A232 );
 a55640a <=( A203  and  a55639a );
 a55643a <=( A235  and  A234 );
 a55646a <=( (not A299)  and  (not A298) );
 a55647a <=( a55646a  and  a55643a );
 a55648a <=( a55647a  and  a55640a );
 a55652a <=( A167  and  (not A168) );
 a55653a <=( (not A169)  and  a55652a );
 a55656a <=( A199  and  A166 );
 a55659a <=( A201  and  (not A200) );
 a55660a <=( a55659a  and  a55656a );
 a55661a <=( a55660a  and  a55653a );
 a55665a <=( (not A233)  and  A232 );
 a55666a <=( A203  and  a55665a );
 a55669a <=( A235  and  A234 );
 a55672a <=( A266  and  (not A265) );
 a55673a <=( a55672a  and  a55669a );
 a55674a <=( a55673a  and  a55666a );
 a55678a <=( A167  and  (not A168) );
 a55679a <=( (not A169)  and  a55678a );
 a55682a <=( A199  and  A166 );
 a55685a <=( A201  and  (not A200) );
 a55686a <=( a55685a  and  a55682a );
 a55687a <=( a55686a  and  a55679a );
 a55691a <=( (not A233)  and  A232 );
 a55692a <=( A203  and  a55691a );
 a55695a <=( A236  and  A234 );
 a55698a <=( (not A300)  and  A298 );
 a55699a <=( a55698a  and  a55695a );
 a55700a <=( a55699a  and  a55692a );
 a55704a <=( A167  and  (not A168) );
 a55705a <=( (not A169)  and  a55704a );
 a55708a <=( A199  and  A166 );
 a55711a <=( A201  and  (not A200) );
 a55712a <=( a55711a  and  a55708a );
 a55713a <=( a55712a  and  a55705a );
 a55717a <=( (not A233)  and  A232 );
 a55718a <=( A203  and  a55717a );
 a55721a <=( A236  and  A234 );
 a55724a <=( A299  and  A298 );
 a55725a <=( a55724a  and  a55721a );
 a55726a <=( a55725a  and  a55718a );
 a55730a <=( A167  and  (not A168) );
 a55731a <=( (not A169)  and  a55730a );
 a55734a <=( A199  and  A166 );
 a55737a <=( A201  and  (not A200) );
 a55738a <=( a55737a  and  a55734a );
 a55739a <=( a55738a  and  a55731a );
 a55743a <=( (not A233)  and  A232 );
 a55744a <=( A203  and  a55743a );
 a55747a <=( A236  and  A234 );
 a55750a <=( (not A299)  and  (not A298) );
 a55751a <=( a55750a  and  a55747a );
 a55752a <=( a55751a  and  a55744a );
 a55756a <=( A167  and  (not A168) );
 a55757a <=( (not A169)  and  a55756a );
 a55760a <=( A199  and  A166 );
 a55763a <=( A201  and  (not A200) );
 a55764a <=( a55763a  and  a55760a );
 a55765a <=( a55764a  and  a55757a );
 a55769a <=( (not A233)  and  A232 );
 a55770a <=( A203  and  a55769a );
 a55773a <=( A236  and  A234 );
 a55776a <=( A266  and  (not A265) );
 a55777a <=( a55776a  and  a55773a );
 a55778a <=( a55777a  and  a55770a );
 a55782a <=( A167  and  (not A168) );
 a55783a <=( (not A169)  and  a55782a );
 a55786a <=( A199  and  A166 );
 a55789a <=( A201  and  (not A200) );
 a55790a <=( a55789a  and  a55786a );
 a55791a <=( a55790a  and  a55783a );
 a55795a <=( (not A233)  and  (not A232) );
 a55796a <=( A203  and  a55795a );
 a55799a <=( A266  and  A265 );
 a55802a <=( A299  and  (not A298) );
 a55803a <=( a55802a  and  a55799a );
 a55804a <=( a55803a  and  a55796a );
 a55808a <=( A167  and  (not A168) );
 a55809a <=( (not A169)  and  a55808a );
 a55812a <=( A199  and  A166 );
 a55815a <=( A201  and  (not A200) );
 a55816a <=( a55815a  and  a55812a );
 a55817a <=( a55816a  and  a55809a );
 a55821a <=( (not A233)  and  (not A232) );
 a55822a <=( A203  and  a55821a );
 a55825a <=( (not A267)  and  (not A266) );
 a55828a <=( A299  and  (not A298) );
 a55829a <=( a55828a  and  a55825a );
 a55830a <=( a55829a  and  a55822a );
 a55834a <=( A167  and  (not A168) );
 a55835a <=( (not A169)  and  a55834a );
 a55838a <=( A199  and  A166 );
 a55841a <=( A201  and  (not A200) );
 a55842a <=( a55841a  and  a55838a );
 a55843a <=( a55842a  and  a55835a );
 a55847a <=( (not A233)  and  (not A232) );
 a55848a <=( A203  and  a55847a );
 a55851a <=( (not A266)  and  (not A265) );
 a55854a <=( A299  and  (not A298) );
 a55855a <=( a55854a  and  a55851a );
 a55856a <=( a55855a  and  a55848a );
 a55860a <=( A167  and  (not A169) );
 a55861a <=( A170  and  a55860a );
 a55864a <=( A199  and  (not A166) );
 a55867a <=( A232  and  A200 );
 a55868a <=( a55867a  and  a55864a );
 a55869a <=( a55868a  and  a55861a );
 a55873a <=( (not A267)  and  A265 );
 a55874a <=( A233  and  a55873a );
 a55877a <=( (not A299)  and  A298 );
 a55880a <=( A301  and  A300 );
 a55881a <=( a55880a  and  a55877a );
 a55882a <=( a55881a  and  a55874a );
 a55886a <=( A167  and  (not A169) );
 a55887a <=( A170  and  a55886a );
 a55890a <=( A199  and  (not A166) );
 a55893a <=( A232  and  A200 );
 a55894a <=( a55893a  and  a55890a );
 a55895a <=( a55894a  and  a55887a );
 a55899a <=( (not A267)  and  A265 );
 a55900a <=( A233  and  a55899a );
 a55903a <=( (not A299)  and  A298 );
 a55906a <=( A302  and  A300 );
 a55907a <=( a55906a  and  a55903a );
 a55908a <=( a55907a  and  a55900a );
 a55912a <=( A167  and  (not A169) );
 a55913a <=( A170  and  a55912a );
 a55916a <=( A199  and  (not A166) );
 a55919a <=( A232  and  A200 );
 a55920a <=( a55919a  and  a55916a );
 a55921a <=( a55920a  and  a55913a );
 a55925a <=( A266  and  A265 );
 a55926a <=( A233  and  a55925a );
 a55929a <=( (not A299)  and  A298 );
 a55932a <=( A301  and  A300 );
 a55933a <=( a55932a  and  a55929a );
 a55934a <=( a55933a  and  a55926a );
 a55938a <=( A167  and  (not A169) );
 a55939a <=( A170  and  a55938a );
 a55942a <=( A199  and  (not A166) );
 a55945a <=( A232  and  A200 );
 a55946a <=( a55945a  and  a55942a );
 a55947a <=( a55946a  and  a55939a );
 a55951a <=( A266  and  A265 );
 a55952a <=( A233  and  a55951a );
 a55955a <=( (not A299)  and  A298 );
 a55958a <=( A302  and  A300 );
 a55959a <=( a55958a  and  a55955a );
 a55960a <=( a55959a  and  a55952a );
 a55964a <=( A167  and  (not A169) );
 a55965a <=( A170  and  a55964a );
 a55968a <=( A199  and  (not A166) );
 a55971a <=( A232  and  A200 );
 a55972a <=( a55971a  and  a55968a );
 a55973a <=( a55972a  and  a55965a );
 a55977a <=( (not A266)  and  (not A265) );
 a55978a <=( A233  and  a55977a );
 a55981a <=( (not A299)  and  A298 );
 a55984a <=( A301  and  A300 );
 a55985a <=( a55984a  and  a55981a );
 a55986a <=( a55985a  and  a55978a );
 a55990a <=( A167  and  (not A169) );
 a55991a <=( A170  and  a55990a );
 a55994a <=( A199  and  (not A166) );
 a55997a <=( A232  and  A200 );
 a55998a <=( a55997a  and  a55994a );
 a55999a <=( a55998a  and  a55991a );
 a56003a <=( (not A266)  and  (not A265) );
 a56004a <=( A233  and  a56003a );
 a56007a <=( (not A299)  and  A298 );
 a56010a <=( A302  and  A300 );
 a56011a <=( a56010a  and  a56007a );
 a56012a <=( a56011a  and  a56004a );
 a56016a <=( A167  and  (not A169) );
 a56017a <=( A170  and  a56016a );
 a56020a <=( A199  and  (not A166) );
 a56023a <=( (not A233)  and  A200 );
 a56024a <=( a56023a  and  a56020a );
 a56025a <=( a56024a  and  a56017a );
 a56029a <=( (not A266)  and  (not A236) );
 a56030a <=( (not A235)  and  a56029a );
 a56033a <=( (not A269)  and  (not A268) );
 a56036a <=( A299  and  (not A298) );
 a56037a <=( a56036a  and  a56033a );
 a56038a <=( a56037a  and  a56030a );
 a56042a <=( A167  and  (not A169) );
 a56043a <=( A170  and  a56042a );
 a56046a <=( A199  and  (not A166) );
 a56049a <=( (not A233)  and  A200 );
 a56050a <=( a56049a  and  a56046a );
 a56051a <=( a56050a  and  a56043a );
 a56055a <=( A266  and  A265 );
 a56056a <=( (not A234)  and  a56055a );
 a56059a <=( (not A299)  and  A298 );
 a56062a <=( A301  and  A300 );
 a56063a <=( a56062a  and  a56059a );
 a56064a <=( a56063a  and  a56056a );
 a56068a <=( A167  and  (not A169) );
 a56069a <=( A170  and  a56068a );
 a56072a <=( A199  and  (not A166) );
 a56075a <=( (not A233)  and  A200 );
 a56076a <=( a56075a  and  a56072a );
 a56077a <=( a56076a  and  a56069a );
 a56081a <=( A266  and  A265 );
 a56082a <=( (not A234)  and  a56081a );
 a56085a <=( (not A299)  and  A298 );
 a56088a <=( A302  and  A300 );
 a56089a <=( a56088a  and  a56085a );
 a56090a <=( a56089a  and  a56082a );
 a56094a <=( A167  and  (not A169) );
 a56095a <=( A170  and  a56094a );
 a56098a <=( A199  and  (not A166) );
 a56101a <=( (not A233)  and  A200 );
 a56102a <=( a56101a  and  a56098a );
 a56103a <=( a56102a  and  a56095a );
 a56107a <=( (not A267)  and  (not A266) );
 a56108a <=( (not A234)  and  a56107a );
 a56111a <=( (not A299)  and  A298 );
 a56114a <=( A301  and  A300 );
 a56115a <=( a56114a  and  a56111a );
 a56116a <=( a56115a  and  a56108a );
 a56120a <=( A167  and  (not A169) );
 a56121a <=( A170  and  a56120a );
 a56124a <=( A199  and  (not A166) );
 a56127a <=( (not A233)  and  A200 );
 a56128a <=( a56127a  and  a56124a );
 a56129a <=( a56128a  and  a56121a );
 a56133a <=( (not A267)  and  (not A266) );
 a56134a <=( (not A234)  and  a56133a );
 a56137a <=( (not A299)  and  A298 );
 a56140a <=( A302  and  A300 );
 a56141a <=( a56140a  and  a56137a );
 a56142a <=( a56141a  and  a56134a );
 a56146a <=( A167  and  (not A169) );
 a56147a <=( A170  and  a56146a );
 a56150a <=( A199  and  (not A166) );
 a56153a <=( (not A233)  and  A200 );
 a56154a <=( a56153a  and  a56150a );
 a56155a <=( a56154a  and  a56147a );
 a56159a <=( (not A266)  and  (not A265) );
 a56160a <=( (not A234)  and  a56159a );
 a56163a <=( (not A299)  and  A298 );
 a56166a <=( A301  and  A300 );
 a56167a <=( a56166a  and  a56163a );
 a56168a <=( a56167a  and  a56160a );
 a56172a <=( A167  and  (not A169) );
 a56173a <=( A170  and  a56172a );
 a56176a <=( A199  and  (not A166) );
 a56179a <=( (not A233)  and  A200 );
 a56180a <=( a56179a  and  a56176a );
 a56181a <=( a56180a  and  a56173a );
 a56185a <=( (not A266)  and  (not A265) );
 a56186a <=( (not A234)  and  a56185a );
 a56189a <=( (not A299)  and  A298 );
 a56192a <=( A302  and  A300 );
 a56193a <=( a56192a  and  a56189a );
 a56194a <=( a56193a  and  a56186a );
 a56198a <=( A167  and  (not A169) );
 a56199a <=( A170  and  a56198a );
 a56202a <=( A199  and  (not A166) );
 a56205a <=( A232  and  A200 );
 a56206a <=( a56205a  and  a56202a );
 a56207a <=( a56206a  and  a56199a );
 a56211a <=( A235  and  A234 );
 a56212a <=( (not A233)  and  a56211a );
 a56215a <=( (not A266)  and  A265 );
 a56218a <=( A268  and  A267 );
 a56219a <=( a56218a  and  a56215a );
 a56220a <=( a56219a  and  a56212a );
 a56224a <=( A167  and  (not A169) );
 a56225a <=( A170  and  a56224a );
 a56228a <=( A199  and  (not A166) );
 a56231a <=( A232  and  A200 );
 a56232a <=( a56231a  and  a56228a );
 a56233a <=( a56232a  and  a56225a );
 a56237a <=( A235  and  A234 );
 a56238a <=( (not A233)  and  a56237a );
 a56241a <=( (not A266)  and  A265 );
 a56244a <=( A269  and  A267 );
 a56245a <=( a56244a  and  a56241a );
 a56246a <=( a56245a  and  a56238a );
 a56250a <=( A167  and  (not A169) );
 a56251a <=( A170  and  a56250a );
 a56254a <=( A199  and  (not A166) );
 a56257a <=( A232  and  A200 );
 a56258a <=( a56257a  and  a56254a );
 a56259a <=( a56258a  and  a56251a );
 a56263a <=( A236  and  A234 );
 a56264a <=( (not A233)  and  a56263a );
 a56267a <=( (not A266)  and  A265 );
 a56270a <=( A268  and  A267 );
 a56271a <=( a56270a  and  a56267a );
 a56272a <=( a56271a  and  a56264a );
 a56276a <=( A167  and  (not A169) );
 a56277a <=( A170  and  a56276a );
 a56280a <=( A199  and  (not A166) );
 a56283a <=( A232  and  A200 );
 a56284a <=( a56283a  and  a56280a );
 a56285a <=( a56284a  and  a56277a );
 a56289a <=( A236  and  A234 );
 a56290a <=( (not A233)  and  a56289a );
 a56293a <=( (not A266)  and  A265 );
 a56296a <=( A269  and  A267 );
 a56297a <=( a56296a  and  a56293a );
 a56298a <=( a56297a  and  a56290a );
 a56302a <=( A167  and  (not A169) );
 a56303a <=( A170  and  a56302a );
 a56306a <=( A199  and  (not A166) );
 a56309a <=( (not A232)  and  A200 );
 a56310a <=( a56309a  and  a56306a );
 a56311a <=( a56310a  and  a56303a );
 a56315a <=( A266  and  A265 );
 a56316a <=( (not A233)  and  a56315a );
 a56319a <=( (not A299)  and  A298 );
 a56322a <=( A301  and  A300 );
 a56323a <=( a56322a  and  a56319a );
 a56324a <=( a56323a  and  a56316a );
 a56328a <=( A167  and  (not A169) );
 a56329a <=( A170  and  a56328a );
 a56332a <=( A199  and  (not A166) );
 a56335a <=( (not A232)  and  A200 );
 a56336a <=( a56335a  and  a56332a );
 a56337a <=( a56336a  and  a56329a );
 a56341a <=( A266  and  A265 );
 a56342a <=( (not A233)  and  a56341a );
 a56345a <=( (not A299)  and  A298 );
 a56348a <=( A302  and  A300 );
 a56349a <=( a56348a  and  a56345a );
 a56350a <=( a56349a  and  a56342a );
 a56354a <=( A167  and  (not A169) );
 a56355a <=( A170  and  a56354a );
 a56358a <=( A199  and  (not A166) );
 a56361a <=( (not A232)  and  A200 );
 a56362a <=( a56361a  and  a56358a );
 a56363a <=( a56362a  and  a56355a );
 a56367a <=( (not A267)  and  (not A266) );
 a56368a <=( (not A233)  and  a56367a );
 a56371a <=( (not A299)  and  A298 );
 a56374a <=( A301  and  A300 );
 a56375a <=( a56374a  and  a56371a );
 a56376a <=( a56375a  and  a56368a );
 a56380a <=( A167  and  (not A169) );
 a56381a <=( A170  and  a56380a );
 a56384a <=( A199  and  (not A166) );
 a56387a <=( (not A232)  and  A200 );
 a56388a <=( a56387a  and  a56384a );
 a56389a <=( a56388a  and  a56381a );
 a56393a <=( (not A267)  and  (not A266) );
 a56394a <=( (not A233)  and  a56393a );
 a56397a <=( (not A299)  and  A298 );
 a56400a <=( A302  and  A300 );
 a56401a <=( a56400a  and  a56397a );
 a56402a <=( a56401a  and  a56394a );
 a56406a <=( A167  and  (not A169) );
 a56407a <=( A170  and  a56406a );
 a56410a <=( A199  and  (not A166) );
 a56413a <=( (not A232)  and  A200 );
 a56414a <=( a56413a  and  a56410a );
 a56415a <=( a56414a  and  a56407a );
 a56419a <=( (not A266)  and  (not A265) );
 a56420a <=( (not A233)  and  a56419a );
 a56423a <=( (not A299)  and  A298 );
 a56426a <=( A301  and  A300 );
 a56427a <=( a56426a  and  a56423a );
 a56428a <=( a56427a  and  a56420a );
 a56432a <=( A167  and  (not A169) );
 a56433a <=( A170  and  a56432a );
 a56436a <=( A199  and  (not A166) );
 a56439a <=( (not A232)  and  A200 );
 a56440a <=( a56439a  and  a56436a );
 a56441a <=( a56440a  and  a56433a );
 a56445a <=( (not A266)  and  (not A265) );
 a56446a <=( (not A233)  and  a56445a );
 a56449a <=( (not A299)  and  A298 );
 a56452a <=( A302  and  A300 );
 a56453a <=( a56452a  and  a56449a );
 a56454a <=( a56453a  and  a56446a );
 a56458a <=( A167  and  (not A169) );
 a56459a <=( A170  and  a56458a );
 a56462a <=( (not A200)  and  (not A166) );
 a56465a <=( (not A203)  and  (not A202) );
 a56466a <=( a56465a  and  a56462a );
 a56467a <=( a56466a  and  a56459a );
 a56471a <=( A265  and  A233 );
 a56472a <=( A232  and  a56471a );
 a56475a <=( (not A269)  and  (not A268) );
 a56478a <=( A299  and  (not A298) );
 a56479a <=( a56478a  and  a56475a );
 a56480a <=( a56479a  and  a56472a );
 a56484a <=( A167  and  (not A169) );
 a56485a <=( A170  and  a56484a );
 a56488a <=( (not A200)  and  (not A166) );
 a56491a <=( (not A203)  and  (not A202) );
 a56492a <=( a56491a  and  a56488a );
 a56493a <=( a56492a  and  a56485a );
 a56497a <=( (not A236)  and  (not A235) );
 a56498a <=( (not A233)  and  a56497a );
 a56501a <=( A266  and  A265 );
 a56504a <=( A299  and  (not A298) );
 a56505a <=( a56504a  and  a56501a );
 a56506a <=( a56505a  and  a56498a );
 a56510a <=( A167  and  (not A169) );
 a56511a <=( A170  and  a56510a );
 a56514a <=( (not A200)  and  (not A166) );
 a56517a <=( (not A203)  and  (not A202) );
 a56518a <=( a56517a  and  a56514a );
 a56519a <=( a56518a  and  a56511a );
 a56523a <=( (not A236)  and  (not A235) );
 a56524a <=( (not A233)  and  a56523a );
 a56527a <=( (not A267)  and  (not A266) );
 a56530a <=( A299  and  (not A298) );
 a56531a <=( a56530a  and  a56527a );
 a56532a <=( a56531a  and  a56524a );
 a56536a <=( A167  and  (not A169) );
 a56537a <=( A170  and  a56536a );
 a56540a <=( (not A200)  and  (not A166) );
 a56543a <=( (not A203)  and  (not A202) );
 a56544a <=( a56543a  and  a56540a );
 a56545a <=( a56544a  and  a56537a );
 a56549a <=( (not A236)  and  (not A235) );
 a56550a <=( (not A233)  and  a56549a );
 a56553a <=( (not A266)  and  (not A265) );
 a56556a <=( A299  and  (not A298) );
 a56557a <=( a56556a  and  a56553a );
 a56558a <=( a56557a  and  a56550a );
 a56562a <=( A167  and  (not A169) );
 a56563a <=( A170  and  a56562a );
 a56566a <=( (not A200)  and  (not A166) );
 a56569a <=( (not A203)  and  (not A202) );
 a56570a <=( a56569a  and  a56566a );
 a56571a <=( a56570a  and  a56563a );
 a56575a <=( (not A266)  and  (not A234) );
 a56576a <=( (not A233)  and  a56575a );
 a56579a <=( (not A269)  and  (not A268) );
 a56582a <=( A299  and  (not A298) );
 a56583a <=( a56582a  and  a56579a );
 a56584a <=( a56583a  and  a56576a );
 a56588a <=( A167  and  (not A169) );
 a56589a <=( A170  and  a56588a );
 a56592a <=( (not A200)  and  (not A166) );
 a56595a <=( (not A203)  and  (not A202) );
 a56596a <=( a56595a  and  a56592a );
 a56597a <=( a56596a  and  a56589a );
 a56601a <=( A234  and  (not A233) );
 a56602a <=( A232  and  a56601a );
 a56605a <=( A298  and  A235 );
 a56608a <=( (not A302)  and  (not A301) );
 a56609a <=( a56608a  and  a56605a );
 a56610a <=( a56609a  and  a56602a );
 a56614a <=( A167  and  (not A169) );
 a56615a <=( A170  and  a56614a );
 a56618a <=( (not A200)  and  (not A166) );
 a56621a <=( (not A203)  and  (not A202) );
 a56622a <=( a56621a  and  a56618a );
 a56623a <=( a56622a  and  a56615a );
 a56627a <=( A234  and  (not A233) );
 a56628a <=( A232  and  a56627a );
 a56631a <=( A298  and  A236 );
 a56634a <=( (not A302)  and  (not A301) );
 a56635a <=( a56634a  and  a56631a );
 a56636a <=( a56635a  and  a56628a );
 a56640a <=( A167  and  (not A169) );
 a56641a <=( A170  and  a56640a );
 a56644a <=( (not A200)  and  (not A166) );
 a56647a <=( (not A203)  and  (not A202) );
 a56648a <=( a56647a  and  a56644a );
 a56649a <=( a56648a  and  a56641a );
 a56653a <=( (not A266)  and  (not A233) );
 a56654a <=( (not A232)  and  a56653a );
 a56657a <=( (not A269)  and  (not A268) );
 a56660a <=( A299  and  (not A298) );
 a56661a <=( a56660a  and  a56657a );
 a56662a <=( a56661a  and  a56654a );
 a56666a <=( A167  and  (not A169) );
 a56667a <=( A170  and  a56666a );
 a56670a <=( (not A200)  and  (not A166) );
 a56673a <=( A232  and  (not A201) );
 a56674a <=( a56673a  and  a56670a );
 a56675a <=( a56674a  and  a56667a );
 a56679a <=( (not A267)  and  A265 );
 a56680a <=( A233  and  a56679a );
 a56683a <=( (not A299)  and  A298 );
 a56686a <=( A301  and  A300 );
 a56687a <=( a56686a  and  a56683a );
 a56688a <=( a56687a  and  a56680a );
 a56692a <=( A167  and  (not A169) );
 a56693a <=( A170  and  a56692a );
 a56696a <=( (not A200)  and  (not A166) );
 a56699a <=( A232  and  (not A201) );
 a56700a <=( a56699a  and  a56696a );
 a56701a <=( a56700a  and  a56693a );
 a56705a <=( (not A267)  and  A265 );
 a56706a <=( A233  and  a56705a );
 a56709a <=( (not A299)  and  A298 );
 a56712a <=( A302  and  A300 );
 a56713a <=( a56712a  and  a56709a );
 a56714a <=( a56713a  and  a56706a );
 a56718a <=( A167  and  (not A169) );
 a56719a <=( A170  and  a56718a );
 a56722a <=( (not A200)  and  (not A166) );
 a56725a <=( A232  and  (not A201) );
 a56726a <=( a56725a  and  a56722a );
 a56727a <=( a56726a  and  a56719a );
 a56731a <=( A266  and  A265 );
 a56732a <=( A233  and  a56731a );
 a56735a <=( (not A299)  and  A298 );
 a56738a <=( A301  and  A300 );
 a56739a <=( a56738a  and  a56735a );
 a56740a <=( a56739a  and  a56732a );
 a56744a <=( A167  and  (not A169) );
 a56745a <=( A170  and  a56744a );
 a56748a <=( (not A200)  and  (not A166) );
 a56751a <=( A232  and  (not A201) );
 a56752a <=( a56751a  and  a56748a );
 a56753a <=( a56752a  and  a56745a );
 a56757a <=( A266  and  A265 );
 a56758a <=( A233  and  a56757a );
 a56761a <=( (not A299)  and  A298 );
 a56764a <=( A302  and  A300 );
 a56765a <=( a56764a  and  a56761a );
 a56766a <=( a56765a  and  a56758a );
 a56770a <=( A167  and  (not A169) );
 a56771a <=( A170  and  a56770a );
 a56774a <=( (not A200)  and  (not A166) );
 a56777a <=( A232  and  (not A201) );
 a56778a <=( a56777a  and  a56774a );
 a56779a <=( a56778a  and  a56771a );
 a56783a <=( (not A266)  and  (not A265) );
 a56784a <=( A233  and  a56783a );
 a56787a <=( (not A299)  and  A298 );
 a56790a <=( A301  and  A300 );
 a56791a <=( a56790a  and  a56787a );
 a56792a <=( a56791a  and  a56784a );
 a56796a <=( A167  and  (not A169) );
 a56797a <=( A170  and  a56796a );
 a56800a <=( (not A200)  and  (not A166) );
 a56803a <=( A232  and  (not A201) );
 a56804a <=( a56803a  and  a56800a );
 a56805a <=( a56804a  and  a56797a );
 a56809a <=( (not A266)  and  (not A265) );
 a56810a <=( A233  and  a56809a );
 a56813a <=( (not A299)  and  A298 );
 a56816a <=( A302  and  A300 );
 a56817a <=( a56816a  and  a56813a );
 a56818a <=( a56817a  and  a56810a );
 a56822a <=( A167  and  (not A169) );
 a56823a <=( A170  and  a56822a );
 a56826a <=( (not A200)  and  (not A166) );
 a56829a <=( (not A233)  and  (not A201) );
 a56830a <=( a56829a  and  a56826a );
 a56831a <=( a56830a  and  a56823a );
 a56835a <=( (not A266)  and  (not A236) );
 a56836a <=( (not A235)  and  a56835a );
 a56839a <=( (not A269)  and  (not A268) );
 a56842a <=( A299  and  (not A298) );
 a56843a <=( a56842a  and  a56839a );
 a56844a <=( a56843a  and  a56836a );
 a56848a <=( A167  and  (not A169) );
 a56849a <=( A170  and  a56848a );
 a56852a <=( (not A200)  and  (not A166) );
 a56855a <=( (not A233)  and  (not A201) );
 a56856a <=( a56855a  and  a56852a );
 a56857a <=( a56856a  and  a56849a );
 a56861a <=( A266  and  A265 );
 a56862a <=( (not A234)  and  a56861a );
 a56865a <=( (not A299)  and  A298 );
 a56868a <=( A301  and  A300 );
 a56869a <=( a56868a  and  a56865a );
 a56870a <=( a56869a  and  a56862a );
 a56874a <=( A167  and  (not A169) );
 a56875a <=( A170  and  a56874a );
 a56878a <=( (not A200)  and  (not A166) );
 a56881a <=( (not A233)  and  (not A201) );
 a56882a <=( a56881a  and  a56878a );
 a56883a <=( a56882a  and  a56875a );
 a56887a <=( A266  and  A265 );
 a56888a <=( (not A234)  and  a56887a );
 a56891a <=( (not A299)  and  A298 );
 a56894a <=( A302  and  A300 );
 a56895a <=( a56894a  and  a56891a );
 a56896a <=( a56895a  and  a56888a );
 a56900a <=( A167  and  (not A169) );
 a56901a <=( A170  and  a56900a );
 a56904a <=( (not A200)  and  (not A166) );
 a56907a <=( (not A233)  and  (not A201) );
 a56908a <=( a56907a  and  a56904a );
 a56909a <=( a56908a  and  a56901a );
 a56913a <=( (not A267)  and  (not A266) );
 a56914a <=( (not A234)  and  a56913a );
 a56917a <=( (not A299)  and  A298 );
 a56920a <=( A301  and  A300 );
 a56921a <=( a56920a  and  a56917a );
 a56922a <=( a56921a  and  a56914a );
 a56926a <=( A167  and  (not A169) );
 a56927a <=( A170  and  a56926a );
 a56930a <=( (not A200)  and  (not A166) );
 a56933a <=( (not A233)  and  (not A201) );
 a56934a <=( a56933a  and  a56930a );
 a56935a <=( a56934a  and  a56927a );
 a56939a <=( (not A267)  and  (not A266) );
 a56940a <=( (not A234)  and  a56939a );
 a56943a <=( (not A299)  and  A298 );
 a56946a <=( A302  and  A300 );
 a56947a <=( a56946a  and  a56943a );
 a56948a <=( a56947a  and  a56940a );
 a56952a <=( A167  and  (not A169) );
 a56953a <=( A170  and  a56952a );
 a56956a <=( (not A200)  and  (not A166) );
 a56959a <=( (not A233)  and  (not A201) );
 a56960a <=( a56959a  and  a56956a );
 a56961a <=( a56960a  and  a56953a );
 a56965a <=( (not A266)  and  (not A265) );
 a56966a <=( (not A234)  and  a56965a );
 a56969a <=( (not A299)  and  A298 );
 a56972a <=( A301  and  A300 );
 a56973a <=( a56972a  and  a56969a );
 a56974a <=( a56973a  and  a56966a );
 a56978a <=( A167  and  (not A169) );
 a56979a <=( A170  and  a56978a );
 a56982a <=( (not A200)  and  (not A166) );
 a56985a <=( (not A233)  and  (not A201) );
 a56986a <=( a56985a  and  a56982a );
 a56987a <=( a56986a  and  a56979a );
 a56991a <=( (not A266)  and  (not A265) );
 a56992a <=( (not A234)  and  a56991a );
 a56995a <=( (not A299)  and  A298 );
 a56998a <=( A302  and  A300 );
 a56999a <=( a56998a  and  a56995a );
 a57000a <=( a56999a  and  a56992a );
 a57004a <=( A167  and  (not A169) );
 a57005a <=( A170  and  a57004a );
 a57008a <=( (not A200)  and  (not A166) );
 a57011a <=( A232  and  (not A201) );
 a57012a <=( a57011a  and  a57008a );
 a57013a <=( a57012a  and  a57005a );
 a57017a <=( A235  and  A234 );
 a57018a <=( (not A233)  and  a57017a );
 a57021a <=( (not A266)  and  A265 );
 a57024a <=( A268  and  A267 );
 a57025a <=( a57024a  and  a57021a );
 a57026a <=( a57025a  and  a57018a );
 a57030a <=( A167  and  (not A169) );
 a57031a <=( A170  and  a57030a );
 a57034a <=( (not A200)  and  (not A166) );
 a57037a <=( A232  and  (not A201) );
 a57038a <=( a57037a  and  a57034a );
 a57039a <=( a57038a  and  a57031a );
 a57043a <=( A235  and  A234 );
 a57044a <=( (not A233)  and  a57043a );
 a57047a <=( (not A266)  and  A265 );
 a57050a <=( A269  and  A267 );
 a57051a <=( a57050a  and  a57047a );
 a57052a <=( a57051a  and  a57044a );
 a57056a <=( A167  and  (not A169) );
 a57057a <=( A170  and  a57056a );
 a57060a <=( (not A200)  and  (not A166) );
 a57063a <=( A232  and  (not A201) );
 a57064a <=( a57063a  and  a57060a );
 a57065a <=( a57064a  and  a57057a );
 a57069a <=( A236  and  A234 );
 a57070a <=( (not A233)  and  a57069a );
 a57073a <=( (not A266)  and  A265 );
 a57076a <=( A268  and  A267 );
 a57077a <=( a57076a  and  a57073a );
 a57078a <=( a57077a  and  a57070a );
 a57082a <=( A167  and  (not A169) );
 a57083a <=( A170  and  a57082a );
 a57086a <=( (not A200)  and  (not A166) );
 a57089a <=( A232  and  (not A201) );
 a57090a <=( a57089a  and  a57086a );
 a57091a <=( a57090a  and  a57083a );
 a57095a <=( A236  and  A234 );
 a57096a <=( (not A233)  and  a57095a );
 a57099a <=( (not A266)  and  A265 );
 a57102a <=( A269  and  A267 );
 a57103a <=( a57102a  and  a57099a );
 a57104a <=( a57103a  and  a57096a );
 a57108a <=( A167  and  (not A169) );
 a57109a <=( A170  and  a57108a );
 a57112a <=( (not A200)  and  (not A166) );
 a57115a <=( (not A232)  and  (not A201) );
 a57116a <=( a57115a  and  a57112a );
 a57117a <=( a57116a  and  a57109a );
 a57121a <=( A266  and  A265 );
 a57122a <=( (not A233)  and  a57121a );
 a57125a <=( (not A299)  and  A298 );
 a57128a <=( A301  and  A300 );
 a57129a <=( a57128a  and  a57125a );
 a57130a <=( a57129a  and  a57122a );
 a57134a <=( A167  and  (not A169) );
 a57135a <=( A170  and  a57134a );
 a57138a <=( (not A200)  and  (not A166) );
 a57141a <=( (not A232)  and  (not A201) );
 a57142a <=( a57141a  and  a57138a );
 a57143a <=( a57142a  and  a57135a );
 a57147a <=( A266  and  A265 );
 a57148a <=( (not A233)  and  a57147a );
 a57151a <=( (not A299)  and  A298 );
 a57154a <=( A302  and  A300 );
 a57155a <=( a57154a  and  a57151a );
 a57156a <=( a57155a  and  a57148a );
 a57160a <=( A167  and  (not A169) );
 a57161a <=( A170  and  a57160a );
 a57164a <=( (not A200)  and  (not A166) );
 a57167a <=( (not A232)  and  (not A201) );
 a57168a <=( a57167a  and  a57164a );
 a57169a <=( a57168a  and  a57161a );
 a57173a <=( (not A267)  and  (not A266) );
 a57174a <=( (not A233)  and  a57173a );
 a57177a <=( (not A299)  and  A298 );
 a57180a <=( A301  and  A300 );
 a57181a <=( a57180a  and  a57177a );
 a57182a <=( a57181a  and  a57174a );
 a57186a <=( A167  and  (not A169) );
 a57187a <=( A170  and  a57186a );
 a57190a <=( (not A200)  and  (not A166) );
 a57193a <=( (not A232)  and  (not A201) );
 a57194a <=( a57193a  and  a57190a );
 a57195a <=( a57194a  and  a57187a );
 a57199a <=( (not A267)  and  (not A266) );
 a57200a <=( (not A233)  and  a57199a );
 a57203a <=( (not A299)  and  A298 );
 a57206a <=( A302  and  A300 );
 a57207a <=( a57206a  and  a57203a );
 a57208a <=( a57207a  and  a57200a );
 a57212a <=( A167  and  (not A169) );
 a57213a <=( A170  and  a57212a );
 a57216a <=( (not A200)  and  (not A166) );
 a57219a <=( (not A232)  and  (not A201) );
 a57220a <=( a57219a  and  a57216a );
 a57221a <=( a57220a  and  a57213a );
 a57225a <=( (not A266)  and  (not A265) );
 a57226a <=( (not A233)  and  a57225a );
 a57229a <=( (not A299)  and  A298 );
 a57232a <=( A301  and  A300 );
 a57233a <=( a57232a  and  a57229a );
 a57234a <=( a57233a  and  a57226a );
 a57238a <=( A167  and  (not A169) );
 a57239a <=( A170  and  a57238a );
 a57242a <=( (not A200)  and  (not A166) );
 a57245a <=( (not A232)  and  (not A201) );
 a57246a <=( a57245a  and  a57242a );
 a57247a <=( a57246a  and  a57239a );
 a57251a <=( (not A266)  and  (not A265) );
 a57252a <=( (not A233)  and  a57251a );
 a57255a <=( (not A299)  and  A298 );
 a57258a <=( A302  and  A300 );
 a57259a <=( a57258a  and  a57255a );
 a57260a <=( a57259a  and  a57252a );
 a57264a <=( A167  and  (not A169) );
 a57265a <=( A170  and  a57264a );
 a57268a <=( (not A199)  and  (not A166) );
 a57271a <=( A232  and  (not A200) );
 a57272a <=( a57271a  and  a57268a );
 a57273a <=( a57272a  and  a57265a );
 a57277a <=( (not A267)  and  A265 );
 a57278a <=( A233  and  a57277a );
 a57281a <=( (not A299)  and  A298 );
 a57284a <=( A301  and  A300 );
 a57285a <=( a57284a  and  a57281a );
 a57286a <=( a57285a  and  a57278a );
 a57290a <=( A167  and  (not A169) );
 a57291a <=( A170  and  a57290a );
 a57294a <=( (not A199)  and  (not A166) );
 a57297a <=( A232  and  (not A200) );
 a57298a <=( a57297a  and  a57294a );
 a57299a <=( a57298a  and  a57291a );
 a57303a <=( (not A267)  and  A265 );
 a57304a <=( A233  and  a57303a );
 a57307a <=( (not A299)  and  A298 );
 a57310a <=( A302  and  A300 );
 a57311a <=( a57310a  and  a57307a );
 a57312a <=( a57311a  and  a57304a );
 a57316a <=( A167  and  (not A169) );
 a57317a <=( A170  and  a57316a );
 a57320a <=( (not A199)  and  (not A166) );
 a57323a <=( A232  and  (not A200) );
 a57324a <=( a57323a  and  a57320a );
 a57325a <=( a57324a  and  a57317a );
 a57329a <=( A266  and  A265 );
 a57330a <=( A233  and  a57329a );
 a57333a <=( (not A299)  and  A298 );
 a57336a <=( A301  and  A300 );
 a57337a <=( a57336a  and  a57333a );
 a57338a <=( a57337a  and  a57330a );
 a57342a <=( A167  and  (not A169) );
 a57343a <=( A170  and  a57342a );
 a57346a <=( (not A199)  and  (not A166) );
 a57349a <=( A232  and  (not A200) );
 a57350a <=( a57349a  and  a57346a );
 a57351a <=( a57350a  and  a57343a );
 a57355a <=( A266  and  A265 );
 a57356a <=( A233  and  a57355a );
 a57359a <=( (not A299)  and  A298 );
 a57362a <=( A302  and  A300 );
 a57363a <=( a57362a  and  a57359a );
 a57364a <=( a57363a  and  a57356a );
 a57368a <=( A167  and  (not A169) );
 a57369a <=( A170  and  a57368a );
 a57372a <=( (not A199)  and  (not A166) );
 a57375a <=( A232  and  (not A200) );
 a57376a <=( a57375a  and  a57372a );
 a57377a <=( a57376a  and  a57369a );
 a57381a <=( (not A266)  and  (not A265) );
 a57382a <=( A233  and  a57381a );
 a57385a <=( (not A299)  and  A298 );
 a57388a <=( A301  and  A300 );
 a57389a <=( a57388a  and  a57385a );
 a57390a <=( a57389a  and  a57382a );
 a57394a <=( A167  and  (not A169) );
 a57395a <=( A170  and  a57394a );
 a57398a <=( (not A199)  and  (not A166) );
 a57401a <=( A232  and  (not A200) );
 a57402a <=( a57401a  and  a57398a );
 a57403a <=( a57402a  and  a57395a );
 a57407a <=( (not A266)  and  (not A265) );
 a57408a <=( A233  and  a57407a );
 a57411a <=( (not A299)  and  A298 );
 a57414a <=( A302  and  A300 );
 a57415a <=( a57414a  and  a57411a );
 a57416a <=( a57415a  and  a57408a );
 a57420a <=( A167  and  (not A169) );
 a57421a <=( A170  and  a57420a );
 a57424a <=( (not A199)  and  (not A166) );
 a57427a <=( (not A233)  and  (not A200) );
 a57428a <=( a57427a  and  a57424a );
 a57429a <=( a57428a  and  a57421a );
 a57433a <=( (not A266)  and  (not A236) );
 a57434a <=( (not A235)  and  a57433a );
 a57437a <=( (not A269)  and  (not A268) );
 a57440a <=( A299  and  (not A298) );
 a57441a <=( a57440a  and  a57437a );
 a57442a <=( a57441a  and  a57434a );
 a57446a <=( A167  and  (not A169) );
 a57447a <=( A170  and  a57446a );
 a57450a <=( (not A199)  and  (not A166) );
 a57453a <=( (not A233)  and  (not A200) );
 a57454a <=( a57453a  and  a57450a );
 a57455a <=( a57454a  and  a57447a );
 a57459a <=( A266  and  A265 );
 a57460a <=( (not A234)  and  a57459a );
 a57463a <=( (not A299)  and  A298 );
 a57466a <=( A301  and  A300 );
 a57467a <=( a57466a  and  a57463a );
 a57468a <=( a57467a  and  a57460a );
 a57472a <=( A167  and  (not A169) );
 a57473a <=( A170  and  a57472a );
 a57476a <=( (not A199)  and  (not A166) );
 a57479a <=( (not A233)  and  (not A200) );
 a57480a <=( a57479a  and  a57476a );
 a57481a <=( a57480a  and  a57473a );
 a57485a <=( A266  and  A265 );
 a57486a <=( (not A234)  and  a57485a );
 a57489a <=( (not A299)  and  A298 );
 a57492a <=( A302  and  A300 );
 a57493a <=( a57492a  and  a57489a );
 a57494a <=( a57493a  and  a57486a );
 a57498a <=( A167  and  (not A169) );
 a57499a <=( A170  and  a57498a );
 a57502a <=( (not A199)  and  (not A166) );
 a57505a <=( (not A233)  and  (not A200) );
 a57506a <=( a57505a  and  a57502a );
 a57507a <=( a57506a  and  a57499a );
 a57511a <=( (not A267)  and  (not A266) );
 a57512a <=( (not A234)  and  a57511a );
 a57515a <=( (not A299)  and  A298 );
 a57518a <=( A301  and  A300 );
 a57519a <=( a57518a  and  a57515a );
 a57520a <=( a57519a  and  a57512a );
 a57524a <=( A167  and  (not A169) );
 a57525a <=( A170  and  a57524a );
 a57528a <=( (not A199)  and  (not A166) );
 a57531a <=( (not A233)  and  (not A200) );
 a57532a <=( a57531a  and  a57528a );
 a57533a <=( a57532a  and  a57525a );
 a57537a <=( (not A267)  and  (not A266) );
 a57538a <=( (not A234)  and  a57537a );
 a57541a <=( (not A299)  and  A298 );
 a57544a <=( A302  and  A300 );
 a57545a <=( a57544a  and  a57541a );
 a57546a <=( a57545a  and  a57538a );
 a57550a <=( A167  and  (not A169) );
 a57551a <=( A170  and  a57550a );
 a57554a <=( (not A199)  and  (not A166) );
 a57557a <=( (not A233)  and  (not A200) );
 a57558a <=( a57557a  and  a57554a );
 a57559a <=( a57558a  and  a57551a );
 a57563a <=( (not A266)  and  (not A265) );
 a57564a <=( (not A234)  and  a57563a );
 a57567a <=( (not A299)  and  A298 );
 a57570a <=( A301  and  A300 );
 a57571a <=( a57570a  and  a57567a );
 a57572a <=( a57571a  and  a57564a );
 a57576a <=( A167  and  (not A169) );
 a57577a <=( A170  and  a57576a );
 a57580a <=( (not A199)  and  (not A166) );
 a57583a <=( (not A233)  and  (not A200) );
 a57584a <=( a57583a  and  a57580a );
 a57585a <=( a57584a  and  a57577a );
 a57589a <=( (not A266)  and  (not A265) );
 a57590a <=( (not A234)  and  a57589a );
 a57593a <=( (not A299)  and  A298 );
 a57596a <=( A302  and  A300 );
 a57597a <=( a57596a  and  a57593a );
 a57598a <=( a57597a  and  a57590a );
 a57602a <=( A167  and  (not A169) );
 a57603a <=( A170  and  a57602a );
 a57606a <=( (not A199)  and  (not A166) );
 a57609a <=( A232  and  (not A200) );
 a57610a <=( a57609a  and  a57606a );
 a57611a <=( a57610a  and  a57603a );
 a57615a <=( A235  and  A234 );
 a57616a <=( (not A233)  and  a57615a );
 a57619a <=( (not A266)  and  A265 );
 a57622a <=( A268  and  A267 );
 a57623a <=( a57622a  and  a57619a );
 a57624a <=( a57623a  and  a57616a );
 a57628a <=( A167  and  (not A169) );
 a57629a <=( A170  and  a57628a );
 a57632a <=( (not A199)  and  (not A166) );
 a57635a <=( A232  and  (not A200) );
 a57636a <=( a57635a  and  a57632a );
 a57637a <=( a57636a  and  a57629a );
 a57641a <=( A235  and  A234 );
 a57642a <=( (not A233)  and  a57641a );
 a57645a <=( (not A266)  and  A265 );
 a57648a <=( A269  and  A267 );
 a57649a <=( a57648a  and  a57645a );
 a57650a <=( a57649a  and  a57642a );
 a57654a <=( A167  and  (not A169) );
 a57655a <=( A170  and  a57654a );
 a57658a <=( (not A199)  and  (not A166) );
 a57661a <=( A232  and  (not A200) );
 a57662a <=( a57661a  and  a57658a );
 a57663a <=( a57662a  and  a57655a );
 a57667a <=( A236  and  A234 );
 a57668a <=( (not A233)  and  a57667a );
 a57671a <=( (not A266)  and  A265 );
 a57674a <=( A268  and  A267 );
 a57675a <=( a57674a  and  a57671a );
 a57676a <=( a57675a  and  a57668a );
 a57680a <=( A167  and  (not A169) );
 a57681a <=( A170  and  a57680a );
 a57684a <=( (not A199)  and  (not A166) );
 a57687a <=( A232  and  (not A200) );
 a57688a <=( a57687a  and  a57684a );
 a57689a <=( a57688a  and  a57681a );
 a57693a <=( A236  and  A234 );
 a57694a <=( (not A233)  and  a57693a );
 a57697a <=( (not A266)  and  A265 );
 a57700a <=( A269  and  A267 );
 a57701a <=( a57700a  and  a57697a );
 a57702a <=( a57701a  and  a57694a );
 a57706a <=( A167  and  (not A169) );
 a57707a <=( A170  and  a57706a );
 a57710a <=( (not A199)  and  (not A166) );
 a57713a <=( (not A232)  and  (not A200) );
 a57714a <=( a57713a  and  a57710a );
 a57715a <=( a57714a  and  a57707a );
 a57719a <=( A266  and  A265 );
 a57720a <=( (not A233)  and  a57719a );
 a57723a <=( (not A299)  and  A298 );
 a57726a <=( A301  and  A300 );
 a57727a <=( a57726a  and  a57723a );
 a57728a <=( a57727a  and  a57720a );
 a57732a <=( A167  and  (not A169) );
 a57733a <=( A170  and  a57732a );
 a57736a <=( (not A199)  and  (not A166) );
 a57739a <=( (not A232)  and  (not A200) );
 a57740a <=( a57739a  and  a57736a );
 a57741a <=( a57740a  and  a57733a );
 a57745a <=( A266  and  A265 );
 a57746a <=( (not A233)  and  a57745a );
 a57749a <=( (not A299)  and  A298 );
 a57752a <=( A302  and  A300 );
 a57753a <=( a57752a  and  a57749a );
 a57754a <=( a57753a  and  a57746a );
 a57758a <=( A167  and  (not A169) );
 a57759a <=( A170  and  a57758a );
 a57762a <=( (not A199)  and  (not A166) );
 a57765a <=( (not A232)  and  (not A200) );
 a57766a <=( a57765a  and  a57762a );
 a57767a <=( a57766a  and  a57759a );
 a57771a <=( (not A267)  and  (not A266) );
 a57772a <=( (not A233)  and  a57771a );
 a57775a <=( (not A299)  and  A298 );
 a57778a <=( A301  and  A300 );
 a57779a <=( a57778a  and  a57775a );
 a57780a <=( a57779a  and  a57772a );
 a57784a <=( A167  and  (not A169) );
 a57785a <=( A170  and  a57784a );
 a57788a <=( (not A199)  and  (not A166) );
 a57791a <=( (not A232)  and  (not A200) );
 a57792a <=( a57791a  and  a57788a );
 a57793a <=( a57792a  and  a57785a );
 a57797a <=( (not A267)  and  (not A266) );
 a57798a <=( (not A233)  and  a57797a );
 a57801a <=( (not A299)  and  A298 );
 a57804a <=( A302  and  A300 );
 a57805a <=( a57804a  and  a57801a );
 a57806a <=( a57805a  and  a57798a );
 a57810a <=( A167  and  (not A169) );
 a57811a <=( A170  and  a57810a );
 a57814a <=( (not A199)  and  (not A166) );
 a57817a <=( (not A232)  and  (not A200) );
 a57818a <=( a57817a  and  a57814a );
 a57819a <=( a57818a  and  a57811a );
 a57823a <=( (not A266)  and  (not A265) );
 a57824a <=( (not A233)  and  a57823a );
 a57827a <=( (not A299)  and  A298 );
 a57830a <=( A301  and  A300 );
 a57831a <=( a57830a  and  a57827a );
 a57832a <=( a57831a  and  a57824a );
 a57836a <=( A167  and  (not A169) );
 a57837a <=( A170  and  a57836a );
 a57840a <=( (not A199)  and  (not A166) );
 a57843a <=( (not A232)  and  (not A200) );
 a57844a <=( a57843a  and  a57840a );
 a57845a <=( a57844a  and  a57837a );
 a57849a <=( (not A266)  and  (not A265) );
 a57850a <=( (not A233)  and  a57849a );
 a57853a <=( (not A299)  and  A298 );
 a57856a <=( A302  and  A300 );
 a57857a <=( a57856a  and  a57853a );
 a57858a <=( a57857a  and  a57850a );
 a57862a <=( (not A167)  and  (not A169) );
 a57863a <=( A170  and  a57862a );
 a57866a <=( A199  and  A166 );
 a57869a <=( A232  and  A200 );
 a57870a <=( a57869a  and  a57866a );
 a57871a <=( a57870a  and  a57863a );
 a57875a <=( (not A267)  and  A265 );
 a57876a <=( A233  and  a57875a );
 a57879a <=( (not A299)  and  A298 );
 a57882a <=( A301  and  A300 );
 a57883a <=( a57882a  and  a57879a );
 a57884a <=( a57883a  and  a57876a );
 a57888a <=( (not A167)  and  (not A169) );
 a57889a <=( A170  and  a57888a );
 a57892a <=( A199  and  A166 );
 a57895a <=( A232  and  A200 );
 a57896a <=( a57895a  and  a57892a );
 a57897a <=( a57896a  and  a57889a );
 a57901a <=( (not A267)  and  A265 );
 a57902a <=( A233  and  a57901a );
 a57905a <=( (not A299)  and  A298 );
 a57908a <=( A302  and  A300 );
 a57909a <=( a57908a  and  a57905a );
 a57910a <=( a57909a  and  a57902a );
 a57914a <=( (not A167)  and  (not A169) );
 a57915a <=( A170  and  a57914a );
 a57918a <=( A199  and  A166 );
 a57921a <=( A232  and  A200 );
 a57922a <=( a57921a  and  a57918a );
 a57923a <=( a57922a  and  a57915a );
 a57927a <=( A266  and  A265 );
 a57928a <=( A233  and  a57927a );
 a57931a <=( (not A299)  and  A298 );
 a57934a <=( A301  and  A300 );
 a57935a <=( a57934a  and  a57931a );
 a57936a <=( a57935a  and  a57928a );
 a57940a <=( (not A167)  and  (not A169) );
 a57941a <=( A170  and  a57940a );
 a57944a <=( A199  and  A166 );
 a57947a <=( A232  and  A200 );
 a57948a <=( a57947a  and  a57944a );
 a57949a <=( a57948a  and  a57941a );
 a57953a <=( A266  and  A265 );
 a57954a <=( A233  and  a57953a );
 a57957a <=( (not A299)  and  A298 );
 a57960a <=( A302  and  A300 );
 a57961a <=( a57960a  and  a57957a );
 a57962a <=( a57961a  and  a57954a );
 a57966a <=( (not A167)  and  (not A169) );
 a57967a <=( A170  and  a57966a );
 a57970a <=( A199  and  A166 );
 a57973a <=( A232  and  A200 );
 a57974a <=( a57973a  and  a57970a );
 a57975a <=( a57974a  and  a57967a );
 a57979a <=( (not A266)  and  (not A265) );
 a57980a <=( A233  and  a57979a );
 a57983a <=( (not A299)  and  A298 );
 a57986a <=( A301  and  A300 );
 a57987a <=( a57986a  and  a57983a );
 a57988a <=( a57987a  and  a57980a );
 a57992a <=( (not A167)  and  (not A169) );
 a57993a <=( A170  and  a57992a );
 a57996a <=( A199  and  A166 );
 a57999a <=( A232  and  A200 );
 a58000a <=( a57999a  and  a57996a );
 a58001a <=( a58000a  and  a57993a );
 a58005a <=( (not A266)  and  (not A265) );
 a58006a <=( A233  and  a58005a );
 a58009a <=( (not A299)  and  A298 );
 a58012a <=( A302  and  A300 );
 a58013a <=( a58012a  and  a58009a );
 a58014a <=( a58013a  and  a58006a );
 a58018a <=( (not A167)  and  (not A169) );
 a58019a <=( A170  and  a58018a );
 a58022a <=( A199  and  A166 );
 a58025a <=( (not A233)  and  A200 );
 a58026a <=( a58025a  and  a58022a );
 a58027a <=( a58026a  and  a58019a );
 a58031a <=( (not A266)  and  (not A236) );
 a58032a <=( (not A235)  and  a58031a );
 a58035a <=( (not A269)  and  (not A268) );
 a58038a <=( A299  and  (not A298) );
 a58039a <=( a58038a  and  a58035a );
 a58040a <=( a58039a  and  a58032a );
 a58044a <=( (not A167)  and  (not A169) );
 a58045a <=( A170  and  a58044a );
 a58048a <=( A199  and  A166 );
 a58051a <=( (not A233)  and  A200 );
 a58052a <=( a58051a  and  a58048a );
 a58053a <=( a58052a  and  a58045a );
 a58057a <=( A266  and  A265 );
 a58058a <=( (not A234)  and  a58057a );
 a58061a <=( (not A299)  and  A298 );
 a58064a <=( A301  and  A300 );
 a58065a <=( a58064a  and  a58061a );
 a58066a <=( a58065a  and  a58058a );
 a58070a <=( (not A167)  and  (not A169) );
 a58071a <=( A170  and  a58070a );
 a58074a <=( A199  and  A166 );
 a58077a <=( (not A233)  and  A200 );
 a58078a <=( a58077a  and  a58074a );
 a58079a <=( a58078a  and  a58071a );
 a58083a <=( A266  and  A265 );
 a58084a <=( (not A234)  and  a58083a );
 a58087a <=( (not A299)  and  A298 );
 a58090a <=( A302  and  A300 );
 a58091a <=( a58090a  and  a58087a );
 a58092a <=( a58091a  and  a58084a );
 a58096a <=( (not A167)  and  (not A169) );
 a58097a <=( A170  and  a58096a );
 a58100a <=( A199  and  A166 );
 a58103a <=( (not A233)  and  A200 );
 a58104a <=( a58103a  and  a58100a );
 a58105a <=( a58104a  and  a58097a );
 a58109a <=( (not A267)  and  (not A266) );
 a58110a <=( (not A234)  and  a58109a );
 a58113a <=( (not A299)  and  A298 );
 a58116a <=( A301  and  A300 );
 a58117a <=( a58116a  and  a58113a );
 a58118a <=( a58117a  and  a58110a );
 a58122a <=( (not A167)  and  (not A169) );
 a58123a <=( A170  and  a58122a );
 a58126a <=( A199  and  A166 );
 a58129a <=( (not A233)  and  A200 );
 a58130a <=( a58129a  and  a58126a );
 a58131a <=( a58130a  and  a58123a );
 a58135a <=( (not A267)  and  (not A266) );
 a58136a <=( (not A234)  and  a58135a );
 a58139a <=( (not A299)  and  A298 );
 a58142a <=( A302  and  A300 );
 a58143a <=( a58142a  and  a58139a );
 a58144a <=( a58143a  and  a58136a );
 a58148a <=( (not A167)  and  (not A169) );
 a58149a <=( A170  and  a58148a );
 a58152a <=( A199  and  A166 );
 a58155a <=( (not A233)  and  A200 );
 a58156a <=( a58155a  and  a58152a );
 a58157a <=( a58156a  and  a58149a );
 a58161a <=( (not A266)  and  (not A265) );
 a58162a <=( (not A234)  and  a58161a );
 a58165a <=( (not A299)  and  A298 );
 a58168a <=( A301  and  A300 );
 a58169a <=( a58168a  and  a58165a );
 a58170a <=( a58169a  and  a58162a );
 a58174a <=( (not A167)  and  (not A169) );
 a58175a <=( A170  and  a58174a );
 a58178a <=( A199  and  A166 );
 a58181a <=( (not A233)  and  A200 );
 a58182a <=( a58181a  and  a58178a );
 a58183a <=( a58182a  and  a58175a );
 a58187a <=( (not A266)  and  (not A265) );
 a58188a <=( (not A234)  and  a58187a );
 a58191a <=( (not A299)  and  A298 );
 a58194a <=( A302  and  A300 );
 a58195a <=( a58194a  and  a58191a );
 a58196a <=( a58195a  and  a58188a );
 a58200a <=( (not A167)  and  (not A169) );
 a58201a <=( A170  and  a58200a );
 a58204a <=( A199  and  A166 );
 a58207a <=( A232  and  A200 );
 a58208a <=( a58207a  and  a58204a );
 a58209a <=( a58208a  and  a58201a );
 a58213a <=( A235  and  A234 );
 a58214a <=( (not A233)  and  a58213a );
 a58217a <=( (not A266)  and  A265 );
 a58220a <=( A268  and  A267 );
 a58221a <=( a58220a  and  a58217a );
 a58222a <=( a58221a  and  a58214a );
 a58226a <=( (not A167)  and  (not A169) );
 a58227a <=( A170  and  a58226a );
 a58230a <=( A199  and  A166 );
 a58233a <=( A232  and  A200 );
 a58234a <=( a58233a  and  a58230a );
 a58235a <=( a58234a  and  a58227a );
 a58239a <=( A235  and  A234 );
 a58240a <=( (not A233)  and  a58239a );
 a58243a <=( (not A266)  and  A265 );
 a58246a <=( A269  and  A267 );
 a58247a <=( a58246a  and  a58243a );
 a58248a <=( a58247a  and  a58240a );
 a58252a <=( (not A167)  and  (not A169) );
 a58253a <=( A170  and  a58252a );
 a58256a <=( A199  and  A166 );
 a58259a <=( A232  and  A200 );
 a58260a <=( a58259a  and  a58256a );
 a58261a <=( a58260a  and  a58253a );
 a58265a <=( A236  and  A234 );
 a58266a <=( (not A233)  and  a58265a );
 a58269a <=( (not A266)  and  A265 );
 a58272a <=( A268  and  A267 );
 a58273a <=( a58272a  and  a58269a );
 a58274a <=( a58273a  and  a58266a );
 a58278a <=( (not A167)  and  (not A169) );
 a58279a <=( A170  and  a58278a );
 a58282a <=( A199  and  A166 );
 a58285a <=( A232  and  A200 );
 a58286a <=( a58285a  and  a58282a );
 a58287a <=( a58286a  and  a58279a );
 a58291a <=( A236  and  A234 );
 a58292a <=( (not A233)  and  a58291a );
 a58295a <=( (not A266)  and  A265 );
 a58298a <=( A269  and  A267 );
 a58299a <=( a58298a  and  a58295a );
 a58300a <=( a58299a  and  a58292a );
 a58304a <=( (not A167)  and  (not A169) );
 a58305a <=( A170  and  a58304a );
 a58308a <=( A199  and  A166 );
 a58311a <=( (not A232)  and  A200 );
 a58312a <=( a58311a  and  a58308a );
 a58313a <=( a58312a  and  a58305a );
 a58317a <=( A266  and  A265 );
 a58318a <=( (not A233)  and  a58317a );
 a58321a <=( (not A299)  and  A298 );
 a58324a <=( A301  and  A300 );
 a58325a <=( a58324a  and  a58321a );
 a58326a <=( a58325a  and  a58318a );
 a58330a <=( (not A167)  and  (not A169) );
 a58331a <=( A170  and  a58330a );
 a58334a <=( A199  and  A166 );
 a58337a <=( (not A232)  and  A200 );
 a58338a <=( a58337a  and  a58334a );
 a58339a <=( a58338a  and  a58331a );
 a58343a <=( A266  and  A265 );
 a58344a <=( (not A233)  and  a58343a );
 a58347a <=( (not A299)  and  A298 );
 a58350a <=( A302  and  A300 );
 a58351a <=( a58350a  and  a58347a );
 a58352a <=( a58351a  and  a58344a );
 a58356a <=( (not A167)  and  (not A169) );
 a58357a <=( A170  and  a58356a );
 a58360a <=( A199  and  A166 );
 a58363a <=( (not A232)  and  A200 );
 a58364a <=( a58363a  and  a58360a );
 a58365a <=( a58364a  and  a58357a );
 a58369a <=( (not A267)  and  (not A266) );
 a58370a <=( (not A233)  and  a58369a );
 a58373a <=( (not A299)  and  A298 );
 a58376a <=( A301  and  A300 );
 a58377a <=( a58376a  and  a58373a );
 a58378a <=( a58377a  and  a58370a );
 a58382a <=( (not A167)  and  (not A169) );
 a58383a <=( A170  and  a58382a );
 a58386a <=( A199  and  A166 );
 a58389a <=( (not A232)  and  A200 );
 a58390a <=( a58389a  and  a58386a );
 a58391a <=( a58390a  and  a58383a );
 a58395a <=( (not A267)  and  (not A266) );
 a58396a <=( (not A233)  and  a58395a );
 a58399a <=( (not A299)  and  A298 );
 a58402a <=( A302  and  A300 );
 a58403a <=( a58402a  and  a58399a );
 a58404a <=( a58403a  and  a58396a );
 a58408a <=( (not A167)  and  (not A169) );
 a58409a <=( A170  and  a58408a );
 a58412a <=( A199  and  A166 );
 a58415a <=( (not A232)  and  A200 );
 a58416a <=( a58415a  and  a58412a );
 a58417a <=( a58416a  and  a58409a );
 a58421a <=( (not A266)  and  (not A265) );
 a58422a <=( (not A233)  and  a58421a );
 a58425a <=( (not A299)  and  A298 );
 a58428a <=( A301  and  A300 );
 a58429a <=( a58428a  and  a58425a );
 a58430a <=( a58429a  and  a58422a );
 a58434a <=( (not A167)  and  (not A169) );
 a58435a <=( A170  and  a58434a );
 a58438a <=( A199  and  A166 );
 a58441a <=( (not A232)  and  A200 );
 a58442a <=( a58441a  and  a58438a );
 a58443a <=( a58442a  and  a58435a );
 a58447a <=( (not A266)  and  (not A265) );
 a58448a <=( (not A233)  and  a58447a );
 a58451a <=( (not A299)  and  A298 );
 a58454a <=( A302  and  A300 );
 a58455a <=( a58454a  and  a58451a );
 a58456a <=( a58455a  and  a58448a );
 a58460a <=( (not A167)  and  (not A169) );
 a58461a <=( A170  and  a58460a );
 a58464a <=( (not A200)  and  A166 );
 a58467a <=( (not A203)  and  (not A202) );
 a58468a <=( a58467a  and  a58464a );
 a58469a <=( a58468a  and  a58461a );
 a58473a <=( A265  and  A233 );
 a58474a <=( A232  and  a58473a );
 a58477a <=( (not A269)  and  (not A268) );
 a58480a <=( A299  and  (not A298) );
 a58481a <=( a58480a  and  a58477a );
 a58482a <=( a58481a  and  a58474a );
 a58486a <=( (not A167)  and  (not A169) );
 a58487a <=( A170  and  a58486a );
 a58490a <=( (not A200)  and  A166 );
 a58493a <=( (not A203)  and  (not A202) );
 a58494a <=( a58493a  and  a58490a );
 a58495a <=( a58494a  and  a58487a );
 a58499a <=( (not A236)  and  (not A235) );
 a58500a <=( (not A233)  and  a58499a );
 a58503a <=( A266  and  A265 );
 a58506a <=( A299  and  (not A298) );
 a58507a <=( a58506a  and  a58503a );
 a58508a <=( a58507a  and  a58500a );
 a58512a <=( (not A167)  and  (not A169) );
 a58513a <=( A170  and  a58512a );
 a58516a <=( (not A200)  and  A166 );
 a58519a <=( (not A203)  and  (not A202) );
 a58520a <=( a58519a  and  a58516a );
 a58521a <=( a58520a  and  a58513a );
 a58525a <=( (not A236)  and  (not A235) );
 a58526a <=( (not A233)  and  a58525a );
 a58529a <=( (not A267)  and  (not A266) );
 a58532a <=( A299  and  (not A298) );
 a58533a <=( a58532a  and  a58529a );
 a58534a <=( a58533a  and  a58526a );
 a58538a <=( (not A167)  and  (not A169) );
 a58539a <=( A170  and  a58538a );
 a58542a <=( (not A200)  and  A166 );
 a58545a <=( (not A203)  and  (not A202) );
 a58546a <=( a58545a  and  a58542a );
 a58547a <=( a58546a  and  a58539a );
 a58551a <=( (not A236)  and  (not A235) );
 a58552a <=( (not A233)  and  a58551a );
 a58555a <=( (not A266)  and  (not A265) );
 a58558a <=( A299  and  (not A298) );
 a58559a <=( a58558a  and  a58555a );
 a58560a <=( a58559a  and  a58552a );
 a58564a <=( (not A167)  and  (not A169) );
 a58565a <=( A170  and  a58564a );
 a58568a <=( (not A200)  and  A166 );
 a58571a <=( (not A203)  and  (not A202) );
 a58572a <=( a58571a  and  a58568a );
 a58573a <=( a58572a  and  a58565a );
 a58577a <=( (not A266)  and  (not A234) );
 a58578a <=( (not A233)  and  a58577a );
 a58581a <=( (not A269)  and  (not A268) );
 a58584a <=( A299  and  (not A298) );
 a58585a <=( a58584a  and  a58581a );
 a58586a <=( a58585a  and  a58578a );
 a58590a <=( (not A167)  and  (not A169) );
 a58591a <=( A170  and  a58590a );
 a58594a <=( (not A200)  and  A166 );
 a58597a <=( (not A203)  and  (not A202) );
 a58598a <=( a58597a  and  a58594a );
 a58599a <=( a58598a  and  a58591a );
 a58603a <=( A234  and  (not A233) );
 a58604a <=( A232  and  a58603a );
 a58607a <=( A298  and  A235 );
 a58610a <=( (not A302)  and  (not A301) );
 a58611a <=( a58610a  and  a58607a );
 a58612a <=( a58611a  and  a58604a );
 a58616a <=( (not A167)  and  (not A169) );
 a58617a <=( A170  and  a58616a );
 a58620a <=( (not A200)  and  A166 );
 a58623a <=( (not A203)  and  (not A202) );
 a58624a <=( a58623a  and  a58620a );
 a58625a <=( a58624a  and  a58617a );
 a58629a <=( A234  and  (not A233) );
 a58630a <=( A232  and  a58629a );
 a58633a <=( A298  and  A236 );
 a58636a <=( (not A302)  and  (not A301) );
 a58637a <=( a58636a  and  a58633a );
 a58638a <=( a58637a  and  a58630a );
 a58642a <=( (not A167)  and  (not A169) );
 a58643a <=( A170  and  a58642a );
 a58646a <=( (not A200)  and  A166 );
 a58649a <=( (not A203)  and  (not A202) );
 a58650a <=( a58649a  and  a58646a );
 a58651a <=( a58650a  and  a58643a );
 a58655a <=( (not A266)  and  (not A233) );
 a58656a <=( (not A232)  and  a58655a );
 a58659a <=( (not A269)  and  (not A268) );
 a58662a <=( A299  and  (not A298) );
 a58663a <=( a58662a  and  a58659a );
 a58664a <=( a58663a  and  a58656a );
 a58668a <=( (not A167)  and  (not A169) );
 a58669a <=( A170  and  a58668a );
 a58672a <=( (not A200)  and  A166 );
 a58675a <=( A232  and  (not A201) );
 a58676a <=( a58675a  and  a58672a );
 a58677a <=( a58676a  and  a58669a );
 a58681a <=( (not A267)  and  A265 );
 a58682a <=( A233  and  a58681a );
 a58685a <=( (not A299)  and  A298 );
 a58688a <=( A301  and  A300 );
 a58689a <=( a58688a  and  a58685a );
 a58690a <=( a58689a  and  a58682a );
 a58694a <=( (not A167)  and  (not A169) );
 a58695a <=( A170  and  a58694a );
 a58698a <=( (not A200)  and  A166 );
 a58701a <=( A232  and  (not A201) );
 a58702a <=( a58701a  and  a58698a );
 a58703a <=( a58702a  and  a58695a );
 a58707a <=( (not A267)  and  A265 );
 a58708a <=( A233  and  a58707a );
 a58711a <=( (not A299)  and  A298 );
 a58714a <=( A302  and  A300 );
 a58715a <=( a58714a  and  a58711a );
 a58716a <=( a58715a  and  a58708a );
 a58720a <=( (not A167)  and  (not A169) );
 a58721a <=( A170  and  a58720a );
 a58724a <=( (not A200)  and  A166 );
 a58727a <=( A232  and  (not A201) );
 a58728a <=( a58727a  and  a58724a );
 a58729a <=( a58728a  and  a58721a );
 a58733a <=( A266  and  A265 );
 a58734a <=( A233  and  a58733a );
 a58737a <=( (not A299)  and  A298 );
 a58740a <=( A301  and  A300 );
 a58741a <=( a58740a  and  a58737a );
 a58742a <=( a58741a  and  a58734a );
 a58746a <=( (not A167)  and  (not A169) );
 a58747a <=( A170  and  a58746a );
 a58750a <=( (not A200)  and  A166 );
 a58753a <=( A232  and  (not A201) );
 a58754a <=( a58753a  and  a58750a );
 a58755a <=( a58754a  and  a58747a );
 a58759a <=( A266  and  A265 );
 a58760a <=( A233  and  a58759a );
 a58763a <=( (not A299)  and  A298 );
 a58766a <=( A302  and  A300 );
 a58767a <=( a58766a  and  a58763a );
 a58768a <=( a58767a  and  a58760a );
 a58772a <=( (not A167)  and  (not A169) );
 a58773a <=( A170  and  a58772a );
 a58776a <=( (not A200)  and  A166 );
 a58779a <=( A232  and  (not A201) );
 a58780a <=( a58779a  and  a58776a );
 a58781a <=( a58780a  and  a58773a );
 a58785a <=( (not A266)  and  (not A265) );
 a58786a <=( A233  and  a58785a );
 a58789a <=( (not A299)  and  A298 );
 a58792a <=( A301  and  A300 );
 a58793a <=( a58792a  and  a58789a );
 a58794a <=( a58793a  and  a58786a );
 a58798a <=( (not A167)  and  (not A169) );
 a58799a <=( A170  and  a58798a );
 a58802a <=( (not A200)  and  A166 );
 a58805a <=( A232  and  (not A201) );
 a58806a <=( a58805a  and  a58802a );
 a58807a <=( a58806a  and  a58799a );
 a58811a <=( (not A266)  and  (not A265) );
 a58812a <=( A233  and  a58811a );
 a58815a <=( (not A299)  and  A298 );
 a58818a <=( A302  and  A300 );
 a58819a <=( a58818a  and  a58815a );
 a58820a <=( a58819a  and  a58812a );
 a58824a <=( (not A167)  and  (not A169) );
 a58825a <=( A170  and  a58824a );
 a58828a <=( (not A200)  and  A166 );
 a58831a <=( (not A233)  and  (not A201) );
 a58832a <=( a58831a  and  a58828a );
 a58833a <=( a58832a  and  a58825a );
 a58837a <=( (not A266)  and  (not A236) );
 a58838a <=( (not A235)  and  a58837a );
 a58841a <=( (not A269)  and  (not A268) );
 a58844a <=( A299  and  (not A298) );
 a58845a <=( a58844a  and  a58841a );
 a58846a <=( a58845a  and  a58838a );
 a58850a <=( (not A167)  and  (not A169) );
 a58851a <=( A170  and  a58850a );
 a58854a <=( (not A200)  and  A166 );
 a58857a <=( (not A233)  and  (not A201) );
 a58858a <=( a58857a  and  a58854a );
 a58859a <=( a58858a  and  a58851a );
 a58863a <=( A266  and  A265 );
 a58864a <=( (not A234)  and  a58863a );
 a58867a <=( (not A299)  and  A298 );
 a58870a <=( A301  and  A300 );
 a58871a <=( a58870a  and  a58867a );
 a58872a <=( a58871a  and  a58864a );
 a58876a <=( (not A167)  and  (not A169) );
 a58877a <=( A170  and  a58876a );
 a58880a <=( (not A200)  and  A166 );
 a58883a <=( (not A233)  and  (not A201) );
 a58884a <=( a58883a  and  a58880a );
 a58885a <=( a58884a  and  a58877a );
 a58889a <=( A266  and  A265 );
 a58890a <=( (not A234)  and  a58889a );
 a58893a <=( (not A299)  and  A298 );
 a58896a <=( A302  and  A300 );
 a58897a <=( a58896a  and  a58893a );
 a58898a <=( a58897a  and  a58890a );
 a58902a <=( (not A167)  and  (not A169) );
 a58903a <=( A170  and  a58902a );
 a58906a <=( (not A200)  and  A166 );
 a58909a <=( (not A233)  and  (not A201) );
 a58910a <=( a58909a  and  a58906a );
 a58911a <=( a58910a  and  a58903a );
 a58915a <=( (not A267)  and  (not A266) );
 a58916a <=( (not A234)  and  a58915a );
 a58919a <=( (not A299)  and  A298 );
 a58922a <=( A301  and  A300 );
 a58923a <=( a58922a  and  a58919a );
 a58924a <=( a58923a  and  a58916a );
 a58928a <=( (not A167)  and  (not A169) );
 a58929a <=( A170  and  a58928a );
 a58932a <=( (not A200)  and  A166 );
 a58935a <=( (not A233)  and  (not A201) );
 a58936a <=( a58935a  and  a58932a );
 a58937a <=( a58936a  and  a58929a );
 a58941a <=( (not A267)  and  (not A266) );
 a58942a <=( (not A234)  and  a58941a );
 a58945a <=( (not A299)  and  A298 );
 a58948a <=( A302  and  A300 );
 a58949a <=( a58948a  and  a58945a );
 a58950a <=( a58949a  and  a58942a );
 a58954a <=( (not A167)  and  (not A169) );
 a58955a <=( A170  and  a58954a );
 a58958a <=( (not A200)  and  A166 );
 a58961a <=( (not A233)  and  (not A201) );
 a58962a <=( a58961a  and  a58958a );
 a58963a <=( a58962a  and  a58955a );
 a58967a <=( (not A266)  and  (not A265) );
 a58968a <=( (not A234)  and  a58967a );
 a58971a <=( (not A299)  and  A298 );
 a58974a <=( A301  and  A300 );
 a58975a <=( a58974a  and  a58971a );
 a58976a <=( a58975a  and  a58968a );
 a58980a <=( (not A167)  and  (not A169) );
 a58981a <=( A170  and  a58980a );
 a58984a <=( (not A200)  and  A166 );
 a58987a <=( (not A233)  and  (not A201) );
 a58988a <=( a58987a  and  a58984a );
 a58989a <=( a58988a  and  a58981a );
 a58993a <=( (not A266)  and  (not A265) );
 a58994a <=( (not A234)  and  a58993a );
 a58997a <=( (not A299)  and  A298 );
 a59000a <=( A302  and  A300 );
 a59001a <=( a59000a  and  a58997a );
 a59002a <=( a59001a  and  a58994a );
 a59006a <=( (not A167)  and  (not A169) );
 a59007a <=( A170  and  a59006a );
 a59010a <=( (not A200)  and  A166 );
 a59013a <=( A232  and  (not A201) );
 a59014a <=( a59013a  and  a59010a );
 a59015a <=( a59014a  and  a59007a );
 a59019a <=( A235  and  A234 );
 a59020a <=( (not A233)  and  a59019a );
 a59023a <=( (not A266)  and  A265 );
 a59026a <=( A268  and  A267 );
 a59027a <=( a59026a  and  a59023a );
 a59028a <=( a59027a  and  a59020a );
 a59032a <=( (not A167)  and  (not A169) );
 a59033a <=( A170  and  a59032a );
 a59036a <=( (not A200)  and  A166 );
 a59039a <=( A232  and  (not A201) );
 a59040a <=( a59039a  and  a59036a );
 a59041a <=( a59040a  and  a59033a );
 a59045a <=( A235  and  A234 );
 a59046a <=( (not A233)  and  a59045a );
 a59049a <=( (not A266)  and  A265 );
 a59052a <=( A269  and  A267 );
 a59053a <=( a59052a  and  a59049a );
 a59054a <=( a59053a  and  a59046a );
 a59058a <=( (not A167)  and  (not A169) );
 a59059a <=( A170  and  a59058a );
 a59062a <=( (not A200)  and  A166 );
 a59065a <=( A232  and  (not A201) );
 a59066a <=( a59065a  and  a59062a );
 a59067a <=( a59066a  and  a59059a );
 a59071a <=( A236  and  A234 );
 a59072a <=( (not A233)  and  a59071a );
 a59075a <=( (not A266)  and  A265 );
 a59078a <=( A268  and  A267 );
 a59079a <=( a59078a  and  a59075a );
 a59080a <=( a59079a  and  a59072a );
 a59084a <=( (not A167)  and  (not A169) );
 a59085a <=( A170  and  a59084a );
 a59088a <=( (not A200)  and  A166 );
 a59091a <=( A232  and  (not A201) );
 a59092a <=( a59091a  and  a59088a );
 a59093a <=( a59092a  and  a59085a );
 a59097a <=( A236  and  A234 );
 a59098a <=( (not A233)  and  a59097a );
 a59101a <=( (not A266)  and  A265 );
 a59104a <=( A269  and  A267 );
 a59105a <=( a59104a  and  a59101a );
 a59106a <=( a59105a  and  a59098a );
 a59110a <=( (not A167)  and  (not A169) );
 a59111a <=( A170  and  a59110a );
 a59114a <=( (not A200)  and  A166 );
 a59117a <=( (not A232)  and  (not A201) );
 a59118a <=( a59117a  and  a59114a );
 a59119a <=( a59118a  and  a59111a );
 a59123a <=( A266  and  A265 );
 a59124a <=( (not A233)  and  a59123a );
 a59127a <=( (not A299)  and  A298 );
 a59130a <=( A301  and  A300 );
 a59131a <=( a59130a  and  a59127a );
 a59132a <=( a59131a  and  a59124a );
 a59136a <=( (not A167)  and  (not A169) );
 a59137a <=( A170  and  a59136a );
 a59140a <=( (not A200)  and  A166 );
 a59143a <=( (not A232)  and  (not A201) );
 a59144a <=( a59143a  and  a59140a );
 a59145a <=( a59144a  and  a59137a );
 a59149a <=( A266  and  A265 );
 a59150a <=( (not A233)  and  a59149a );
 a59153a <=( (not A299)  and  A298 );
 a59156a <=( A302  and  A300 );
 a59157a <=( a59156a  and  a59153a );
 a59158a <=( a59157a  and  a59150a );
 a59162a <=( (not A167)  and  (not A169) );
 a59163a <=( A170  and  a59162a );
 a59166a <=( (not A200)  and  A166 );
 a59169a <=( (not A232)  and  (not A201) );
 a59170a <=( a59169a  and  a59166a );
 a59171a <=( a59170a  and  a59163a );
 a59175a <=( (not A267)  and  (not A266) );
 a59176a <=( (not A233)  and  a59175a );
 a59179a <=( (not A299)  and  A298 );
 a59182a <=( A301  and  A300 );
 a59183a <=( a59182a  and  a59179a );
 a59184a <=( a59183a  and  a59176a );
 a59188a <=( (not A167)  and  (not A169) );
 a59189a <=( A170  and  a59188a );
 a59192a <=( (not A200)  and  A166 );
 a59195a <=( (not A232)  and  (not A201) );
 a59196a <=( a59195a  and  a59192a );
 a59197a <=( a59196a  and  a59189a );
 a59201a <=( (not A267)  and  (not A266) );
 a59202a <=( (not A233)  and  a59201a );
 a59205a <=( (not A299)  and  A298 );
 a59208a <=( A302  and  A300 );
 a59209a <=( a59208a  and  a59205a );
 a59210a <=( a59209a  and  a59202a );
 a59214a <=( (not A167)  and  (not A169) );
 a59215a <=( A170  and  a59214a );
 a59218a <=( (not A200)  and  A166 );
 a59221a <=( (not A232)  and  (not A201) );
 a59222a <=( a59221a  and  a59218a );
 a59223a <=( a59222a  and  a59215a );
 a59227a <=( (not A266)  and  (not A265) );
 a59228a <=( (not A233)  and  a59227a );
 a59231a <=( (not A299)  and  A298 );
 a59234a <=( A301  and  A300 );
 a59235a <=( a59234a  and  a59231a );
 a59236a <=( a59235a  and  a59228a );
 a59240a <=( (not A167)  and  (not A169) );
 a59241a <=( A170  and  a59240a );
 a59244a <=( (not A200)  and  A166 );
 a59247a <=( (not A232)  and  (not A201) );
 a59248a <=( a59247a  and  a59244a );
 a59249a <=( a59248a  and  a59241a );
 a59253a <=( (not A266)  and  (not A265) );
 a59254a <=( (not A233)  and  a59253a );
 a59257a <=( (not A299)  and  A298 );
 a59260a <=( A302  and  A300 );
 a59261a <=( a59260a  and  a59257a );
 a59262a <=( a59261a  and  a59254a );
 a59266a <=( (not A167)  and  (not A169) );
 a59267a <=( A170  and  a59266a );
 a59270a <=( (not A199)  and  A166 );
 a59273a <=( A232  and  (not A200) );
 a59274a <=( a59273a  and  a59270a );
 a59275a <=( a59274a  and  a59267a );
 a59279a <=( (not A267)  and  A265 );
 a59280a <=( A233  and  a59279a );
 a59283a <=( (not A299)  and  A298 );
 a59286a <=( A301  and  A300 );
 a59287a <=( a59286a  and  a59283a );
 a59288a <=( a59287a  and  a59280a );
 a59292a <=( (not A167)  and  (not A169) );
 a59293a <=( A170  and  a59292a );
 a59296a <=( (not A199)  and  A166 );
 a59299a <=( A232  and  (not A200) );
 a59300a <=( a59299a  and  a59296a );
 a59301a <=( a59300a  and  a59293a );
 a59305a <=( (not A267)  and  A265 );
 a59306a <=( A233  and  a59305a );
 a59309a <=( (not A299)  and  A298 );
 a59312a <=( A302  and  A300 );
 a59313a <=( a59312a  and  a59309a );
 a59314a <=( a59313a  and  a59306a );
 a59318a <=( (not A167)  and  (not A169) );
 a59319a <=( A170  and  a59318a );
 a59322a <=( (not A199)  and  A166 );
 a59325a <=( A232  and  (not A200) );
 a59326a <=( a59325a  and  a59322a );
 a59327a <=( a59326a  and  a59319a );
 a59331a <=( A266  and  A265 );
 a59332a <=( A233  and  a59331a );
 a59335a <=( (not A299)  and  A298 );
 a59338a <=( A301  and  A300 );
 a59339a <=( a59338a  and  a59335a );
 a59340a <=( a59339a  and  a59332a );
 a59344a <=( (not A167)  and  (not A169) );
 a59345a <=( A170  and  a59344a );
 a59348a <=( (not A199)  and  A166 );
 a59351a <=( A232  and  (not A200) );
 a59352a <=( a59351a  and  a59348a );
 a59353a <=( a59352a  and  a59345a );
 a59357a <=( A266  and  A265 );
 a59358a <=( A233  and  a59357a );
 a59361a <=( (not A299)  and  A298 );
 a59364a <=( A302  and  A300 );
 a59365a <=( a59364a  and  a59361a );
 a59366a <=( a59365a  and  a59358a );
 a59370a <=( (not A167)  and  (not A169) );
 a59371a <=( A170  and  a59370a );
 a59374a <=( (not A199)  and  A166 );
 a59377a <=( A232  and  (not A200) );
 a59378a <=( a59377a  and  a59374a );
 a59379a <=( a59378a  and  a59371a );
 a59383a <=( (not A266)  and  (not A265) );
 a59384a <=( A233  and  a59383a );
 a59387a <=( (not A299)  and  A298 );
 a59390a <=( A301  and  A300 );
 a59391a <=( a59390a  and  a59387a );
 a59392a <=( a59391a  and  a59384a );
 a59396a <=( (not A167)  and  (not A169) );
 a59397a <=( A170  and  a59396a );
 a59400a <=( (not A199)  and  A166 );
 a59403a <=( A232  and  (not A200) );
 a59404a <=( a59403a  and  a59400a );
 a59405a <=( a59404a  and  a59397a );
 a59409a <=( (not A266)  and  (not A265) );
 a59410a <=( A233  and  a59409a );
 a59413a <=( (not A299)  and  A298 );
 a59416a <=( A302  and  A300 );
 a59417a <=( a59416a  and  a59413a );
 a59418a <=( a59417a  and  a59410a );
 a59422a <=( (not A167)  and  (not A169) );
 a59423a <=( A170  and  a59422a );
 a59426a <=( (not A199)  and  A166 );
 a59429a <=( (not A233)  and  (not A200) );
 a59430a <=( a59429a  and  a59426a );
 a59431a <=( a59430a  and  a59423a );
 a59435a <=( (not A266)  and  (not A236) );
 a59436a <=( (not A235)  and  a59435a );
 a59439a <=( (not A269)  and  (not A268) );
 a59442a <=( A299  and  (not A298) );
 a59443a <=( a59442a  and  a59439a );
 a59444a <=( a59443a  and  a59436a );
 a59448a <=( (not A167)  and  (not A169) );
 a59449a <=( A170  and  a59448a );
 a59452a <=( (not A199)  and  A166 );
 a59455a <=( (not A233)  and  (not A200) );
 a59456a <=( a59455a  and  a59452a );
 a59457a <=( a59456a  and  a59449a );
 a59461a <=( A266  and  A265 );
 a59462a <=( (not A234)  and  a59461a );
 a59465a <=( (not A299)  and  A298 );
 a59468a <=( A301  and  A300 );
 a59469a <=( a59468a  and  a59465a );
 a59470a <=( a59469a  and  a59462a );
 a59474a <=( (not A167)  and  (not A169) );
 a59475a <=( A170  and  a59474a );
 a59478a <=( (not A199)  and  A166 );
 a59481a <=( (not A233)  and  (not A200) );
 a59482a <=( a59481a  and  a59478a );
 a59483a <=( a59482a  and  a59475a );
 a59487a <=( A266  and  A265 );
 a59488a <=( (not A234)  and  a59487a );
 a59491a <=( (not A299)  and  A298 );
 a59494a <=( A302  and  A300 );
 a59495a <=( a59494a  and  a59491a );
 a59496a <=( a59495a  and  a59488a );
 a59500a <=( (not A167)  and  (not A169) );
 a59501a <=( A170  and  a59500a );
 a59504a <=( (not A199)  and  A166 );
 a59507a <=( (not A233)  and  (not A200) );
 a59508a <=( a59507a  and  a59504a );
 a59509a <=( a59508a  and  a59501a );
 a59513a <=( (not A267)  and  (not A266) );
 a59514a <=( (not A234)  and  a59513a );
 a59517a <=( (not A299)  and  A298 );
 a59520a <=( A301  and  A300 );
 a59521a <=( a59520a  and  a59517a );
 a59522a <=( a59521a  and  a59514a );
 a59526a <=( (not A167)  and  (not A169) );
 a59527a <=( A170  and  a59526a );
 a59530a <=( (not A199)  and  A166 );
 a59533a <=( (not A233)  and  (not A200) );
 a59534a <=( a59533a  and  a59530a );
 a59535a <=( a59534a  and  a59527a );
 a59539a <=( (not A267)  and  (not A266) );
 a59540a <=( (not A234)  and  a59539a );
 a59543a <=( (not A299)  and  A298 );
 a59546a <=( A302  and  A300 );
 a59547a <=( a59546a  and  a59543a );
 a59548a <=( a59547a  and  a59540a );
 a59552a <=( (not A167)  and  (not A169) );
 a59553a <=( A170  and  a59552a );
 a59556a <=( (not A199)  and  A166 );
 a59559a <=( (not A233)  and  (not A200) );
 a59560a <=( a59559a  and  a59556a );
 a59561a <=( a59560a  and  a59553a );
 a59565a <=( (not A266)  and  (not A265) );
 a59566a <=( (not A234)  and  a59565a );
 a59569a <=( (not A299)  and  A298 );
 a59572a <=( A301  and  A300 );
 a59573a <=( a59572a  and  a59569a );
 a59574a <=( a59573a  and  a59566a );
 a59578a <=( (not A167)  and  (not A169) );
 a59579a <=( A170  and  a59578a );
 a59582a <=( (not A199)  and  A166 );
 a59585a <=( (not A233)  and  (not A200) );
 a59586a <=( a59585a  and  a59582a );
 a59587a <=( a59586a  and  a59579a );
 a59591a <=( (not A266)  and  (not A265) );
 a59592a <=( (not A234)  and  a59591a );
 a59595a <=( (not A299)  and  A298 );
 a59598a <=( A302  and  A300 );
 a59599a <=( a59598a  and  a59595a );
 a59600a <=( a59599a  and  a59592a );
 a59604a <=( (not A167)  and  (not A169) );
 a59605a <=( A170  and  a59604a );
 a59608a <=( (not A199)  and  A166 );
 a59611a <=( A232  and  (not A200) );
 a59612a <=( a59611a  and  a59608a );
 a59613a <=( a59612a  and  a59605a );
 a59617a <=( A235  and  A234 );
 a59618a <=( (not A233)  and  a59617a );
 a59621a <=( (not A266)  and  A265 );
 a59624a <=( A268  and  A267 );
 a59625a <=( a59624a  and  a59621a );
 a59626a <=( a59625a  and  a59618a );
 a59630a <=( (not A167)  and  (not A169) );
 a59631a <=( A170  and  a59630a );
 a59634a <=( (not A199)  and  A166 );
 a59637a <=( A232  and  (not A200) );
 a59638a <=( a59637a  and  a59634a );
 a59639a <=( a59638a  and  a59631a );
 a59643a <=( A235  and  A234 );
 a59644a <=( (not A233)  and  a59643a );
 a59647a <=( (not A266)  and  A265 );
 a59650a <=( A269  and  A267 );
 a59651a <=( a59650a  and  a59647a );
 a59652a <=( a59651a  and  a59644a );
 a59656a <=( (not A167)  and  (not A169) );
 a59657a <=( A170  and  a59656a );
 a59660a <=( (not A199)  and  A166 );
 a59663a <=( A232  and  (not A200) );
 a59664a <=( a59663a  and  a59660a );
 a59665a <=( a59664a  and  a59657a );
 a59669a <=( A236  and  A234 );
 a59670a <=( (not A233)  and  a59669a );
 a59673a <=( (not A266)  and  A265 );
 a59676a <=( A268  and  A267 );
 a59677a <=( a59676a  and  a59673a );
 a59678a <=( a59677a  and  a59670a );
 a59682a <=( (not A167)  and  (not A169) );
 a59683a <=( A170  and  a59682a );
 a59686a <=( (not A199)  and  A166 );
 a59689a <=( A232  and  (not A200) );
 a59690a <=( a59689a  and  a59686a );
 a59691a <=( a59690a  and  a59683a );
 a59695a <=( A236  and  A234 );
 a59696a <=( (not A233)  and  a59695a );
 a59699a <=( (not A266)  and  A265 );
 a59702a <=( A269  and  A267 );
 a59703a <=( a59702a  and  a59699a );
 a59704a <=( a59703a  and  a59696a );
 a59708a <=( (not A167)  and  (not A169) );
 a59709a <=( A170  and  a59708a );
 a59712a <=( (not A199)  and  A166 );
 a59715a <=( (not A232)  and  (not A200) );
 a59716a <=( a59715a  and  a59712a );
 a59717a <=( a59716a  and  a59709a );
 a59721a <=( A266  and  A265 );
 a59722a <=( (not A233)  and  a59721a );
 a59725a <=( (not A299)  and  A298 );
 a59728a <=( A301  and  A300 );
 a59729a <=( a59728a  and  a59725a );
 a59730a <=( a59729a  and  a59722a );
 a59734a <=( (not A167)  and  (not A169) );
 a59735a <=( A170  and  a59734a );
 a59738a <=( (not A199)  and  A166 );
 a59741a <=( (not A232)  and  (not A200) );
 a59742a <=( a59741a  and  a59738a );
 a59743a <=( a59742a  and  a59735a );
 a59747a <=( A266  and  A265 );
 a59748a <=( (not A233)  and  a59747a );
 a59751a <=( (not A299)  and  A298 );
 a59754a <=( A302  and  A300 );
 a59755a <=( a59754a  and  a59751a );
 a59756a <=( a59755a  and  a59748a );
 a59760a <=( (not A167)  and  (not A169) );
 a59761a <=( A170  and  a59760a );
 a59764a <=( (not A199)  and  A166 );
 a59767a <=( (not A232)  and  (not A200) );
 a59768a <=( a59767a  and  a59764a );
 a59769a <=( a59768a  and  a59761a );
 a59773a <=( (not A267)  and  (not A266) );
 a59774a <=( (not A233)  and  a59773a );
 a59777a <=( (not A299)  and  A298 );
 a59780a <=( A301  and  A300 );
 a59781a <=( a59780a  and  a59777a );
 a59782a <=( a59781a  and  a59774a );
 a59786a <=( (not A167)  and  (not A169) );
 a59787a <=( A170  and  a59786a );
 a59790a <=( (not A199)  and  A166 );
 a59793a <=( (not A232)  and  (not A200) );
 a59794a <=( a59793a  and  a59790a );
 a59795a <=( a59794a  and  a59787a );
 a59799a <=( (not A267)  and  (not A266) );
 a59800a <=( (not A233)  and  a59799a );
 a59803a <=( (not A299)  and  A298 );
 a59806a <=( A302  and  A300 );
 a59807a <=( a59806a  and  a59803a );
 a59808a <=( a59807a  and  a59800a );
 a59812a <=( (not A167)  and  (not A169) );
 a59813a <=( A170  and  a59812a );
 a59816a <=( (not A199)  and  A166 );
 a59819a <=( (not A232)  and  (not A200) );
 a59820a <=( a59819a  and  a59816a );
 a59821a <=( a59820a  and  a59813a );
 a59825a <=( (not A266)  and  (not A265) );
 a59826a <=( (not A233)  and  a59825a );
 a59829a <=( (not A299)  and  A298 );
 a59832a <=( A301  and  A300 );
 a59833a <=( a59832a  and  a59829a );
 a59834a <=( a59833a  and  a59826a );
 a59838a <=( (not A167)  and  (not A169) );
 a59839a <=( A170  and  a59838a );
 a59842a <=( (not A199)  and  A166 );
 a59845a <=( (not A232)  and  (not A200) );
 a59846a <=( a59845a  and  a59842a );
 a59847a <=( a59846a  and  a59839a );
 a59851a <=( (not A266)  and  (not A265) );
 a59852a <=( (not A233)  and  a59851a );
 a59855a <=( (not A299)  and  A298 );
 a59858a <=( A302  and  A300 );
 a59859a <=( a59858a  and  a59855a );
 a59860a <=( a59859a  and  a59852a );
 a59864a <=( (not A168)  and  (not A169) );
 a59865a <=( (not A170)  and  a59864a );
 a59868a <=( (not A200)  and  A199 );
 a59871a <=( A202  and  A201 );
 a59872a <=( a59871a  and  a59868a );
 a59873a <=( a59872a  and  a59865a );
 a59877a <=( A265  and  A233 );
 a59878a <=( A232  and  a59877a );
 a59881a <=( (not A269)  and  (not A268) );
 a59884a <=( A299  and  (not A298) );
 a59885a <=( a59884a  and  a59881a );
 a59886a <=( a59885a  and  a59878a );
 a59890a <=( (not A168)  and  (not A169) );
 a59891a <=( (not A170)  and  a59890a );
 a59894a <=( (not A200)  and  A199 );
 a59897a <=( A202  and  A201 );
 a59898a <=( a59897a  and  a59894a );
 a59899a <=( a59898a  and  a59891a );
 a59903a <=( (not A236)  and  (not A235) );
 a59904a <=( (not A233)  and  a59903a );
 a59907a <=( A266  and  A265 );
 a59910a <=( A299  and  (not A298) );
 a59911a <=( a59910a  and  a59907a );
 a59912a <=( a59911a  and  a59904a );
 a59916a <=( (not A168)  and  (not A169) );
 a59917a <=( (not A170)  and  a59916a );
 a59920a <=( (not A200)  and  A199 );
 a59923a <=( A202  and  A201 );
 a59924a <=( a59923a  and  a59920a );
 a59925a <=( a59924a  and  a59917a );
 a59929a <=( (not A236)  and  (not A235) );
 a59930a <=( (not A233)  and  a59929a );
 a59933a <=( (not A267)  and  (not A266) );
 a59936a <=( A299  and  (not A298) );
 a59937a <=( a59936a  and  a59933a );
 a59938a <=( a59937a  and  a59930a );
 a59942a <=( (not A168)  and  (not A169) );
 a59943a <=( (not A170)  and  a59942a );
 a59946a <=( (not A200)  and  A199 );
 a59949a <=( A202  and  A201 );
 a59950a <=( a59949a  and  a59946a );
 a59951a <=( a59950a  and  a59943a );
 a59955a <=( (not A236)  and  (not A235) );
 a59956a <=( (not A233)  and  a59955a );
 a59959a <=( (not A266)  and  (not A265) );
 a59962a <=( A299  and  (not A298) );
 a59963a <=( a59962a  and  a59959a );
 a59964a <=( a59963a  and  a59956a );
 a59968a <=( (not A168)  and  (not A169) );
 a59969a <=( (not A170)  and  a59968a );
 a59972a <=( (not A200)  and  A199 );
 a59975a <=( A202  and  A201 );
 a59976a <=( a59975a  and  a59972a );
 a59977a <=( a59976a  and  a59969a );
 a59981a <=( (not A266)  and  (not A234) );
 a59982a <=( (not A233)  and  a59981a );
 a59985a <=( (not A269)  and  (not A268) );
 a59988a <=( A299  and  (not A298) );
 a59989a <=( a59988a  and  a59985a );
 a59990a <=( a59989a  and  a59982a );
 a59994a <=( (not A168)  and  (not A169) );
 a59995a <=( (not A170)  and  a59994a );
 a59998a <=( (not A200)  and  A199 );
 a60001a <=( A202  and  A201 );
 a60002a <=( a60001a  and  a59998a );
 a60003a <=( a60002a  and  a59995a );
 a60007a <=( A234  and  (not A233) );
 a60008a <=( A232  and  a60007a );
 a60011a <=( A298  and  A235 );
 a60014a <=( (not A302)  and  (not A301) );
 a60015a <=( a60014a  and  a60011a );
 a60016a <=( a60015a  and  a60008a );
 a60020a <=( (not A168)  and  (not A169) );
 a60021a <=( (not A170)  and  a60020a );
 a60024a <=( (not A200)  and  A199 );
 a60027a <=( A202  and  A201 );
 a60028a <=( a60027a  and  a60024a );
 a60029a <=( a60028a  and  a60021a );
 a60033a <=( A234  and  (not A233) );
 a60034a <=( A232  and  a60033a );
 a60037a <=( A298  and  A236 );
 a60040a <=( (not A302)  and  (not A301) );
 a60041a <=( a60040a  and  a60037a );
 a60042a <=( a60041a  and  a60034a );
 a60046a <=( (not A168)  and  (not A169) );
 a60047a <=( (not A170)  and  a60046a );
 a60050a <=( (not A200)  and  A199 );
 a60053a <=( A202  and  A201 );
 a60054a <=( a60053a  and  a60050a );
 a60055a <=( a60054a  and  a60047a );
 a60059a <=( (not A266)  and  (not A233) );
 a60060a <=( (not A232)  and  a60059a );
 a60063a <=( (not A269)  and  (not A268) );
 a60066a <=( A299  and  (not A298) );
 a60067a <=( a60066a  and  a60063a );
 a60068a <=( a60067a  and  a60060a );
 a60072a <=( (not A168)  and  (not A169) );
 a60073a <=( (not A170)  and  a60072a );
 a60076a <=( (not A200)  and  A199 );
 a60079a <=( A203  and  A201 );
 a60080a <=( a60079a  and  a60076a );
 a60081a <=( a60080a  and  a60073a );
 a60085a <=( A265  and  A233 );
 a60086a <=( A232  and  a60085a );
 a60089a <=( (not A269)  and  (not A268) );
 a60092a <=( A299  and  (not A298) );
 a60093a <=( a60092a  and  a60089a );
 a60094a <=( a60093a  and  a60086a );
 a60098a <=( (not A168)  and  (not A169) );
 a60099a <=( (not A170)  and  a60098a );
 a60102a <=( (not A200)  and  A199 );
 a60105a <=( A203  and  A201 );
 a60106a <=( a60105a  and  a60102a );
 a60107a <=( a60106a  and  a60099a );
 a60111a <=( (not A236)  and  (not A235) );
 a60112a <=( (not A233)  and  a60111a );
 a60115a <=( A266  and  A265 );
 a60118a <=( A299  and  (not A298) );
 a60119a <=( a60118a  and  a60115a );
 a60120a <=( a60119a  and  a60112a );
 a60124a <=( (not A168)  and  (not A169) );
 a60125a <=( (not A170)  and  a60124a );
 a60128a <=( (not A200)  and  A199 );
 a60131a <=( A203  and  A201 );
 a60132a <=( a60131a  and  a60128a );
 a60133a <=( a60132a  and  a60125a );
 a60137a <=( (not A236)  and  (not A235) );
 a60138a <=( (not A233)  and  a60137a );
 a60141a <=( (not A267)  and  (not A266) );
 a60144a <=( A299  and  (not A298) );
 a60145a <=( a60144a  and  a60141a );
 a60146a <=( a60145a  and  a60138a );
 a60150a <=( (not A168)  and  (not A169) );
 a60151a <=( (not A170)  and  a60150a );
 a60154a <=( (not A200)  and  A199 );
 a60157a <=( A203  and  A201 );
 a60158a <=( a60157a  and  a60154a );
 a60159a <=( a60158a  and  a60151a );
 a60163a <=( (not A236)  and  (not A235) );
 a60164a <=( (not A233)  and  a60163a );
 a60167a <=( (not A266)  and  (not A265) );
 a60170a <=( A299  and  (not A298) );
 a60171a <=( a60170a  and  a60167a );
 a60172a <=( a60171a  and  a60164a );
 a60176a <=( (not A168)  and  (not A169) );
 a60177a <=( (not A170)  and  a60176a );
 a60180a <=( (not A200)  and  A199 );
 a60183a <=( A203  and  A201 );
 a60184a <=( a60183a  and  a60180a );
 a60185a <=( a60184a  and  a60177a );
 a60189a <=( (not A266)  and  (not A234) );
 a60190a <=( (not A233)  and  a60189a );
 a60193a <=( (not A269)  and  (not A268) );
 a60196a <=( A299  and  (not A298) );
 a60197a <=( a60196a  and  a60193a );
 a60198a <=( a60197a  and  a60190a );
 a60202a <=( (not A168)  and  (not A169) );
 a60203a <=( (not A170)  and  a60202a );
 a60206a <=( (not A200)  and  A199 );
 a60209a <=( A203  and  A201 );
 a60210a <=( a60209a  and  a60206a );
 a60211a <=( a60210a  and  a60203a );
 a60215a <=( A234  and  (not A233) );
 a60216a <=( A232  and  a60215a );
 a60219a <=( A298  and  A235 );
 a60222a <=( (not A302)  and  (not A301) );
 a60223a <=( a60222a  and  a60219a );
 a60224a <=( a60223a  and  a60216a );
 a60228a <=( (not A168)  and  (not A169) );
 a60229a <=( (not A170)  and  a60228a );
 a60232a <=( (not A200)  and  A199 );
 a60235a <=( A203  and  A201 );
 a60236a <=( a60235a  and  a60232a );
 a60237a <=( a60236a  and  a60229a );
 a60241a <=( A234  and  (not A233) );
 a60242a <=( A232  and  a60241a );
 a60245a <=( A298  and  A236 );
 a60248a <=( (not A302)  and  (not A301) );
 a60249a <=( a60248a  and  a60245a );
 a60250a <=( a60249a  and  a60242a );
 a60254a <=( (not A168)  and  (not A169) );
 a60255a <=( (not A170)  and  a60254a );
 a60258a <=( (not A200)  and  A199 );
 a60261a <=( A203  and  A201 );
 a60262a <=( a60261a  and  a60258a );
 a60263a <=( a60262a  and  a60255a );
 a60267a <=( (not A266)  and  (not A233) );
 a60268a <=( (not A232)  and  a60267a );
 a60271a <=( (not A269)  and  (not A268) );
 a60274a <=( A299  and  (not A298) );
 a60275a <=( a60274a  and  a60271a );
 a60276a <=( a60275a  and  a60268a );
 a60280a <=( (not A200)  and  A166 );
 a60281a <=( A168  and  a60280a );
 a60284a <=( (not A203)  and  (not A202) );
 a60287a <=( (not A235)  and  (not A233) );
 a60288a <=( a60287a  and  a60284a );
 a60289a <=( a60288a  and  a60281a );
 a60292a <=( (not A266)  and  (not A236) );
 a60295a <=( (not A269)  and  (not A268) );
 a60296a <=( a60295a  and  a60292a );
 a60299a <=( (not A299)  and  A298 );
 a60302a <=( A301  and  A300 );
 a60303a <=( a60302a  and  a60299a );
 a60304a <=( a60303a  and  a60296a );
 a60308a <=( (not A200)  and  A166 );
 a60309a <=( A168  and  a60308a );
 a60312a <=( (not A203)  and  (not A202) );
 a60315a <=( (not A235)  and  (not A233) );
 a60316a <=( a60315a  and  a60312a );
 a60317a <=( a60316a  and  a60309a );
 a60320a <=( (not A266)  and  (not A236) );
 a60323a <=( (not A269)  and  (not A268) );
 a60324a <=( a60323a  and  a60320a );
 a60327a <=( (not A299)  and  A298 );
 a60330a <=( A302  and  A300 );
 a60331a <=( a60330a  and  a60327a );
 a60332a <=( a60331a  and  a60324a );
 a60336a <=( (not A200)  and  A167 );
 a60337a <=( A168  and  a60336a );
 a60340a <=( (not A203)  and  (not A202) );
 a60343a <=( (not A235)  and  (not A233) );
 a60344a <=( a60343a  and  a60340a );
 a60345a <=( a60344a  and  a60337a );
 a60348a <=( (not A266)  and  (not A236) );
 a60351a <=( (not A269)  and  (not A268) );
 a60352a <=( a60351a  and  a60348a );
 a60355a <=( (not A299)  and  A298 );
 a60358a <=( A301  and  A300 );
 a60359a <=( a60358a  and  a60355a );
 a60360a <=( a60359a  and  a60352a );
 a60364a <=( (not A200)  and  A167 );
 a60365a <=( A168  and  a60364a );
 a60368a <=( (not A203)  and  (not A202) );
 a60371a <=( (not A235)  and  (not A233) );
 a60372a <=( a60371a  and  a60368a );
 a60373a <=( a60372a  and  a60365a );
 a60376a <=( (not A266)  and  (not A236) );
 a60379a <=( (not A269)  and  (not A268) );
 a60380a <=( a60379a  and  a60376a );
 a60383a <=( (not A299)  and  A298 );
 a60386a <=( A302  and  A300 );
 a60387a <=( a60386a  and  a60383a );
 a60388a <=( a60387a  and  a60380a );
 a60392a <=( (not A166)  and  (not A167) );
 a60393a <=( A170  and  a60392a );
 a60396a <=( A200  and  (not A199) );
 a60399a <=( (not A235)  and  (not A233) );
 a60400a <=( a60399a  and  a60396a );
 a60401a <=( a60400a  and  a60393a );
 a60404a <=( (not A266)  and  (not A236) );
 a60407a <=( (not A269)  and  (not A268) );
 a60408a <=( a60407a  and  a60404a );
 a60411a <=( (not A299)  and  A298 );
 a60414a <=( A301  and  A300 );
 a60415a <=( a60414a  and  a60411a );
 a60416a <=( a60415a  and  a60408a );
 a60420a <=( (not A166)  and  (not A167) );
 a60421a <=( A170  and  a60420a );
 a60424a <=( A200  and  (not A199) );
 a60427a <=( (not A235)  and  (not A233) );
 a60428a <=( a60427a  and  a60424a );
 a60429a <=( a60428a  and  a60421a );
 a60432a <=( (not A266)  and  (not A236) );
 a60435a <=( (not A269)  and  (not A268) );
 a60436a <=( a60435a  and  a60432a );
 a60439a <=( (not A299)  and  A298 );
 a60442a <=( A302  and  A300 );
 a60443a <=( a60442a  and  a60439a );
 a60444a <=( a60443a  and  a60436a );
 a60448a <=( (not A166)  and  (not A167) );
 a60449a <=( A170  and  a60448a );
 a60452a <=( (not A200)  and  A199 );
 a60455a <=( A202  and  A201 );
 a60456a <=( a60455a  and  a60452a );
 a60457a <=( a60456a  and  a60449a );
 a60460a <=( A233  and  A232 );
 a60463a <=( (not A267)  and  A265 );
 a60464a <=( a60463a  and  a60460a );
 a60467a <=( (not A299)  and  A298 );
 a60470a <=( A301  and  A300 );
 a60471a <=( a60470a  and  a60467a );
 a60472a <=( a60471a  and  a60464a );
 a60476a <=( (not A166)  and  (not A167) );
 a60477a <=( A170  and  a60476a );
 a60480a <=( (not A200)  and  A199 );
 a60483a <=( A202  and  A201 );
 a60484a <=( a60483a  and  a60480a );
 a60485a <=( a60484a  and  a60477a );
 a60488a <=( A233  and  A232 );
 a60491a <=( (not A267)  and  A265 );
 a60492a <=( a60491a  and  a60488a );
 a60495a <=( (not A299)  and  A298 );
 a60498a <=( A302  and  A300 );
 a60499a <=( a60498a  and  a60495a );
 a60500a <=( a60499a  and  a60492a );
 a60504a <=( (not A166)  and  (not A167) );
 a60505a <=( A170  and  a60504a );
 a60508a <=( (not A200)  and  A199 );
 a60511a <=( A202  and  A201 );
 a60512a <=( a60511a  and  a60508a );
 a60513a <=( a60512a  and  a60505a );
 a60516a <=( A233  and  A232 );
 a60519a <=( A266  and  A265 );
 a60520a <=( a60519a  and  a60516a );
 a60523a <=( (not A299)  and  A298 );
 a60526a <=( A301  and  A300 );
 a60527a <=( a60526a  and  a60523a );
 a60528a <=( a60527a  and  a60520a );
 a60532a <=( (not A166)  and  (not A167) );
 a60533a <=( A170  and  a60532a );
 a60536a <=( (not A200)  and  A199 );
 a60539a <=( A202  and  A201 );
 a60540a <=( a60539a  and  a60536a );
 a60541a <=( a60540a  and  a60533a );
 a60544a <=( A233  and  A232 );
 a60547a <=( A266  and  A265 );
 a60548a <=( a60547a  and  a60544a );
 a60551a <=( (not A299)  and  A298 );
 a60554a <=( A302  and  A300 );
 a60555a <=( a60554a  and  a60551a );
 a60556a <=( a60555a  and  a60548a );
 a60560a <=( (not A166)  and  (not A167) );
 a60561a <=( A170  and  a60560a );
 a60564a <=( (not A200)  and  A199 );
 a60567a <=( A202  and  A201 );
 a60568a <=( a60567a  and  a60564a );
 a60569a <=( a60568a  and  a60561a );
 a60572a <=( A233  and  A232 );
 a60575a <=( (not A266)  and  (not A265) );
 a60576a <=( a60575a  and  a60572a );
 a60579a <=( (not A299)  and  A298 );
 a60582a <=( A301  and  A300 );
 a60583a <=( a60582a  and  a60579a );
 a60584a <=( a60583a  and  a60576a );
 a60588a <=( (not A166)  and  (not A167) );
 a60589a <=( A170  and  a60588a );
 a60592a <=( (not A200)  and  A199 );
 a60595a <=( A202  and  A201 );
 a60596a <=( a60595a  and  a60592a );
 a60597a <=( a60596a  and  a60589a );
 a60600a <=( A233  and  A232 );
 a60603a <=( (not A266)  and  (not A265) );
 a60604a <=( a60603a  and  a60600a );
 a60607a <=( (not A299)  and  A298 );
 a60610a <=( A302  and  A300 );
 a60611a <=( a60610a  and  a60607a );
 a60612a <=( a60611a  and  a60604a );
 a60616a <=( (not A166)  and  (not A167) );
 a60617a <=( A170  and  a60616a );
 a60620a <=( (not A200)  and  A199 );
 a60623a <=( A202  and  A201 );
 a60624a <=( a60623a  and  a60620a );
 a60625a <=( a60624a  and  a60617a );
 a60628a <=( (not A235)  and  (not A233) );
 a60631a <=( (not A266)  and  (not A236) );
 a60632a <=( a60631a  and  a60628a );
 a60635a <=( (not A269)  and  (not A268) );
 a60638a <=( A299  and  (not A298) );
 a60639a <=( a60638a  and  a60635a );
 a60640a <=( a60639a  and  a60632a );
 a60644a <=( (not A166)  and  (not A167) );
 a60645a <=( A170  and  a60644a );
 a60648a <=( (not A200)  and  A199 );
 a60651a <=( A202  and  A201 );
 a60652a <=( a60651a  and  a60648a );
 a60653a <=( a60652a  and  a60645a );
 a60656a <=( (not A234)  and  (not A233) );
 a60659a <=( A266  and  A265 );
 a60660a <=( a60659a  and  a60656a );
 a60663a <=( (not A299)  and  A298 );
 a60666a <=( A301  and  A300 );
 a60667a <=( a60666a  and  a60663a );
 a60668a <=( a60667a  and  a60660a );
 a60672a <=( (not A166)  and  (not A167) );
 a60673a <=( A170  and  a60672a );
 a60676a <=( (not A200)  and  A199 );
 a60679a <=( A202  and  A201 );
 a60680a <=( a60679a  and  a60676a );
 a60681a <=( a60680a  and  a60673a );
 a60684a <=( (not A234)  and  (not A233) );
 a60687a <=( A266  and  A265 );
 a60688a <=( a60687a  and  a60684a );
 a60691a <=( (not A299)  and  A298 );
 a60694a <=( A302  and  A300 );
 a60695a <=( a60694a  and  a60691a );
 a60696a <=( a60695a  and  a60688a );
 a60700a <=( (not A166)  and  (not A167) );
 a60701a <=( A170  and  a60700a );
 a60704a <=( (not A200)  and  A199 );
 a60707a <=( A202  and  A201 );
 a60708a <=( a60707a  and  a60704a );
 a60709a <=( a60708a  and  a60701a );
 a60712a <=( (not A234)  and  (not A233) );
 a60715a <=( (not A267)  and  (not A266) );
 a60716a <=( a60715a  and  a60712a );
 a60719a <=( (not A299)  and  A298 );
 a60722a <=( A301  and  A300 );
 a60723a <=( a60722a  and  a60719a );
 a60724a <=( a60723a  and  a60716a );
 a60728a <=( (not A166)  and  (not A167) );
 a60729a <=( A170  and  a60728a );
 a60732a <=( (not A200)  and  A199 );
 a60735a <=( A202  and  A201 );
 a60736a <=( a60735a  and  a60732a );
 a60737a <=( a60736a  and  a60729a );
 a60740a <=( (not A234)  and  (not A233) );
 a60743a <=( (not A267)  and  (not A266) );
 a60744a <=( a60743a  and  a60740a );
 a60747a <=( (not A299)  and  A298 );
 a60750a <=( A302  and  A300 );
 a60751a <=( a60750a  and  a60747a );
 a60752a <=( a60751a  and  a60744a );
 a60756a <=( (not A166)  and  (not A167) );
 a60757a <=( A170  and  a60756a );
 a60760a <=( (not A200)  and  A199 );
 a60763a <=( A202  and  A201 );
 a60764a <=( a60763a  and  a60760a );
 a60765a <=( a60764a  and  a60757a );
 a60768a <=( (not A234)  and  (not A233) );
 a60771a <=( (not A266)  and  (not A265) );
 a60772a <=( a60771a  and  a60768a );
 a60775a <=( (not A299)  and  A298 );
 a60778a <=( A301  and  A300 );
 a60779a <=( a60778a  and  a60775a );
 a60780a <=( a60779a  and  a60772a );
 a60784a <=( (not A166)  and  (not A167) );
 a60785a <=( A170  and  a60784a );
 a60788a <=( (not A200)  and  A199 );
 a60791a <=( A202  and  A201 );
 a60792a <=( a60791a  and  a60788a );
 a60793a <=( a60792a  and  a60785a );
 a60796a <=( (not A234)  and  (not A233) );
 a60799a <=( (not A266)  and  (not A265) );
 a60800a <=( a60799a  and  a60796a );
 a60803a <=( (not A299)  and  A298 );
 a60806a <=( A302  and  A300 );
 a60807a <=( a60806a  and  a60803a );
 a60808a <=( a60807a  and  a60800a );
 a60812a <=( (not A166)  and  (not A167) );
 a60813a <=( A170  and  a60812a );
 a60816a <=( (not A200)  and  A199 );
 a60819a <=( A202  and  A201 );
 a60820a <=( a60819a  and  a60816a );
 a60821a <=( a60820a  and  a60813a );
 a60824a <=( (not A233)  and  A232 );
 a60827a <=( A235  and  A234 );
 a60828a <=( a60827a  and  a60824a );
 a60831a <=( (not A266)  and  A265 );
 a60834a <=( A268  and  A267 );
 a60835a <=( a60834a  and  a60831a );
 a60836a <=( a60835a  and  a60828a );
 a60840a <=( (not A166)  and  (not A167) );
 a60841a <=( A170  and  a60840a );
 a60844a <=( (not A200)  and  A199 );
 a60847a <=( A202  and  A201 );
 a60848a <=( a60847a  and  a60844a );
 a60849a <=( a60848a  and  a60841a );
 a60852a <=( (not A233)  and  A232 );
 a60855a <=( A235  and  A234 );
 a60856a <=( a60855a  and  a60852a );
 a60859a <=( (not A266)  and  A265 );
 a60862a <=( A269  and  A267 );
 a60863a <=( a60862a  and  a60859a );
 a60864a <=( a60863a  and  a60856a );
 a60868a <=( (not A166)  and  (not A167) );
 a60869a <=( A170  and  a60868a );
 a60872a <=( (not A200)  and  A199 );
 a60875a <=( A202  and  A201 );
 a60876a <=( a60875a  and  a60872a );
 a60877a <=( a60876a  and  a60869a );
 a60880a <=( (not A233)  and  A232 );
 a60883a <=( A236  and  A234 );
 a60884a <=( a60883a  and  a60880a );
 a60887a <=( (not A266)  and  A265 );
 a60890a <=( A268  and  A267 );
 a60891a <=( a60890a  and  a60887a );
 a60892a <=( a60891a  and  a60884a );
 a60896a <=( (not A166)  and  (not A167) );
 a60897a <=( A170  and  a60896a );
 a60900a <=( (not A200)  and  A199 );
 a60903a <=( A202  and  A201 );
 a60904a <=( a60903a  and  a60900a );
 a60905a <=( a60904a  and  a60897a );
 a60908a <=( (not A233)  and  A232 );
 a60911a <=( A236  and  A234 );
 a60912a <=( a60911a  and  a60908a );
 a60915a <=( (not A266)  and  A265 );
 a60918a <=( A269  and  A267 );
 a60919a <=( a60918a  and  a60915a );
 a60920a <=( a60919a  and  a60912a );
 a60924a <=( (not A166)  and  (not A167) );
 a60925a <=( A170  and  a60924a );
 a60928a <=( (not A200)  and  A199 );
 a60931a <=( A202  and  A201 );
 a60932a <=( a60931a  and  a60928a );
 a60933a <=( a60932a  and  a60925a );
 a60936a <=( (not A233)  and  (not A232) );
 a60939a <=( A266  and  A265 );
 a60940a <=( a60939a  and  a60936a );
 a60943a <=( (not A299)  and  A298 );
 a60946a <=( A301  and  A300 );
 a60947a <=( a60946a  and  a60943a );
 a60948a <=( a60947a  and  a60940a );
 a60952a <=( (not A166)  and  (not A167) );
 a60953a <=( A170  and  a60952a );
 a60956a <=( (not A200)  and  A199 );
 a60959a <=( A202  and  A201 );
 a60960a <=( a60959a  and  a60956a );
 a60961a <=( a60960a  and  a60953a );
 a60964a <=( (not A233)  and  (not A232) );
 a60967a <=( A266  and  A265 );
 a60968a <=( a60967a  and  a60964a );
 a60971a <=( (not A299)  and  A298 );
 a60974a <=( A302  and  A300 );
 a60975a <=( a60974a  and  a60971a );
 a60976a <=( a60975a  and  a60968a );
 a60980a <=( (not A166)  and  (not A167) );
 a60981a <=( A170  and  a60980a );
 a60984a <=( (not A200)  and  A199 );
 a60987a <=( A202  and  A201 );
 a60988a <=( a60987a  and  a60984a );
 a60989a <=( a60988a  and  a60981a );
 a60992a <=( (not A233)  and  (not A232) );
 a60995a <=( (not A267)  and  (not A266) );
 a60996a <=( a60995a  and  a60992a );
 a60999a <=( (not A299)  and  A298 );
 a61002a <=( A301  and  A300 );
 a61003a <=( a61002a  and  a60999a );
 a61004a <=( a61003a  and  a60996a );
 a61008a <=( (not A166)  and  (not A167) );
 a61009a <=( A170  and  a61008a );
 a61012a <=( (not A200)  and  A199 );
 a61015a <=( A202  and  A201 );
 a61016a <=( a61015a  and  a61012a );
 a61017a <=( a61016a  and  a61009a );
 a61020a <=( (not A233)  and  (not A232) );
 a61023a <=( (not A267)  and  (not A266) );
 a61024a <=( a61023a  and  a61020a );
 a61027a <=( (not A299)  and  A298 );
 a61030a <=( A302  and  A300 );
 a61031a <=( a61030a  and  a61027a );
 a61032a <=( a61031a  and  a61024a );
 a61036a <=( (not A166)  and  (not A167) );
 a61037a <=( A170  and  a61036a );
 a61040a <=( (not A200)  and  A199 );
 a61043a <=( A202  and  A201 );
 a61044a <=( a61043a  and  a61040a );
 a61045a <=( a61044a  and  a61037a );
 a61048a <=( (not A233)  and  (not A232) );
 a61051a <=( (not A266)  and  (not A265) );
 a61052a <=( a61051a  and  a61048a );
 a61055a <=( (not A299)  and  A298 );
 a61058a <=( A301  and  A300 );
 a61059a <=( a61058a  and  a61055a );
 a61060a <=( a61059a  and  a61052a );
 a61064a <=( (not A166)  and  (not A167) );
 a61065a <=( A170  and  a61064a );
 a61068a <=( (not A200)  and  A199 );
 a61071a <=( A202  and  A201 );
 a61072a <=( a61071a  and  a61068a );
 a61073a <=( a61072a  and  a61065a );
 a61076a <=( (not A233)  and  (not A232) );
 a61079a <=( (not A266)  and  (not A265) );
 a61080a <=( a61079a  and  a61076a );
 a61083a <=( (not A299)  and  A298 );
 a61086a <=( A302  and  A300 );
 a61087a <=( a61086a  and  a61083a );
 a61088a <=( a61087a  and  a61080a );
 a61092a <=( (not A166)  and  (not A167) );
 a61093a <=( A170  and  a61092a );
 a61096a <=( (not A200)  and  A199 );
 a61099a <=( A203  and  A201 );
 a61100a <=( a61099a  and  a61096a );
 a61101a <=( a61100a  and  a61093a );
 a61104a <=( A233  and  A232 );
 a61107a <=( (not A267)  and  A265 );
 a61108a <=( a61107a  and  a61104a );
 a61111a <=( (not A299)  and  A298 );
 a61114a <=( A301  and  A300 );
 a61115a <=( a61114a  and  a61111a );
 a61116a <=( a61115a  and  a61108a );
 a61120a <=( (not A166)  and  (not A167) );
 a61121a <=( A170  and  a61120a );
 a61124a <=( (not A200)  and  A199 );
 a61127a <=( A203  and  A201 );
 a61128a <=( a61127a  and  a61124a );
 a61129a <=( a61128a  and  a61121a );
 a61132a <=( A233  and  A232 );
 a61135a <=( (not A267)  and  A265 );
 a61136a <=( a61135a  and  a61132a );
 a61139a <=( (not A299)  and  A298 );
 a61142a <=( A302  and  A300 );
 a61143a <=( a61142a  and  a61139a );
 a61144a <=( a61143a  and  a61136a );
 a61148a <=( (not A166)  and  (not A167) );
 a61149a <=( A170  and  a61148a );
 a61152a <=( (not A200)  and  A199 );
 a61155a <=( A203  and  A201 );
 a61156a <=( a61155a  and  a61152a );
 a61157a <=( a61156a  and  a61149a );
 a61160a <=( A233  and  A232 );
 a61163a <=( A266  and  A265 );
 a61164a <=( a61163a  and  a61160a );
 a61167a <=( (not A299)  and  A298 );
 a61170a <=( A301  and  A300 );
 a61171a <=( a61170a  and  a61167a );
 a61172a <=( a61171a  and  a61164a );
 a61176a <=( (not A166)  and  (not A167) );
 a61177a <=( A170  and  a61176a );
 a61180a <=( (not A200)  and  A199 );
 a61183a <=( A203  and  A201 );
 a61184a <=( a61183a  and  a61180a );
 a61185a <=( a61184a  and  a61177a );
 a61188a <=( A233  and  A232 );
 a61191a <=( A266  and  A265 );
 a61192a <=( a61191a  and  a61188a );
 a61195a <=( (not A299)  and  A298 );
 a61198a <=( A302  and  A300 );
 a61199a <=( a61198a  and  a61195a );
 a61200a <=( a61199a  and  a61192a );
 a61204a <=( (not A166)  and  (not A167) );
 a61205a <=( A170  and  a61204a );
 a61208a <=( (not A200)  and  A199 );
 a61211a <=( A203  and  A201 );
 a61212a <=( a61211a  and  a61208a );
 a61213a <=( a61212a  and  a61205a );
 a61216a <=( A233  and  A232 );
 a61219a <=( (not A266)  and  (not A265) );
 a61220a <=( a61219a  and  a61216a );
 a61223a <=( (not A299)  and  A298 );
 a61226a <=( A301  and  A300 );
 a61227a <=( a61226a  and  a61223a );
 a61228a <=( a61227a  and  a61220a );
 a61232a <=( (not A166)  and  (not A167) );
 a61233a <=( A170  and  a61232a );
 a61236a <=( (not A200)  and  A199 );
 a61239a <=( A203  and  A201 );
 a61240a <=( a61239a  and  a61236a );
 a61241a <=( a61240a  and  a61233a );
 a61244a <=( A233  and  A232 );
 a61247a <=( (not A266)  and  (not A265) );
 a61248a <=( a61247a  and  a61244a );
 a61251a <=( (not A299)  and  A298 );
 a61254a <=( A302  and  A300 );
 a61255a <=( a61254a  and  a61251a );
 a61256a <=( a61255a  and  a61248a );
 a61260a <=( (not A166)  and  (not A167) );
 a61261a <=( A170  and  a61260a );
 a61264a <=( (not A200)  and  A199 );
 a61267a <=( A203  and  A201 );
 a61268a <=( a61267a  and  a61264a );
 a61269a <=( a61268a  and  a61261a );
 a61272a <=( (not A235)  and  (not A233) );
 a61275a <=( (not A266)  and  (not A236) );
 a61276a <=( a61275a  and  a61272a );
 a61279a <=( (not A269)  and  (not A268) );
 a61282a <=( A299  and  (not A298) );
 a61283a <=( a61282a  and  a61279a );
 a61284a <=( a61283a  and  a61276a );
 a61288a <=( (not A166)  and  (not A167) );
 a61289a <=( A170  and  a61288a );
 a61292a <=( (not A200)  and  A199 );
 a61295a <=( A203  and  A201 );
 a61296a <=( a61295a  and  a61292a );
 a61297a <=( a61296a  and  a61289a );
 a61300a <=( (not A234)  and  (not A233) );
 a61303a <=( A266  and  A265 );
 a61304a <=( a61303a  and  a61300a );
 a61307a <=( (not A299)  and  A298 );
 a61310a <=( A301  and  A300 );
 a61311a <=( a61310a  and  a61307a );
 a61312a <=( a61311a  and  a61304a );
 a61316a <=( (not A166)  and  (not A167) );
 a61317a <=( A170  and  a61316a );
 a61320a <=( (not A200)  and  A199 );
 a61323a <=( A203  and  A201 );
 a61324a <=( a61323a  and  a61320a );
 a61325a <=( a61324a  and  a61317a );
 a61328a <=( (not A234)  and  (not A233) );
 a61331a <=( A266  and  A265 );
 a61332a <=( a61331a  and  a61328a );
 a61335a <=( (not A299)  and  A298 );
 a61338a <=( A302  and  A300 );
 a61339a <=( a61338a  and  a61335a );
 a61340a <=( a61339a  and  a61332a );
 a61344a <=( (not A166)  and  (not A167) );
 a61345a <=( A170  and  a61344a );
 a61348a <=( (not A200)  and  A199 );
 a61351a <=( A203  and  A201 );
 a61352a <=( a61351a  and  a61348a );
 a61353a <=( a61352a  and  a61345a );
 a61356a <=( (not A234)  and  (not A233) );
 a61359a <=( (not A267)  and  (not A266) );
 a61360a <=( a61359a  and  a61356a );
 a61363a <=( (not A299)  and  A298 );
 a61366a <=( A301  and  A300 );
 a61367a <=( a61366a  and  a61363a );
 a61368a <=( a61367a  and  a61360a );
 a61372a <=( (not A166)  and  (not A167) );
 a61373a <=( A170  and  a61372a );
 a61376a <=( (not A200)  and  A199 );
 a61379a <=( A203  and  A201 );
 a61380a <=( a61379a  and  a61376a );
 a61381a <=( a61380a  and  a61373a );
 a61384a <=( (not A234)  and  (not A233) );
 a61387a <=( (not A267)  and  (not A266) );
 a61388a <=( a61387a  and  a61384a );
 a61391a <=( (not A299)  and  A298 );
 a61394a <=( A302  and  A300 );
 a61395a <=( a61394a  and  a61391a );
 a61396a <=( a61395a  and  a61388a );
 a61400a <=( (not A166)  and  (not A167) );
 a61401a <=( A170  and  a61400a );
 a61404a <=( (not A200)  and  A199 );
 a61407a <=( A203  and  A201 );
 a61408a <=( a61407a  and  a61404a );
 a61409a <=( a61408a  and  a61401a );
 a61412a <=( (not A234)  and  (not A233) );
 a61415a <=( (not A266)  and  (not A265) );
 a61416a <=( a61415a  and  a61412a );
 a61419a <=( (not A299)  and  A298 );
 a61422a <=( A301  and  A300 );
 a61423a <=( a61422a  and  a61419a );
 a61424a <=( a61423a  and  a61416a );
 a61428a <=( (not A166)  and  (not A167) );
 a61429a <=( A170  and  a61428a );
 a61432a <=( (not A200)  and  A199 );
 a61435a <=( A203  and  A201 );
 a61436a <=( a61435a  and  a61432a );
 a61437a <=( a61436a  and  a61429a );
 a61440a <=( (not A234)  and  (not A233) );
 a61443a <=( (not A266)  and  (not A265) );
 a61444a <=( a61443a  and  a61440a );
 a61447a <=( (not A299)  and  A298 );
 a61450a <=( A302  and  A300 );
 a61451a <=( a61450a  and  a61447a );
 a61452a <=( a61451a  and  a61444a );
 a61456a <=( (not A166)  and  (not A167) );
 a61457a <=( A170  and  a61456a );
 a61460a <=( (not A200)  and  A199 );
 a61463a <=( A203  and  A201 );
 a61464a <=( a61463a  and  a61460a );
 a61465a <=( a61464a  and  a61457a );
 a61468a <=( (not A233)  and  A232 );
 a61471a <=( A235  and  A234 );
 a61472a <=( a61471a  and  a61468a );
 a61475a <=( (not A266)  and  A265 );
 a61478a <=( A268  and  A267 );
 a61479a <=( a61478a  and  a61475a );
 a61480a <=( a61479a  and  a61472a );
 a61484a <=( (not A166)  and  (not A167) );
 a61485a <=( A170  and  a61484a );
 a61488a <=( (not A200)  and  A199 );
 a61491a <=( A203  and  A201 );
 a61492a <=( a61491a  and  a61488a );
 a61493a <=( a61492a  and  a61485a );
 a61496a <=( (not A233)  and  A232 );
 a61499a <=( A235  and  A234 );
 a61500a <=( a61499a  and  a61496a );
 a61503a <=( (not A266)  and  A265 );
 a61506a <=( A269  and  A267 );
 a61507a <=( a61506a  and  a61503a );
 a61508a <=( a61507a  and  a61500a );
 a61512a <=( (not A166)  and  (not A167) );
 a61513a <=( A170  and  a61512a );
 a61516a <=( (not A200)  and  A199 );
 a61519a <=( A203  and  A201 );
 a61520a <=( a61519a  and  a61516a );
 a61521a <=( a61520a  and  a61513a );
 a61524a <=( (not A233)  and  A232 );
 a61527a <=( A236  and  A234 );
 a61528a <=( a61527a  and  a61524a );
 a61531a <=( (not A266)  and  A265 );
 a61534a <=( A268  and  A267 );
 a61535a <=( a61534a  and  a61531a );
 a61536a <=( a61535a  and  a61528a );
 a61540a <=( (not A166)  and  (not A167) );
 a61541a <=( A170  and  a61540a );
 a61544a <=( (not A200)  and  A199 );
 a61547a <=( A203  and  A201 );
 a61548a <=( a61547a  and  a61544a );
 a61549a <=( a61548a  and  a61541a );
 a61552a <=( (not A233)  and  A232 );
 a61555a <=( A236  and  A234 );
 a61556a <=( a61555a  and  a61552a );
 a61559a <=( (not A266)  and  A265 );
 a61562a <=( A269  and  A267 );
 a61563a <=( a61562a  and  a61559a );
 a61564a <=( a61563a  and  a61556a );
 a61568a <=( (not A166)  and  (not A167) );
 a61569a <=( A170  and  a61568a );
 a61572a <=( (not A200)  and  A199 );
 a61575a <=( A203  and  A201 );
 a61576a <=( a61575a  and  a61572a );
 a61577a <=( a61576a  and  a61569a );
 a61580a <=( (not A233)  and  (not A232) );
 a61583a <=( A266  and  A265 );
 a61584a <=( a61583a  and  a61580a );
 a61587a <=( (not A299)  and  A298 );
 a61590a <=( A301  and  A300 );
 a61591a <=( a61590a  and  a61587a );
 a61592a <=( a61591a  and  a61584a );
 a61596a <=( (not A166)  and  (not A167) );
 a61597a <=( A170  and  a61596a );
 a61600a <=( (not A200)  and  A199 );
 a61603a <=( A203  and  A201 );
 a61604a <=( a61603a  and  a61600a );
 a61605a <=( a61604a  and  a61597a );
 a61608a <=( (not A233)  and  (not A232) );
 a61611a <=( A266  and  A265 );
 a61612a <=( a61611a  and  a61608a );
 a61615a <=( (not A299)  and  A298 );
 a61618a <=( A302  and  A300 );
 a61619a <=( a61618a  and  a61615a );
 a61620a <=( a61619a  and  a61612a );
 a61624a <=( (not A166)  and  (not A167) );
 a61625a <=( A170  and  a61624a );
 a61628a <=( (not A200)  and  A199 );
 a61631a <=( A203  and  A201 );
 a61632a <=( a61631a  and  a61628a );
 a61633a <=( a61632a  and  a61625a );
 a61636a <=( (not A233)  and  (not A232) );
 a61639a <=( (not A267)  and  (not A266) );
 a61640a <=( a61639a  and  a61636a );
 a61643a <=( (not A299)  and  A298 );
 a61646a <=( A301  and  A300 );
 a61647a <=( a61646a  and  a61643a );
 a61648a <=( a61647a  and  a61640a );
 a61652a <=( (not A166)  and  (not A167) );
 a61653a <=( A170  and  a61652a );
 a61656a <=( (not A200)  and  A199 );
 a61659a <=( A203  and  A201 );
 a61660a <=( a61659a  and  a61656a );
 a61661a <=( a61660a  and  a61653a );
 a61664a <=( (not A233)  and  (not A232) );
 a61667a <=( (not A267)  and  (not A266) );
 a61668a <=( a61667a  and  a61664a );
 a61671a <=( (not A299)  and  A298 );
 a61674a <=( A302  and  A300 );
 a61675a <=( a61674a  and  a61671a );
 a61676a <=( a61675a  and  a61668a );
 a61680a <=( (not A166)  and  (not A167) );
 a61681a <=( A170  and  a61680a );
 a61684a <=( (not A200)  and  A199 );
 a61687a <=( A203  and  A201 );
 a61688a <=( a61687a  and  a61684a );
 a61689a <=( a61688a  and  a61681a );
 a61692a <=( (not A233)  and  (not A232) );
 a61695a <=( (not A266)  and  (not A265) );
 a61696a <=( a61695a  and  a61692a );
 a61699a <=( (not A299)  and  A298 );
 a61702a <=( A301  and  A300 );
 a61703a <=( a61702a  and  a61699a );
 a61704a <=( a61703a  and  a61696a );
 a61708a <=( (not A166)  and  (not A167) );
 a61709a <=( A170  and  a61708a );
 a61712a <=( (not A200)  and  A199 );
 a61715a <=( A203  and  A201 );
 a61716a <=( a61715a  and  a61712a );
 a61717a <=( a61716a  and  a61709a );
 a61720a <=( (not A233)  and  (not A232) );
 a61723a <=( (not A266)  and  (not A265) );
 a61724a <=( a61723a  and  a61720a );
 a61727a <=( (not A299)  and  A298 );
 a61730a <=( A302  and  A300 );
 a61731a <=( a61730a  and  a61727a );
 a61732a <=( a61731a  and  a61724a );
 a61736a <=( A167  and  (not A168) );
 a61737a <=( A170  and  a61736a );
 a61740a <=( (not A199)  and  A166 );
 a61743a <=( A232  and  A200 );
 a61744a <=( a61743a  and  a61740a );
 a61745a <=( a61744a  and  a61737a );
 a61748a <=( A265  and  A233 );
 a61751a <=( (not A269)  and  (not A268) );
 a61752a <=( a61751a  and  a61748a );
 a61755a <=( (not A299)  and  A298 );
 a61758a <=( A301  and  A300 );
 a61759a <=( a61758a  and  a61755a );
 a61760a <=( a61759a  and  a61752a );
 a61764a <=( A167  and  (not A168) );
 a61765a <=( A170  and  a61764a );
 a61768a <=( (not A199)  and  A166 );
 a61771a <=( A232  and  A200 );
 a61772a <=( a61771a  and  a61768a );
 a61773a <=( a61772a  and  a61765a );
 a61776a <=( A265  and  A233 );
 a61779a <=( (not A269)  and  (not A268) );
 a61780a <=( a61779a  and  a61776a );
 a61783a <=( (not A299)  and  A298 );
 a61786a <=( A302  and  A300 );
 a61787a <=( a61786a  and  a61783a );
 a61788a <=( a61787a  and  a61780a );
 a61792a <=( A167  and  (not A168) );
 a61793a <=( A170  and  a61792a );
 a61796a <=( (not A199)  and  A166 );
 a61799a <=( (not A233)  and  A200 );
 a61800a <=( a61799a  and  a61796a );
 a61801a <=( a61800a  and  a61793a );
 a61804a <=( (not A236)  and  (not A235) );
 a61807a <=( A266  and  A265 );
 a61808a <=( a61807a  and  a61804a );
 a61811a <=( (not A299)  and  A298 );
 a61814a <=( A301  and  A300 );
 a61815a <=( a61814a  and  a61811a );
 a61816a <=( a61815a  and  a61808a );
 a61820a <=( A167  and  (not A168) );
 a61821a <=( A170  and  a61820a );
 a61824a <=( (not A199)  and  A166 );
 a61827a <=( (not A233)  and  A200 );
 a61828a <=( a61827a  and  a61824a );
 a61829a <=( a61828a  and  a61821a );
 a61832a <=( (not A236)  and  (not A235) );
 a61835a <=( A266  and  A265 );
 a61836a <=( a61835a  and  a61832a );
 a61839a <=( (not A299)  and  A298 );
 a61842a <=( A302  and  A300 );
 a61843a <=( a61842a  and  a61839a );
 a61844a <=( a61843a  and  a61836a );
 a61848a <=( A167  and  (not A168) );
 a61849a <=( A170  and  a61848a );
 a61852a <=( (not A199)  and  A166 );
 a61855a <=( (not A233)  and  A200 );
 a61856a <=( a61855a  and  a61852a );
 a61857a <=( a61856a  and  a61849a );
 a61860a <=( (not A236)  and  (not A235) );
 a61863a <=( (not A267)  and  (not A266) );
 a61864a <=( a61863a  and  a61860a );
 a61867a <=( (not A299)  and  A298 );
 a61870a <=( A301  and  A300 );
 a61871a <=( a61870a  and  a61867a );
 a61872a <=( a61871a  and  a61864a );
 a61876a <=( A167  and  (not A168) );
 a61877a <=( A170  and  a61876a );
 a61880a <=( (not A199)  and  A166 );
 a61883a <=( (not A233)  and  A200 );
 a61884a <=( a61883a  and  a61880a );
 a61885a <=( a61884a  and  a61877a );
 a61888a <=( (not A236)  and  (not A235) );
 a61891a <=( (not A267)  and  (not A266) );
 a61892a <=( a61891a  and  a61888a );
 a61895a <=( (not A299)  and  A298 );
 a61898a <=( A302  and  A300 );
 a61899a <=( a61898a  and  a61895a );
 a61900a <=( a61899a  and  a61892a );
 a61904a <=( A167  and  (not A168) );
 a61905a <=( A170  and  a61904a );
 a61908a <=( (not A199)  and  A166 );
 a61911a <=( (not A233)  and  A200 );
 a61912a <=( a61911a  and  a61908a );
 a61913a <=( a61912a  and  a61905a );
 a61916a <=( (not A236)  and  (not A235) );
 a61919a <=( (not A266)  and  (not A265) );
 a61920a <=( a61919a  and  a61916a );
 a61923a <=( (not A299)  and  A298 );
 a61926a <=( A301  and  A300 );
 a61927a <=( a61926a  and  a61923a );
 a61928a <=( a61927a  and  a61920a );
 a61932a <=( A167  and  (not A168) );
 a61933a <=( A170  and  a61932a );
 a61936a <=( (not A199)  and  A166 );
 a61939a <=( (not A233)  and  A200 );
 a61940a <=( a61939a  and  a61936a );
 a61941a <=( a61940a  and  a61933a );
 a61944a <=( (not A236)  and  (not A235) );
 a61947a <=( (not A266)  and  (not A265) );
 a61948a <=( a61947a  and  a61944a );
 a61951a <=( (not A299)  and  A298 );
 a61954a <=( A302  and  A300 );
 a61955a <=( a61954a  and  a61951a );
 a61956a <=( a61955a  and  a61948a );
 a61960a <=( A167  and  (not A168) );
 a61961a <=( A170  and  a61960a );
 a61964a <=( (not A199)  and  A166 );
 a61967a <=( (not A233)  and  A200 );
 a61968a <=( a61967a  and  a61964a );
 a61969a <=( a61968a  and  a61961a );
 a61972a <=( (not A266)  and  (not A234) );
 a61975a <=( (not A269)  and  (not A268) );
 a61976a <=( a61975a  and  a61972a );
 a61979a <=( (not A299)  and  A298 );
 a61982a <=( A301  and  A300 );
 a61983a <=( a61982a  and  a61979a );
 a61984a <=( a61983a  and  a61976a );
 a61988a <=( A167  and  (not A168) );
 a61989a <=( A170  and  a61988a );
 a61992a <=( (not A199)  and  A166 );
 a61995a <=( (not A233)  and  A200 );
 a61996a <=( a61995a  and  a61992a );
 a61997a <=( a61996a  and  a61989a );
 a62000a <=( (not A266)  and  (not A234) );
 a62003a <=( (not A269)  and  (not A268) );
 a62004a <=( a62003a  and  a62000a );
 a62007a <=( (not A299)  and  A298 );
 a62010a <=( A302  and  A300 );
 a62011a <=( a62010a  and  a62007a );
 a62012a <=( a62011a  and  a62004a );
 a62016a <=( A167  and  (not A168) );
 a62017a <=( A170  and  a62016a );
 a62020a <=( (not A199)  and  A166 );
 a62023a <=( (not A232)  and  A200 );
 a62024a <=( a62023a  and  a62020a );
 a62025a <=( a62024a  and  a62017a );
 a62028a <=( (not A266)  and  (not A233) );
 a62031a <=( (not A269)  and  (not A268) );
 a62032a <=( a62031a  and  a62028a );
 a62035a <=( (not A299)  and  A298 );
 a62038a <=( A301  and  A300 );
 a62039a <=( a62038a  and  a62035a );
 a62040a <=( a62039a  and  a62032a );
 a62044a <=( A167  and  (not A168) );
 a62045a <=( A170  and  a62044a );
 a62048a <=( (not A199)  and  A166 );
 a62051a <=( (not A232)  and  A200 );
 a62052a <=( a62051a  and  a62048a );
 a62053a <=( a62052a  and  a62045a );
 a62056a <=( (not A266)  and  (not A233) );
 a62059a <=( (not A269)  and  (not A268) );
 a62060a <=( a62059a  and  a62056a );
 a62063a <=( (not A299)  and  A298 );
 a62066a <=( A302  and  A300 );
 a62067a <=( a62066a  and  a62063a );
 a62068a <=( a62067a  and  a62060a );
 a62072a <=( A167  and  (not A168) );
 a62073a <=( (not A170)  and  a62072a );
 a62076a <=( (not A199)  and  (not A166) );
 a62079a <=( A232  and  A200 );
 a62080a <=( a62079a  and  a62076a );
 a62081a <=( a62080a  and  a62073a );
 a62084a <=( A265  and  A233 );
 a62087a <=( (not A269)  and  (not A268) );
 a62088a <=( a62087a  and  a62084a );
 a62091a <=( (not A299)  and  A298 );
 a62094a <=( A301  and  A300 );
 a62095a <=( a62094a  and  a62091a );
 a62096a <=( a62095a  and  a62088a );
 a62100a <=( A167  and  (not A168) );
 a62101a <=( (not A170)  and  a62100a );
 a62104a <=( (not A199)  and  (not A166) );
 a62107a <=( A232  and  A200 );
 a62108a <=( a62107a  and  a62104a );
 a62109a <=( a62108a  and  a62101a );
 a62112a <=( A265  and  A233 );
 a62115a <=( (not A269)  and  (not A268) );
 a62116a <=( a62115a  and  a62112a );
 a62119a <=( (not A299)  and  A298 );
 a62122a <=( A302  and  A300 );
 a62123a <=( a62122a  and  a62119a );
 a62124a <=( a62123a  and  a62116a );
 a62128a <=( A167  and  (not A168) );
 a62129a <=( (not A170)  and  a62128a );
 a62132a <=( (not A199)  and  (not A166) );
 a62135a <=( (not A233)  and  A200 );
 a62136a <=( a62135a  and  a62132a );
 a62137a <=( a62136a  and  a62129a );
 a62140a <=( (not A236)  and  (not A235) );
 a62143a <=( A266  and  A265 );
 a62144a <=( a62143a  and  a62140a );
 a62147a <=( (not A299)  and  A298 );
 a62150a <=( A301  and  A300 );
 a62151a <=( a62150a  and  a62147a );
 a62152a <=( a62151a  and  a62144a );
 a62156a <=( A167  and  (not A168) );
 a62157a <=( (not A170)  and  a62156a );
 a62160a <=( (not A199)  and  (not A166) );
 a62163a <=( (not A233)  and  A200 );
 a62164a <=( a62163a  and  a62160a );
 a62165a <=( a62164a  and  a62157a );
 a62168a <=( (not A236)  and  (not A235) );
 a62171a <=( A266  and  A265 );
 a62172a <=( a62171a  and  a62168a );
 a62175a <=( (not A299)  and  A298 );
 a62178a <=( A302  and  A300 );
 a62179a <=( a62178a  and  a62175a );
 a62180a <=( a62179a  and  a62172a );
 a62184a <=( A167  and  (not A168) );
 a62185a <=( (not A170)  and  a62184a );
 a62188a <=( (not A199)  and  (not A166) );
 a62191a <=( (not A233)  and  A200 );
 a62192a <=( a62191a  and  a62188a );
 a62193a <=( a62192a  and  a62185a );
 a62196a <=( (not A236)  and  (not A235) );
 a62199a <=( (not A267)  and  (not A266) );
 a62200a <=( a62199a  and  a62196a );
 a62203a <=( (not A299)  and  A298 );
 a62206a <=( A301  and  A300 );
 a62207a <=( a62206a  and  a62203a );
 a62208a <=( a62207a  and  a62200a );
 a62212a <=( A167  and  (not A168) );
 a62213a <=( (not A170)  and  a62212a );
 a62216a <=( (not A199)  and  (not A166) );
 a62219a <=( (not A233)  and  A200 );
 a62220a <=( a62219a  and  a62216a );
 a62221a <=( a62220a  and  a62213a );
 a62224a <=( (not A236)  and  (not A235) );
 a62227a <=( (not A267)  and  (not A266) );
 a62228a <=( a62227a  and  a62224a );
 a62231a <=( (not A299)  and  A298 );
 a62234a <=( A302  and  A300 );
 a62235a <=( a62234a  and  a62231a );
 a62236a <=( a62235a  and  a62228a );
 a62240a <=( A167  and  (not A168) );
 a62241a <=( (not A170)  and  a62240a );
 a62244a <=( (not A199)  and  (not A166) );
 a62247a <=( (not A233)  and  A200 );
 a62248a <=( a62247a  and  a62244a );
 a62249a <=( a62248a  and  a62241a );
 a62252a <=( (not A236)  and  (not A235) );
 a62255a <=( (not A266)  and  (not A265) );
 a62256a <=( a62255a  and  a62252a );
 a62259a <=( (not A299)  and  A298 );
 a62262a <=( A301  and  A300 );
 a62263a <=( a62262a  and  a62259a );
 a62264a <=( a62263a  and  a62256a );
 a62268a <=( A167  and  (not A168) );
 a62269a <=( (not A170)  and  a62268a );
 a62272a <=( (not A199)  and  (not A166) );
 a62275a <=( (not A233)  and  A200 );
 a62276a <=( a62275a  and  a62272a );
 a62277a <=( a62276a  and  a62269a );
 a62280a <=( (not A236)  and  (not A235) );
 a62283a <=( (not A266)  and  (not A265) );
 a62284a <=( a62283a  and  a62280a );
 a62287a <=( (not A299)  and  A298 );
 a62290a <=( A302  and  A300 );
 a62291a <=( a62290a  and  a62287a );
 a62292a <=( a62291a  and  a62284a );
 a62296a <=( A167  and  (not A168) );
 a62297a <=( (not A170)  and  a62296a );
 a62300a <=( (not A199)  and  (not A166) );
 a62303a <=( (not A233)  and  A200 );
 a62304a <=( a62303a  and  a62300a );
 a62305a <=( a62304a  and  a62297a );
 a62308a <=( (not A266)  and  (not A234) );
 a62311a <=( (not A269)  and  (not A268) );
 a62312a <=( a62311a  and  a62308a );
 a62315a <=( (not A299)  and  A298 );
 a62318a <=( A301  and  A300 );
 a62319a <=( a62318a  and  a62315a );
 a62320a <=( a62319a  and  a62312a );
 a62324a <=( A167  and  (not A168) );
 a62325a <=( (not A170)  and  a62324a );
 a62328a <=( (not A199)  and  (not A166) );
 a62331a <=( (not A233)  and  A200 );
 a62332a <=( a62331a  and  a62328a );
 a62333a <=( a62332a  and  a62325a );
 a62336a <=( (not A266)  and  (not A234) );
 a62339a <=( (not A269)  and  (not A268) );
 a62340a <=( a62339a  and  a62336a );
 a62343a <=( (not A299)  and  A298 );
 a62346a <=( A302  and  A300 );
 a62347a <=( a62346a  and  a62343a );
 a62348a <=( a62347a  and  a62340a );
 a62352a <=( A167  and  (not A168) );
 a62353a <=( (not A170)  and  a62352a );
 a62356a <=( (not A199)  and  (not A166) );
 a62359a <=( (not A232)  and  A200 );
 a62360a <=( a62359a  and  a62356a );
 a62361a <=( a62360a  and  a62353a );
 a62364a <=( (not A266)  and  (not A233) );
 a62367a <=( (not A269)  and  (not A268) );
 a62368a <=( a62367a  and  a62364a );
 a62371a <=( (not A299)  and  A298 );
 a62374a <=( A301  and  A300 );
 a62375a <=( a62374a  and  a62371a );
 a62376a <=( a62375a  and  a62368a );
 a62380a <=( A167  and  (not A168) );
 a62381a <=( (not A170)  and  a62380a );
 a62384a <=( (not A199)  and  (not A166) );
 a62387a <=( (not A232)  and  A200 );
 a62388a <=( a62387a  and  a62384a );
 a62389a <=( a62388a  and  a62381a );
 a62392a <=( (not A266)  and  (not A233) );
 a62395a <=( (not A269)  and  (not A268) );
 a62396a <=( a62395a  and  a62392a );
 a62399a <=( (not A299)  and  A298 );
 a62402a <=( A302  and  A300 );
 a62403a <=( a62402a  and  a62399a );
 a62404a <=( a62403a  and  a62396a );
 a62408a <=( (not A167)  and  (not A168) );
 a62409a <=( (not A170)  and  a62408a );
 a62412a <=( (not A199)  and  A166 );
 a62415a <=( A232  and  A200 );
 a62416a <=( a62415a  and  a62412a );
 a62417a <=( a62416a  and  a62409a );
 a62420a <=( A265  and  A233 );
 a62423a <=( (not A269)  and  (not A268) );
 a62424a <=( a62423a  and  a62420a );
 a62427a <=( (not A299)  and  A298 );
 a62430a <=( A301  and  A300 );
 a62431a <=( a62430a  and  a62427a );
 a62432a <=( a62431a  and  a62424a );
 a62436a <=( (not A167)  and  (not A168) );
 a62437a <=( (not A170)  and  a62436a );
 a62440a <=( (not A199)  and  A166 );
 a62443a <=( A232  and  A200 );
 a62444a <=( a62443a  and  a62440a );
 a62445a <=( a62444a  and  a62437a );
 a62448a <=( A265  and  A233 );
 a62451a <=( (not A269)  and  (not A268) );
 a62452a <=( a62451a  and  a62448a );
 a62455a <=( (not A299)  and  A298 );
 a62458a <=( A302  and  A300 );
 a62459a <=( a62458a  and  a62455a );
 a62460a <=( a62459a  and  a62452a );
 a62464a <=( (not A167)  and  (not A168) );
 a62465a <=( (not A170)  and  a62464a );
 a62468a <=( (not A199)  and  A166 );
 a62471a <=( (not A233)  and  A200 );
 a62472a <=( a62471a  and  a62468a );
 a62473a <=( a62472a  and  a62465a );
 a62476a <=( (not A236)  and  (not A235) );
 a62479a <=( A266  and  A265 );
 a62480a <=( a62479a  and  a62476a );
 a62483a <=( (not A299)  and  A298 );
 a62486a <=( A301  and  A300 );
 a62487a <=( a62486a  and  a62483a );
 a62488a <=( a62487a  and  a62480a );
 a62492a <=( (not A167)  and  (not A168) );
 a62493a <=( (not A170)  and  a62492a );
 a62496a <=( (not A199)  and  A166 );
 a62499a <=( (not A233)  and  A200 );
 a62500a <=( a62499a  and  a62496a );
 a62501a <=( a62500a  and  a62493a );
 a62504a <=( (not A236)  and  (not A235) );
 a62507a <=( A266  and  A265 );
 a62508a <=( a62507a  and  a62504a );
 a62511a <=( (not A299)  and  A298 );
 a62514a <=( A302  and  A300 );
 a62515a <=( a62514a  and  a62511a );
 a62516a <=( a62515a  and  a62508a );
 a62520a <=( (not A167)  and  (not A168) );
 a62521a <=( (not A170)  and  a62520a );
 a62524a <=( (not A199)  and  A166 );
 a62527a <=( (not A233)  and  A200 );
 a62528a <=( a62527a  and  a62524a );
 a62529a <=( a62528a  and  a62521a );
 a62532a <=( (not A236)  and  (not A235) );
 a62535a <=( (not A267)  and  (not A266) );
 a62536a <=( a62535a  and  a62532a );
 a62539a <=( (not A299)  and  A298 );
 a62542a <=( A301  and  A300 );
 a62543a <=( a62542a  and  a62539a );
 a62544a <=( a62543a  and  a62536a );
 a62548a <=( (not A167)  and  (not A168) );
 a62549a <=( (not A170)  and  a62548a );
 a62552a <=( (not A199)  and  A166 );
 a62555a <=( (not A233)  and  A200 );
 a62556a <=( a62555a  and  a62552a );
 a62557a <=( a62556a  and  a62549a );
 a62560a <=( (not A236)  and  (not A235) );
 a62563a <=( (not A267)  and  (not A266) );
 a62564a <=( a62563a  and  a62560a );
 a62567a <=( (not A299)  and  A298 );
 a62570a <=( A302  and  A300 );
 a62571a <=( a62570a  and  a62567a );
 a62572a <=( a62571a  and  a62564a );
 a62576a <=( (not A167)  and  (not A168) );
 a62577a <=( (not A170)  and  a62576a );
 a62580a <=( (not A199)  and  A166 );
 a62583a <=( (not A233)  and  A200 );
 a62584a <=( a62583a  and  a62580a );
 a62585a <=( a62584a  and  a62577a );
 a62588a <=( (not A236)  and  (not A235) );
 a62591a <=( (not A266)  and  (not A265) );
 a62592a <=( a62591a  and  a62588a );
 a62595a <=( (not A299)  and  A298 );
 a62598a <=( A301  and  A300 );
 a62599a <=( a62598a  and  a62595a );
 a62600a <=( a62599a  and  a62592a );
 a62604a <=( (not A167)  and  (not A168) );
 a62605a <=( (not A170)  and  a62604a );
 a62608a <=( (not A199)  and  A166 );
 a62611a <=( (not A233)  and  A200 );
 a62612a <=( a62611a  and  a62608a );
 a62613a <=( a62612a  and  a62605a );
 a62616a <=( (not A236)  and  (not A235) );
 a62619a <=( (not A266)  and  (not A265) );
 a62620a <=( a62619a  and  a62616a );
 a62623a <=( (not A299)  and  A298 );
 a62626a <=( A302  and  A300 );
 a62627a <=( a62626a  and  a62623a );
 a62628a <=( a62627a  and  a62620a );
 a62632a <=( (not A167)  and  (not A168) );
 a62633a <=( (not A170)  and  a62632a );
 a62636a <=( (not A199)  and  A166 );
 a62639a <=( (not A233)  and  A200 );
 a62640a <=( a62639a  and  a62636a );
 a62641a <=( a62640a  and  a62633a );
 a62644a <=( (not A266)  and  (not A234) );
 a62647a <=( (not A269)  and  (not A268) );
 a62648a <=( a62647a  and  a62644a );
 a62651a <=( (not A299)  and  A298 );
 a62654a <=( A301  and  A300 );
 a62655a <=( a62654a  and  a62651a );
 a62656a <=( a62655a  and  a62648a );
 a62660a <=( (not A167)  and  (not A168) );
 a62661a <=( (not A170)  and  a62660a );
 a62664a <=( (not A199)  and  A166 );
 a62667a <=( (not A233)  and  A200 );
 a62668a <=( a62667a  and  a62664a );
 a62669a <=( a62668a  and  a62661a );
 a62672a <=( (not A266)  and  (not A234) );
 a62675a <=( (not A269)  and  (not A268) );
 a62676a <=( a62675a  and  a62672a );
 a62679a <=( (not A299)  and  A298 );
 a62682a <=( A302  and  A300 );
 a62683a <=( a62682a  and  a62679a );
 a62684a <=( a62683a  and  a62676a );
 a62688a <=( (not A167)  and  (not A168) );
 a62689a <=( (not A170)  and  a62688a );
 a62692a <=( (not A199)  and  A166 );
 a62695a <=( (not A232)  and  A200 );
 a62696a <=( a62695a  and  a62692a );
 a62697a <=( a62696a  and  a62689a );
 a62700a <=( (not A266)  and  (not A233) );
 a62703a <=( (not A269)  and  (not A268) );
 a62704a <=( a62703a  and  a62700a );
 a62707a <=( (not A299)  and  A298 );
 a62710a <=( A301  and  A300 );
 a62711a <=( a62710a  and  a62707a );
 a62712a <=( a62711a  and  a62704a );
 a62716a <=( (not A167)  and  (not A168) );
 a62717a <=( (not A170)  and  a62716a );
 a62720a <=( (not A199)  and  A166 );
 a62723a <=( (not A232)  and  A200 );
 a62724a <=( a62723a  and  a62720a );
 a62725a <=( a62724a  and  a62717a );
 a62728a <=( (not A266)  and  (not A233) );
 a62731a <=( (not A269)  and  (not A268) );
 a62732a <=( a62731a  and  a62728a );
 a62735a <=( (not A299)  and  A298 );
 a62738a <=( A302  and  A300 );
 a62739a <=( a62738a  and  a62735a );
 a62740a <=( a62739a  and  a62732a );
 a62744a <=( A167  and  (not A168) );
 a62745a <=( A169  and  a62744a );
 a62748a <=( (not A199)  and  (not A166) );
 a62751a <=( A232  and  A200 );
 a62752a <=( a62751a  and  a62748a );
 a62753a <=( a62752a  and  a62745a );
 a62756a <=( A265  and  A233 );
 a62759a <=( (not A269)  and  (not A268) );
 a62760a <=( a62759a  and  a62756a );
 a62763a <=( (not A299)  and  A298 );
 a62766a <=( A301  and  A300 );
 a62767a <=( a62766a  and  a62763a );
 a62768a <=( a62767a  and  a62760a );
 a62772a <=( A167  and  (not A168) );
 a62773a <=( A169  and  a62772a );
 a62776a <=( (not A199)  and  (not A166) );
 a62779a <=( A232  and  A200 );
 a62780a <=( a62779a  and  a62776a );
 a62781a <=( a62780a  and  a62773a );
 a62784a <=( A265  and  A233 );
 a62787a <=( (not A269)  and  (not A268) );
 a62788a <=( a62787a  and  a62784a );
 a62791a <=( (not A299)  and  A298 );
 a62794a <=( A302  and  A300 );
 a62795a <=( a62794a  and  a62791a );
 a62796a <=( a62795a  and  a62788a );
 a62800a <=( A167  and  (not A168) );
 a62801a <=( A169  and  a62800a );
 a62804a <=( (not A199)  and  (not A166) );
 a62807a <=( (not A233)  and  A200 );
 a62808a <=( a62807a  and  a62804a );
 a62809a <=( a62808a  and  a62801a );
 a62812a <=( (not A236)  and  (not A235) );
 a62815a <=( A266  and  A265 );
 a62816a <=( a62815a  and  a62812a );
 a62819a <=( (not A299)  and  A298 );
 a62822a <=( A301  and  A300 );
 a62823a <=( a62822a  and  a62819a );
 a62824a <=( a62823a  and  a62816a );
 a62828a <=( A167  and  (not A168) );
 a62829a <=( A169  and  a62828a );
 a62832a <=( (not A199)  and  (not A166) );
 a62835a <=( (not A233)  and  A200 );
 a62836a <=( a62835a  and  a62832a );
 a62837a <=( a62836a  and  a62829a );
 a62840a <=( (not A236)  and  (not A235) );
 a62843a <=( A266  and  A265 );
 a62844a <=( a62843a  and  a62840a );
 a62847a <=( (not A299)  and  A298 );
 a62850a <=( A302  and  A300 );
 a62851a <=( a62850a  and  a62847a );
 a62852a <=( a62851a  and  a62844a );
 a62856a <=( A167  and  (not A168) );
 a62857a <=( A169  and  a62856a );
 a62860a <=( (not A199)  and  (not A166) );
 a62863a <=( (not A233)  and  A200 );
 a62864a <=( a62863a  and  a62860a );
 a62865a <=( a62864a  and  a62857a );
 a62868a <=( (not A236)  and  (not A235) );
 a62871a <=( (not A267)  and  (not A266) );
 a62872a <=( a62871a  and  a62868a );
 a62875a <=( (not A299)  and  A298 );
 a62878a <=( A301  and  A300 );
 a62879a <=( a62878a  and  a62875a );
 a62880a <=( a62879a  and  a62872a );
 a62884a <=( A167  and  (not A168) );
 a62885a <=( A169  and  a62884a );
 a62888a <=( (not A199)  and  (not A166) );
 a62891a <=( (not A233)  and  A200 );
 a62892a <=( a62891a  and  a62888a );
 a62893a <=( a62892a  and  a62885a );
 a62896a <=( (not A236)  and  (not A235) );
 a62899a <=( (not A267)  and  (not A266) );
 a62900a <=( a62899a  and  a62896a );
 a62903a <=( (not A299)  and  A298 );
 a62906a <=( A302  and  A300 );
 a62907a <=( a62906a  and  a62903a );
 a62908a <=( a62907a  and  a62900a );
 a62912a <=( A167  and  (not A168) );
 a62913a <=( A169  and  a62912a );
 a62916a <=( (not A199)  and  (not A166) );
 a62919a <=( (not A233)  and  A200 );
 a62920a <=( a62919a  and  a62916a );
 a62921a <=( a62920a  and  a62913a );
 a62924a <=( (not A236)  and  (not A235) );
 a62927a <=( (not A266)  and  (not A265) );
 a62928a <=( a62927a  and  a62924a );
 a62931a <=( (not A299)  and  A298 );
 a62934a <=( A301  and  A300 );
 a62935a <=( a62934a  and  a62931a );
 a62936a <=( a62935a  and  a62928a );
 a62940a <=( A167  and  (not A168) );
 a62941a <=( A169  and  a62940a );
 a62944a <=( (not A199)  and  (not A166) );
 a62947a <=( (not A233)  and  A200 );
 a62948a <=( a62947a  and  a62944a );
 a62949a <=( a62948a  and  a62941a );
 a62952a <=( (not A236)  and  (not A235) );
 a62955a <=( (not A266)  and  (not A265) );
 a62956a <=( a62955a  and  a62952a );
 a62959a <=( (not A299)  and  A298 );
 a62962a <=( A302  and  A300 );
 a62963a <=( a62962a  and  a62959a );
 a62964a <=( a62963a  and  a62956a );
 a62968a <=( A167  and  (not A168) );
 a62969a <=( A169  and  a62968a );
 a62972a <=( (not A199)  and  (not A166) );
 a62975a <=( (not A233)  and  A200 );
 a62976a <=( a62975a  and  a62972a );
 a62977a <=( a62976a  and  a62969a );
 a62980a <=( (not A266)  and  (not A234) );
 a62983a <=( (not A269)  and  (not A268) );
 a62984a <=( a62983a  and  a62980a );
 a62987a <=( (not A299)  and  A298 );
 a62990a <=( A301  and  A300 );
 a62991a <=( a62990a  and  a62987a );
 a62992a <=( a62991a  and  a62984a );
 a62996a <=( A167  and  (not A168) );
 a62997a <=( A169  and  a62996a );
 a63000a <=( (not A199)  and  (not A166) );
 a63003a <=( (not A233)  and  A200 );
 a63004a <=( a63003a  and  a63000a );
 a63005a <=( a63004a  and  a62997a );
 a63008a <=( (not A266)  and  (not A234) );
 a63011a <=( (not A269)  and  (not A268) );
 a63012a <=( a63011a  and  a63008a );
 a63015a <=( (not A299)  and  A298 );
 a63018a <=( A302  and  A300 );
 a63019a <=( a63018a  and  a63015a );
 a63020a <=( a63019a  and  a63012a );
 a63024a <=( A167  and  (not A168) );
 a63025a <=( A169  and  a63024a );
 a63028a <=( (not A199)  and  (not A166) );
 a63031a <=( (not A232)  and  A200 );
 a63032a <=( a63031a  and  a63028a );
 a63033a <=( a63032a  and  a63025a );
 a63036a <=( (not A266)  and  (not A233) );
 a63039a <=( (not A269)  and  (not A268) );
 a63040a <=( a63039a  and  a63036a );
 a63043a <=( (not A299)  and  A298 );
 a63046a <=( A301  and  A300 );
 a63047a <=( a63046a  and  a63043a );
 a63048a <=( a63047a  and  a63040a );
 a63052a <=( A167  and  (not A168) );
 a63053a <=( A169  and  a63052a );
 a63056a <=( (not A199)  and  (not A166) );
 a63059a <=( (not A232)  and  A200 );
 a63060a <=( a63059a  and  a63056a );
 a63061a <=( a63060a  and  a63053a );
 a63064a <=( (not A266)  and  (not A233) );
 a63067a <=( (not A269)  and  (not A268) );
 a63068a <=( a63067a  and  a63064a );
 a63071a <=( (not A299)  and  A298 );
 a63074a <=( A302  and  A300 );
 a63075a <=( a63074a  and  a63071a );
 a63076a <=( a63075a  and  a63068a );
 a63080a <=( A167  and  (not A168) );
 a63081a <=( A169  and  a63080a );
 a63084a <=( A199  and  (not A166) );
 a63087a <=( A201  and  (not A200) );
 a63088a <=( a63087a  and  a63084a );
 a63089a <=( a63088a  and  a63081a );
 a63092a <=( A232  and  A202 );
 a63095a <=( A265  and  A233 );
 a63096a <=( a63095a  and  a63092a );
 a63099a <=( (not A269)  and  (not A268) );
 a63102a <=( A299  and  (not A298) );
 a63103a <=( a63102a  and  a63099a );
 a63104a <=( a63103a  and  a63096a );
 a63108a <=( A167  and  (not A168) );
 a63109a <=( A169  and  a63108a );
 a63112a <=( A199  and  (not A166) );
 a63115a <=( A201  and  (not A200) );
 a63116a <=( a63115a  and  a63112a );
 a63117a <=( a63116a  and  a63109a );
 a63120a <=( (not A233)  and  A202 );
 a63123a <=( (not A236)  and  (not A235) );
 a63124a <=( a63123a  and  a63120a );
 a63127a <=( A266  and  A265 );
 a63130a <=( A299  and  (not A298) );
 a63131a <=( a63130a  and  a63127a );
 a63132a <=( a63131a  and  a63124a );
 a63136a <=( A167  and  (not A168) );
 a63137a <=( A169  and  a63136a );
 a63140a <=( A199  and  (not A166) );
 a63143a <=( A201  and  (not A200) );
 a63144a <=( a63143a  and  a63140a );
 a63145a <=( a63144a  and  a63137a );
 a63148a <=( (not A233)  and  A202 );
 a63151a <=( (not A236)  and  (not A235) );
 a63152a <=( a63151a  and  a63148a );
 a63155a <=( (not A267)  and  (not A266) );
 a63158a <=( A299  and  (not A298) );
 a63159a <=( a63158a  and  a63155a );
 a63160a <=( a63159a  and  a63152a );
 a63164a <=( A167  and  (not A168) );
 a63165a <=( A169  and  a63164a );
 a63168a <=( A199  and  (not A166) );
 a63171a <=( A201  and  (not A200) );
 a63172a <=( a63171a  and  a63168a );
 a63173a <=( a63172a  and  a63165a );
 a63176a <=( (not A233)  and  A202 );
 a63179a <=( (not A236)  and  (not A235) );
 a63180a <=( a63179a  and  a63176a );
 a63183a <=( (not A266)  and  (not A265) );
 a63186a <=( A299  and  (not A298) );
 a63187a <=( a63186a  and  a63183a );
 a63188a <=( a63187a  and  a63180a );
 a63192a <=( A167  and  (not A168) );
 a63193a <=( A169  and  a63192a );
 a63196a <=( A199  and  (not A166) );
 a63199a <=( A201  and  (not A200) );
 a63200a <=( a63199a  and  a63196a );
 a63201a <=( a63200a  and  a63193a );
 a63204a <=( (not A233)  and  A202 );
 a63207a <=( (not A266)  and  (not A234) );
 a63208a <=( a63207a  and  a63204a );
 a63211a <=( (not A269)  and  (not A268) );
 a63214a <=( A299  and  (not A298) );
 a63215a <=( a63214a  and  a63211a );
 a63216a <=( a63215a  and  a63208a );
 a63220a <=( A167  and  (not A168) );
 a63221a <=( A169  and  a63220a );
 a63224a <=( A199  and  (not A166) );
 a63227a <=( A201  and  (not A200) );
 a63228a <=( a63227a  and  a63224a );
 a63229a <=( a63228a  and  a63221a );
 a63232a <=( A232  and  A202 );
 a63235a <=( A234  and  (not A233) );
 a63236a <=( a63235a  and  a63232a );
 a63239a <=( A298  and  A235 );
 a63242a <=( (not A302)  and  (not A301) );
 a63243a <=( a63242a  and  a63239a );
 a63244a <=( a63243a  and  a63236a );
 a63248a <=( A167  and  (not A168) );
 a63249a <=( A169  and  a63248a );
 a63252a <=( A199  and  (not A166) );
 a63255a <=( A201  and  (not A200) );
 a63256a <=( a63255a  and  a63252a );
 a63257a <=( a63256a  and  a63249a );
 a63260a <=( A232  and  A202 );
 a63263a <=( A234  and  (not A233) );
 a63264a <=( a63263a  and  a63260a );
 a63267a <=( A298  and  A236 );
 a63270a <=( (not A302)  and  (not A301) );
 a63271a <=( a63270a  and  a63267a );
 a63272a <=( a63271a  and  a63264a );
 a63276a <=( A167  and  (not A168) );
 a63277a <=( A169  and  a63276a );
 a63280a <=( A199  and  (not A166) );
 a63283a <=( A201  and  (not A200) );
 a63284a <=( a63283a  and  a63280a );
 a63285a <=( a63284a  and  a63277a );
 a63288a <=( (not A232)  and  A202 );
 a63291a <=( (not A266)  and  (not A233) );
 a63292a <=( a63291a  and  a63288a );
 a63295a <=( (not A269)  and  (not A268) );
 a63298a <=( A299  and  (not A298) );
 a63299a <=( a63298a  and  a63295a );
 a63300a <=( a63299a  and  a63292a );
 a63304a <=( A167  and  (not A168) );
 a63305a <=( A169  and  a63304a );
 a63308a <=( A199  and  (not A166) );
 a63311a <=( A201  and  (not A200) );
 a63312a <=( a63311a  and  a63308a );
 a63313a <=( a63312a  and  a63305a );
 a63316a <=( A232  and  A203 );
 a63319a <=( A265  and  A233 );
 a63320a <=( a63319a  and  a63316a );
 a63323a <=( (not A269)  and  (not A268) );
 a63326a <=( A299  and  (not A298) );
 a63327a <=( a63326a  and  a63323a );
 a63328a <=( a63327a  and  a63320a );
 a63332a <=( A167  and  (not A168) );
 a63333a <=( A169  and  a63332a );
 a63336a <=( A199  and  (not A166) );
 a63339a <=( A201  and  (not A200) );
 a63340a <=( a63339a  and  a63336a );
 a63341a <=( a63340a  and  a63333a );
 a63344a <=( (not A233)  and  A203 );
 a63347a <=( (not A236)  and  (not A235) );
 a63348a <=( a63347a  and  a63344a );
 a63351a <=( A266  and  A265 );
 a63354a <=( A299  and  (not A298) );
 a63355a <=( a63354a  and  a63351a );
 a63356a <=( a63355a  and  a63348a );
 a63360a <=( A167  and  (not A168) );
 a63361a <=( A169  and  a63360a );
 a63364a <=( A199  and  (not A166) );
 a63367a <=( A201  and  (not A200) );
 a63368a <=( a63367a  and  a63364a );
 a63369a <=( a63368a  and  a63361a );
 a63372a <=( (not A233)  and  A203 );
 a63375a <=( (not A236)  and  (not A235) );
 a63376a <=( a63375a  and  a63372a );
 a63379a <=( (not A267)  and  (not A266) );
 a63382a <=( A299  and  (not A298) );
 a63383a <=( a63382a  and  a63379a );
 a63384a <=( a63383a  and  a63376a );
 a63388a <=( A167  and  (not A168) );
 a63389a <=( A169  and  a63388a );
 a63392a <=( A199  and  (not A166) );
 a63395a <=( A201  and  (not A200) );
 a63396a <=( a63395a  and  a63392a );
 a63397a <=( a63396a  and  a63389a );
 a63400a <=( (not A233)  and  A203 );
 a63403a <=( (not A236)  and  (not A235) );
 a63404a <=( a63403a  and  a63400a );
 a63407a <=( (not A266)  and  (not A265) );
 a63410a <=( A299  and  (not A298) );
 a63411a <=( a63410a  and  a63407a );
 a63412a <=( a63411a  and  a63404a );
 a63416a <=( A167  and  (not A168) );
 a63417a <=( A169  and  a63416a );
 a63420a <=( A199  and  (not A166) );
 a63423a <=( A201  and  (not A200) );
 a63424a <=( a63423a  and  a63420a );
 a63425a <=( a63424a  and  a63417a );
 a63428a <=( (not A233)  and  A203 );
 a63431a <=( (not A266)  and  (not A234) );
 a63432a <=( a63431a  and  a63428a );
 a63435a <=( (not A269)  and  (not A268) );
 a63438a <=( A299  and  (not A298) );
 a63439a <=( a63438a  and  a63435a );
 a63440a <=( a63439a  and  a63432a );
 a63444a <=( A167  and  (not A168) );
 a63445a <=( A169  and  a63444a );
 a63448a <=( A199  and  (not A166) );
 a63451a <=( A201  and  (not A200) );
 a63452a <=( a63451a  and  a63448a );
 a63453a <=( a63452a  and  a63445a );
 a63456a <=( A232  and  A203 );
 a63459a <=( A234  and  (not A233) );
 a63460a <=( a63459a  and  a63456a );
 a63463a <=( A298  and  A235 );
 a63466a <=( (not A302)  and  (not A301) );
 a63467a <=( a63466a  and  a63463a );
 a63468a <=( a63467a  and  a63460a );
 a63472a <=( A167  and  (not A168) );
 a63473a <=( A169  and  a63472a );
 a63476a <=( A199  and  (not A166) );
 a63479a <=( A201  and  (not A200) );
 a63480a <=( a63479a  and  a63476a );
 a63481a <=( a63480a  and  a63473a );
 a63484a <=( A232  and  A203 );
 a63487a <=( A234  and  (not A233) );
 a63488a <=( a63487a  and  a63484a );
 a63491a <=( A298  and  A236 );
 a63494a <=( (not A302)  and  (not A301) );
 a63495a <=( a63494a  and  a63491a );
 a63496a <=( a63495a  and  a63488a );
 a63500a <=( A167  and  (not A168) );
 a63501a <=( A169  and  a63500a );
 a63504a <=( A199  and  (not A166) );
 a63507a <=( A201  and  (not A200) );
 a63508a <=( a63507a  and  a63504a );
 a63509a <=( a63508a  and  a63501a );
 a63512a <=( (not A232)  and  A203 );
 a63515a <=( (not A266)  and  (not A233) );
 a63516a <=( a63515a  and  a63512a );
 a63519a <=( (not A269)  and  (not A268) );
 a63522a <=( A299  and  (not A298) );
 a63523a <=( a63522a  and  a63519a );
 a63524a <=( a63523a  and  a63516a );
 a63528a <=( (not A167)  and  (not A168) );
 a63529a <=( A169  and  a63528a );
 a63532a <=( (not A199)  and  A166 );
 a63535a <=( A232  and  A200 );
 a63536a <=( a63535a  and  a63532a );
 a63537a <=( a63536a  and  a63529a );
 a63540a <=( A265  and  A233 );
 a63543a <=( (not A269)  and  (not A268) );
 a63544a <=( a63543a  and  a63540a );
 a63547a <=( (not A299)  and  A298 );
 a63550a <=( A301  and  A300 );
 a63551a <=( a63550a  and  a63547a );
 a63552a <=( a63551a  and  a63544a );
 a63556a <=( (not A167)  and  (not A168) );
 a63557a <=( A169  and  a63556a );
 a63560a <=( (not A199)  and  A166 );
 a63563a <=( A232  and  A200 );
 a63564a <=( a63563a  and  a63560a );
 a63565a <=( a63564a  and  a63557a );
 a63568a <=( A265  and  A233 );
 a63571a <=( (not A269)  and  (not A268) );
 a63572a <=( a63571a  and  a63568a );
 a63575a <=( (not A299)  and  A298 );
 a63578a <=( A302  and  A300 );
 a63579a <=( a63578a  and  a63575a );
 a63580a <=( a63579a  and  a63572a );
 a63584a <=( (not A167)  and  (not A168) );
 a63585a <=( A169  and  a63584a );
 a63588a <=( (not A199)  and  A166 );
 a63591a <=( (not A233)  and  A200 );
 a63592a <=( a63591a  and  a63588a );
 a63593a <=( a63592a  and  a63585a );
 a63596a <=( (not A236)  and  (not A235) );
 a63599a <=( A266  and  A265 );
 a63600a <=( a63599a  and  a63596a );
 a63603a <=( (not A299)  and  A298 );
 a63606a <=( A301  and  A300 );
 a63607a <=( a63606a  and  a63603a );
 a63608a <=( a63607a  and  a63600a );
 a63612a <=( (not A167)  and  (not A168) );
 a63613a <=( A169  and  a63612a );
 a63616a <=( (not A199)  and  A166 );
 a63619a <=( (not A233)  and  A200 );
 a63620a <=( a63619a  and  a63616a );
 a63621a <=( a63620a  and  a63613a );
 a63624a <=( (not A236)  and  (not A235) );
 a63627a <=( A266  and  A265 );
 a63628a <=( a63627a  and  a63624a );
 a63631a <=( (not A299)  and  A298 );
 a63634a <=( A302  and  A300 );
 a63635a <=( a63634a  and  a63631a );
 a63636a <=( a63635a  and  a63628a );
 a63640a <=( (not A167)  and  (not A168) );
 a63641a <=( A169  and  a63640a );
 a63644a <=( (not A199)  and  A166 );
 a63647a <=( (not A233)  and  A200 );
 a63648a <=( a63647a  and  a63644a );
 a63649a <=( a63648a  and  a63641a );
 a63652a <=( (not A236)  and  (not A235) );
 a63655a <=( (not A267)  and  (not A266) );
 a63656a <=( a63655a  and  a63652a );
 a63659a <=( (not A299)  and  A298 );
 a63662a <=( A301  and  A300 );
 a63663a <=( a63662a  and  a63659a );
 a63664a <=( a63663a  and  a63656a );
 a63668a <=( (not A167)  and  (not A168) );
 a63669a <=( A169  and  a63668a );
 a63672a <=( (not A199)  and  A166 );
 a63675a <=( (not A233)  and  A200 );
 a63676a <=( a63675a  and  a63672a );
 a63677a <=( a63676a  and  a63669a );
 a63680a <=( (not A236)  and  (not A235) );
 a63683a <=( (not A267)  and  (not A266) );
 a63684a <=( a63683a  and  a63680a );
 a63687a <=( (not A299)  and  A298 );
 a63690a <=( A302  and  A300 );
 a63691a <=( a63690a  and  a63687a );
 a63692a <=( a63691a  and  a63684a );
 a63696a <=( (not A167)  and  (not A168) );
 a63697a <=( A169  and  a63696a );
 a63700a <=( (not A199)  and  A166 );
 a63703a <=( (not A233)  and  A200 );
 a63704a <=( a63703a  and  a63700a );
 a63705a <=( a63704a  and  a63697a );
 a63708a <=( (not A236)  and  (not A235) );
 a63711a <=( (not A266)  and  (not A265) );
 a63712a <=( a63711a  and  a63708a );
 a63715a <=( (not A299)  and  A298 );
 a63718a <=( A301  and  A300 );
 a63719a <=( a63718a  and  a63715a );
 a63720a <=( a63719a  and  a63712a );
 a63724a <=( (not A167)  and  (not A168) );
 a63725a <=( A169  and  a63724a );
 a63728a <=( (not A199)  and  A166 );
 a63731a <=( (not A233)  and  A200 );
 a63732a <=( a63731a  and  a63728a );
 a63733a <=( a63732a  and  a63725a );
 a63736a <=( (not A236)  and  (not A235) );
 a63739a <=( (not A266)  and  (not A265) );
 a63740a <=( a63739a  and  a63736a );
 a63743a <=( (not A299)  and  A298 );
 a63746a <=( A302  and  A300 );
 a63747a <=( a63746a  and  a63743a );
 a63748a <=( a63747a  and  a63740a );
 a63752a <=( (not A167)  and  (not A168) );
 a63753a <=( A169  and  a63752a );
 a63756a <=( (not A199)  and  A166 );
 a63759a <=( (not A233)  and  A200 );
 a63760a <=( a63759a  and  a63756a );
 a63761a <=( a63760a  and  a63753a );
 a63764a <=( (not A266)  and  (not A234) );
 a63767a <=( (not A269)  and  (not A268) );
 a63768a <=( a63767a  and  a63764a );
 a63771a <=( (not A299)  and  A298 );
 a63774a <=( A301  and  A300 );
 a63775a <=( a63774a  and  a63771a );
 a63776a <=( a63775a  and  a63768a );
 a63780a <=( (not A167)  and  (not A168) );
 a63781a <=( A169  and  a63780a );
 a63784a <=( (not A199)  and  A166 );
 a63787a <=( (not A233)  and  A200 );
 a63788a <=( a63787a  and  a63784a );
 a63789a <=( a63788a  and  a63781a );
 a63792a <=( (not A266)  and  (not A234) );
 a63795a <=( (not A269)  and  (not A268) );
 a63796a <=( a63795a  and  a63792a );
 a63799a <=( (not A299)  and  A298 );
 a63802a <=( A302  and  A300 );
 a63803a <=( a63802a  and  a63799a );
 a63804a <=( a63803a  and  a63796a );
 a63808a <=( (not A167)  and  (not A168) );
 a63809a <=( A169  and  a63808a );
 a63812a <=( (not A199)  and  A166 );
 a63815a <=( (not A232)  and  A200 );
 a63816a <=( a63815a  and  a63812a );
 a63817a <=( a63816a  and  a63809a );
 a63820a <=( (not A266)  and  (not A233) );
 a63823a <=( (not A269)  and  (not A268) );
 a63824a <=( a63823a  and  a63820a );
 a63827a <=( (not A299)  and  A298 );
 a63830a <=( A301  and  A300 );
 a63831a <=( a63830a  and  a63827a );
 a63832a <=( a63831a  and  a63824a );
 a63836a <=( (not A167)  and  (not A168) );
 a63837a <=( A169  and  a63836a );
 a63840a <=( (not A199)  and  A166 );
 a63843a <=( (not A232)  and  A200 );
 a63844a <=( a63843a  and  a63840a );
 a63845a <=( a63844a  and  a63837a );
 a63848a <=( (not A266)  and  (not A233) );
 a63851a <=( (not A269)  and  (not A268) );
 a63852a <=( a63851a  and  a63848a );
 a63855a <=( (not A299)  and  A298 );
 a63858a <=( A302  and  A300 );
 a63859a <=( a63858a  and  a63855a );
 a63860a <=( a63859a  and  a63852a );
 a63864a <=( (not A167)  and  (not A168) );
 a63865a <=( A169  and  a63864a );
 a63868a <=( A199  and  A166 );
 a63871a <=( A201  and  (not A200) );
 a63872a <=( a63871a  and  a63868a );
 a63873a <=( a63872a  and  a63865a );
 a63876a <=( A232  and  A202 );
 a63879a <=( A265  and  A233 );
 a63880a <=( a63879a  and  a63876a );
 a63883a <=( (not A269)  and  (not A268) );
 a63886a <=( A299  and  (not A298) );
 a63887a <=( a63886a  and  a63883a );
 a63888a <=( a63887a  and  a63880a );
 a63892a <=( (not A167)  and  (not A168) );
 a63893a <=( A169  and  a63892a );
 a63896a <=( A199  and  A166 );
 a63899a <=( A201  and  (not A200) );
 a63900a <=( a63899a  and  a63896a );
 a63901a <=( a63900a  and  a63893a );
 a63904a <=( (not A233)  and  A202 );
 a63907a <=( (not A236)  and  (not A235) );
 a63908a <=( a63907a  and  a63904a );
 a63911a <=( A266  and  A265 );
 a63914a <=( A299  and  (not A298) );
 a63915a <=( a63914a  and  a63911a );
 a63916a <=( a63915a  and  a63908a );
 a63920a <=( (not A167)  and  (not A168) );
 a63921a <=( A169  and  a63920a );
 a63924a <=( A199  and  A166 );
 a63927a <=( A201  and  (not A200) );
 a63928a <=( a63927a  and  a63924a );
 a63929a <=( a63928a  and  a63921a );
 a63932a <=( (not A233)  and  A202 );
 a63935a <=( (not A236)  and  (not A235) );
 a63936a <=( a63935a  and  a63932a );
 a63939a <=( (not A267)  and  (not A266) );
 a63942a <=( A299  and  (not A298) );
 a63943a <=( a63942a  and  a63939a );
 a63944a <=( a63943a  and  a63936a );
 a63948a <=( (not A167)  and  (not A168) );
 a63949a <=( A169  and  a63948a );
 a63952a <=( A199  and  A166 );
 a63955a <=( A201  and  (not A200) );
 a63956a <=( a63955a  and  a63952a );
 a63957a <=( a63956a  and  a63949a );
 a63960a <=( (not A233)  and  A202 );
 a63963a <=( (not A236)  and  (not A235) );
 a63964a <=( a63963a  and  a63960a );
 a63967a <=( (not A266)  and  (not A265) );
 a63970a <=( A299  and  (not A298) );
 a63971a <=( a63970a  and  a63967a );
 a63972a <=( a63971a  and  a63964a );
 a63976a <=( (not A167)  and  (not A168) );
 a63977a <=( A169  and  a63976a );
 a63980a <=( A199  and  A166 );
 a63983a <=( A201  and  (not A200) );
 a63984a <=( a63983a  and  a63980a );
 a63985a <=( a63984a  and  a63977a );
 a63988a <=( (not A233)  and  A202 );
 a63991a <=( (not A266)  and  (not A234) );
 a63992a <=( a63991a  and  a63988a );
 a63995a <=( (not A269)  and  (not A268) );
 a63998a <=( A299  and  (not A298) );
 a63999a <=( a63998a  and  a63995a );
 a64000a <=( a63999a  and  a63992a );
 a64004a <=( (not A167)  and  (not A168) );
 a64005a <=( A169  and  a64004a );
 a64008a <=( A199  and  A166 );
 a64011a <=( A201  and  (not A200) );
 a64012a <=( a64011a  and  a64008a );
 a64013a <=( a64012a  and  a64005a );
 a64016a <=( A232  and  A202 );
 a64019a <=( A234  and  (not A233) );
 a64020a <=( a64019a  and  a64016a );
 a64023a <=( A298  and  A235 );
 a64026a <=( (not A302)  and  (not A301) );
 a64027a <=( a64026a  and  a64023a );
 a64028a <=( a64027a  and  a64020a );
 a64032a <=( (not A167)  and  (not A168) );
 a64033a <=( A169  and  a64032a );
 a64036a <=( A199  and  A166 );
 a64039a <=( A201  and  (not A200) );
 a64040a <=( a64039a  and  a64036a );
 a64041a <=( a64040a  and  a64033a );
 a64044a <=( A232  and  A202 );
 a64047a <=( A234  and  (not A233) );
 a64048a <=( a64047a  and  a64044a );
 a64051a <=( A298  and  A236 );
 a64054a <=( (not A302)  and  (not A301) );
 a64055a <=( a64054a  and  a64051a );
 a64056a <=( a64055a  and  a64048a );
 a64060a <=( (not A167)  and  (not A168) );
 a64061a <=( A169  and  a64060a );
 a64064a <=( A199  and  A166 );
 a64067a <=( A201  and  (not A200) );
 a64068a <=( a64067a  and  a64064a );
 a64069a <=( a64068a  and  a64061a );
 a64072a <=( (not A232)  and  A202 );
 a64075a <=( (not A266)  and  (not A233) );
 a64076a <=( a64075a  and  a64072a );
 a64079a <=( (not A269)  and  (not A268) );
 a64082a <=( A299  and  (not A298) );
 a64083a <=( a64082a  and  a64079a );
 a64084a <=( a64083a  and  a64076a );
 a64088a <=( (not A167)  and  (not A168) );
 a64089a <=( A169  and  a64088a );
 a64092a <=( A199  and  A166 );
 a64095a <=( A201  and  (not A200) );
 a64096a <=( a64095a  and  a64092a );
 a64097a <=( a64096a  and  a64089a );
 a64100a <=( A232  and  A203 );
 a64103a <=( A265  and  A233 );
 a64104a <=( a64103a  and  a64100a );
 a64107a <=( (not A269)  and  (not A268) );
 a64110a <=( A299  and  (not A298) );
 a64111a <=( a64110a  and  a64107a );
 a64112a <=( a64111a  and  a64104a );
 a64116a <=( (not A167)  and  (not A168) );
 a64117a <=( A169  and  a64116a );
 a64120a <=( A199  and  A166 );
 a64123a <=( A201  and  (not A200) );
 a64124a <=( a64123a  and  a64120a );
 a64125a <=( a64124a  and  a64117a );
 a64128a <=( (not A233)  and  A203 );
 a64131a <=( (not A236)  and  (not A235) );
 a64132a <=( a64131a  and  a64128a );
 a64135a <=( A266  and  A265 );
 a64138a <=( A299  and  (not A298) );
 a64139a <=( a64138a  and  a64135a );
 a64140a <=( a64139a  and  a64132a );
 a64144a <=( (not A167)  and  (not A168) );
 a64145a <=( A169  and  a64144a );
 a64148a <=( A199  and  A166 );
 a64151a <=( A201  and  (not A200) );
 a64152a <=( a64151a  and  a64148a );
 a64153a <=( a64152a  and  a64145a );
 a64156a <=( (not A233)  and  A203 );
 a64159a <=( (not A236)  and  (not A235) );
 a64160a <=( a64159a  and  a64156a );
 a64163a <=( (not A267)  and  (not A266) );
 a64166a <=( A299  and  (not A298) );
 a64167a <=( a64166a  and  a64163a );
 a64168a <=( a64167a  and  a64160a );
 a64172a <=( (not A167)  and  (not A168) );
 a64173a <=( A169  and  a64172a );
 a64176a <=( A199  and  A166 );
 a64179a <=( A201  and  (not A200) );
 a64180a <=( a64179a  and  a64176a );
 a64181a <=( a64180a  and  a64173a );
 a64184a <=( (not A233)  and  A203 );
 a64187a <=( (not A236)  and  (not A235) );
 a64188a <=( a64187a  and  a64184a );
 a64191a <=( (not A266)  and  (not A265) );
 a64194a <=( A299  and  (not A298) );
 a64195a <=( a64194a  and  a64191a );
 a64196a <=( a64195a  and  a64188a );
 a64200a <=( (not A167)  and  (not A168) );
 a64201a <=( A169  and  a64200a );
 a64204a <=( A199  and  A166 );
 a64207a <=( A201  and  (not A200) );
 a64208a <=( a64207a  and  a64204a );
 a64209a <=( a64208a  and  a64201a );
 a64212a <=( (not A233)  and  A203 );
 a64215a <=( (not A266)  and  (not A234) );
 a64216a <=( a64215a  and  a64212a );
 a64219a <=( (not A269)  and  (not A268) );
 a64222a <=( A299  and  (not A298) );
 a64223a <=( a64222a  and  a64219a );
 a64224a <=( a64223a  and  a64216a );
 a64228a <=( (not A167)  and  (not A168) );
 a64229a <=( A169  and  a64228a );
 a64232a <=( A199  and  A166 );
 a64235a <=( A201  and  (not A200) );
 a64236a <=( a64235a  and  a64232a );
 a64237a <=( a64236a  and  a64229a );
 a64240a <=( A232  and  A203 );
 a64243a <=( A234  and  (not A233) );
 a64244a <=( a64243a  and  a64240a );
 a64247a <=( A298  and  A235 );
 a64250a <=( (not A302)  and  (not A301) );
 a64251a <=( a64250a  and  a64247a );
 a64252a <=( a64251a  and  a64244a );
 a64256a <=( (not A167)  and  (not A168) );
 a64257a <=( A169  and  a64256a );
 a64260a <=( A199  and  A166 );
 a64263a <=( A201  and  (not A200) );
 a64264a <=( a64263a  and  a64260a );
 a64265a <=( a64264a  and  a64257a );
 a64268a <=( A232  and  A203 );
 a64271a <=( A234  and  (not A233) );
 a64272a <=( a64271a  and  a64268a );
 a64275a <=( A298  and  A236 );
 a64278a <=( (not A302)  and  (not A301) );
 a64279a <=( a64278a  and  a64275a );
 a64280a <=( a64279a  and  a64272a );
 a64284a <=( (not A167)  and  (not A168) );
 a64285a <=( A169  and  a64284a );
 a64288a <=( A199  and  A166 );
 a64291a <=( A201  and  (not A200) );
 a64292a <=( a64291a  and  a64288a );
 a64293a <=( a64292a  and  a64285a );
 a64296a <=( (not A232)  and  A203 );
 a64299a <=( (not A266)  and  (not A233) );
 a64300a <=( a64299a  and  a64296a );
 a64303a <=( (not A269)  and  (not A268) );
 a64306a <=( A299  and  (not A298) );
 a64307a <=( a64306a  and  a64303a );
 a64308a <=( a64307a  and  a64300a );
 a64312a <=( (not A168)  and  A169 );
 a64313a <=( A170  and  a64312a );
 a64316a <=( (not A200)  and  A199 );
 a64319a <=( A202  and  A201 );
 a64320a <=( a64319a  and  a64316a );
 a64321a <=( a64320a  and  a64313a );
 a64324a <=( A233  and  A232 );
 a64327a <=( (not A267)  and  A265 );
 a64328a <=( a64327a  and  a64324a );
 a64331a <=( (not A299)  and  A298 );
 a64334a <=( A301  and  A300 );
 a64335a <=( a64334a  and  a64331a );
 a64336a <=( a64335a  and  a64328a );
 a64340a <=( (not A168)  and  A169 );
 a64341a <=( A170  and  a64340a );
 a64344a <=( (not A200)  and  A199 );
 a64347a <=( A202  and  A201 );
 a64348a <=( a64347a  and  a64344a );
 a64349a <=( a64348a  and  a64341a );
 a64352a <=( A233  and  A232 );
 a64355a <=( (not A267)  and  A265 );
 a64356a <=( a64355a  and  a64352a );
 a64359a <=( (not A299)  and  A298 );
 a64362a <=( A302  and  A300 );
 a64363a <=( a64362a  and  a64359a );
 a64364a <=( a64363a  and  a64356a );
 a64368a <=( (not A168)  and  A169 );
 a64369a <=( A170  and  a64368a );
 a64372a <=( (not A200)  and  A199 );
 a64375a <=( A202  and  A201 );
 a64376a <=( a64375a  and  a64372a );
 a64377a <=( a64376a  and  a64369a );
 a64380a <=( A233  and  A232 );
 a64383a <=( A266  and  A265 );
 a64384a <=( a64383a  and  a64380a );
 a64387a <=( (not A299)  and  A298 );
 a64390a <=( A301  and  A300 );
 a64391a <=( a64390a  and  a64387a );
 a64392a <=( a64391a  and  a64384a );
 a64396a <=( (not A168)  and  A169 );
 a64397a <=( A170  and  a64396a );
 a64400a <=( (not A200)  and  A199 );
 a64403a <=( A202  and  A201 );
 a64404a <=( a64403a  and  a64400a );
 a64405a <=( a64404a  and  a64397a );
 a64408a <=( A233  and  A232 );
 a64411a <=( A266  and  A265 );
 a64412a <=( a64411a  and  a64408a );
 a64415a <=( (not A299)  and  A298 );
 a64418a <=( A302  and  A300 );
 a64419a <=( a64418a  and  a64415a );
 a64420a <=( a64419a  and  a64412a );
 a64424a <=( (not A168)  and  A169 );
 a64425a <=( A170  and  a64424a );
 a64428a <=( (not A200)  and  A199 );
 a64431a <=( A202  and  A201 );
 a64432a <=( a64431a  and  a64428a );
 a64433a <=( a64432a  and  a64425a );
 a64436a <=( A233  and  A232 );
 a64439a <=( (not A266)  and  (not A265) );
 a64440a <=( a64439a  and  a64436a );
 a64443a <=( (not A299)  and  A298 );
 a64446a <=( A301  and  A300 );
 a64447a <=( a64446a  and  a64443a );
 a64448a <=( a64447a  and  a64440a );
 a64452a <=( (not A168)  and  A169 );
 a64453a <=( A170  and  a64452a );
 a64456a <=( (not A200)  and  A199 );
 a64459a <=( A202  and  A201 );
 a64460a <=( a64459a  and  a64456a );
 a64461a <=( a64460a  and  a64453a );
 a64464a <=( A233  and  A232 );
 a64467a <=( (not A266)  and  (not A265) );
 a64468a <=( a64467a  and  a64464a );
 a64471a <=( (not A299)  and  A298 );
 a64474a <=( A302  and  A300 );
 a64475a <=( a64474a  and  a64471a );
 a64476a <=( a64475a  and  a64468a );
 a64480a <=( (not A168)  and  A169 );
 a64481a <=( A170  and  a64480a );
 a64484a <=( (not A200)  and  A199 );
 a64487a <=( A202  and  A201 );
 a64488a <=( a64487a  and  a64484a );
 a64489a <=( a64488a  and  a64481a );
 a64492a <=( (not A235)  and  (not A233) );
 a64495a <=( (not A266)  and  (not A236) );
 a64496a <=( a64495a  and  a64492a );
 a64499a <=( (not A269)  and  (not A268) );
 a64502a <=( A299  and  (not A298) );
 a64503a <=( a64502a  and  a64499a );
 a64504a <=( a64503a  and  a64496a );
 a64508a <=( (not A168)  and  A169 );
 a64509a <=( A170  and  a64508a );
 a64512a <=( (not A200)  and  A199 );
 a64515a <=( A202  and  A201 );
 a64516a <=( a64515a  and  a64512a );
 a64517a <=( a64516a  and  a64509a );
 a64520a <=( (not A234)  and  (not A233) );
 a64523a <=( A266  and  A265 );
 a64524a <=( a64523a  and  a64520a );
 a64527a <=( (not A299)  and  A298 );
 a64530a <=( A301  and  A300 );
 a64531a <=( a64530a  and  a64527a );
 a64532a <=( a64531a  and  a64524a );
 a64536a <=( (not A168)  and  A169 );
 a64537a <=( A170  and  a64536a );
 a64540a <=( (not A200)  and  A199 );
 a64543a <=( A202  and  A201 );
 a64544a <=( a64543a  and  a64540a );
 a64545a <=( a64544a  and  a64537a );
 a64548a <=( (not A234)  and  (not A233) );
 a64551a <=( A266  and  A265 );
 a64552a <=( a64551a  and  a64548a );
 a64555a <=( (not A299)  and  A298 );
 a64558a <=( A302  and  A300 );
 a64559a <=( a64558a  and  a64555a );
 a64560a <=( a64559a  and  a64552a );
 a64564a <=( (not A168)  and  A169 );
 a64565a <=( A170  and  a64564a );
 a64568a <=( (not A200)  and  A199 );
 a64571a <=( A202  and  A201 );
 a64572a <=( a64571a  and  a64568a );
 a64573a <=( a64572a  and  a64565a );
 a64576a <=( (not A233)  and  A232 );
 a64579a <=( A235  and  A234 );
 a64580a <=( a64579a  and  a64576a );
 a64583a <=( (not A266)  and  A265 );
 a64586a <=( A268  and  A267 );
 a64587a <=( a64586a  and  a64583a );
 a64588a <=( a64587a  and  a64580a );
 a64592a <=( (not A168)  and  A169 );
 a64593a <=( A170  and  a64592a );
 a64596a <=( (not A200)  and  A199 );
 a64599a <=( A202  and  A201 );
 a64600a <=( a64599a  and  a64596a );
 a64601a <=( a64600a  and  a64593a );
 a64604a <=( (not A233)  and  A232 );
 a64607a <=( A235  and  A234 );
 a64608a <=( a64607a  and  a64604a );
 a64611a <=( (not A266)  and  A265 );
 a64614a <=( A269  and  A267 );
 a64615a <=( a64614a  and  a64611a );
 a64616a <=( a64615a  and  a64608a );
 a64620a <=( (not A168)  and  A169 );
 a64621a <=( A170  and  a64620a );
 a64624a <=( (not A200)  and  A199 );
 a64627a <=( A202  and  A201 );
 a64628a <=( a64627a  and  a64624a );
 a64629a <=( a64628a  and  a64621a );
 a64632a <=( (not A233)  and  A232 );
 a64635a <=( A236  and  A234 );
 a64636a <=( a64635a  and  a64632a );
 a64639a <=( (not A266)  and  A265 );
 a64642a <=( A268  and  A267 );
 a64643a <=( a64642a  and  a64639a );
 a64644a <=( a64643a  and  a64636a );
 a64648a <=( (not A168)  and  A169 );
 a64649a <=( A170  and  a64648a );
 a64652a <=( (not A200)  and  A199 );
 a64655a <=( A202  and  A201 );
 a64656a <=( a64655a  and  a64652a );
 a64657a <=( a64656a  and  a64649a );
 a64660a <=( (not A233)  and  A232 );
 a64663a <=( A236  and  A234 );
 a64664a <=( a64663a  and  a64660a );
 a64667a <=( (not A266)  and  A265 );
 a64670a <=( A269  and  A267 );
 a64671a <=( a64670a  and  a64667a );
 a64672a <=( a64671a  and  a64664a );
 a64676a <=( (not A168)  and  A169 );
 a64677a <=( A170  and  a64676a );
 a64680a <=( (not A200)  and  A199 );
 a64683a <=( A202  and  A201 );
 a64684a <=( a64683a  and  a64680a );
 a64685a <=( a64684a  and  a64677a );
 a64688a <=( (not A233)  and  (not A232) );
 a64691a <=( A266  and  A265 );
 a64692a <=( a64691a  and  a64688a );
 a64695a <=( (not A299)  and  A298 );
 a64698a <=( A301  and  A300 );
 a64699a <=( a64698a  and  a64695a );
 a64700a <=( a64699a  and  a64692a );
 a64704a <=( (not A168)  and  A169 );
 a64705a <=( A170  and  a64704a );
 a64708a <=( (not A200)  and  A199 );
 a64711a <=( A202  and  A201 );
 a64712a <=( a64711a  and  a64708a );
 a64713a <=( a64712a  and  a64705a );
 a64716a <=( (not A233)  and  (not A232) );
 a64719a <=( A266  and  A265 );
 a64720a <=( a64719a  and  a64716a );
 a64723a <=( (not A299)  and  A298 );
 a64726a <=( A302  and  A300 );
 a64727a <=( a64726a  and  a64723a );
 a64728a <=( a64727a  and  a64720a );
 a64732a <=( (not A168)  and  A169 );
 a64733a <=( A170  and  a64732a );
 a64736a <=( (not A200)  and  A199 );
 a64739a <=( A203  and  A201 );
 a64740a <=( a64739a  and  a64736a );
 a64741a <=( a64740a  and  a64733a );
 a64744a <=( A233  and  A232 );
 a64747a <=( (not A267)  and  A265 );
 a64748a <=( a64747a  and  a64744a );
 a64751a <=( (not A299)  and  A298 );
 a64754a <=( A301  and  A300 );
 a64755a <=( a64754a  and  a64751a );
 a64756a <=( a64755a  and  a64748a );
 a64760a <=( (not A168)  and  A169 );
 a64761a <=( A170  and  a64760a );
 a64764a <=( (not A200)  and  A199 );
 a64767a <=( A203  and  A201 );
 a64768a <=( a64767a  and  a64764a );
 a64769a <=( a64768a  and  a64761a );
 a64772a <=( A233  and  A232 );
 a64775a <=( (not A267)  and  A265 );
 a64776a <=( a64775a  and  a64772a );
 a64779a <=( (not A299)  and  A298 );
 a64782a <=( A302  and  A300 );
 a64783a <=( a64782a  and  a64779a );
 a64784a <=( a64783a  and  a64776a );
 a64788a <=( (not A168)  and  A169 );
 a64789a <=( A170  and  a64788a );
 a64792a <=( (not A200)  and  A199 );
 a64795a <=( A203  and  A201 );
 a64796a <=( a64795a  and  a64792a );
 a64797a <=( a64796a  and  a64789a );
 a64800a <=( A233  and  A232 );
 a64803a <=( A266  and  A265 );
 a64804a <=( a64803a  and  a64800a );
 a64807a <=( (not A299)  and  A298 );
 a64810a <=( A301  and  A300 );
 a64811a <=( a64810a  and  a64807a );
 a64812a <=( a64811a  and  a64804a );
 a64816a <=( (not A168)  and  A169 );
 a64817a <=( A170  and  a64816a );
 a64820a <=( (not A200)  and  A199 );
 a64823a <=( A203  and  A201 );
 a64824a <=( a64823a  and  a64820a );
 a64825a <=( a64824a  and  a64817a );
 a64828a <=( A233  and  A232 );
 a64831a <=( A266  and  A265 );
 a64832a <=( a64831a  and  a64828a );
 a64835a <=( (not A299)  and  A298 );
 a64838a <=( A302  and  A300 );
 a64839a <=( a64838a  and  a64835a );
 a64840a <=( a64839a  and  a64832a );
 a64844a <=( (not A168)  and  A169 );
 a64845a <=( A170  and  a64844a );
 a64848a <=( (not A200)  and  A199 );
 a64851a <=( A203  and  A201 );
 a64852a <=( a64851a  and  a64848a );
 a64853a <=( a64852a  and  a64845a );
 a64856a <=( A233  and  A232 );
 a64859a <=( (not A266)  and  (not A265) );
 a64860a <=( a64859a  and  a64856a );
 a64863a <=( (not A299)  and  A298 );
 a64866a <=( A301  and  A300 );
 a64867a <=( a64866a  and  a64863a );
 a64868a <=( a64867a  and  a64860a );
 a64872a <=( (not A168)  and  A169 );
 a64873a <=( A170  and  a64872a );
 a64876a <=( (not A200)  and  A199 );
 a64879a <=( A203  and  A201 );
 a64880a <=( a64879a  and  a64876a );
 a64881a <=( a64880a  and  a64873a );
 a64884a <=( A233  and  A232 );
 a64887a <=( (not A266)  and  (not A265) );
 a64888a <=( a64887a  and  a64884a );
 a64891a <=( (not A299)  and  A298 );
 a64894a <=( A302  and  A300 );
 a64895a <=( a64894a  and  a64891a );
 a64896a <=( a64895a  and  a64888a );
 a64900a <=( (not A168)  and  A169 );
 a64901a <=( A170  and  a64900a );
 a64904a <=( (not A200)  and  A199 );
 a64907a <=( A203  and  A201 );
 a64908a <=( a64907a  and  a64904a );
 a64909a <=( a64908a  and  a64901a );
 a64912a <=( (not A235)  and  (not A233) );
 a64915a <=( (not A266)  and  (not A236) );
 a64916a <=( a64915a  and  a64912a );
 a64919a <=( (not A269)  and  (not A268) );
 a64922a <=( A299  and  (not A298) );
 a64923a <=( a64922a  and  a64919a );
 a64924a <=( a64923a  and  a64916a );
 a64928a <=( (not A168)  and  A169 );
 a64929a <=( A170  and  a64928a );
 a64932a <=( (not A200)  and  A199 );
 a64935a <=( A203  and  A201 );
 a64936a <=( a64935a  and  a64932a );
 a64937a <=( a64936a  and  a64929a );
 a64940a <=( (not A234)  and  (not A233) );
 a64943a <=( A266  and  A265 );
 a64944a <=( a64943a  and  a64940a );
 a64947a <=( (not A299)  and  A298 );
 a64950a <=( A301  and  A300 );
 a64951a <=( a64950a  and  a64947a );
 a64952a <=( a64951a  and  a64944a );
 a64956a <=( (not A168)  and  A169 );
 a64957a <=( A170  and  a64956a );
 a64960a <=( (not A200)  and  A199 );
 a64963a <=( A203  and  A201 );
 a64964a <=( a64963a  and  a64960a );
 a64965a <=( a64964a  and  a64957a );
 a64968a <=( (not A234)  and  (not A233) );
 a64971a <=( A266  and  A265 );
 a64972a <=( a64971a  and  a64968a );
 a64975a <=( (not A299)  and  A298 );
 a64978a <=( A302  and  A300 );
 a64979a <=( a64978a  and  a64975a );
 a64980a <=( a64979a  and  a64972a );
 a64984a <=( (not A168)  and  A169 );
 a64985a <=( A170  and  a64984a );
 a64988a <=( (not A200)  and  A199 );
 a64991a <=( A203  and  A201 );
 a64992a <=( a64991a  and  a64988a );
 a64993a <=( a64992a  and  a64985a );
 a64996a <=( (not A233)  and  A232 );
 a64999a <=( A235  and  A234 );
 a65000a <=( a64999a  and  a64996a );
 a65003a <=( (not A266)  and  A265 );
 a65006a <=( A268  and  A267 );
 a65007a <=( a65006a  and  a65003a );
 a65008a <=( a65007a  and  a65000a );
 a65012a <=( (not A168)  and  A169 );
 a65013a <=( A170  and  a65012a );
 a65016a <=( (not A200)  and  A199 );
 a65019a <=( A203  and  A201 );
 a65020a <=( a65019a  and  a65016a );
 a65021a <=( a65020a  and  a65013a );
 a65024a <=( (not A233)  and  A232 );
 a65027a <=( A235  and  A234 );
 a65028a <=( a65027a  and  a65024a );
 a65031a <=( (not A266)  and  A265 );
 a65034a <=( A269  and  A267 );
 a65035a <=( a65034a  and  a65031a );
 a65036a <=( a65035a  and  a65028a );
 a65040a <=( (not A168)  and  A169 );
 a65041a <=( A170  and  a65040a );
 a65044a <=( (not A200)  and  A199 );
 a65047a <=( A203  and  A201 );
 a65048a <=( a65047a  and  a65044a );
 a65049a <=( a65048a  and  a65041a );
 a65052a <=( (not A233)  and  A232 );
 a65055a <=( A236  and  A234 );
 a65056a <=( a65055a  and  a65052a );
 a65059a <=( (not A266)  and  A265 );
 a65062a <=( A268  and  A267 );
 a65063a <=( a65062a  and  a65059a );
 a65064a <=( a65063a  and  a65056a );
 a65068a <=( (not A168)  and  A169 );
 a65069a <=( A170  and  a65068a );
 a65072a <=( (not A200)  and  A199 );
 a65075a <=( A203  and  A201 );
 a65076a <=( a65075a  and  a65072a );
 a65077a <=( a65076a  and  a65069a );
 a65080a <=( (not A233)  and  A232 );
 a65083a <=( A236  and  A234 );
 a65084a <=( a65083a  and  a65080a );
 a65087a <=( (not A266)  and  A265 );
 a65090a <=( A269  and  A267 );
 a65091a <=( a65090a  and  a65087a );
 a65092a <=( a65091a  and  a65084a );
 a65096a <=( (not A168)  and  A169 );
 a65097a <=( A170  and  a65096a );
 a65100a <=( (not A200)  and  A199 );
 a65103a <=( A203  and  A201 );
 a65104a <=( a65103a  and  a65100a );
 a65105a <=( a65104a  and  a65097a );
 a65108a <=( (not A233)  and  (not A232) );
 a65111a <=( A266  and  A265 );
 a65112a <=( a65111a  and  a65108a );
 a65115a <=( (not A299)  and  A298 );
 a65118a <=( A301  and  A300 );
 a65119a <=( a65118a  and  a65115a );
 a65120a <=( a65119a  and  a65112a );
 a65124a <=( (not A168)  and  A169 );
 a65125a <=( A170  and  a65124a );
 a65128a <=( (not A200)  and  A199 );
 a65131a <=( A203  and  A201 );
 a65132a <=( a65131a  and  a65128a );
 a65133a <=( a65132a  and  a65125a );
 a65136a <=( (not A233)  and  (not A232) );
 a65139a <=( A266  and  A265 );
 a65140a <=( a65139a  and  a65136a );
 a65143a <=( (not A299)  and  A298 );
 a65146a <=( A302  and  A300 );
 a65147a <=( a65146a  and  a65143a );
 a65148a <=( a65147a  and  a65140a );
 a65152a <=( A167  and  A169 );
 a65153a <=( (not A170)  and  a65152a );
 a65156a <=( A199  and  A166 );
 a65159a <=( A232  and  A200 );
 a65160a <=( a65159a  and  a65156a );
 a65161a <=( a65160a  and  a65153a );
 a65164a <=( A265  and  A233 );
 a65167a <=( (not A269)  and  (not A268) );
 a65168a <=( a65167a  and  a65164a );
 a65171a <=( (not A299)  and  A298 );
 a65174a <=( A301  and  A300 );
 a65175a <=( a65174a  and  a65171a );
 a65176a <=( a65175a  and  a65168a );
 a65180a <=( A167  and  A169 );
 a65181a <=( (not A170)  and  a65180a );
 a65184a <=( A199  and  A166 );
 a65187a <=( A232  and  A200 );
 a65188a <=( a65187a  and  a65184a );
 a65189a <=( a65188a  and  a65181a );
 a65192a <=( A265  and  A233 );
 a65195a <=( (not A269)  and  (not A268) );
 a65196a <=( a65195a  and  a65192a );
 a65199a <=( (not A299)  and  A298 );
 a65202a <=( A302  and  A300 );
 a65203a <=( a65202a  and  a65199a );
 a65204a <=( a65203a  and  a65196a );
 a65208a <=( A167  and  A169 );
 a65209a <=( (not A170)  and  a65208a );
 a65212a <=( A199  and  A166 );
 a65215a <=( (not A233)  and  A200 );
 a65216a <=( a65215a  and  a65212a );
 a65217a <=( a65216a  and  a65209a );
 a65220a <=( (not A236)  and  (not A235) );
 a65223a <=( A266  and  A265 );
 a65224a <=( a65223a  and  a65220a );
 a65227a <=( (not A299)  and  A298 );
 a65230a <=( A301  and  A300 );
 a65231a <=( a65230a  and  a65227a );
 a65232a <=( a65231a  and  a65224a );
 a65236a <=( A167  and  A169 );
 a65237a <=( (not A170)  and  a65236a );
 a65240a <=( A199  and  A166 );
 a65243a <=( (not A233)  and  A200 );
 a65244a <=( a65243a  and  a65240a );
 a65245a <=( a65244a  and  a65237a );
 a65248a <=( (not A236)  and  (not A235) );
 a65251a <=( A266  and  A265 );
 a65252a <=( a65251a  and  a65248a );
 a65255a <=( (not A299)  and  A298 );
 a65258a <=( A302  and  A300 );
 a65259a <=( a65258a  and  a65255a );
 a65260a <=( a65259a  and  a65252a );
 a65264a <=( A167  and  A169 );
 a65265a <=( (not A170)  and  a65264a );
 a65268a <=( A199  and  A166 );
 a65271a <=( (not A233)  and  A200 );
 a65272a <=( a65271a  and  a65268a );
 a65273a <=( a65272a  and  a65265a );
 a65276a <=( (not A236)  and  (not A235) );
 a65279a <=( (not A267)  and  (not A266) );
 a65280a <=( a65279a  and  a65276a );
 a65283a <=( (not A299)  and  A298 );
 a65286a <=( A301  and  A300 );
 a65287a <=( a65286a  and  a65283a );
 a65288a <=( a65287a  and  a65280a );
 a65292a <=( A167  and  A169 );
 a65293a <=( (not A170)  and  a65292a );
 a65296a <=( A199  and  A166 );
 a65299a <=( (not A233)  and  A200 );
 a65300a <=( a65299a  and  a65296a );
 a65301a <=( a65300a  and  a65293a );
 a65304a <=( (not A236)  and  (not A235) );
 a65307a <=( (not A267)  and  (not A266) );
 a65308a <=( a65307a  and  a65304a );
 a65311a <=( (not A299)  and  A298 );
 a65314a <=( A302  and  A300 );
 a65315a <=( a65314a  and  a65311a );
 a65316a <=( a65315a  and  a65308a );
 a65320a <=( A167  and  A169 );
 a65321a <=( (not A170)  and  a65320a );
 a65324a <=( A199  and  A166 );
 a65327a <=( (not A233)  and  A200 );
 a65328a <=( a65327a  and  a65324a );
 a65329a <=( a65328a  and  a65321a );
 a65332a <=( (not A236)  and  (not A235) );
 a65335a <=( (not A266)  and  (not A265) );
 a65336a <=( a65335a  and  a65332a );
 a65339a <=( (not A299)  and  A298 );
 a65342a <=( A301  and  A300 );
 a65343a <=( a65342a  and  a65339a );
 a65344a <=( a65343a  and  a65336a );
 a65348a <=( A167  and  A169 );
 a65349a <=( (not A170)  and  a65348a );
 a65352a <=( A199  and  A166 );
 a65355a <=( (not A233)  and  A200 );
 a65356a <=( a65355a  and  a65352a );
 a65357a <=( a65356a  and  a65349a );
 a65360a <=( (not A236)  and  (not A235) );
 a65363a <=( (not A266)  and  (not A265) );
 a65364a <=( a65363a  and  a65360a );
 a65367a <=( (not A299)  and  A298 );
 a65370a <=( A302  and  A300 );
 a65371a <=( a65370a  and  a65367a );
 a65372a <=( a65371a  and  a65364a );
 a65376a <=( A167  and  A169 );
 a65377a <=( (not A170)  and  a65376a );
 a65380a <=( A199  and  A166 );
 a65383a <=( (not A233)  and  A200 );
 a65384a <=( a65383a  and  a65380a );
 a65385a <=( a65384a  and  a65377a );
 a65388a <=( (not A266)  and  (not A234) );
 a65391a <=( (not A269)  and  (not A268) );
 a65392a <=( a65391a  and  a65388a );
 a65395a <=( (not A299)  and  A298 );
 a65398a <=( A301  and  A300 );
 a65399a <=( a65398a  and  a65395a );
 a65400a <=( a65399a  and  a65392a );
 a65404a <=( A167  and  A169 );
 a65405a <=( (not A170)  and  a65404a );
 a65408a <=( A199  and  A166 );
 a65411a <=( (not A233)  and  A200 );
 a65412a <=( a65411a  and  a65408a );
 a65413a <=( a65412a  and  a65405a );
 a65416a <=( (not A266)  and  (not A234) );
 a65419a <=( (not A269)  and  (not A268) );
 a65420a <=( a65419a  and  a65416a );
 a65423a <=( (not A299)  and  A298 );
 a65426a <=( A302  and  A300 );
 a65427a <=( a65426a  and  a65423a );
 a65428a <=( a65427a  and  a65420a );
 a65432a <=( A167  and  A169 );
 a65433a <=( (not A170)  and  a65432a );
 a65436a <=( A199  and  A166 );
 a65439a <=( (not A232)  and  A200 );
 a65440a <=( a65439a  and  a65436a );
 a65441a <=( a65440a  and  a65433a );
 a65444a <=( (not A266)  and  (not A233) );
 a65447a <=( (not A269)  and  (not A268) );
 a65448a <=( a65447a  and  a65444a );
 a65451a <=( (not A299)  and  A298 );
 a65454a <=( A301  and  A300 );
 a65455a <=( a65454a  and  a65451a );
 a65456a <=( a65455a  and  a65448a );
 a65460a <=( A167  and  A169 );
 a65461a <=( (not A170)  and  a65460a );
 a65464a <=( A199  and  A166 );
 a65467a <=( (not A232)  and  A200 );
 a65468a <=( a65467a  and  a65464a );
 a65469a <=( a65468a  and  a65461a );
 a65472a <=( (not A266)  and  (not A233) );
 a65475a <=( (not A269)  and  (not A268) );
 a65476a <=( a65475a  and  a65472a );
 a65479a <=( (not A299)  and  A298 );
 a65482a <=( A302  and  A300 );
 a65483a <=( a65482a  and  a65479a );
 a65484a <=( a65483a  and  a65476a );
 a65488a <=( A167  and  A169 );
 a65489a <=( (not A170)  and  a65488a );
 a65492a <=( (not A200)  and  A166 );
 a65495a <=( (not A203)  and  (not A202) );
 a65496a <=( a65495a  and  a65492a );
 a65497a <=( a65496a  and  a65489a );
 a65500a <=( A233  and  A232 );
 a65503a <=( (not A267)  and  A265 );
 a65504a <=( a65503a  and  a65500a );
 a65507a <=( (not A299)  and  A298 );
 a65510a <=( A301  and  A300 );
 a65511a <=( a65510a  and  a65507a );
 a65512a <=( a65511a  and  a65504a );
 a65516a <=( A167  and  A169 );
 a65517a <=( (not A170)  and  a65516a );
 a65520a <=( (not A200)  and  A166 );
 a65523a <=( (not A203)  and  (not A202) );
 a65524a <=( a65523a  and  a65520a );
 a65525a <=( a65524a  and  a65517a );
 a65528a <=( A233  and  A232 );
 a65531a <=( (not A267)  and  A265 );
 a65532a <=( a65531a  and  a65528a );
 a65535a <=( (not A299)  and  A298 );
 a65538a <=( A302  and  A300 );
 a65539a <=( a65538a  and  a65535a );
 a65540a <=( a65539a  and  a65532a );
 a65544a <=( A167  and  A169 );
 a65545a <=( (not A170)  and  a65544a );
 a65548a <=( (not A200)  and  A166 );
 a65551a <=( (not A203)  and  (not A202) );
 a65552a <=( a65551a  and  a65548a );
 a65553a <=( a65552a  and  a65545a );
 a65556a <=( A233  and  A232 );
 a65559a <=( A266  and  A265 );
 a65560a <=( a65559a  and  a65556a );
 a65563a <=( (not A299)  and  A298 );
 a65566a <=( A301  and  A300 );
 a65567a <=( a65566a  and  a65563a );
 a65568a <=( a65567a  and  a65560a );
 a65572a <=( A167  and  A169 );
 a65573a <=( (not A170)  and  a65572a );
 a65576a <=( (not A200)  and  A166 );
 a65579a <=( (not A203)  and  (not A202) );
 a65580a <=( a65579a  and  a65576a );
 a65581a <=( a65580a  and  a65573a );
 a65584a <=( A233  and  A232 );
 a65587a <=( A266  and  A265 );
 a65588a <=( a65587a  and  a65584a );
 a65591a <=( (not A299)  and  A298 );
 a65594a <=( A302  and  A300 );
 a65595a <=( a65594a  and  a65591a );
 a65596a <=( a65595a  and  a65588a );
 a65600a <=( A167  and  A169 );
 a65601a <=( (not A170)  and  a65600a );
 a65604a <=( (not A200)  and  A166 );
 a65607a <=( (not A203)  and  (not A202) );
 a65608a <=( a65607a  and  a65604a );
 a65609a <=( a65608a  and  a65601a );
 a65612a <=( A233  and  A232 );
 a65615a <=( (not A266)  and  (not A265) );
 a65616a <=( a65615a  and  a65612a );
 a65619a <=( (not A299)  and  A298 );
 a65622a <=( A301  and  A300 );
 a65623a <=( a65622a  and  a65619a );
 a65624a <=( a65623a  and  a65616a );
 a65628a <=( A167  and  A169 );
 a65629a <=( (not A170)  and  a65628a );
 a65632a <=( (not A200)  and  A166 );
 a65635a <=( (not A203)  and  (not A202) );
 a65636a <=( a65635a  and  a65632a );
 a65637a <=( a65636a  and  a65629a );
 a65640a <=( A233  and  A232 );
 a65643a <=( (not A266)  and  (not A265) );
 a65644a <=( a65643a  and  a65640a );
 a65647a <=( (not A299)  and  A298 );
 a65650a <=( A302  and  A300 );
 a65651a <=( a65650a  and  a65647a );
 a65652a <=( a65651a  and  a65644a );
 a65656a <=( A167  and  A169 );
 a65657a <=( (not A170)  and  a65656a );
 a65660a <=( (not A200)  and  A166 );
 a65663a <=( (not A203)  and  (not A202) );
 a65664a <=( a65663a  and  a65660a );
 a65665a <=( a65664a  and  a65657a );
 a65668a <=( (not A235)  and  (not A233) );
 a65671a <=( (not A266)  and  (not A236) );
 a65672a <=( a65671a  and  a65668a );
 a65675a <=( (not A269)  and  (not A268) );
 a65678a <=( A299  and  (not A298) );
 a65679a <=( a65678a  and  a65675a );
 a65680a <=( a65679a  and  a65672a );
 a65684a <=( A167  and  A169 );
 a65685a <=( (not A170)  and  a65684a );
 a65688a <=( (not A200)  and  A166 );
 a65691a <=( (not A203)  and  (not A202) );
 a65692a <=( a65691a  and  a65688a );
 a65693a <=( a65692a  and  a65685a );
 a65696a <=( (not A234)  and  (not A233) );
 a65699a <=( A266  and  A265 );
 a65700a <=( a65699a  and  a65696a );
 a65703a <=( (not A299)  and  A298 );
 a65706a <=( A301  and  A300 );
 a65707a <=( a65706a  and  a65703a );
 a65708a <=( a65707a  and  a65700a );
 a65712a <=( A167  and  A169 );
 a65713a <=( (not A170)  and  a65712a );
 a65716a <=( (not A200)  and  A166 );
 a65719a <=( (not A203)  and  (not A202) );
 a65720a <=( a65719a  and  a65716a );
 a65721a <=( a65720a  and  a65713a );
 a65724a <=( (not A234)  and  (not A233) );
 a65727a <=( A266  and  A265 );
 a65728a <=( a65727a  and  a65724a );
 a65731a <=( (not A299)  and  A298 );
 a65734a <=( A302  and  A300 );
 a65735a <=( a65734a  and  a65731a );
 a65736a <=( a65735a  and  a65728a );
 a65740a <=( A167  and  A169 );
 a65741a <=( (not A170)  and  a65740a );
 a65744a <=( (not A200)  and  A166 );
 a65747a <=( (not A203)  and  (not A202) );
 a65748a <=( a65747a  and  a65744a );
 a65749a <=( a65748a  and  a65741a );
 a65752a <=( (not A234)  and  (not A233) );
 a65755a <=( (not A267)  and  (not A266) );
 a65756a <=( a65755a  and  a65752a );
 a65759a <=( (not A299)  and  A298 );
 a65762a <=( A301  and  A300 );
 a65763a <=( a65762a  and  a65759a );
 a65764a <=( a65763a  and  a65756a );
 a65768a <=( A167  and  A169 );
 a65769a <=( (not A170)  and  a65768a );
 a65772a <=( (not A200)  and  A166 );
 a65775a <=( (not A203)  and  (not A202) );
 a65776a <=( a65775a  and  a65772a );
 a65777a <=( a65776a  and  a65769a );
 a65780a <=( (not A234)  and  (not A233) );
 a65783a <=( (not A267)  and  (not A266) );
 a65784a <=( a65783a  and  a65780a );
 a65787a <=( (not A299)  and  A298 );
 a65790a <=( A302  and  A300 );
 a65791a <=( a65790a  and  a65787a );
 a65792a <=( a65791a  and  a65784a );
 a65796a <=( A167  and  A169 );
 a65797a <=( (not A170)  and  a65796a );
 a65800a <=( (not A200)  and  A166 );
 a65803a <=( (not A203)  and  (not A202) );
 a65804a <=( a65803a  and  a65800a );
 a65805a <=( a65804a  and  a65797a );
 a65808a <=( (not A234)  and  (not A233) );
 a65811a <=( (not A266)  and  (not A265) );
 a65812a <=( a65811a  and  a65808a );
 a65815a <=( (not A299)  and  A298 );
 a65818a <=( A301  and  A300 );
 a65819a <=( a65818a  and  a65815a );
 a65820a <=( a65819a  and  a65812a );
 a65824a <=( A167  and  A169 );
 a65825a <=( (not A170)  and  a65824a );
 a65828a <=( (not A200)  and  A166 );
 a65831a <=( (not A203)  and  (not A202) );
 a65832a <=( a65831a  and  a65828a );
 a65833a <=( a65832a  and  a65825a );
 a65836a <=( (not A234)  and  (not A233) );
 a65839a <=( (not A266)  and  (not A265) );
 a65840a <=( a65839a  and  a65836a );
 a65843a <=( (not A299)  and  A298 );
 a65846a <=( A302  and  A300 );
 a65847a <=( a65846a  and  a65843a );
 a65848a <=( a65847a  and  a65840a );
 a65852a <=( A167  and  A169 );
 a65853a <=( (not A170)  and  a65852a );
 a65856a <=( (not A200)  and  A166 );
 a65859a <=( (not A203)  and  (not A202) );
 a65860a <=( a65859a  and  a65856a );
 a65861a <=( a65860a  and  a65853a );
 a65864a <=( (not A233)  and  A232 );
 a65867a <=( A235  and  A234 );
 a65868a <=( a65867a  and  a65864a );
 a65871a <=( (not A266)  and  A265 );
 a65874a <=( A268  and  A267 );
 a65875a <=( a65874a  and  a65871a );
 a65876a <=( a65875a  and  a65868a );
 a65880a <=( A167  and  A169 );
 a65881a <=( (not A170)  and  a65880a );
 a65884a <=( (not A200)  and  A166 );
 a65887a <=( (not A203)  and  (not A202) );
 a65888a <=( a65887a  and  a65884a );
 a65889a <=( a65888a  and  a65881a );
 a65892a <=( (not A233)  and  A232 );
 a65895a <=( A235  and  A234 );
 a65896a <=( a65895a  and  a65892a );
 a65899a <=( (not A266)  and  A265 );
 a65902a <=( A269  and  A267 );
 a65903a <=( a65902a  and  a65899a );
 a65904a <=( a65903a  and  a65896a );
 a65908a <=( A167  and  A169 );
 a65909a <=( (not A170)  and  a65908a );
 a65912a <=( (not A200)  and  A166 );
 a65915a <=( (not A203)  and  (not A202) );
 a65916a <=( a65915a  and  a65912a );
 a65917a <=( a65916a  and  a65909a );
 a65920a <=( (not A233)  and  A232 );
 a65923a <=( A236  and  A234 );
 a65924a <=( a65923a  and  a65920a );
 a65927a <=( (not A266)  and  A265 );
 a65930a <=( A268  and  A267 );
 a65931a <=( a65930a  and  a65927a );
 a65932a <=( a65931a  and  a65924a );
 a65936a <=( A167  and  A169 );
 a65937a <=( (not A170)  and  a65936a );
 a65940a <=( (not A200)  and  A166 );
 a65943a <=( (not A203)  and  (not A202) );
 a65944a <=( a65943a  and  a65940a );
 a65945a <=( a65944a  and  a65937a );
 a65948a <=( (not A233)  and  A232 );
 a65951a <=( A236  and  A234 );
 a65952a <=( a65951a  and  a65948a );
 a65955a <=( (not A266)  and  A265 );
 a65958a <=( A269  and  A267 );
 a65959a <=( a65958a  and  a65955a );
 a65960a <=( a65959a  and  a65952a );
 a65964a <=( A167  and  A169 );
 a65965a <=( (not A170)  and  a65964a );
 a65968a <=( (not A200)  and  A166 );
 a65971a <=( (not A203)  and  (not A202) );
 a65972a <=( a65971a  and  a65968a );
 a65973a <=( a65972a  and  a65965a );
 a65976a <=( (not A233)  and  (not A232) );
 a65979a <=( A266  and  A265 );
 a65980a <=( a65979a  and  a65976a );
 a65983a <=( (not A299)  and  A298 );
 a65986a <=( A301  and  A300 );
 a65987a <=( a65986a  and  a65983a );
 a65988a <=( a65987a  and  a65980a );
 a65992a <=( A167  and  A169 );
 a65993a <=( (not A170)  and  a65992a );
 a65996a <=( (not A200)  and  A166 );
 a65999a <=( (not A203)  and  (not A202) );
 a66000a <=( a65999a  and  a65996a );
 a66001a <=( a66000a  and  a65993a );
 a66004a <=( (not A233)  and  (not A232) );
 a66007a <=( A266  and  A265 );
 a66008a <=( a66007a  and  a66004a );
 a66011a <=( (not A299)  and  A298 );
 a66014a <=( A302  and  A300 );
 a66015a <=( a66014a  and  a66011a );
 a66016a <=( a66015a  and  a66008a );
 a66020a <=( A167  and  A169 );
 a66021a <=( (not A170)  and  a66020a );
 a66024a <=( (not A200)  and  A166 );
 a66027a <=( (not A203)  and  (not A202) );
 a66028a <=( a66027a  and  a66024a );
 a66029a <=( a66028a  and  a66021a );
 a66032a <=( (not A233)  and  (not A232) );
 a66035a <=( (not A267)  and  (not A266) );
 a66036a <=( a66035a  and  a66032a );
 a66039a <=( (not A299)  and  A298 );
 a66042a <=( A301  and  A300 );
 a66043a <=( a66042a  and  a66039a );
 a66044a <=( a66043a  and  a66036a );
 a66048a <=( A167  and  A169 );
 a66049a <=( (not A170)  and  a66048a );
 a66052a <=( (not A200)  and  A166 );
 a66055a <=( (not A203)  and  (not A202) );
 a66056a <=( a66055a  and  a66052a );
 a66057a <=( a66056a  and  a66049a );
 a66060a <=( (not A233)  and  (not A232) );
 a66063a <=( (not A267)  and  (not A266) );
 a66064a <=( a66063a  and  a66060a );
 a66067a <=( (not A299)  and  A298 );
 a66070a <=( A302  and  A300 );
 a66071a <=( a66070a  and  a66067a );
 a66072a <=( a66071a  and  a66064a );
 a66076a <=( A167  and  A169 );
 a66077a <=( (not A170)  and  a66076a );
 a66080a <=( (not A200)  and  A166 );
 a66083a <=( (not A203)  and  (not A202) );
 a66084a <=( a66083a  and  a66080a );
 a66085a <=( a66084a  and  a66077a );
 a66088a <=( (not A233)  and  (not A232) );
 a66091a <=( (not A266)  and  (not A265) );
 a66092a <=( a66091a  and  a66088a );
 a66095a <=( (not A299)  and  A298 );
 a66098a <=( A301  and  A300 );
 a66099a <=( a66098a  and  a66095a );
 a66100a <=( a66099a  and  a66092a );
 a66104a <=( A167  and  A169 );
 a66105a <=( (not A170)  and  a66104a );
 a66108a <=( (not A200)  and  A166 );
 a66111a <=( (not A203)  and  (not A202) );
 a66112a <=( a66111a  and  a66108a );
 a66113a <=( a66112a  and  a66105a );
 a66116a <=( (not A233)  and  (not A232) );
 a66119a <=( (not A266)  and  (not A265) );
 a66120a <=( a66119a  and  a66116a );
 a66123a <=( (not A299)  and  A298 );
 a66126a <=( A302  and  A300 );
 a66127a <=( a66126a  and  a66123a );
 a66128a <=( a66127a  and  a66120a );
 a66132a <=( A167  and  A169 );
 a66133a <=( (not A170)  and  a66132a );
 a66136a <=( (not A200)  and  A166 );
 a66139a <=( A232  and  (not A201) );
 a66140a <=( a66139a  and  a66136a );
 a66141a <=( a66140a  and  a66133a );
 a66144a <=( A265  and  A233 );
 a66147a <=( (not A269)  and  (not A268) );
 a66148a <=( a66147a  and  a66144a );
 a66151a <=( (not A299)  and  A298 );
 a66154a <=( A301  and  A300 );
 a66155a <=( a66154a  and  a66151a );
 a66156a <=( a66155a  and  a66148a );
 a66160a <=( A167  and  A169 );
 a66161a <=( (not A170)  and  a66160a );
 a66164a <=( (not A200)  and  A166 );
 a66167a <=( A232  and  (not A201) );
 a66168a <=( a66167a  and  a66164a );
 a66169a <=( a66168a  and  a66161a );
 a66172a <=( A265  and  A233 );
 a66175a <=( (not A269)  and  (not A268) );
 a66176a <=( a66175a  and  a66172a );
 a66179a <=( (not A299)  and  A298 );
 a66182a <=( A302  and  A300 );
 a66183a <=( a66182a  and  a66179a );
 a66184a <=( a66183a  and  a66176a );
 a66188a <=( A167  and  A169 );
 a66189a <=( (not A170)  and  a66188a );
 a66192a <=( (not A200)  and  A166 );
 a66195a <=( (not A233)  and  (not A201) );
 a66196a <=( a66195a  and  a66192a );
 a66197a <=( a66196a  and  a66189a );
 a66200a <=( (not A236)  and  (not A235) );
 a66203a <=( A266  and  A265 );
 a66204a <=( a66203a  and  a66200a );
 a66207a <=( (not A299)  and  A298 );
 a66210a <=( A301  and  A300 );
 a66211a <=( a66210a  and  a66207a );
 a66212a <=( a66211a  and  a66204a );
 a66216a <=( A167  and  A169 );
 a66217a <=( (not A170)  and  a66216a );
 a66220a <=( (not A200)  and  A166 );
 a66223a <=( (not A233)  and  (not A201) );
 a66224a <=( a66223a  and  a66220a );
 a66225a <=( a66224a  and  a66217a );
 a66228a <=( (not A236)  and  (not A235) );
 a66231a <=( A266  and  A265 );
 a66232a <=( a66231a  and  a66228a );
 a66235a <=( (not A299)  and  A298 );
 a66238a <=( A302  and  A300 );
 a66239a <=( a66238a  and  a66235a );
 a66240a <=( a66239a  and  a66232a );
 a66244a <=( A167  and  A169 );
 a66245a <=( (not A170)  and  a66244a );
 a66248a <=( (not A200)  and  A166 );
 a66251a <=( (not A233)  and  (not A201) );
 a66252a <=( a66251a  and  a66248a );
 a66253a <=( a66252a  and  a66245a );
 a66256a <=( (not A236)  and  (not A235) );
 a66259a <=( (not A267)  and  (not A266) );
 a66260a <=( a66259a  and  a66256a );
 a66263a <=( (not A299)  and  A298 );
 a66266a <=( A301  and  A300 );
 a66267a <=( a66266a  and  a66263a );
 a66268a <=( a66267a  and  a66260a );
 a66272a <=( A167  and  A169 );
 a66273a <=( (not A170)  and  a66272a );
 a66276a <=( (not A200)  and  A166 );
 a66279a <=( (not A233)  and  (not A201) );
 a66280a <=( a66279a  and  a66276a );
 a66281a <=( a66280a  and  a66273a );
 a66284a <=( (not A236)  and  (not A235) );
 a66287a <=( (not A267)  and  (not A266) );
 a66288a <=( a66287a  and  a66284a );
 a66291a <=( (not A299)  and  A298 );
 a66294a <=( A302  and  A300 );
 a66295a <=( a66294a  and  a66291a );
 a66296a <=( a66295a  and  a66288a );
 a66300a <=( A167  and  A169 );
 a66301a <=( (not A170)  and  a66300a );
 a66304a <=( (not A200)  and  A166 );
 a66307a <=( (not A233)  and  (not A201) );
 a66308a <=( a66307a  and  a66304a );
 a66309a <=( a66308a  and  a66301a );
 a66312a <=( (not A236)  and  (not A235) );
 a66315a <=( (not A266)  and  (not A265) );
 a66316a <=( a66315a  and  a66312a );
 a66319a <=( (not A299)  and  A298 );
 a66322a <=( A301  and  A300 );
 a66323a <=( a66322a  and  a66319a );
 a66324a <=( a66323a  and  a66316a );
 a66328a <=( A167  and  A169 );
 a66329a <=( (not A170)  and  a66328a );
 a66332a <=( (not A200)  and  A166 );
 a66335a <=( (not A233)  and  (not A201) );
 a66336a <=( a66335a  and  a66332a );
 a66337a <=( a66336a  and  a66329a );
 a66340a <=( (not A236)  and  (not A235) );
 a66343a <=( (not A266)  and  (not A265) );
 a66344a <=( a66343a  and  a66340a );
 a66347a <=( (not A299)  and  A298 );
 a66350a <=( A302  and  A300 );
 a66351a <=( a66350a  and  a66347a );
 a66352a <=( a66351a  and  a66344a );
 a66356a <=( A167  and  A169 );
 a66357a <=( (not A170)  and  a66356a );
 a66360a <=( (not A200)  and  A166 );
 a66363a <=( (not A233)  and  (not A201) );
 a66364a <=( a66363a  and  a66360a );
 a66365a <=( a66364a  and  a66357a );
 a66368a <=( (not A266)  and  (not A234) );
 a66371a <=( (not A269)  and  (not A268) );
 a66372a <=( a66371a  and  a66368a );
 a66375a <=( (not A299)  and  A298 );
 a66378a <=( A301  and  A300 );
 a66379a <=( a66378a  and  a66375a );
 a66380a <=( a66379a  and  a66372a );
 a66384a <=( A167  and  A169 );
 a66385a <=( (not A170)  and  a66384a );
 a66388a <=( (not A200)  and  A166 );
 a66391a <=( (not A233)  and  (not A201) );
 a66392a <=( a66391a  and  a66388a );
 a66393a <=( a66392a  and  a66385a );
 a66396a <=( (not A266)  and  (not A234) );
 a66399a <=( (not A269)  and  (not A268) );
 a66400a <=( a66399a  and  a66396a );
 a66403a <=( (not A299)  and  A298 );
 a66406a <=( A302  and  A300 );
 a66407a <=( a66406a  and  a66403a );
 a66408a <=( a66407a  and  a66400a );
 a66412a <=( A167  and  A169 );
 a66413a <=( (not A170)  and  a66412a );
 a66416a <=( (not A200)  and  A166 );
 a66419a <=( (not A232)  and  (not A201) );
 a66420a <=( a66419a  and  a66416a );
 a66421a <=( a66420a  and  a66413a );
 a66424a <=( (not A266)  and  (not A233) );
 a66427a <=( (not A269)  and  (not A268) );
 a66428a <=( a66427a  and  a66424a );
 a66431a <=( (not A299)  and  A298 );
 a66434a <=( A301  and  A300 );
 a66435a <=( a66434a  and  a66431a );
 a66436a <=( a66435a  and  a66428a );
 a66440a <=( A167  and  A169 );
 a66441a <=( (not A170)  and  a66440a );
 a66444a <=( (not A200)  and  A166 );
 a66447a <=( (not A232)  and  (not A201) );
 a66448a <=( a66447a  and  a66444a );
 a66449a <=( a66448a  and  a66441a );
 a66452a <=( (not A266)  and  (not A233) );
 a66455a <=( (not A269)  and  (not A268) );
 a66456a <=( a66455a  and  a66452a );
 a66459a <=( (not A299)  and  A298 );
 a66462a <=( A302  and  A300 );
 a66463a <=( a66462a  and  a66459a );
 a66464a <=( a66463a  and  a66456a );
 a66468a <=( A167  and  A169 );
 a66469a <=( (not A170)  and  a66468a );
 a66472a <=( (not A199)  and  A166 );
 a66475a <=( A232  and  (not A200) );
 a66476a <=( a66475a  and  a66472a );
 a66477a <=( a66476a  and  a66469a );
 a66480a <=( A265  and  A233 );
 a66483a <=( (not A269)  and  (not A268) );
 a66484a <=( a66483a  and  a66480a );
 a66487a <=( (not A299)  and  A298 );
 a66490a <=( A301  and  A300 );
 a66491a <=( a66490a  and  a66487a );
 a66492a <=( a66491a  and  a66484a );
 a66496a <=( A167  and  A169 );
 a66497a <=( (not A170)  and  a66496a );
 a66500a <=( (not A199)  and  A166 );
 a66503a <=( A232  and  (not A200) );
 a66504a <=( a66503a  and  a66500a );
 a66505a <=( a66504a  and  a66497a );
 a66508a <=( A265  and  A233 );
 a66511a <=( (not A269)  and  (not A268) );
 a66512a <=( a66511a  and  a66508a );
 a66515a <=( (not A299)  and  A298 );
 a66518a <=( A302  and  A300 );
 a66519a <=( a66518a  and  a66515a );
 a66520a <=( a66519a  and  a66512a );
 a66524a <=( A167  and  A169 );
 a66525a <=( (not A170)  and  a66524a );
 a66528a <=( (not A199)  and  A166 );
 a66531a <=( (not A233)  and  (not A200) );
 a66532a <=( a66531a  and  a66528a );
 a66533a <=( a66532a  and  a66525a );
 a66536a <=( (not A236)  and  (not A235) );
 a66539a <=( A266  and  A265 );
 a66540a <=( a66539a  and  a66536a );
 a66543a <=( (not A299)  and  A298 );
 a66546a <=( A301  and  A300 );
 a66547a <=( a66546a  and  a66543a );
 a66548a <=( a66547a  and  a66540a );
 a66552a <=( A167  and  A169 );
 a66553a <=( (not A170)  and  a66552a );
 a66556a <=( (not A199)  and  A166 );
 a66559a <=( (not A233)  and  (not A200) );
 a66560a <=( a66559a  and  a66556a );
 a66561a <=( a66560a  and  a66553a );
 a66564a <=( (not A236)  and  (not A235) );
 a66567a <=( A266  and  A265 );
 a66568a <=( a66567a  and  a66564a );
 a66571a <=( (not A299)  and  A298 );
 a66574a <=( A302  and  A300 );
 a66575a <=( a66574a  and  a66571a );
 a66576a <=( a66575a  and  a66568a );
 a66580a <=( A167  and  A169 );
 a66581a <=( (not A170)  and  a66580a );
 a66584a <=( (not A199)  and  A166 );
 a66587a <=( (not A233)  and  (not A200) );
 a66588a <=( a66587a  and  a66584a );
 a66589a <=( a66588a  and  a66581a );
 a66592a <=( (not A236)  and  (not A235) );
 a66595a <=( (not A267)  and  (not A266) );
 a66596a <=( a66595a  and  a66592a );
 a66599a <=( (not A299)  and  A298 );
 a66602a <=( A301  and  A300 );
 a66603a <=( a66602a  and  a66599a );
 a66604a <=( a66603a  and  a66596a );
 a66608a <=( A167  and  A169 );
 a66609a <=( (not A170)  and  a66608a );
 a66612a <=( (not A199)  and  A166 );
 a66615a <=( (not A233)  and  (not A200) );
 a66616a <=( a66615a  and  a66612a );
 a66617a <=( a66616a  and  a66609a );
 a66620a <=( (not A236)  and  (not A235) );
 a66623a <=( (not A267)  and  (not A266) );
 a66624a <=( a66623a  and  a66620a );
 a66627a <=( (not A299)  and  A298 );
 a66630a <=( A302  and  A300 );
 a66631a <=( a66630a  and  a66627a );
 a66632a <=( a66631a  and  a66624a );
 a66636a <=( A167  and  A169 );
 a66637a <=( (not A170)  and  a66636a );
 a66640a <=( (not A199)  and  A166 );
 a66643a <=( (not A233)  and  (not A200) );
 a66644a <=( a66643a  and  a66640a );
 a66645a <=( a66644a  and  a66637a );
 a66648a <=( (not A236)  and  (not A235) );
 a66651a <=( (not A266)  and  (not A265) );
 a66652a <=( a66651a  and  a66648a );
 a66655a <=( (not A299)  and  A298 );
 a66658a <=( A301  and  A300 );
 a66659a <=( a66658a  and  a66655a );
 a66660a <=( a66659a  and  a66652a );
 a66664a <=( A167  and  A169 );
 a66665a <=( (not A170)  and  a66664a );
 a66668a <=( (not A199)  and  A166 );
 a66671a <=( (not A233)  and  (not A200) );
 a66672a <=( a66671a  and  a66668a );
 a66673a <=( a66672a  and  a66665a );
 a66676a <=( (not A236)  and  (not A235) );
 a66679a <=( (not A266)  and  (not A265) );
 a66680a <=( a66679a  and  a66676a );
 a66683a <=( (not A299)  and  A298 );
 a66686a <=( A302  and  A300 );
 a66687a <=( a66686a  and  a66683a );
 a66688a <=( a66687a  and  a66680a );
 a66692a <=( A167  and  A169 );
 a66693a <=( (not A170)  and  a66692a );
 a66696a <=( (not A199)  and  A166 );
 a66699a <=( (not A233)  and  (not A200) );
 a66700a <=( a66699a  and  a66696a );
 a66701a <=( a66700a  and  a66693a );
 a66704a <=( (not A266)  and  (not A234) );
 a66707a <=( (not A269)  and  (not A268) );
 a66708a <=( a66707a  and  a66704a );
 a66711a <=( (not A299)  and  A298 );
 a66714a <=( A301  and  A300 );
 a66715a <=( a66714a  and  a66711a );
 a66716a <=( a66715a  and  a66708a );
 a66720a <=( A167  and  A169 );
 a66721a <=( (not A170)  and  a66720a );
 a66724a <=( (not A199)  and  A166 );
 a66727a <=( (not A233)  and  (not A200) );
 a66728a <=( a66727a  and  a66724a );
 a66729a <=( a66728a  and  a66721a );
 a66732a <=( (not A266)  and  (not A234) );
 a66735a <=( (not A269)  and  (not A268) );
 a66736a <=( a66735a  and  a66732a );
 a66739a <=( (not A299)  and  A298 );
 a66742a <=( A302  and  A300 );
 a66743a <=( a66742a  and  a66739a );
 a66744a <=( a66743a  and  a66736a );
 a66748a <=( A167  and  A169 );
 a66749a <=( (not A170)  and  a66748a );
 a66752a <=( (not A199)  and  A166 );
 a66755a <=( (not A232)  and  (not A200) );
 a66756a <=( a66755a  and  a66752a );
 a66757a <=( a66756a  and  a66749a );
 a66760a <=( (not A266)  and  (not A233) );
 a66763a <=( (not A269)  and  (not A268) );
 a66764a <=( a66763a  and  a66760a );
 a66767a <=( (not A299)  and  A298 );
 a66770a <=( A301  and  A300 );
 a66771a <=( a66770a  and  a66767a );
 a66772a <=( a66771a  and  a66764a );
 a66776a <=( A167  and  A169 );
 a66777a <=( (not A170)  and  a66776a );
 a66780a <=( (not A199)  and  A166 );
 a66783a <=( (not A232)  and  (not A200) );
 a66784a <=( a66783a  and  a66780a );
 a66785a <=( a66784a  and  a66777a );
 a66788a <=( (not A266)  and  (not A233) );
 a66791a <=( (not A269)  and  (not A268) );
 a66792a <=( a66791a  and  a66788a );
 a66795a <=( (not A299)  and  A298 );
 a66798a <=( A302  and  A300 );
 a66799a <=( a66798a  and  a66795a );
 a66800a <=( a66799a  and  a66792a );
 a66804a <=( (not A167)  and  A169 );
 a66805a <=( (not A170)  and  a66804a );
 a66808a <=( A199  and  (not A166) );
 a66811a <=( A232  and  A200 );
 a66812a <=( a66811a  and  a66808a );
 a66813a <=( a66812a  and  a66805a );
 a66816a <=( A265  and  A233 );
 a66819a <=( (not A269)  and  (not A268) );
 a66820a <=( a66819a  and  a66816a );
 a66823a <=( (not A299)  and  A298 );
 a66826a <=( A301  and  A300 );
 a66827a <=( a66826a  and  a66823a );
 a66828a <=( a66827a  and  a66820a );
 a66832a <=( (not A167)  and  A169 );
 a66833a <=( (not A170)  and  a66832a );
 a66836a <=( A199  and  (not A166) );
 a66839a <=( A232  and  A200 );
 a66840a <=( a66839a  and  a66836a );
 a66841a <=( a66840a  and  a66833a );
 a66844a <=( A265  and  A233 );
 a66847a <=( (not A269)  and  (not A268) );
 a66848a <=( a66847a  and  a66844a );
 a66851a <=( (not A299)  and  A298 );
 a66854a <=( A302  and  A300 );
 a66855a <=( a66854a  and  a66851a );
 a66856a <=( a66855a  and  a66848a );
 a66860a <=( (not A167)  and  A169 );
 a66861a <=( (not A170)  and  a66860a );
 a66864a <=( A199  and  (not A166) );
 a66867a <=( (not A233)  and  A200 );
 a66868a <=( a66867a  and  a66864a );
 a66869a <=( a66868a  and  a66861a );
 a66872a <=( (not A236)  and  (not A235) );
 a66875a <=( A266  and  A265 );
 a66876a <=( a66875a  and  a66872a );
 a66879a <=( (not A299)  and  A298 );
 a66882a <=( A301  and  A300 );
 a66883a <=( a66882a  and  a66879a );
 a66884a <=( a66883a  and  a66876a );
 a66888a <=( (not A167)  and  A169 );
 a66889a <=( (not A170)  and  a66888a );
 a66892a <=( A199  and  (not A166) );
 a66895a <=( (not A233)  and  A200 );
 a66896a <=( a66895a  and  a66892a );
 a66897a <=( a66896a  and  a66889a );
 a66900a <=( (not A236)  and  (not A235) );
 a66903a <=( A266  and  A265 );
 a66904a <=( a66903a  and  a66900a );
 a66907a <=( (not A299)  and  A298 );
 a66910a <=( A302  and  A300 );
 a66911a <=( a66910a  and  a66907a );
 a66912a <=( a66911a  and  a66904a );
 a66916a <=( (not A167)  and  A169 );
 a66917a <=( (not A170)  and  a66916a );
 a66920a <=( A199  and  (not A166) );
 a66923a <=( (not A233)  and  A200 );
 a66924a <=( a66923a  and  a66920a );
 a66925a <=( a66924a  and  a66917a );
 a66928a <=( (not A236)  and  (not A235) );
 a66931a <=( (not A267)  and  (not A266) );
 a66932a <=( a66931a  and  a66928a );
 a66935a <=( (not A299)  and  A298 );
 a66938a <=( A301  and  A300 );
 a66939a <=( a66938a  and  a66935a );
 a66940a <=( a66939a  and  a66932a );
 a66944a <=( (not A167)  and  A169 );
 a66945a <=( (not A170)  and  a66944a );
 a66948a <=( A199  and  (not A166) );
 a66951a <=( (not A233)  and  A200 );
 a66952a <=( a66951a  and  a66948a );
 a66953a <=( a66952a  and  a66945a );
 a66956a <=( (not A236)  and  (not A235) );
 a66959a <=( (not A267)  and  (not A266) );
 a66960a <=( a66959a  and  a66956a );
 a66963a <=( (not A299)  and  A298 );
 a66966a <=( A302  and  A300 );
 a66967a <=( a66966a  and  a66963a );
 a66968a <=( a66967a  and  a66960a );
 a66972a <=( (not A167)  and  A169 );
 a66973a <=( (not A170)  and  a66972a );
 a66976a <=( A199  and  (not A166) );
 a66979a <=( (not A233)  and  A200 );
 a66980a <=( a66979a  and  a66976a );
 a66981a <=( a66980a  and  a66973a );
 a66984a <=( (not A236)  and  (not A235) );
 a66987a <=( (not A266)  and  (not A265) );
 a66988a <=( a66987a  and  a66984a );
 a66991a <=( (not A299)  and  A298 );
 a66994a <=( A301  and  A300 );
 a66995a <=( a66994a  and  a66991a );
 a66996a <=( a66995a  and  a66988a );
 a67000a <=( (not A167)  and  A169 );
 a67001a <=( (not A170)  and  a67000a );
 a67004a <=( A199  and  (not A166) );
 a67007a <=( (not A233)  and  A200 );
 a67008a <=( a67007a  and  a67004a );
 a67009a <=( a67008a  and  a67001a );
 a67012a <=( (not A236)  and  (not A235) );
 a67015a <=( (not A266)  and  (not A265) );
 a67016a <=( a67015a  and  a67012a );
 a67019a <=( (not A299)  and  A298 );
 a67022a <=( A302  and  A300 );
 a67023a <=( a67022a  and  a67019a );
 a67024a <=( a67023a  and  a67016a );
 a67028a <=( (not A167)  and  A169 );
 a67029a <=( (not A170)  and  a67028a );
 a67032a <=( A199  and  (not A166) );
 a67035a <=( (not A233)  and  A200 );
 a67036a <=( a67035a  and  a67032a );
 a67037a <=( a67036a  and  a67029a );
 a67040a <=( (not A266)  and  (not A234) );
 a67043a <=( (not A269)  and  (not A268) );
 a67044a <=( a67043a  and  a67040a );
 a67047a <=( (not A299)  and  A298 );
 a67050a <=( A301  and  A300 );
 a67051a <=( a67050a  and  a67047a );
 a67052a <=( a67051a  and  a67044a );
 a67056a <=( (not A167)  and  A169 );
 a67057a <=( (not A170)  and  a67056a );
 a67060a <=( A199  and  (not A166) );
 a67063a <=( (not A233)  and  A200 );
 a67064a <=( a67063a  and  a67060a );
 a67065a <=( a67064a  and  a67057a );
 a67068a <=( (not A266)  and  (not A234) );
 a67071a <=( (not A269)  and  (not A268) );
 a67072a <=( a67071a  and  a67068a );
 a67075a <=( (not A299)  and  A298 );
 a67078a <=( A302  and  A300 );
 a67079a <=( a67078a  and  a67075a );
 a67080a <=( a67079a  and  a67072a );
 a67084a <=( (not A167)  and  A169 );
 a67085a <=( (not A170)  and  a67084a );
 a67088a <=( A199  and  (not A166) );
 a67091a <=( (not A232)  and  A200 );
 a67092a <=( a67091a  and  a67088a );
 a67093a <=( a67092a  and  a67085a );
 a67096a <=( (not A266)  and  (not A233) );
 a67099a <=( (not A269)  and  (not A268) );
 a67100a <=( a67099a  and  a67096a );
 a67103a <=( (not A299)  and  A298 );
 a67106a <=( A301  and  A300 );
 a67107a <=( a67106a  and  a67103a );
 a67108a <=( a67107a  and  a67100a );
 a67112a <=( (not A167)  and  A169 );
 a67113a <=( (not A170)  and  a67112a );
 a67116a <=( A199  and  (not A166) );
 a67119a <=( (not A232)  and  A200 );
 a67120a <=( a67119a  and  a67116a );
 a67121a <=( a67120a  and  a67113a );
 a67124a <=( (not A266)  and  (not A233) );
 a67127a <=( (not A269)  and  (not A268) );
 a67128a <=( a67127a  and  a67124a );
 a67131a <=( (not A299)  and  A298 );
 a67134a <=( A302  and  A300 );
 a67135a <=( a67134a  and  a67131a );
 a67136a <=( a67135a  and  a67128a );
 a67140a <=( (not A167)  and  A169 );
 a67141a <=( (not A170)  and  a67140a );
 a67144a <=( (not A200)  and  (not A166) );
 a67147a <=( (not A203)  and  (not A202) );
 a67148a <=( a67147a  and  a67144a );
 a67149a <=( a67148a  and  a67141a );
 a67152a <=( A233  and  A232 );
 a67155a <=( (not A267)  and  A265 );
 a67156a <=( a67155a  and  a67152a );
 a67159a <=( (not A299)  and  A298 );
 a67162a <=( A301  and  A300 );
 a67163a <=( a67162a  and  a67159a );
 a67164a <=( a67163a  and  a67156a );
 a67168a <=( (not A167)  and  A169 );
 a67169a <=( (not A170)  and  a67168a );
 a67172a <=( (not A200)  and  (not A166) );
 a67175a <=( (not A203)  and  (not A202) );
 a67176a <=( a67175a  and  a67172a );
 a67177a <=( a67176a  and  a67169a );
 a67180a <=( A233  and  A232 );
 a67183a <=( (not A267)  and  A265 );
 a67184a <=( a67183a  and  a67180a );
 a67187a <=( (not A299)  and  A298 );
 a67190a <=( A302  and  A300 );
 a67191a <=( a67190a  and  a67187a );
 a67192a <=( a67191a  and  a67184a );
 a67196a <=( (not A167)  and  A169 );
 a67197a <=( (not A170)  and  a67196a );
 a67200a <=( (not A200)  and  (not A166) );
 a67203a <=( (not A203)  and  (not A202) );
 a67204a <=( a67203a  and  a67200a );
 a67205a <=( a67204a  and  a67197a );
 a67208a <=( A233  and  A232 );
 a67211a <=( A266  and  A265 );
 a67212a <=( a67211a  and  a67208a );
 a67215a <=( (not A299)  and  A298 );
 a67218a <=( A301  and  A300 );
 a67219a <=( a67218a  and  a67215a );
 a67220a <=( a67219a  and  a67212a );
 a67224a <=( (not A167)  and  A169 );
 a67225a <=( (not A170)  and  a67224a );
 a67228a <=( (not A200)  and  (not A166) );
 a67231a <=( (not A203)  and  (not A202) );
 a67232a <=( a67231a  and  a67228a );
 a67233a <=( a67232a  and  a67225a );
 a67236a <=( A233  and  A232 );
 a67239a <=( A266  and  A265 );
 a67240a <=( a67239a  and  a67236a );
 a67243a <=( (not A299)  and  A298 );
 a67246a <=( A302  and  A300 );
 a67247a <=( a67246a  and  a67243a );
 a67248a <=( a67247a  and  a67240a );
 a67252a <=( (not A167)  and  A169 );
 a67253a <=( (not A170)  and  a67252a );
 a67256a <=( (not A200)  and  (not A166) );
 a67259a <=( (not A203)  and  (not A202) );
 a67260a <=( a67259a  and  a67256a );
 a67261a <=( a67260a  and  a67253a );
 a67264a <=( A233  and  A232 );
 a67267a <=( (not A266)  and  (not A265) );
 a67268a <=( a67267a  and  a67264a );
 a67271a <=( (not A299)  and  A298 );
 a67274a <=( A301  and  A300 );
 a67275a <=( a67274a  and  a67271a );
 a67276a <=( a67275a  and  a67268a );
 a67280a <=( (not A167)  and  A169 );
 a67281a <=( (not A170)  and  a67280a );
 a67284a <=( (not A200)  and  (not A166) );
 a67287a <=( (not A203)  and  (not A202) );
 a67288a <=( a67287a  and  a67284a );
 a67289a <=( a67288a  and  a67281a );
 a67292a <=( A233  and  A232 );
 a67295a <=( (not A266)  and  (not A265) );
 a67296a <=( a67295a  and  a67292a );
 a67299a <=( (not A299)  and  A298 );
 a67302a <=( A302  and  A300 );
 a67303a <=( a67302a  and  a67299a );
 a67304a <=( a67303a  and  a67296a );
 a67308a <=( (not A167)  and  A169 );
 a67309a <=( (not A170)  and  a67308a );
 a67312a <=( (not A200)  and  (not A166) );
 a67315a <=( (not A203)  and  (not A202) );
 a67316a <=( a67315a  and  a67312a );
 a67317a <=( a67316a  and  a67309a );
 a67320a <=( (not A235)  and  (not A233) );
 a67323a <=( (not A266)  and  (not A236) );
 a67324a <=( a67323a  and  a67320a );
 a67327a <=( (not A269)  and  (not A268) );
 a67330a <=( A299  and  (not A298) );
 a67331a <=( a67330a  and  a67327a );
 a67332a <=( a67331a  and  a67324a );
 a67336a <=( (not A167)  and  A169 );
 a67337a <=( (not A170)  and  a67336a );
 a67340a <=( (not A200)  and  (not A166) );
 a67343a <=( (not A203)  and  (not A202) );
 a67344a <=( a67343a  and  a67340a );
 a67345a <=( a67344a  and  a67337a );
 a67348a <=( (not A234)  and  (not A233) );
 a67351a <=( A266  and  A265 );
 a67352a <=( a67351a  and  a67348a );
 a67355a <=( (not A299)  and  A298 );
 a67358a <=( A301  and  A300 );
 a67359a <=( a67358a  and  a67355a );
 a67360a <=( a67359a  and  a67352a );
 a67364a <=( (not A167)  and  A169 );
 a67365a <=( (not A170)  and  a67364a );
 a67368a <=( (not A200)  and  (not A166) );
 a67371a <=( (not A203)  and  (not A202) );
 a67372a <=( a67371a  and  a67368a );
 a67373a <=( a67372a  and  a67365a );
 a67376a <=( (not A234)  and  (not A233) );
 a67379a <=( A266  and  A265 );
 a67380a <=( a67379a  and  a67376a );
 a67383a <=( (not A299)  and  A298 );
 a67386a <=( A302  and  A300 );
 a67387a <=( a67386a  and  a67383a );
 a67388a <=( a67387a  and  a67380a );
 a67392a <=( (not A167)  and  A169 );
 a67393a <=( (not A170)  and  a67392a );
 a67396a <=( (not A200)  and  (not A166) );
 a67399a <=( (not A203)  and  (not A202) );
 a67400a <=( a67399a  and  a67396a );
 a67401a <=( a67400a  and  a67393a );
 a67404a <=( (not A234)  and  (not A233) );
 a67407a <=( (not A267)  and  (not A266) );
 a67408a <=( a67407a  and  a67404a );
 a67411a <=( (not A299)  and  A298 );
 a67414a <=( A301  and  A300 );
 a67415a <=( a67414a  and  a67411a );
 a67416a <=( a67415a  and  a67408a );
 a67420a <=( (not A167)  and  A169 );
 a67421a <=( (not A170)  and  a67420a );
 a67424a <=( (not A200)  and  (not A166) );
 a67427a <=( (not A203)  and  (not A202) );
 a67428a <=( a67427a  and  a67424a );
 a67429a <=( a67428a  and  a67421a );
 a67432a <=( (not A234)  and  (not A233) );
 a67435a <=( (not A267)  and  (not A266) );
 a67436a <=( a67435a  and  a67432a );
 a67439a <=( (not A299)  and  A298 );
 a67442a <=( A302  and  A300 );
 a67443a <=( a67442a  and  a67439a );
 a67444a <=( a67443a  and  a67436a );
 a67448a <=( (not A167)  and  A169 );
 a67449a <=( (not A170)  and  a67448a );
 a67452a <=( (not A200)  and  (not A166) );
 a67455a <=( (not A203)  and  (not A202) );
 a67456a <=( a67455a  and  a67452a );
 a67457a <=( a67456a  and  a67449a );
 a67460a <=( (not A234)  and  (not A233) );
 a67463a <=( (not A266)  and  (not A265) );
 a67464a <=( a67463a  and  a67460a );
 a67467a <=( (not A299)  and  A298 );
 a67470a <=( A301  and  A300 );
 a67471a <=( a67470a  and  a67467a );
 a67472a <=( a67471a  and  a67464a );
 a67476a <=( (not A167)  and  A169 );
 a67477a <=( (not A170)  and  a67476a );
 a67480a <=( (not A200)  and  (not A166) );
 a67483a <=( (not A203)  and  (not A202) );
 a67484a <=( a67483a  and  a67480a );
 a67485a <=( a67484a  and  a67477a );
 a67488a <=( (not A234)  and  (not A233) );
 a67491a <=( (not A266)  and  (not A265) );
 a67492a <=( a67491a  and  a67488a );
 a67495a <=( (not A299)  and  A298 );
 a67498a <=( A302  and  A300 );
 a67499a <=( a67498a  and  a67495a );
 a67500a <=( a67499a  and  a67492a );
 a67504a <=( (not A167)  and  A169 );
 a67505a <=( (not A170)  and  a67504a );
 a67508a <=( (not A200)  and  (not A166) );
 a67511a <=( (not A203)  and  (not A202) );
 a67512a <=( a67511a  and  a67508a );
 a67513a <=( a67512a  and  a67505a );
 a67516a <=( (not A233)  and  A232 );
 a67519a <=( A235  and  A234 );
 a67520a <=( a67519a  and  a67516a );
 a67523a <=( (not A266)  and  A265 );
 a67526a <=( A268  and  A267 );
 a67527a <=( a67526a  and  a67523a );
 a67528a <=( a67527a  and  a67520a );
 a67532a <=( (not A167)  and  A169 );
 a67533a <=( (not A170)  and  a67532a );
 a67536a <=( (not A200)  and  (not A166) );
 a67539a <=( (not A203)  and  (not A202) );
 a67540a <=( a67539a  and  a67536a );
 a67541a <=( a67540a  and  a67533a );
 a67544a <=( (not A233)  and  A232 );
 a67547a <=( A235  and  A234 );
 a67548a <=( a67547a  and  a67544a );
 a67551a <=( (not A266)  and  A265 );
 a67554a <=( A269  and  A267 );
 a67555a <=( a67554a  and  a67551a );
 a67556a <=( a67555a  and  a67548a );
 a67560a <=( (not A167)  and  A169 );
 a67561a <=( (not A170)  and  a67560a );
 a67564a <=( (not A200)  and  (not A166) );
 a67567a <=( (not A203)  and  (not A202) );
 a67568a <=( a67567a  and  a67564a );
 a67569a <=( a67568a  and  a67561a );
 a67572a <=( (not A233)  and  A232 );
 a67575a <=( A236  and  A234 );
 a67576a <=( a67575a  and  a67572a );
 a67579a <=( (not A266)  and  A265 );
 a67582a <=( A268  and  A267 );
 a67583a <=( a67582a  and  a67579a );
 a67584a <=( a67583a  and  a67576a );
 a67588a <=( (not A167)  and  A169 );
 a67589a <=( (not A170)  and  a67588a );
 a67592a <=( (not A200)  and  (not A166) );
 a67595a <=( (not A203)  and  (not A202) );
 a67596a <=( a67595a  and  a67592a );
 a67597a <=( a67596a  and  a67589a );
 a67600a <=( (not A233)  and  A232 );
 a67603a <=( A236  and  A234 );
 a67604a <=( a67603a  and  a67600a );
 a67607a <=( (not A266)  and  A265 );
 a67610a <=( A269  and  A267 );
 a67611a <=( a67610a  and  a67607a );
 a67612a <=( a67611a  and  a67604a );
 a67616a <=( (not A167)  and  A169 );
 a67617a <=( (not A170)  and  a67616a );
 a67620a <=( (not A200)  and  (not A166) );
 a67623a <=( (not A203)  and  (not A202) );
 a67624a <=( a67623a  and  a67620a );
 a67625a <=( a67624a  and  a67617a );
 a67628a <=( (not A233)  and  (not A232) );
 a67631a <=( A266  and  A265 );
 a67632a <=( a67631a  and  a67628a );
 a67635a <=( (not A299)  and  A298 );
 a67638a <=( A301  and  A300 );
 a67639a <=( a67638a  and  a67635a );
 a67640a <=( a67639a  and  a67632a );
 a67644a <=( (not A167)  and  A169 );
 a67645a <=( (not A170)  and  a67644a );
 a67648a <=( (not A200)  and  (not A166) );
 a67651a <=( (not A203)  and  (not A202) );
 a67652a <=( a67651a  and  a67648a );
 a67653a <=( a67652a  and  a67645a );
 a67656a <=( (not A233)  and  (not A232) );
 a67659a <=( A266  and  A265 );
 a67660a <=( a67659a  and  a67656a );
 a67663a <=( (not A299)  and  A298 );
 a67666a <=( A302  and  A300 );
 a67667a <=( a67666a  and  a67663a );
 a67668a <=( a67667a  and  a67660a );
 a67672a <=( (not A167)  and  A169 );
 a67673a <=( (not A170)  and  a67672a );
 a67676a <=( (not A200)  and  (not A166) );
 a67679a <=( (not A203)  and  (not A202) );
 a67680a <=( a67679a  and  a67676a );
 a67681a <=( a67680a  and  a67673a );
 a67684a <=( (not A233)  and  (not A232) );
 a67687a <=( (not A267)  and  (not A266) );
 a67688a <=( a67687a  and  a67684a );
 a67691a <=( (not A299)  and  A298 );
 a67694a <=( A301  and  A300 );
 a67695a <=( a67694a  and  a67691a );
 a67696a <=( a67695a  and  a67688a );
 a67700a <=( (not A167)  and  A169 );
 a67701a <=( (not A170)  and  a67700a );
 a67704a <=( (not A200)  and  (not A166) );
 a67707a <=( (not A203)  and  (not A202) );
 a67708a <=( a67707a  and  a67704a );
 a67709a <=( a67708a  and  a67701a );
 a67712a <=( (not A233)  and  (not A232) );
 a67715a <=( (not A267)  and  (not A266) );
 a67716a <=( a67715a  and  a67712a );
 a67719a <=( (not A299)  and  A298 );
 a67722a <=( A302  and  A300 );
 a67723a <=( a67722a  and  a67719a );
 a67724a <=( a67723a  and  a67716a );
 a67728a <=( (not A167)  and  A169 );
 a67729a <=( (not A170)  and  a67728a );
 a67732a <=( (not A200)  and  (not A166) );
 a67735a <=( (not A203)  and  (not A202) );
 a67736a <=( a67735a  and  a67732a );
 a67737a <=( a67736a  and  a67729a );
 a67740a <=( (not A233)  and  (not A232) );
 a67743a <=( (not A266)  and  (not A265) );
 a67744a <=( a67743a  and  a67740a );
 a67747a <=( (not A299)  and  A298 );
 a67750a <=( A301  and  A300 );
 a67751a <=( a67750a  and  a67747a );
 a67752a <=( a67751a  and  a67744a );
 a67756a <=( (not A167)  and  A169 );
 a67757a <=( (not A170)  and  a67756a );
 a67760a <=( (not A200)  and  (not A166) );
 a67763a <=( (not A203)  and  (not A202) );
 a67764a <=( a67763a  and  a67760a );
 a67765a <=( a67764a  and  a67757a );
 a67768a <=( (not A233)  and  (not A232) );
 a67771a <=( (not A266)  and  (not A265) );
 a67772a <=( a67771a  and  a67768a );
 a67775a <=( (not A299)  and  A298 );
 a67778a <=( A302  and  A300 );
 a67779a <=( a67778a  and  a67775a );
 a67780a <=( a67779a  and  a67772a );
 a67784a <=( (not A167)  and  A169 );
 a67785a <=( (not A170)  and  a67784a );
 a67788a <=( (not A200)  and  (not A166) );
 a67791a <=( A232  and  (not A201) );
 a67792a <=( a67791a  and  a67788a );
 a67793a <=( a67792a  and  a67785a );
 a67796a <=( A265  and  A233 );
 a67799a <=( (not A269)  and  (not A268) );
 a67800a <=( a67799a  and  a67796a );
 a67803a <=( (not A299)  and  A298 );
 a67806a <=( A301  and  A300 );
 a67807a <=( a67806a  and  a67803a );
 a67808a <=( a67807a  and  a67800a );
 a67812a <=( (not A167)  and  A169 );
 a67813a <=( (not A170)  and  a67812a );
 a67816a <=( (not A200)  and  (not A166) );
 a67819a <=( A232  and  (not A201) );
 a67820a <=( a67819a  and  a67816a );
 a67821a <=( a67820a  and  a67813a );
 a67824a <=( A265  and  A233 );
 a67827a <=( (not A269)  and  (not A268) );
 a67828a <=( a67827a  and  a67824a );
 a67831a <=( (not A299)  and  A298 );
 a67834a <=( A302  and  A300 );
 a67835a <=( a67834a  and  a67831a );
 a67836a <=( a67835a  and  a67828a );
 a67840a <=( (not A167)  and  A169 );
 a67841a <=( (not A170)  and  a67840a );
 a67844a <=( (not A200)  and  (not A166) );
 a67847a <=( (not A233)  and  (not A201) );
 a67848a <=( a67847a  and  a67844a );
 a67849a <=( a67848a  and  a67841a );
 a67852a <=( (not A236)  and  (not A235) );
 a67855a <=( A266  and  A265 );
 a67856a <=( a67855a  and  a67852a );
 a67859a <=( (not A299)  and  A298 );
 a67862a <=( A301  and  A300 );
 a67863a <=( a67862a  and  a67859a );
 a67864a <=( a67863a  and  a67856a );
 a67868a <=( (not A167)  and  A169 );
 a67869a <=( (not A170)  and  a67868a );
 a67872a <=( (not A200)  and  (not A166) );
 a67875a <=( (not A233)  and  (not A201) );
 a67876a <=( a67875a  and  a67872a );
 a67877a <=( a67876a  and  a67869a );
 a67880a <=( (not A236)  and  (not A235) );
 a67883a <=( A266  and  A265 );
 a67884a <=( a67883a  and  a67880a );
 a67887a <=( (not A299)  and  A298 );
 a67890a <=( A302  and  A300 );
 a67891a <=( a67890a  and  a67887a );
 a67892a <=( a67891a  and  a67884a );
 a67896a <=( (not A167)  and  A169 );
 a67897a <=( (not A170)  and  a67896a );
 a67900a <=( (not A200)  and  (not A166) );
 a67903a <=( (not A233)  and  (not A201) );
 a67904a <=( a67903a  and  a67900a );
 a67905a <=( a67904a  and  a67897a );
 a67908a <=( (not A236)  and  (not A235) );
 a67911a <=( (not A267)  and  (not A266) );
 a67912a <=( a67911a  and  a67908a );
 a67915a <=( (not A299)  and  A298 );
 a67918a <=( A301  and  A300 );
 a67919a <=( a67918a  and  a67915a );
 a67920a <=( a67919a  and  a67912a );
 a67924a <=( (not A167)  and  A169 );
 a67925a <=( (not A170)  and  a67924a );
 a67928a <=( (not A200)  and  (not A166) );
 a67931a <=( (not A233)  and  (not A201) );
 a67932a <=( a67931a  and  a67928a );
 a67933a <=( a67932a  and  a67925a );
 a67936a <=( (not A236)  and  (not A235) );
 a67939a <=( (not A267)  and  (not A266) );
 a67940a <=( a67939a  and  a67936a );
 a67943a <=( (not A299)  and  A298 );
 a67946a <=( A302  and  A300 );
 a67947a <=( a67946a  and  a67943a );
 a67948a <=( a67947a  and  a67940a );
 a67952a <=( (not A167)  and  A169 );
 a67953a <=( (not A170)  and  a67952a );
 a67956a <=( (not A200)  and  (not A166) );
 a67959a <=( (not A233)  and  (not A201) );
 a67960a <=( a67959a  and  a67956a );
 a67961a <=( a67960a  and  a67953a );
 a67964a <=( (not A236)  and  (not A235) );
 a67967a <=( (not A266)  and  (not A265) );
 a67968a <=( a67967a  and  a67964a );
 a67971a <=( (not A299)  and  A298 );
 a67974a <=( A301  and  A300 );
 a67975a <=( a67974a  and  a67971a );
 a67976a <=( a67975a  and  a67968a );
 a67980a <=( (not A167)  and  A169 );
 a67981a <=( (not A170)  and  a67980a );
 a67984a <=( (not A200)  and  (not A166) );
 a67987a <=( (not A233)  and  (not A201) );
 a67988a <=( a67987a  and  a67984a );
 a67989a <=( a67988a  and  a67981a );
 a67992a <=( (not A236)  and  (not A235) );
 a67995a <=( (not A266)  and  (not A265) );
 a67996a <=( a67995a  and  a67992a );
 a67999a <=( (not A299)  and  A298 );
 a68002a <=( A302  and  A300 );
 a68003a <=( a68002a  and  a67999a );
 a68004a <=( a68003a  and  a67996a );
 a68008a <=( (not A167)  and  A169 );
 a68009a <=( (not A170)  and  a68008a );
 a68012a <=( (not A200)  and  (not A166) );
 a68015a <=( (not A233)  and  (not A201) );
 a68016a <=( a68015a  and  a68012a );
 a68017a <=( a68016a  and  a68009a );
 a68020a <=( (not A266)  and  (not A234) );
 a68023a <=( (not A269)  and  (not A268) );
 a68024a <=( a68023a  and  a68020a );
 a68027a <=( (not A299)  and  A298 );
 a68030a <=( A301  and  A300 );
 a68031a <=( a68030a  and  a68027a );
 a68032a <=( a68031a  and  a68024a );
 a68036a <=( (not A167)  and  A169 );
 a68037a <=( (not A170)  and  a68036a );
 a68040a <=( (not A200)  and  (not A166) );
 a68043a <=( (not A233)  and  (not A201) );
 a68044a <=( a68043a  and  a68040a );
 a68045a <=( a68044a  and  a68037a );
 a68048a <=( (not A266)  and  (not A234) );
 a68051a <=( (not A269)  and  (not A268) );
 a68052a <=( a68051a  and  a68048a );
 a68055a <=( (not A299)  and  A298 );
 a68058a <=( A302  and  A300 );
 a68059a <=( a68058a  and  a68055a );
 a68060a <=( a68059a  and  a68052a );
 a68064a <=( (not A167)  and  A169 );
 a68065a <=( (not A170)  and  a68064a );
 a68068a <=( (not A200)  and  (not A166) );
 a68071a <=( (not A232)  and  (not A201) );
 a68072a <=( a68071a  and  a68068a );
 a68073a <=( a68072a  and  a68065a );
 a68076a <=( (not A266)  and  (not A233) );
 a68079a <=( (not A269)  and  (not A268) );
 a68080a <=( a68079a  and  a68076a );
 a68083a <=( (not A299)  and  A298 );
 a68086a <=( A301  and  A300 );
 a68087a <=( a68086a  and  a68083a );
 a68088a <=( a68087a  and  a68080a );
 a68092a <=( (not A167)  and  A169 );
 a68093a <=( (not A170)  and  a68092a );
 a68096a <=( (not A200)  and  (not A166) );
 a68099a <=( (not A232)  and  (not A201) );
 a68100a <=( a68099a  and  a68096a );
 a68101a <=( a68100a  and  a68093a );
 a68104a <=( (not A266)  and  (not A233) );
 a68107a <=( (not A269)  and  (not A268) );
 a68108a <=( a68107a  and  a68104a );
 a68111a <=( (not A299)  and  A298 );
 a68114a <=( A302  and  A300 );
 a68115a <=( a68114a  and  a68111a );
 a68116a <=( a68115a  and  a68108a );
 a68120a <=( (not A167)  and  A169 );
 a68121a <=( (not A170)  and  a68120a );
 a68124a <=( (not A199)  and  (not A166) );
 a68127a <=( A232  and  (not A200) );
 a68128a <=( a68127a  and  a68124a );
 a68129a <=( a68128a  and  a68121a );
 a68132a <=( A265  and  A233 );
 a68135a <=( (not A269)  and  (not A268) );
 a68136a <=( a68135a  and  a68132a );
 a68139a <=( (not A299)  and  A298 );
 a68142a <=( A301  and  A300 );
 a68143a <=( a68142a  and  a68139a );
 a68144a <=( a68143a  and  a68136a );
 a68148a <=( (not A167)  and  A169 );
 a68149a <=( (not A170)  and  a68148a );
 a68152a <=( (not A199)  and  (not A166) );
 a68155a <=( A232  and  (not A200) );
 a68156a <=( a68155a  and  a68152a );
 a68157a <=( a68156a  and  a68149a );
 a68160a <=( A265  and  A233 );
 a68163a <=( (not A269)  and  (not A268) );
 a68164a <=( a68163a  and  a68160a );
 a68167a <=( (not A299)  and  A298 );
 a68170a <=( A302  and  A300 );
 a68171a <=( a68170a  and  a68167a );
 a68172a <=( a68171a  and  a68164a );
 a68176a <=( (not A167)  and  A169 );
 a68177a <=( (not A170)  and  a68176a );
 a68180a <=( (not A199)  and  (not A166) );
 a68183a <=( (not A233)  and  (not A200) );
 a68184a <=( a68183a  and  a68180a );
 a68185a <=( a68184a  and  a68177a );
 a68188a <=( (not A236)  and  (not A235) );
 a68191a <=( A266  and  A265 );
 a68192a <=( a68191a  and  a68188a );
 a68195a <=( (not A299)  and  A298 );
 a68198a <=( A301  and  A300 );
 a68199a <=( a68198a  and  a68195a );
 a68200a <=( a68199a  and  a68192a );
 a68204a <=( (not A167)  and  A169 );
 a68205a <=( (not A170)  and  a68204a );
 a68208a <=( (not A199)  and  (not A166) );
 a68211a <=( (not A233)  and  (not A200) );
 a68212a <=( a68211a  and  a68208a );
 a68213a <=( a68212a  and  a68205a );
 a68216a <=( (not A236)  and  (not A235) );
 a68219a <=( A266  and  A265 );
 a68220a <=( a68219a  and  a68216a );
 a68223a <=( (not A299)  and  A298 );
 a68226a <=( A302  and  A300 );
 a68227a <=( a68226a  and  a68223a );
 a68228a <=( a68227a  and  a68220a );
 a68232a <=( (not A167)  and  A169 );
 a68233a <=( (not A170)  and  a68232a );
 a68236a <=( (not A199)  and  (not A166) );
 a68239a <=( (not A233)  and  (not A200) );
 a68240a <=( a68239a  and  a68236a );
 a68241a <=( a68240a  and  a68233a );
 a68244a <=( (not A236)  and  (not A235) );
 a68247a <=( (not A267)  and  (not A266) );
 a68248a <=( a68247a  and  a68244a );
 a68251a <=( (not A299)  and  A298 );
 a68254a <=( A301  and  A300 );
 a68255a <=( a68254a  and  a68251a );
 a68256a <=( a68255a  and  a68248a );
 a68260a <=( (not A167)  and  A169 );
 a68261a <=( (not A170)  and  a68260a );
 a68264a <=( (not A199)  and  (not A166) );
 a68267a <=( (not A233)  and  (not A200) );
 a68268a <=( a68267a  and  a68264a );
 a68269a <=( a68268a  and  a68261a );
 a68272a <=( (not A236)  and  (not A235) );
 a68275a <=( (not A267)  and  (not A266) );
 a68276a <=( a68275a  and  a68272a );
 a68279a <=( (not A299)  and  A298 );
 a68282a <=( A302  and  A300 );
 a68283a <=( a68282a  and  a68279a );
 a68284a <=( a68283a  and  a68276a );
 a68288a <=( (not A167)  and  A169 );
 a68289a <=( (not A170)  and  a68288a );
 a68292a <=( (not A199)  and  (not A166) );
 a68295a <=( (not A233)  and  (not A200) );
 a68296a <=( a68295a  and  a68292a );
 a68297a <=( a68296a  and  a68289a );
 a68300a <=( (not A236)  and  (not A235) );
 a68303a <=( (not A266)  and  (not A265) );
 a68304a <=( a68303a  and  a68300a );
 a68307a <=( (not A299)  and  A298 );
 a68310a <=( A301  and  A300 );
 a68311a <=( a68310a  and  a68307a );
 a68312a <=( a68311a  and  a68304a );
 a68316a <=( (not A167)  and  A169 );
 a68317a <=( (not A170)  and  a68316a );
 a68320a <=( (not A199)  and  (not A166) );
 a68323a <=( (not A233)  and  (not A200) );
 a68324a <=( a68323a  and  a68320a );
 a68325a <=( a68324a  and  a68317a );
 a68328a <=( (not A236)  and  (not A235) );
 a68331a <=( (not A266)  and  (not A265) );
 a68332a <=( a68331a  and  a68328a );
 a68335a <=( (not A299)  and  A298 );
 a68338a <=( A302  and  A300 );
 a68339a <=( a68338a  and  a68335a );
 a68340a <=( a68339a  and  a68332a );
 a68344a <=( (not A167)  and  A169 );
 a68345a <=( (not A170)  and  a68344a );
 a68348a <=( (not A199)  and  (not A166) );
 a68351a <=( (not A233)  and  (not A200) );
 a68352a <=( a68351a  and  a68348a );
 a68353a <=( a68352a  and  a68345a );
 a68356a <=( (not A266)  and  (not A234) );
 a68359a <=( (not A269)  and  (not A268) );
 a68360a <=( a68359a  and  a68356a );
 a68363a <=( (not A299)  and  A298 );
 a68366a <=( A301  and  A300 );
 a68367a <=( a68366a  and  a68363a );
 a68368a <=( a68367a  and  a68360a );
 a68372a <=( (not A167)  and  A169 );
 a68373a <=( (not A170)  and  a68372a );
 a68376a <=( (not A199)  and  (not A166) );
 a68379a <=( (not A233)  and  (not A200) );
 a68380a <=( a68379a  and  a68376a );
 a68381a <=( a68380a  and  a68373a );
 a68384a <=( (not A266)  and  (not A234) );
 a68387a <=( (not A269)  and  (not A268) );
 a68388a <=( a68387a  and  a68384a );
 a68391a <=( (not A299)  and  A298 );
 a68394a <=( A302  and  A300 );
 a68395a <=( a68394a  and  a68391a );
 a68396a <=( a68395a  and  a68388a );
 a68400a <=( (not A167)  and  A169 );
 a68401a <=( (not A170)  and  a68400a );
 a68404a <=( (not A199)  and  (not A166) );
 a68407a <=( (not A232)  and  (not A200) );
 a68408a <=( a68407a  and  a68404a );
 a68409a <=( a68408a  and  a68401a );
 a68412a <=( (not A266)  and  (not A233) );
 a68415a <=( (not A269)  and  (not A268) );
 a68416a <=( a68415a  and  a68412a );
 a68419a <=( (not A299)  and  A298 );
 a68422a <=( A301  and  A300 );
 a68423a <=( a68422a  and  a68419a );
 a68424a <=( a68423a  and  a68416a );
 a68428a <=( (not A167)  and  A169 );
 a68429a <=( (not A170)  and  a68428a );
 a68432a <=( (not A199)  and  (not A166) );
 a68435a <=( (not A232)  and  (not A200) );
 a68436a <=( a68435a  and  a68432a );
 a68437a <=( a68436a  and  a68429a );
 a68440a <=( (not A266)  and  (not A233) );
 a68443a <=( (not A269)  and  (not A268) );
 a68444a <=( a68443a  and  a68440a );
 a68447a <=( (not A299)  and  A298 );
 a68450a <=( A302  and  A300 );
 a68451a <=( a68450a  and  a68447a );
 a68452a <=( a68451a  and  a68444a );
 a68456a <=( (not A166)  and  (not A167) );
 a68457a <=( (not A169)  and  a68456a );
 a68460a <=( A200  and  (not A199) );
 a68463a <=( (not A235)  and  (not A233) );
 a68464a <=( a68463a  and  a68460a );
 a68465a <=( a68464a  and  a68457a );
 a68468a <=( (not A266)  and  (not A236) );
 a68471a <=( (not A269)  and  (not A268) );
 a68472a <=( a68471a  and  a68468a );
 a68475a <=( (not A299)  and  A298 );
 a68478a <=( A301  and  A300 );
 a68479a <=( a68478a  and  a68475a );
 a68480a <=( a68479a  and  a68472a );
 a68484a <=( (not A166)  and  (not A167) );
 a68485a <=( (not A169)  and  a68484a );
 a68488a <=( A200  and  (not A199) );
 a68491a <=( (not A235)  and  (not A233) );
 a68492a <=( a68491a  and  a68488a );
 a68493a <=( a68492a  and  a68485a );
 a68496a <=( (not A266)  and  (not A236) );
 a68499a <=( (not A269)  and  (not A268) );
 a68500a <=( a68499a  and  a68496a );
 a68503a <=( (not A299)  and  A298 );
 a68506a <=( A302  and  A300 );
 a68507a <=( a68506a  and  a68503a );
 a68508a <=( a68507a  and  a68500a );
 a68512a <=( (not A166)  and  (not A167) );
 a68513a <=( (not A169)  and  a68512a );
 a68516a <=( (not A200)  and  A199 );
 a68519a <=( A202  and  A201 );
 a68520a <=( a68519a  and  a68516a );
 a68521a <=( a68520a  and  a68513a );
 a68524a <=( A233  and  A232 );
 a68527a <=( (not A267)  and  A265 );
 a68528a <=( a68527a  and  a68524a );
 a68531a <=( (not A299)  and  A298 );
 a68534a <=( A301  and  A300 );
 a68535a <=( a68534a  and  a68531a );
 a68536a <=( a68535a  and  a68528a );
 a68540a <=( (not A166)  and  (not A167) );
 a68541a <=( (not A169)  and  a68540a );
 a68544a <=( (not A200)  and  A199 );
 a68547a <=( A202  and  A201 );
 a68548a <=( a68547a  and  a68544a );
 a68549a <=( a68548a  and  a68541a );
 a68552a <=( A233  and  A232 );
 a68555a <=( (not A267)  and  A265 );
 a68556a <=( a68555a  and  a68552a );
 a68559a <=( (not A299)  and  A298 );
 a68562a <=( A302  and  A300 );
 a68563a <=( a68562a  and  a68559a );
 a68564a <=( a68563a  and  a68556a );
 a68568a <=( (not A166)  and  (not A167) );
 a68569a <=( (not A169)  and  a68568a );
 a68572a <=( (not A200)  and  A199 );
 a68575a <=( A202  and  A201 );
 a68576a <=( a68575a  and  a68572a );
 a68577a <=( a68576a  and  a68569a );
 a68580a <=( A233  and  A232 );
 a68583a <=( A266  and  A265 );
 a68584a <=( a68583a  and  a68580a );
 a68587a <=( (not A299)  and  A298 );
 a68590a <=( A301  and  A300 );
 a68591a <=( a68590a  and  a68587a );
 a68592a <=( a68591a  and  a68584a );
 a68596a <=( (not A166)  and  (not A167) );
 a68597a <=( (not A169)  and  a68596a );
 a68600a <=( (not A200)  and  A199 );
 a68603a <=( A202  and  A201 );
 a68604a <=( a68603a  and  a68600a );
 a68605a <=( a68604a  and  a68597a );
 a68608a <=( A233  and  A232 );
 a68611a <=( A266  and  A265 );
 a68612a <=( a68611a  and  a68608a );
 a68615a <=( (not A299)  and  A298 );
 a68618a <=( A302  and  A300 );
 a68619a <=( a68618a  and  a68615a );
 a68620a <=( a68619a  and  a68612a );
 a68624a <=( (not A166)  and  (not A167) );
 a68625a <=( (not A169)  and  a68624a );
 a68628a <=( (not A200)  and  A199 );
 a68631a <=( A202  and  A201 );
 a68632a <=( a68631a  and  a68628a );
 a68633a <=( a68632a  and  a68625a );
 a68636a <=( A233  and  A232 );
 a68639a <=( (not A266)  and  (not A265) );
 a68640a <=( a68639a  and  a68636a );
 a68643a <=( (not A299)  and  A298 );
 a68646a <=( A301  and  A300 );
 a68647a <=( a68646a  and  a68643a );
 a68648a <=( a68647a  and  a68640a );
 a68652a <=( (not A166)  and  (not A167) );
 a68653a <=( (not A169)  and  a68652a );
 a68656a <=( (not A200)  and  A199 );
 a68659a <=( A202  and  A201 );
 a68660a <=( a68659a  and  a68656a );
 a68661a <=( a68660a  and  a68653a );
 a68664a <=( A233  and  A232 );
 a68667a <=( (not A266)  and  (not A265) );
 a68668a <=( a68667a  and  a68664a );
 a68671a <=( (not A299)  and  A298 );
 a68674a <=( A302  and  A300 );
 a68675a <=( a68674a  and  a68671a );
 a68676a <=( a68675a  and  a68668a );
 a68680a <=( (not A166)  and  (not A167) );
 a68681a <=( (not A169)  and  a68680a );
 a68684a <=( (not A200)  and  A199 );
 a68687a <=( A202  and  A201 );
 a68688a <=( a68687a  and  a68684a );
 a68689a <=( a68688a  and  a68681a );
 a68692a <=( (not A235)  and  (not A233) );
 a68695a <=( (not A266)  and  (not A236) );
 a68696a <=( a68695a  and  a68692a );
 a68699a <=( (not A269)  and  (not A268) );
 a68702a <=( A299  and  (not A298) );
 a68703a <=( a68702a  and  a68699a );
 a68704a <=( a68703a  and  a68696a );
 a68708a <=( (not A166)  and  (not A167) );
 a68709a <=( (not A169)  and  a68708a );
 a68712a <=( (not A200)  and  A199 );
 a68715a <=( A202  and  A201 );
 a68716a <=( a68715a  and  a68712a );
 a68717a <=( a68716a  and  a68709a );
 a68720a <=( (not A234)  and  (not A233) );
 a68723a <=( A266  and  A265 );
 a68724a <=( a68723a  and  a68720a );
 a68727a <=( (not A299)  and  A298 );
 a68730a <=( A301  and  A300 );
 a68731a <=( a68730a  and  a68727a );
 a68732a <=( a68731a  and  a68724a );
 a68736a <=( (not A166)  and  (not A167) );
 a68737a <=( (not A169)  and  a68736a );
 a68740a <=( (not A200)  and  A199 );
 a68743a <=( A202  and  A201 );
 a68744a <=( a68743a  and  a68740a );
 a68745a <=( a68744a  and  a68737a );
 a68748a <=( (not A234)  and  (not A233) );
 a68751a <=( A266  and  A265 );
 a68752a <=( a68751a  and  a68748a );
 a68755a <=( (not A299)  and  A298 );
 a68758a <=( A302  and  A300 );
 a68759a <=( a68758a  and  a68755a );
 a68760a <=( a68759a  and  a68752a );
 a68764a <=( (not A166)  and  (not A167) );
 a68765a <=( (not A169)  and  a68764a );
 a68768a <=( (not A200)  and  A199 );
 a68771a <=( A202  and  A201 );
 a68772a <=( a68771a  and  a68768a );
 a68773a <=( a68772a  and  a68765a );
 a68776a <=( (not A234)  and  (not A233) );
 a68779a <=( (not A267)  and  (not A266) );
 a68780a <=( a68779a  and  a68776a );
 a68783a <=( (not A299)  and  A298 );
 a68786a <=( A301  and  A300 );
 a68787a <=( a68786a  and  a68783a );
 a68788a <=( a68787a  and  a68780a );
 a68792a <=( (not A166)  and  (not A167) );
 a68793a <=( (not A169)  and  a68792a );
 a68796a <=( (not A200)  and  A199 );
 a68799a <=( A202  and  A201 );
 a68800a <=( a68799a  and  a68796a );
 a68801a <=( a68800a  and  a68793a );
 a68804a <=( (not A234)  and  (not A233) );
 a68807a <=( (not A267)  and  (not A266) );
 a68808a <=( a68807a  and  a68804a );
 a68811a <=( (not A299)  and  A298 );
 a68814a <=( A302  and  A300 );
 a68815a <=( a68814a  and  a68811a );
 a68816a <=( a68815a  and  a68808a );
 a68820a <=( (not A166)  and  (not A167) );
 a68821a <=( (not A169)  and  a68820a );
 a68824a <=( (not A200)  and  A199 );
 a68827a <=( A202  and  A201 );
 a68828a <=( a68827a  and  a68824a );
 a68829a <=( a68828a  and  a68821a );
 a68832a <=( (not A234)  and  (not A233) );
 a68835a <=( (not A266)  and  (not A265) );
 a68836a <=( a68835a  and  a68832a );
 a68839a <=( (not A299)  and  A298 );
 a68842a <=( A301  and  A300 );
 a68843a <=( a68842a  and  a68839a );
 a68844a <=( a68843a  and  a68836a );
 a68848a <=( (not A166)  and  (not A167) );
 a68849a <=( (not A169)  and  a68848a );
 a68852a <=( (not A200)  and  A199 );
 a68855a <=( A202  and  A201 );
 a68856a <=( a68855a  and  a68852a );
 a68857a <=( a68856a  and  a68849a );
 a68860a <=( (not A234)  and  (not A233) );
 a68863a <=( (not A266)  and  (not A265) );
 a68864a <=( a68863a  and  a68860a );
 a68867a <=( (not A299)  and  A298 );
 a68870a <=( A302  and  A300 );
 a68871a <=( a68870a  and  a68867a );
 a68872a <=( a68871a  and  a68864a );
 a68876a <=( (not A166)  and  (not A167) );
 a68877a <=( (not A169)  and  a68876a );
 a68880a <=( (not A200)  and  A199 );
 a68883a <=( A202  and  A201 );
 a68884a <=( a68883a  and  a68880a );
 a68885a <=( a68884a  and  a68877a );
 a68888a <=( (not A233)  and  A232 );
 a68891a <=( A235  and  A234 );
 a68892a <=( a68891a  and  a68888a );
 a68895a <=( (not A266)  and  A265 );
 a68898a <=( A268  and  A267 );
 a68899a <=( a68898a  and  a68895a );
 a68900a <=( a68899a  and  a68892a );
 a68904a <=( (not A166)  and  (not A167) );
 a68905a <=( (not A169)  and  a68904a );
 a68908a <=( (not A200)  and  A199 );
 a68911a <=( A202  and  A201 );
 a68912a <=( a68911a  and  a68908a );
 a68913a <=( a68912a  and  a68905a );
 a68916a <=( (not A233)  and  A232 );
 a68919a <=( A235  and  A234 );
 a68920a <=( a68919a  and  a68916a );
 a68923a <=( (not A266)  and  A265 );
 a68926a <=( A269  and  A267 );
 a68927a <=( a68926a  and  a68923a );
 a68928a <=( a68927a  and  a68920a );
 a68932a <=( (not A166)  and  (not A167) );
 a68933a <=( (not A169)  and  a68932a );
 a68936a <=( (not A200)  and  A199 );
 a68939a <=( A202  and  A201 );
 a68940a <=( a68939a  and  a68936a );
 a68941a <=( a68940a  and  a68933a );
 a68944a <=( (not A233)  and  A232 );
 a68947a <=( A236  and  A234 );
 a68948a <=( a68947a  and  a68944a );
 a68951a <=( (not A266)  and  A265 );
 a68954a <=( A268  and  A267 );
 a68955a <=( a68954a  and  a68951a );
 a68956a <=( a68955a  and  a68948a );
 a68960a <=( (not A166)  and  (not A167) );
 a68961a <=( (not A169)  and  a68960a );
 a68964a <=( (not A200)  and  A199 );
 a68967a <=( A202  and  A201 );
 a68968a <=( a68967a  and  a68964a );
 a68969a <=( a68968a  and  a68961a );
 a68972a <=( (not A233)  and  A232 );
 a68975a <=( A236  and  A234 );
 a68976a <=( a68975a  and  a68972a );
 a68979a <=( (not A266)  and  A265 );
 a68982a <=( A269  and  A267 );
 a68983a <=( a68982a  and  a68979a );
 a68984a <=( a68983a  and  a68976a );
 a68988a <=( (not A166)  and  (not A167) );
 a68989a <=( (not A169)  and  a68988a );
 a68992a <=( (not A200)  and  A199 );
 a68995a <=( A202  and  A201 );
 a68996a <=( a68995a  and  a68992a );
 a68997a <=( a68996a  and  a68989a );
 a69000a <=( (not A233)  and  (not A232) );
 a69003a <=( A266  and  A265 );
 a69004a <=( a69003a  and  a69000a );
 a69007a <=( (not A299)  and  A298 );
 a69010a <=( A301  and  A300 );
 a69011a <=( a69010a  and  a69007a );
 a69012a <=( a69011a  and  a69004a );
 a69016a <=( (not A166)  and  (not A167) );
 a69017a <=( (not A169)  and  a69016a );
 a69020a <=( (not A200)  and  A199 );
 a69023a <=( A202  and  A201 );
 a69024a <=( a69023a  and  a69020a );
 a69025a <=( a69024a  and  a69017a );
 a69028a <=( (not A233)  and  (not A232) );
 a69031a <=( A266  and  A265 );
 a69032a <=( a69031a  and  a69028a );
 a69035a <=( (not A299)  and  A298 );
 a69038a <=( A302  and  A300 );
 a69039a <=( a69038a  and  a69035a );
 a69040a <=( a69039a  and  a69032a );
 a69044a <=( (not A166)  and  (not A167) );
 a69045a <=( (not A169)  and  a69044a );
 a69048a <=( (not A200)  and  A199 );
 a69051a <=( A202  and  A201 );
 a69052a <=( a69051a  and  a69048a );
 a69053a <=( a69052a  and  a69045a );
 a69056a <=( (not A233)  and  (not A232) );
 a69059a <=( (not A267)  and  (not A266) );
 a69060a <=( a69059a  and  a69056a );
 a69063a <=( (not A299)  and  A298 );
 a69066a <=( A301  and  A300 );
 a69067a <=( a69066a  and  a69063a );
 a69068a <=( a69067a  and  a69060a );
 a69072a <=( (not A166)  and  (not A167) );
 a69073a <=( (not A169)  and  a69072a );
 a69076a <=( (not A200)  and  A199 );
 a69079a <=( A202  and  A201 );
 a69080a <=( a69079a  and  a69076a );
 a69081a <=( a69080a  and  a69073a );
 a69084a <=( (not A233)  and  (not A232) );
 a69087a <=( (not A267)  and  (not A266) );
 a69088a <=( a69087a  and  a69084a );
 a69091a <=( (not A299)  and  A298 );
 a69094a <=( A302  and  A300 );
 a69095a <=( a69094a  and  a69091a );
 a69096a <=( a69095a  and  a69088a );
 a69100a <=( (not A166)  and  (not A167) );
 a69101a <=( (not A169)  and  a69100a );
 a69104a <=( (not A200)  and  A199 );
 a69107a <=( A202  and  A201 );
 a69108a <=( a69107a  and  a69104a );
 a69109a <=( a69108a  and  a69101a );
 a69112a <=( (not A233)  and  (not A232) );
 a69115a <=( (not A266)  and  (not A265) );
 a69116a <=( a69115a  and  a69112a );
 a69119a <=( (not A299)  and  A298 );
 a69122a <=( A301  and  A300 );
 a69123a <=( a69122a  and  a69119a );
 a69124a <=( a69123a  and  a69116a );
 a69128a <=( (not A166)  and  (not A167) );
 a69129a <=( (not A169)  and  a69128a );
 a69132a <=( (not A200)  and  A199 );
 a69135a <=( A202  and  A201 );
 a69136a <=( a69135a  and  a69132a );
 a69137a <=( a69136a  and  a69129a );
 a69140a <=( (not A233)  and  (not A232) );
 a69143a <=( (not A266)  and  (not A265) );
 a69144a <=( a69143a  and  a69140a );
 a69147a <=( (not A299)  and  A298 );
 a69150a <=( A302  and  A300 );
 a69151a <=( a69150a  and  a69147a );
 a69152a <=( a69151a  and  a69144a );
 a69156a <=( (not A166)  and  (not A167) );
 a69157a <=( (not A169)  and  a69156a );
 a69160a <=( (not A200)  and  A199 );
 a69163a <=( A203  and  A201 );
 a69164a <=( a69163a  and  a69160a );
 a69165a <=( a69164a  and  a69157a );
 a69168a <=( A233  and  A232 );
 a69171a <=( (not A267)  and  A265 );
 a69172a <=( a69171a  and  a69168a );
 a69175a <=( (not A299)  and  A298 );
 a69178a <=( A301  and  A300 );
 a69179a <=( a69178a  and  a69175a );
 a69180a <=( a69179a  and  a69172a );
 a69184a <=( (not A166)  and  (not A167) );
 a69185a <=( (not A169)  and  a69184a );
 a69188a <=( (not A200)  and  A199 );
 a69191a <=( A203  and  A201 );
 a69192a <=( a69191a  and  a69188a );
 a69193a <=( a69192a  and  a69185a );
 a69196a <=( A233  and  A232 );
 a69199a <=( (not A267)  and  A265 );
 a69200a <=( a69199a  and  a69196a );
 a69203a <=( (not A299)  and  A298 );
 a69206a <=( A302  and  A300 );
 a69207a <=( a69206a  and  a69203a );
 a69208a <=( a69207a  and  a69200a );
 a69212a <=( (not A166)  and  (not A167) );
 a69213a <=( (not A169)  and  a69212a );
 a69216a <=( (not A200)  and  A199 );
 a69219a <=( A203  and  A201 );
 a69220a <=( a69219a  and  a69216a );
 a69221a <=( a69220a  and  a69213a );
 a69224a <=( A233  and  A232 );
 a69227a <=( A266  and  A265 );
 a69228a <=( a69227a  and  a69224a );
 a69231a <=( (not A299)  and  A298 );
 a69234a <=( A301  and  A300 );
 a69235a <=( a69234a  and  a69231a );
 a69236a <=( a69235a  and  a69228a );
 a69240a <=( (not A166)  and  (not A167) );
 a69241a <=( (not A169)  and  a69240a );
 a69244a <=( (not A200)  and  A199 );
 a69247a <=( A203  and  A201 );
 a69248a <=( a69247a  and  a69244a );
 a69249a <=( a69248a  and  a69241a );
 a69252a <=( A233  and  A232 );
 a69255a <=( A266  and  A265 );
 a69256a <=( a69255a  and  a69252a );
 a69259a <=( (not A299)  and  A298 );
 a69262a <=( A302  and  A300 );
 a69263a <=( a69262a  and  a69259a );
 a69264a <=( a69263a  and  a69256a );
 a69268a <=( (not A166)  and  (not A167) );
 a69269a <=( (not A169)  and  a69268a );
 a69272a <=( (not A200)  and  A199 );
 a69275a <=( A203  and  A201 );
 a69276a <=( a69275a  and  a69272a );
 a69277a <=( a69276a  and  a69269a );
 a69280a <=( A233  and  A232 );
 a69283a <=( (not A266)  and  (not A265) );
 a69284a <=( a69283a  and  a69280a );
 a69287a <=( (not A299)  and  A298 );
 a69290a <=( A301  and  A300 );
 a69291a <=( a69290a  and  a69287a );
 a69292a <=( a69291a  and  a69284a );
 a69296a <=( (not A166)  and  (not A167) );
 a69297a <=( (not A169)  and  a69296a );
 a69300a <=( (not A200)  and  A199 );
 a69303a <=( A203  and  A201 );
 a69304a <=( a69303a  and  a69300a );
 a69305a <=( a69304a  and  a69297a );
 a69308a <=( A233  and  A232 );
 a69311a <=( (not A266)  and  (not A265) );
 a69312a <=( a69311a  and  a69308a );
 a69315a <=( (not A299)  and  A298 );
 a69318a <=( A302  and  A300 );
 a69319a <=( a69318a  and  a69315a );
 a69320a <=( a69319a  and  a69312a );
 a69324a <=( (not A166)  and  (not A167) );
 a69325a <=( (not A169)  and  a69324a );
 a69328a <=( (not A200)  and  A199 );
 a69331a <=( A203  and  A201 );
 a69332a <=( a69331a  and  a69328a );
 a69333a <=( a69332a  and  a69325a );
 a69336a <=( (not A235)  and  (not A233) );
 a69339a <=( (not A266)  and  (not A236) );
 a69340a <=( a69339a  and  a69336a );
 a69343a <=( (not A269)  and  (not A268) );
 a69346a <=( A299  and  (not A298) );
 a69347a <=( a69346a  and  a69343a );
 a69348a <=( a69347a  and  a69340a );
 a69352a <=( (not A166)  and  (not A167) );
 a69353a <=( (not A169)  and  a69352a );
 a69356a <=( (not A200)  and  A199 );
 a69359a <=( A203  and  A201 );
 a69360a <=( a69359a  and  a69356a );
 a69361a <=( a69360a  and  a69353a );
 a69364a <=( (not A234)  and  (not A233) );
 a69367a <=( A266  and  A265 );
 a69368a <=( a69367a  and  a69364a );
 a69371a <=( (not A299)  and  A298 );
 a69374a <=( A301  and  A300 );
 a69375a <=( a69374a  and  a69371a );
 a69376a <=( a69375a  and  a69368a );
 a69380a <=( (not A166)  and  (not A167) );
 a69381a <=( (not A169)  and  a69380a );
 a69384a <=( (not A200)  and  A199 );
 a69387a <=( A203  and  A201 );
 a69388a <=( a69387a  and  a69384a );
 a69389a <=( a69388a  and  a69381a );
 a69392a <=( (not A234)  and  (not A233) );
 a69395a <=( A266  and  A265 );
 a69396a <=( a69395a  and  a69392a );
 a69399a <=( (not A299)  and  A298 );
 a69402a <=( A302  and  A300 );
 a69403a <=( a69402a  and  a69399a );
 a69404a <=( a69403a  and  a69396a );
 a69408a <=( (not A166)  and  (not A167) );
 a69409a <=( (not A169)  and  a69408a );
 a69412a <=( (not A200)  and  A199 );
 a69415a <=( A203  and  A201 );
 a69416a <=( a69415a  and  a69412a );
 a69417a <=( a69416a  and  a69409a );
 a69420a <=( (not A234)  and  (not A233) );
 a69423a <=( (not A267)  and  (not A266) );
 a69424a <=( a69423a  and  a69420a );
 a69427a <=( (not A299)  and  A298 );
 a69430a <=( A301  and  A300 );
 a69431a <=( a69430a  and  a69427a );
 a69432a <=( a69431a  and  a69424a );
 a69436a <=( (not A166)  and  (not A167) );
 a69437a <=( (not A169)  and  a69436a );
 a69440a <=( (not A200)  and  A199 );
 a69443a <=( A203  and  A201 );
 a69444a <=( a69443a  and  a69440a );
 a69445a <=( a69444a  and  a69437a );
 a69448a <=( (not A234)  and  (not A233) );
 a69451a <=( (not A267)  and  (not A266) );
 a69452a <=( a69451a  and  a69448a );
 a69455a <=( (not A299)  and  A298 );
 a69458a <=( A302  and  A300 );
 a69459a <=( a69458a  and  a69455a );
 a69460a <=( a69459a  and  a69452a );
 a69464a <=( (not A166)  and  (not A167) );
 a69465a <=( (not A169)  and  a69464a );
 a69468a <=( (not A200)  and  A199 );
 a69471a <=( A203  and  A201 );
 a69472a <=( a69471a  and  a69468a );
 a69473a <=( a69472a  and  a69465a );
 a69476a <=( (not A234)  and  (not A233) );
 a69479a <=( (not A266)  and  (not A265) );
 a69480a <=( a69479a  and  a69476a );
 a69483a <=( (not A299)  and  A298 );
 a69486a <=( A301  and  A300 );
 a69487a <=( a69486a  and  a69483a );
 a69488a <=( a69487a  and  a69480a );
 a69492a <=( (not A166)  and  (not A167) );
 a69493a <=( (not A169)  and  a69492a );
 a69496a <=( (not A200)  and  A199 );
 a69499a <=( A203  and  A201 );
 a69500a <=( a69499a  and  a69496a );
 a69501a <=( a69500a  and  a69493a );
 a69504a <=( (not A234)  and  (not A233) );
 a69507a <=( (not A266)  and  (not A265) );
 a69508a <=( a69507a  and  a69504a );
 a69511a <=( (not A299)  and  A298 );
 a69514a <=( A302  and  A300 );
 a69515a <=( a69514a  and  a69511a );
 a69516a <=( a69515a  and  a69508a );
 a69520a <=( (not A166)  and  (not A167) );
 a69521a <=( (not A169)  and  a69520a );
 a69524a <=( (not A200)  and  A199 );
 a69527a <=( A203  and  A201 );
 a69528a <=( a69527a  and  a69524a );
 a69529a <=( a69528a  and  a69521a );
 a69532a <=( (not A233)  and  A232 );
 a69535a <=( A235  and  A234 );
 a69536a <=( a69535a  and  a69532a );
 a69539a <=( (not A266)  and  A265 );
 a69542a <=( A268  and  A267 );
 a69543a <=( a69542a  and  a69539a );
 a69544a <=( a69543a  and  a69536a );
 a69548a <=( (not A166)  and  (not A167) );
 a69549a <=( (not A169)  and  a69548a );
 a69552a <=( (not A200)  and  A199 );
 a69555a <=( A203  and  A201 );
 a69556a <=( a69555a  and  a69552a );
 a69557a <=( a69556a  and  a69549a );
 a69560a <=( (not A233)  and  A232 );
 a69563a <=( A235  and  A234 );
 a69564a <=( a69563a  and  a69560a );
 a69567a <=( (not A266)  and  A265 );
 a69570a <=( A269  and  A267 );
 a69571a <=( a69570a  and  a69567a );
 a69572a <=( a69571a  and  a69564a );
 a69576a <=( (not A166)  and  (not A167) );
 a69577a <=( (not A169)  and  a69576a );
 a69580a <=( (not A200)  and  A199 );
 a69583a <=( A203  and  A201 );
 a69584a <=( a69583a  and  a69580a );
 a69585a <=( a69584a  and  a69577a );
 a69588a <=( (not A233)  and  A232 );
 a69591a <=( A236  and  A234 );
 a69592a <=( a69591a  and  a69588a );
 a69595a <=( (not A266)  and  A265 );
 a69598a <=( A268  and  A267 );
 a69599a <=( a69598a  and  a69595a );
 a69600a <=( a69599a  and  a69592a );
 a69604a <=( (not A166)  and  (not A167) );
 a69605a <=( (not A169)  and  a69604a );
 a69608a <=( (not A200)  and  A199 );
 a69611a <=( A203  and  A201 );
 a69612a <=( a69611a  and  a69608a );
 a69613a <=( a69612a  and  a69605a );
 a69616a <=( (not A233)  and  A232 );
 a69619a <=( A236  and  A234 );
 a69620a <=( a69619a  and  a69616a );
 a69623a <=( (not A266)  and  A265 );
 a69626a <=( A269  and  A267 );
 a69627a <=( a69626a  and  a69623a );
 a69628a <=( a69627a  and  a69620a );
 a69632a <=( (not A166)  and  (not A167) );
 a69633a <=( (not A169)  and  a69632a );
 a69636a <=( (not A200)  and  A199 );
 a69639a <=( A203  and  A201 );
 a69640a <=( a69639a  and  a69636a );
 a69641a <=( a69640a  and  a69633a );
 a69644a <=( (not A233)  and  (not A232) );
 a69647a <=( A266  and  A265 );
 a69648a <=( a69647a  and  a69644a );
 a69651a <=( (not A299)  and  A298 );
 a69654a <=( A301  and  A300 );
 a69655a <=( a69654a  and  a69651a );
 a69656a <=( a69655a  and  a69648a );
 a69660a <=( (not A166)  and  (not A167) );
 a69661a <=( (not A169)  and  a69660a );
 a69664a <=( (not A200)  and  A199 );
 a69667a <=( A203  and  A201 );
 a69668a <=( a69667a  and  a69664a );
 a69669a <=( a69668a  and  a69661a );
 a69672a <=( (not A233)  and  (not A232) );
 a69675a <=( A266  and  A265 );
 a69676a <=( a69675a  and  a69672a );
 a69679a <=( (not A299)  and  A298 );
 a69682a <=( A302  and  A300 );
 a69683a <=( a69682a  and  a69679a );
 a69684a <=( a69683a  and  a69676a );
 a69688a <=( (not A166)  and  (not A167) );
 a69689a <=( (not A169)  and  a69688a );
 a69692a <=( (not A200)  and  A199 );
 a69695a <=( A203  and  A201 );
 a69696a <=( a69695a  and  a69692a );
 a69697a <=( a69696a  and  a69689a );
 a69700a <=( (not A233)  and  (not A232) );
 a69703a <=( (not A267)  and  (not A266) );
 a69704a <=( a69703a  and  a69700a );
 a69707a <=( (not A299)  and  A298 );
 a69710a <=( A301  and  A300 );
 a69711a <=( a69710a  and  a69707a );
 a69712a <=( a69711a  and  a69704a );
 a69716a <=( (not A166)  and  (not A167) );
 a69717a <=( (not A169)  and  a69716a );
 a69720a <=( (not A200)  and  A199 );
 a69723a <=( A203  and  A201 );
 a69724a <=( a69723a  and  a69720a );
 a69725a <=( a69724a  and  a69717a );
 a69728a <=( (not A233)  and  (not A232) );
 a69731a <=( (not A267)  and  (not A266) );
 a69732a <=( a69731a  and  a69728a );
 a69735a <=( (not A299)  and  A298 );
 a69738a <=( A302  and  A300 );
 a69739a <=( a69738a  and  a69735a );
 a69740a <=( a69739a  and  a69732a );
 a69744a <=( (not A166)  and  (not A167) );
 a69745a <=( (not A169)  and  a69744a );
 a69748a <=( (not A200)  and  A199 );
 a69751a <=( A203  and  A201 );
 a69752a <=( a69751a  and  a69748a );
 a69753a <=( a69752a  and  a69745a );
 a69756a <=( (not A233)  and  (not A232) );
 a69759a <=( (not A266)  and  (not A265) );
 a69760a <=( a69759a  and  a69756a );
 a69763a <=( (not A299)  and  A298 );
 a69766a <=( A301  and  A300 );
 a69767a <=( a69766a  and  a69763a );
 a69768a <=( a69767a  and  a69760a );
 a69772a <=( (not A166)  and  (not A167) );
 a69773a <=( (not A169)  and  a69772a );
 a69776a <=( (not A200)  and  A199 );
 a69779a <=( A203  and  A201 );
 a69780a <=( a69779a  and  a69776a );
 a69781a <=( a69780a  and  a69773a );
 a69784a <=( (not A233)  and  (not A232) );
 a69787a <=( (not A266)  and  (not A265) );
 a69788a <=( a69787a  and  a69784a );
 a69791a <=( (not A299)  and  A298 );
 a69794a <=( A302  and  A300 );
 a69795a <=( a69794a  and  a69791a );
 a69796a <=( a69795a  and  a69788a );
 a69800a <=( A167  and  (not A168) );
 a69801a <=( (not A169)  and  a69800a );
 a69804a <=( (not A199)  and  A166 );
 a69807a <=( A232  and  A200 );
 a69808a <=( a69807a  and  a69804a );
 a69809a <=( a69808a  and  a69801a );
 a69812a <=( A265  and  A233 );
 a69815a <=( (not A269)  and  (not A268) );
 a69816a <=( a69815a  and  a69812a );
 a69819a <=( (not A299)  and  A298 );
 a69822a <=( A301  and  A300 );
 a69823a <=( a69822a  and  a69819a );
 a69824a <=( a69823a  and  a69816a );
 a69828a <=( A167  and  (not A168) );
 a69829a <=( (not A169)  and  a69828a );
 a69832a <=( (not A199)  and  A166 );
 a69835a <=( A232  and  A200 );
 a69836a <=( a69835a  and  a69832a );
 a69837a <=( a69836a  and  a69829a );
 a69840a <=( A265  and  A233 );
 a69843a <=( (not A269)  and  (not A268) );
 a69844a <=( a69843a  and  a69840a );
 a69847a <=( (not A299)  and  A298 );
 a69850a <=( A302  and  A300 );
 a69851a <=( a69850a  and  a69847a );
 a69852a <=( a69851a  and  a69844a );
 a69856a <=( A167  and  (not A168) );
 a69857a <=( (not A169)  and  a69856a );
 a69860a <=( (not A199)  and  A166 );
 a69863a <=( (not A233)  and  A200 );
 a69864a <=( a69863a  and  a69860a );
 a69865a <=( a69864a  and  a69857a );
 a69868a <=( (not A236)  and  (not A235) );
 a69871a <=( A266  and  A265 );
 a69872a <=( a69871a  and  a69868a );
 a69875a <=( (not A299)  and  A298 );
 a69878a <=( A301  and  A300 );
 a69879a <=( a69878a  and  a69875a );
 a69880a <=( a69879a  and  a69872a );
 a69884a <=( A167  and  (not A168) );
 a69885a <=( (not A169)  and  a69884a );
 a69888a <=( (not A199)  and  A166 );
 a69891a <=( (not A233)  and  A200 );
 a69892a <=( a69891a  and  a69888a );
 a69893a <=( a69892a  and  a69885a );
 a69896a <=( (not A236)  and  (not A235) );
 a69899a <=( A266  and  A265 );
 a69900a <=( a69899a  and  a69896a );
 a69903a <=( (not A299)  and  A298 );
 a69906a <=( A302  and  A300 );
 a69907a <=( a69906a  and  a69903a );
 a69908a <=( a69907a  and  a69900a );
 a69912a <=( A167  and  (not A168) );
 a69913a <=( (not A169)  and  a69912a );
 a69916a <=( (not A199)  and  A166 );
 a69919a <=( (not A233)  and  A200 );
 a69920a <=( a69919a  and  a69916a );
 a69921a <=( a69920a  and  a69913a );
 a69924a <=( (not A236)  and  (not A235) );
 a69927a <=( (not A267)  and  (not A266) );
 a69928a <=( a69927a  and  a69924a );
 a69931a <=( (not A299)  and  A298 );
 a69934a <=( A301  and  A300 );
 a69935a <=( a69934a  and  a69931a );
 a69936a <=( a69935a  and  a69928a );
 a69940a <=( A167  and  (not A168) );
 a69941a <=( (not A169)  and  a69940a );
 a69944a <=( (not A199)  and  A166 );
 a69947a <=( (not A233)  and  A200 );
 a69948a <=( a69947a  and  a69944a );
 a69949a <=( a69948a  and  a69941a );
 a69952a <=( (not A236)  and  (not A235) );
 a69955a <=( (not A267)  and  (not A266) );
 a69956a <=( a69955a  and  a69952a );
 a69959a <=( (not A299)  and  A298 );
 a69962a <=( A302  and  A300 );
 a69963a <=( a69962a  and  a69959a );
 a69964a <=( a69963a  and  a69956a );
 a69968a <=( A167  and  (not A168) );
 a69969a <=( (not A169)  and  a69968a );
 a69972a <=( (not A199)  and  A166 );
 a69975a <=( (not A233)  and  A200 );
 a69976a <=( a69975a  and  a69972a );
 a69977a <=( a69976a  and  a69969a );
 a69980a <=( (not A236)  and  (not A235) );
 a69983a <=( (not A266)  and  (not A265) );
 a69984a <=( a69983a  and  a69980a );
 a69987a <=( (not A299)  and  A298 );
 a69990a <=( A301  and  A300 );
 a69991a <=( a69990a  and  a69987a );
 a69992a <=( a69991a  and  a69984a );
 a69996a <=( A167  and  (not A168) );
 a69997a <=( (not A169)  and  a69996a );
 a70000a <=( (not A199)  and  A166 );
 a70003a <=( (not A233)  and  A200 );
 a70004a <=( a70003a  and  a70000a );
 a70005a <=( a70004a  and  a69997a );
 a70008a <=( (not A236)  and  (not A235) );
 a70011a <=( (not A266)  and  (not A265) );
 a70012a <=( a70011a  and  a70008a );
 a70015a <=( (not A299)  and  A298 );
 a70018a <=( A302  and  A300 );
 a70019a <=( a70018a  and  a70015a );
 a70020a <=( a70019a  and  a70012a );
 a70024a <=( A167  and  (not A168) );
 a70025a <=( (not A169)  and  a70024a );
 a70028a <=( (not A199)  and  A166 );
 a70031a <=( (not A233)  and  A200 );
 a70032a <=( a70031a  and  a70028a );
 a70033a <=( a70032a  and  a70025a );
 a70036a <=( (not A266)  and  (not A234) );
 a70039a <=( (not A269)  and  (not A268) );
 a70040a <=( a70039a  and  a70036a );
 a70043a <=( (not A299)  and  A298 );
 a70046a <=( A301  and  A300 );
 a70047a <=( a70046a  and  a70043a );
 a70048a <=( a70047a  and  a70040a );
 a70052a <=( A167  and  (not A168) );
 a70053a <=( (not A169)  and  a70052a );
 a70056a <=( (not A199)  and  A166 );
 a70059a <=( (not A233)  and  A200 );
 a70060a <=( a70059a  and  a70056a );
 a70061a <=( a70060a  and  a70053a );
 a70064a <=( (not A266)  and  (not A234) );
 a70067a <=( (not A269)  and  (not A268) );
 a70068a <=( a70067a  and  a70064a );
 a70071a <=( (not A299)  and  A298 );
 a70074a <=( A302  and  A300 );
 a70075a <=( a70074a  and  a70071a );
 a70076a <=( a70075a  and  a70068a );
 a70080a <=( A167  and  (not A168) );
 a70081a <=( (not A169)  and  a70080a );
 a70084a <=( (not A199)  and  A166 );
 a70087a <=( (not A232)  and  A200 );
 a70088a <=( a70087a  and  a70084a );
 a70089a <=( a70088a  and  a70081a );
 a70092a <=( (not A266)  and  (not A233) );
 a70095a <=( (not A269)  and  (not A268) );
 a70096a <=( a70095a  and  a70092a );
 a70099a <=( (not A299)  and  A298 );
 a70102a <=( A301  and  A300 );
 a70103a <=( a70102a  and  a70099a );
 a70104a <=( a70103a  and  a70096a );
 a70108a <=( A167  and  (not A168) );
 a70109a <=( (not A169)  and  a70108a );
 a70112a <=( (not A199)  and  A166 );
 a70115a <=( (not A232)  and  A200 );
 a70116a <=( a70115a  and  a70112a );
 a70117a <=( a70116a  and  a70109a );
 a70120a <=( (not A266)  and  (not A233) );
 a70123a <=( (not A269)  and  (not A268) );
 a70124a <=( a70123a  and  a70120a );
 a70127a <=( (not A299)  and  A298 );
 a70130a <=( A302  and  A300 );
 a70131a <=( a70130a  and  a70127a );
 a70132a <=( a70131a  and  a70124a );
 a70136a <=( A167  and  (not A168) );
 a70137a <=( (not A169)  and  a70136a );
 a70140a <=( A199  and  A166 );
 a70143a <=( A201  and  (not A200) );
 a70144a <=( a70143a  and  a70140a );
 a70145a <=( a70144a  and  a70137a );
 a70148a <=( A232  and  A202 );
 a70151a <=( A265  and  A233 );
 a70152a <=( a70151a  and  a70148a );
 a70155a <=( (not A269)  and  (not A268) );
 a70158a <=( A299  and  (not A298) );
 a70159a <=( a70158a  and  a70155a );
 a70160a <=( a70159a  and  a70152a );
 a70164a <=( A167  and  (not A168) );
 a70165a <=( (not A169)  and  a70164a );
 a70168a <=( A199  and  A166 );
 a70171a <=( A201  and  (not A200) );
 a70172a <=( a70171a  and  a70168a );
 a70173a <=( a70172a  and  a70165a );
 a70176a <=( (not A233)  and  A202 );
 a70179a <=( (not A236)  and  (not A235) );
 a70180a <=( a70179a  and  a70176a );
 a70183a <=( A266  and  A265 );
 a70186a <=( A299  and  (not A298) );
 a70187a <=( a70186a  and  a70183a );
 a70188a <=( a70187a  and  a70180a );
 a70192a <=( A167  and  (not A168) );
 a70193a <=( (not A169)  and  a70192a );
 a70196a <=( A199  and  A166 );
 a70199a <=( A201  and  (not A200) );
 a70200a <=( a70199a  and  a70196a );
 a70201a <=( a70200a  and  a70193a );
 a70204a <=( (not A233)  and  A202 );
 a70207a <=( (not A236)  and  (not A235) );
 a70208a <=( a70207a  and  a70204a );
 a70211a <=( (not A267)  and  (not A266) );
 a70214a <=( A299  and  (not A298) );
 a70215a <=( a70214a  and  a70211a );
 a70216a <=( a70215a  and  a70208a );
 a70220a <=( A167  and  (not A168) );
 a70221a <=( (not A169)  and  a70220a );
 a70224a <=( A199  and  A166 );
 a70227a <=( A201  and  (not A200) );
 a70228a <=( a70227a  and  a70224a );
 a70229a <=( a70228a  and  a70221a );
 a70232a <=( (not A233)  and  A202 );
 a70235a <=( (not A236)  and  (not A235) );
 a70236a <=( a70235a  and  a70232a );
 a70239a <=( (not A266)  and  (not A265) );
 a70242a <=( A299  and  (not A298) );
 a70243a <=( a70242a  and  a70239a );
 a70244a <=( a70243a  and  a70236a );
 a70248a <=( A167  and  (not A168) );
 a70249a <=( (not A169)  and  a70248a );
 a70252a <=( A199  and  A166 );
 a70255a <=( A201  and  (not A200) );
 a70256a <=( a70255a  and  a70252a );
 a70257a <=( a70256a  and  a70249a );
 a70260a <=( (not A233)  and  A202 );
 a70263a <=( (not A266)  and  (not A234) );
 a70264a <=( a70263a  and  a70260a );
 a70267a <=( (not A269)  and  (not A268) );
 a70270a <=( A299  and  (not A298) );
 a70271a <=( a70270a  and  a70267a );
 a70272a <=( a70271a  and  a70264a );
 a70276a <=( A167  and  (not A168) );
 a70277a <=( (not A169)  and  a70276a );
 a70280a <=( A199  and  A166 );
 a70283a <=( A201  and  (not A200) );
 a70284a <=( a70283a  and  a70280a );
 a70285a <=( a70284a  and  a70277a );
 a70288a <=( A232  and  A202 );
 a70291a <=( A234  and  (not A233) );
 a70292a <=( a70291a  and  a70288a );
 a70295a <=( A298  and  A235 );
 a70298a <=( (not A302)  and  (not A301) );
 a70299a <=( a70298a  and  a70295a );
 a70300a <=( a70299a  and  a70292a );
 a70304a <=( A167  and  (not A168) );
 a70305a <=( (not A169)  and  a70304a );
 a70308a <=( A199  and  A166 );
 a70311a <=( A201  and  (not A200) );
 a70312a <=( a70311a  and  a70308a );
 a70313a <=( a70312a  and  a70305a );
 a70316a <=( A232  and  A202 );
 a70319a <=( A234  and  (not A233) );
 a70320a <=( a70319a  and  a70316a );
 a70323a <=( A298  and  A236 );
 a70326a <=( (not A302)  and  (not A301) );
 a70327a <=( a70326a  and  a70323a );
 a70328a <=( a70327a  and  a70320a );
 a70332a <=( A167  and  (not A168) );
 a70333a <=( (not A169)  and  a70332a );
 a70336a <=( A199  and  A166 );
 a70339a <=( A201  and  (not A200) );
 a70340a <=( a70339a  and  a70336a );
 a70341a <=( a70340a  and  a70333a );
 a70344a <=( (not A232)  and  A202 );
 a70347a <=( (not A266)  and  (not A233) );
 a70348a <=( a70347a  and  a70344a );
 a70351a <=( (not A269)  and  (not A268) );
 a70354a <=( A299  and  (not A298) );
 a70355a <=( a70354a  and  a70351a );
 a70356a <=( a70355a  and  a70348a );
 a70360a <=( A167  and  (not A168) );
 a70361a <=( (not A169)  and  a70360a );
 a70364a <=( A199  and  A166 );
 a70367a <=( A201  and  (not A200) );
 a70368a <=( a70367a  and  a70364a );
 a70369a <=( a70368a  and  a70361a );
 a70372a <=( A232  and  A203 );
 a70375a <=( A265  and  A233 );
 a70376a <=( a70375a  and  a70372a );
 a70379a <=( (not A269)  and  (not A268) );
 a70382a <=( A299  and  (not A298) );
 a70383a <=( a70382a  and  a70379a );
 a70384a <=( a70383a  and  a70376a );
 a70388a <=( A167  and  (not A168) );
 a70389a <=( (not A169)  and  a70388a );
 a70392a <=( A199  and  A166 );
 a70395a <=( A201  and  (not A200) );
 a70396a <=( a70395a  and  a70392a );
 a70397a <=( a70396a  and  a70389a );
 a70400a <=( (not A233)  and  A203 );
 a70403a <=( (not A236)  and  (not A235) );
 a70404a <=( a70403a  and  a70400a );
 a70407a <=( A266  and  A265 );
 a70410a <=( A299  and  (not A298) );
 a70411a <=( a70410a  and  a70407a );
 a70412a <=( a70411a  and  a70404a );
 a70416a <=( A167  and  (not A168) );
 a70417a <=( (not A169)  and  a70416a );
 a70420a <=( A199  and  A166 );
 a70423a <=( A201  and  (not A200) );
 a70424a <=( a70423a  and  a70420a );
 a70425a <=( a70424a  and  a70417a );
 a70428a <=( (not A233)  and  A203 );
 a70431a <=( (not A236)  and  (not A235) );
 a70432a <=( a70431a  and  a70428a );
 a70435a <=( (not A267)  and  (not A266) );
 a70438a <=( A299  and  (not A298) );
 a70439a <=( a70438a  and  a70435a );
 a70440a <=( a70439a  and  a70432a );
 a70444a <=( A167  and  (not A168) );
 a70445a <=( (not A169)  and  a70444a );
 a70448a <=( A199  and  A166 );
 a70451a <=( A201  and  (not A200) );
 a70452a <=( a70451a  and  a70448a );
 a70453a <=( a70452a  and  a70445a );
 a70456a <=( (not A233)  and  A203 );
 a70459a <=( (not A236)  and  (not A235) );
 a70460a <=( a70459a  and  a70456a );
 a70463a <=( (not A266)  and  (not A265) );
 a70466a <=( A299  and  (not A298) );
 a70467a <=( a70466a  and  a70463a );
 a70468a <=( a70467a  and  a70460a );
 a70472a <=( A167  and  (not A168) );
 a70473a <=( (not A169)  and  a70472a );
 a70476a <=( A199  and  A166 );
 a70479a <=( A201  and  (not A200) );
 a70480a <=( a70479a  and  a70476a );
 a70481a <=( a70480a  and  a70473a );
 a70484a <=( (not A233)  and  A203 );
 a70487a <=( (not A266)  and  (not A234) );
 a70488a <=( a70487a  and  a70484a );
 a70491a <=( (not A269)  and  (not A268) );
 a70494a <=( A299  and  (not A298) );
 a70495a <=( a70494a  and  a70491a );
 a70496a <=( a70495a  and  a70488a );
 a70500a <=( A167  and  (not A168) );
 a70501a <=( (not A169)  and  a70500a );
 a70504a <=( A199  and  A166 );
 a70507a <=( A201  and  (not A200) );
 a70508a <=( a70507a  and  a70504a );
 a70509a <=( a70508a  and  a70501a );
 a70512a <=( A232  and  A203 );
 a70515a <=( A234  and  (not A233) );
 a70516a <=( a70515a  and  a70512a );
 a70519a <=( A298  and  A235 );
 a70522a <=( (not A302)  and  (not A301) );
 a70523a <=( a70522a  and  a70519a );
 a70524a <=( a70523a  and  a70516a );
 a70528a <=( A167  and  (not A168) );
 a70529a <=( (not A169)  and  a70528a );
 a70532a <=( A199  and  A166 );
 a70535a <=( A201  and  (not A200) );
 a70536a <=( a70535a  and  a70532a );
 a70537a <=( a70536a  and  a70529a );
 a70540a <=( A232  and  A203 );
 a70543a <=( A234  and  (not A233) );
 a70544a <=( a70543a  and  a70540a );
 a70547a <=( A298  and  A236 );
 a70550a <=( (not A302)  and  (not A301) );
 a70551a <=( a70550a  and  a70547a );
 a70552a <=( a70551a  and  a70544a );
 a70556a <=( A167  and  (not A168) );
 a70557a <=( (not A169)  and  a70556a );
 a70560a <=( A199  and  A166 );
 a70563a <=( A201  and  (not A200) );
 a70564a <=( a70563a  and  a70560a );
 a70565a <=( a70564a  and  a70557a );
 a70568a <=( (not A232)  and  A203 );
 a70571a <=( (not A266)  and  (not A233) );
 a70572a <=( a70571a  and  a70568a );
 a70575a <=( (not A269)  and  (not A268) );
 a70578a <=( A299  and  (not A298) );
 a70579a <=( a70578a  and  a70575a );
 a70580a <=( a70579a  and  a70572a );
 a70584a <=( A167  and  (not A169) );
 a70585a <=( A170  and  a70584a );
 a70588a <=( A199  and  (not A166) );
 a70591a <=( A232  and  A200 );
 a70592a <=( a70591a  and  a70588a );
 a70593a <=( a70592a  and  a70585a );
 a70596a <=( A265  and  A233 );
 a70599a <=( (not A269)  and  (not A268) );
 a70600a <=( a70599a  and  a70596a );
 a70603a <=( (not A299)  and  A298 );
 a70606a <=( A301  and  A300 );
 a70607a <=( a70606a  and  a70603a );
 a70608a <=( a70607a  and  a70600a );
 a70612a <=( A167  and  (not A169) );
 a70613a <=( A170  and  a70612a );
 a70616a <=( A199  and  (not A166) );
 a70619a <=( A232  and  A200 );
 a70620a <=( a70619a  and  a70616a );
 a70621a <=( a70620a  and  a70613a );
 a70624a <=( A265  and  A233 );
 a70627a <=( (not A269)  and  (not A268) );
 a70628a <=( a70627a  and  a70624a );
 a70631a <=( (not A299)  and  A298 );
 a70634a <=( A302  and  A300 );
 a70635a <=( a70634a  and  a70631a );
 a70636a <=( a70635a  and  a70628a );
 a70640a <=( A167  and  (not A169) );
 a70641a <=( A170  and  a70640a );
 a70644a <=( A199  and  (not A166) );
 a70647a <=( (not A233)  and  A200 );
 a70648a <=( a70647a  and  a70644a );
 a70649a <=( a70648a  and  a70641a );
 a70652a <=( (not A236)  and  (not A235) );
 a70655a <=( A266  and  A265 );
 a70656a <=( a70655a  and  a70652a );
 a70659a <=( (not A299)  and  A298 );
 a70662a <=( A301  and  A300 );
 a70663a <=( a70662a  and  a70659a );
 a70664a <=( a70663a  and  a70656a );
 a70668a <=( A167  and  (not A169) );
 a70669a <=( A170  and  a70668a );
 a70672a <=( A199  and  (not A166) );
 a70675a <=( (not A233)  and  A200 );
 a70676a <=( a70675a  and  a70672a );
 a70677a <=( a70676a  and  a70669a );
 a70680a <=( (not A236)  and  (not A235) );
 a70683a <=( A266  and  A265 );
 a70684a <=( a70683a  and  a70680a );
 a70687a <=( (not A299)  and  A298 );
 a70690a <=( A302  and  A300 );
 a70691a <=( a70690a  and  a70687a );
 a70692a <=( a70691a  and  a70684a );
 a70696a <=( A167  and  (not A169) );
 a70697a <=( A170  and  a70696a );
 a70700a <=( A199  and  (not A166) );
 a70703a <=( (not A233)  and  A200 );
 a70704a <=( a70703a  and  a70700a );
 a70705a <=( a70704a  and  a70697a );
 a70708a <=( (not A236)  and  (not A235) );
 a70711a <=( (not A267)  and  (not A266) );
 a70712a <=( a70711a  and  a70708a );
 a70715a <=( (not A299)  and  A298 );
 a70718a <=( A301  and  A300 );
 a70719a <=( a70718a  and  a70715a );
 a70720a <=( a70719a  and  a70712a );
 a70724a <=( A167  and  (not A169) );
 a70725a <=( A170  and  a70724a );
 a70728a <=( A199  and  (not A166) );
 a70731a <=( (not A233)  and  A200 );
 a70732a <=( a70731a  and  a70728a );
 a70733a <=( a70732a  and  a70725a );
 a70736a <=( (not A236)  and  (not A235) );
 a70739a <=( (not A267)  and  (not A266) );
 a70740a <=( a70739a  and  a70736a );
 a70743a <=( (not A299)  and  A298 );
 a70746a <=( A302  and  A300 );
 a70747a <=( a70746a  and  a70743a );
 a70748a <=( a70747a  and  a70740a );
 a70752a <=( A167  and  (not A169) );
 a70753a <=( A170  and  a70752a );
 a70756a <=( A199  and  (not A166) );
 a70759a <=( (not A233)  and  A200 );
 a70760a <=( a70759a  and  a70756a );
 a70761a <=( a70760a  and  a70753a );
 a70764a <=( (not A236)  and  (not A235) );
 a70767a <=( (not A266)  and  (not A265) );
 a70768a <=( a70767a  and  a70764a );
 a70771a <=( (not A299)  and  A298 );
 a70774a <=( A301  and  A300 );
 a70775a <=( a70774a  and  a70771a );
 a70776a <=( a70775a  and  a70768a );
 a70780a <=( A167  and  (not A169) );
 a70781a <=( A170  and  a70780a );
 a70784a <=( A199  and  (not A166) );
 a70787a <=( (not A233)  and  A200 );
 a70788a <=( a70787a  and  a70784a );
 a70789a <=( a70788a  and  a70781a );
 a70792a <=( (not A236)  and  (not A235) );
 a70795a <=( (not A266)  and  (not A265) );
 a70796a <=( a70795a  and  a70792a );
 a70799a <=( (not A299)  and  A298 );
 a70802a <=( A302  and  A300 );
 a70803a <=( a70802a  and  a70799a );
 a70804a <=( a70803a  and  a70796a );
 a70808a <=( A167  and  (not A169) );
 a70809a <=( A170  and  a70808a );
 a70812a <=( A199  and  (not A166) );
 a70815a <=( (not A233)  and  A200 );
 a70816a <=( a70815a  and  a70812a );
 a70817a <=( a70816a  and  a70809a );
 a70820a <=( (not A266)  and  (not A234) );
 a70823a <=( (not A269)  and  (not A268) );
 a70824a <=( a70823a  and  a70820a );
 a70827a <=( (not A299)  and  A298 );
 a70830a <=( A301  and  A300 );
 a70831a <=( a70830a  and  a70827a );
 a70832a <=( a70831a  and  a70824a );
 a70836a <=( A167  and  (not A169) );
 a70837a <=( A170  and  a70836a );
 a70840a <=( A199  and  (not A166) );
 a70843a <=( (not A233)  and  A200 );
 a70844a <=( a70843a  and  a70840a );
 a70845a <=( a70844a  and  a70837a );
 a70848a <=( (not A266)  and  (not A234) );
 a70851a <=( (not A269)  and  (not A268) );
 a70852a <=( a70851a  and  a70848a );
 a70855a <=( (not A299)  and  A298 );
 a70858a <=( A302  and  A300 );
 a70859a <=( a70858a  and  a70855a );
 a70860a <=( a70859a  and  a70852a );
 a70864a <=( A167  and  (not A169) );
 a70865a <=( A170  and  a70864a );
 a70868a <=( A199  and  (not A166) );
 a70871a <=( (not A232)  and  A200 );
 a70872a <=( a70871a  and  a70868a );
 a70873a <=( a70872a  and  a70865a );
 a70876a <=( (not A266)  and  (not A233) );
 a70879a <=( (not A269)  and  (not A268) );
 a70880a <=( a70879a  and  a70876a );
 a70883a <=( (not A299)  and  A298 );
 a70886a <=( A301  and  A300 );
 a70887a <=( a70886a  and  a70883a );
 a70888a <=( a70887a  and  a70880a );
 a70892a <=( A167  and  (not A169) );
 a70893a <=( A170  and  a70892a );
 a70896a <=( A199  and  (not A166) );
 a70899a <=( (not A232)  and  A200 );
 a70900a <=( a70899a  and  a70896a );
 a70901a <=( a70900a  and  a70893a );
 a70904a <=( (not A266)  and  (not A233) );
 a70907a <=( (not A269)  and  (not A268) );
 a70908a <=( a70907a  and  a70904a );
 a70911a <=( (not A299)  and  A298 );
 a70914a <=( A302  and  A300 );
 a70915a <=( a70914a  and  a70911a );
 a70916a <=( a70915a  and  a70908a );
 a70920a <=( A167  and  (not A169) );
 a70921a <=( A170  and  a70920a );
 a70924a <=( (not A200)  and  (not A166) );
 a70927a <=( (not A203)  and  (not A202) );
 a70928a <=( a70927a  and  a70924a );
 a70929a <=( a70928a  and  a70921a );
 a70932a <=( A233  and  A232 );
 a70935a <=( (not A267)  and  A265 );
 a70936a <=( a70935a  and  a70932a );
 a70939a <=( (not A299)  and  A298 );
 a70942a <=( A301  and  A300 );
 a70943a <=( a70942a  and  a70939a );
 a70944a <=( a70943a  and  a70936a );
 a70948a <=( A167  and  (not A169) );
 a70949a <=( A170  and  a70948a );
 a70952a <=( (not A200)  and  (not A166) );
 a70955a <=( (not A203)  and  (not A202) );
 a70956a <=( a70955a  and  a70952a );
 a70957a <=( a70956a  and  a70949a );
 a70960a <=( A233  and  A232 );
 a70963a <=( (not A267)  and  A265 );
 a70964a <=( a70963a  and  a70960a );
 a70967a <=( (not A299)  and  A298 );
 a70970a <=( A302  and  A300 );
 a70971a <=( a70970a  and  a70967a );
 a70972a <=( a70971a  and  a70964a );
 a70976a <=( A167  and  (not A169) );
 a70977a <=( A170  and  a70976a );
 a70980a <=( (not A200)  and  (not A166) );
 a70983a <=( (not A203)  and  (not A202) );
 a70984a <=( a70983a  and  a70980a );
 a70985a <=( a70984a  and  a70977a );
 a70988a <=( A233  and  A232 );
 a70991a <=( A266  and  A265 );
 a70992a <=( a70991a  and  a70988a );
 a70995a <=( (not A299)  and  A298 );
 a70998a <=( A301  and  A300 );
 a70999a <=( a70998a  and  a70995a );
 a71000a <=( a70999a  and  a70992a );
 a71004a <=( A167  and  (not A169) );
 a71005a <=( A170  and  a71004a );
 a71008a <=( (not A200)  and  (not A166) );
 a71011a <=( (not A203)  and  (not A202) );
 a71012a <=( a71011a  and  a71008a );
 a71013a <=( a71012a  and  a71005a );
 a71016a <=( A233  and  A232 );
 a71019a <=( A266  and  A265 );
 a71020a <=( a71019a  and  a71016a );
 a71023a <=( (not A299)  and  A298 );
 a71026a <=( A302  and  A300 );
 a71027a <=( a71026a  and  a71023a );
 a71028a <=( a71027a  and  a71020a );
 a71032a <=( A167  and  (not A169) );
 a71033a <=( A170  and  a71032a );
 a71036a <=( (not A200)  and  (not A166) );
 a71039a <=( (not A203)  and  (not A202) );
 a71040a <=( a71039a  and  a71036a );
 a71041a <=( a71040a  and  a71033a );
 a71044a <=( A233  and  A232 );
 a71047a <=( (not A266)  and  (not A265) );
 a71048a <=( a71047a  and  a71044a );
 a71051a <=( (not A299)  and  A298 );
 a71054a <=( A301  and  A300 );
 a71055a <=( a71054a  and  a71051a );
 a71056a <=( a71055a  and  a71048a );
 a71060a <=( A167  and  (not A169) );
 a71061a <=( A170  and  a71060a );
 a71064a <=( (not A200)  and  (not A166) );
 a71067a <=( (not A203)  and  (not A202) );
 a71068a <=( a71067a  and  a71064a );
 a71069a <=( a71068a  and  a71061a );
 a71072a <=( A233  and  A232 );
 a71075a <=( (not A266)  and  (not A265) );
 a71076a <=( a71075a  and  a71072a );
 a71079a <=( (not A299)  and  A298 );
 a71082a <=( A302  and  A300 );
 a71083a <=( a71082a  and  a71079a );
 a71084a <=( a71083a  and  a71076a );
 a71088a <=( A167  and  (not A169) );
 a71089a <=( A170  and  a71088a );
 a71092a <=( (not A200)  and  (not A166) );
 a71095a <=( (not A203)  and  (not A202) );
 a71096a <=( a71095a  and  a71092a );
 a71097a <=( a71096a  and  a71089a );
 a71100a <=( (not A235)  and  (not A233) );
 a71103a <=( (not A266)  and  (not A236) );
 a71104a <=( a71103a  and  a71100a );
 a71107a <=( (not A269)  and  (not A268) );
 a71110a <=( A299  and  (not A298) );
 a71111a <=( a71110a  and  a71107a );
 a71112a <=( a71111a  and  a71104a );
 a71116a <=( A167  and  (not A169) );
 a71117a <=( A170  and  a71116a );
 a71120a <=( (not A200)  and  (not A166) );
 a71123a <=( (not A203)  and  (not A202) );
 a71124a <=( a71123a  and  a71120a );
 a71125a <=( a71124a  and  a71117a );
 a71128a <=( (not A234)  and  (not A233) );
 a71131a <=( A266  and  A265 );
 a71132a <=( a71131a  and  a71128a );
 a71135a <=( (not A299)  and  A298 );
 a71138a <=( A301  and  A300 );
 a71139a <=( a71138a  and  a71135a );
 a71140a <=( a71139a  and  a71132a );
 a71144a <=( A167  and  (not A169) );
 a71145a <=( A170  and  a71144a );
 a71148a <=( (not A200)  and  (not A166) );
 a71151a <=( (not A203)  and  (not A202) );
 a71152a <=( a71151a  and  a71148a );
 a71153a <=( a71152a  and  a71145a );
 a71156a <=( (not A234)  and  (not A233) );
 a71159a <=( A266  and  A265 );
 a71160a <=( a71159a  and  a71156a );
 a71163a <=( (not A299)  and  A298 );
 a71166a <=( A302  and  A300 );
 a71167a <=( a71166a  and  a71163a );
 a71168a <=( a71167a  and  a71160a );
 a71172a <=( A167  and  (not A169) );
 a71173a <=( A170  and  a71172a );
 a71176a <=( (not A200)  and  (not A166) );
 a71179a <=( (not A203)  and  (not A202) );
 a71180a <=( a71179a  and  a71176a );
 a71181a <=( a71180a  and  a71173a );
 a71184a <=( (not A234)  and  (not A233) );
 a71187a <=( (not A267)  and  (not A266) );
 a71188a <=( a71187a  and  a71184a );
 a71191a <=( (not A299)  and  A298 );
 a71194a <=( A301  and  A300 );
 a71195a <=( a71194a  and  a71191a );
 a71196a <=( a71195a  and  a71188a );
 a71200a <=( A167  and  (not A169) );
 a71201a <=( A170  and  a71200a );
 a71204a <=( (not A200)  and  (not A166) );
 a71207a <=( (not A203)  and  (not A202) );
 a71208a <=( a71207a  and  a71204a );
 a71209a <=( a71208a  and  a71201a );
 a71212a <=( (not A234)  and  (not A233) );
 a71215a <=( (not A267)  and  (not A266) );
 a71216a <=( a71215a  and  a71212a );
 a71219a <=( (not A299)  and  A298 );
 a71222a <=( A302  and  A300 );
 a71223a <=( a71222a  and  a71219a );
 a71224a <=( a71223a  and  a71216a );
 a71228a <=( A167  and  (not A169) );
 a71229a <=( A170  and  a71228a );
 a71232a <=( (not A200)  and  (not A166) );
 a71235a <=( (not A203)  and  (not A202) );
 a71236a <=( a71235a  and  a71232a );
 a71237a <=( a71236a  and  a71229a );
 a71240a <=( (not A234)  and  (not A233) );
 a71243a <=( (not A266)  and  (not A265) );
 a71244a <=( a71243a  and  a71240a );
 a71247a <=( (not A299)  and  A298 );
 a71250a <=( A301  and  A300 );
 a71251a <=( a71250a  and  a71247a );
 a71252a <=( a71251a  and  a71244a );
 a71256a <=( A167  and  (not A169) );
 a71257a <=( A170  and  a71256a );
 a71260a <=( (not A200)  and  (not A166) );
 a71263a <=( (not A203)  and  (not A202) );
 a71264a <=( a71263a  and  a71260a );
 a71265a <=( a71264a  and  a71257a );
 a71268a <=( (not A234)  and  (not A233) );
 a71271a <=( (not A266)  and  (not A265) );
 a71272a <=( a71271a  and  a71268a );
 a71275a <=( (not A299)  and  A298 );
 a71278a <=( A302  and  A300 );
 a71279a <=( a71278a  and  a71275a );
 a71280a <=( a71279a  and  a71272a );
 a71284a <=( A167  and  (not A169) );
 a71285a <=( A170  and  a71284a );
 a71288a <=( (not A200)  and  (not A166) );
 a71291a <=( (not A203)  and  (not A202) );
 a71292a <=( a71291a  and  a71288a );
 a71293a <=( a71292a  and  a71285a );
 a71296a <=( (not A233)  and  A232 );
 a71299a <=( A235  and  A234 );
 a71300a <=( a71299a  and  a71296a );
 a71303a <=( (not A266)  and  A265 );
 a71306a <=( A268  and  A267 );
 a71307a <=( a71306a  and  a71303a );
 a71308a <=( a71307a  and  a71300a );
 a71312a <=( A167  and  (not A169) );
 a71313a <=( A170  and  a71312a );
 a71316a <=( (not A200)  and  (not A166) );
 a71319a <=( (not A203)  and  (not A202) );
 a71320a <=( a71319a  and  a71316a );
 a71321a <=( a71320a  and  a71313a );
 a71324a <=( (not A233)  and  A232 );
 a71327a <=( A235  and  A234 );
 a71328a <=( a71327a  and  a71324a );
 a71331a <=( (not A266)  and  A265 );
 a71334a <=( A269  and  A267 );
 a71335a <=( a71334a  and  a71331a );
 a71336a <=( a71335a  and  a71328a );
 a71340a <=( A167  and  (not A169) );
 a71341a <=( A170  and  a71340a );
 a71344a <=( (not A200)  and  (not A166) );
 a71347a <=( (not A203)  and  (not A202) );
 a71348a <=( a71347a  and  a71344a );
 a71349a <=( a71348a  and  a71341a );
 a71352a <=( (not A233)  and  A232 );
 a71355a <=( A236  and  A234 );
 a71356a <=( a71355a  and  a71352a );
 a71359a <=( (not A266)  and  A265 );
 a71362a <=( A268  and  A267 );
 a71363a <=( a71362a  and  a71359a );
 a71364a <=( a71363a  and  a71356a );
 a71368a <=( A167  and  (not A169) );
 a71369a <=( A170  and  a71368a );
 a71372a <=( (not A200)  and  (not A166) );
 a71375a <=( (not A203)  and  (not A202) );
 a71376a <=( a71375a  and  a71372a );
 a71377a <=( a71376a  and  a71369a );
 a71380a <=( (not A233)  and  A232 );
 a71383a <=( A236  and  A234 );
 a71384a <=( a71383a  and  a71380a );
 a71387a <=( (not A266)  and  A265 );
 a71390a <=( A269  and  A267 );
 a71391a <=( a71390a  and  a71387a );
 a71392a <=( a71391a  and  a71384a );
 a71396a <=( A167  and  (not A169) );
 a71397a <=( A170  and  a71396a );
 a71400a <=( (not A200)  and  (not A166) );
 a71403a <=( (not A203)  and  (not A202) );
 a71404a <=( a71403a  and  a71400a );
 a71405a <=( a71404a  and  a71397a );
 a71408a <=( (not A233)  and  (not A232) );
 a71411a <=( A266  and  A265 );
 a71412a <=( a71411a  and  a71408a );
 a71415a <=( (not A299)  and  A298 );
 a71418a <=( A301  and  A300 );
 a71419a <=( a71418a  and  a71415a );
 a71420a <=( a71419a  and  a71412a );
 a71424a <=( A167  and  (not A169) );
 a71425a <=( A170  and  a71424a );
 a71428a <=( (not A200)  and  (not A166) );
 a71431a <=( (not A203)  and  (not A202) );
 a71432a <=( a71431a  and  a71428a );
 a71433a <=( a71432a  and  a71425a );
 a71436a <=( (not A233)  and  (not A232) );
 a71439a <=( A266  and  A265 );
 a71440a <=( a71439a  and  a71436a );
 a71443a <=( (not A299)  and  A298 );
 a71446a <=( A302  and  A300 );
 a71447a <=( a71446a  and  a71443a );
 a71448a <=( a71447a  and  a71440a );
 a71452a <=( A167  and  (not A169) );
 a71453a <=( A170  and  a71452a );
 a71456a <=( (not A200)  and  (not A166) );
 a71459a <=( (not A203)  and  (not A202) );
 a71460a <=( a71459a  and  a71456a );
 a71461a <=( a71460a  and  a71453a );
 a71464a <=( (not A233)  and  (not A232) );
 a71467a <=( (not A267)  and  (not A266) );
 a71468a <=( a71467a  and  a71464a );
 a71471a <=( (not A299)  and  A298 );
 a71474a <=( A301  and  A300 );
 a71475a <=( a71474a  and  a71471a );
 a71476a <=( a71475a  and  a71468a );
 a71480a <=( A167  and  (not A169) );
 a71481a <=( A170  and  a71480a );
 a71484a <=( (not A200)  and  (not A166) );
 a71487a <=( (not A203)  and  (not A202) );
 a71488a <=( a71487a  and  a71484a );
 a71489a <=( a71488a  and  a71481a );
 a71492a <=( (not A233)  and  (not A232) );
 a71495a <=( (not A267)  and  (not A266) );
 a71496a <=( a71495a  and  a71492a );
 a71499a <=( (not A299)  and  A298 );
 a71502a <=( A302  and  A300 );
 a71503a <=( a71502a  and  a71499a );
 a71504a <=( a71503a  and  a71496a );
 a71508a <=( A167  and  (not A169) );
 a71509a <=( A170  and  a71508a );
 a71512a <=( (not A200)  and  (not A166) );
 a71515a <=( (not A203)  and  (not A202) );
 a71516a <=( a71515a  and  a71512a );
 a71517a <=( a71516a  and  a71509a );
 a71520a <=( (not A233)  and  (not A232) );
 a71523a <=( (not A266)  and  (not A265) );
 a71524a <=( a71523a  and  a71520a );
 a71527a <=( (not A299)  and  A298 );
 a71530a <=( A301  and  A300 );
 a71531a <=( a71530a  and  a71527a );
 a71532a <=( a71531a  and  a71524a );
 a71536a <=( A167  and  (not A169) );
 a71537a <=( A170  and  a71536a );
 a71540a <=( (not A200)  and  (not A166) );
 a71543a <=( (not A203)  and  (not A202) );
 a71544a <=( a71543a  and  a71540a );
 a71545a <=( a71544a  and  a71537a );
 a71548a <=( (not A233)  and  (not A232) );
 a71551a <=( (not A266)  and  (not A265) );
 a71552a <=( a71551a  and  a71548a );
 a71555a <=( (not A299)  and  A298 );
 a71558a <=( A302  and  A300 );
 a71559a <=( a71558a  and  a71555a );
 a71560a <=( a71559a  and  a71552a );
 a71564a <=( A167  and  (not A169) );
 a71565a <=( A170  and  a71564a );
 a71568a <=( (not A200)  and  (not A166) );
 a71571a <=( A232  and  (not A201) );
 a71572a <=( a71571a  and  a71568a );
 a71573a <=( a71572a  and  a71565a );
 a71576a <=( A265  and  A233 );
 a71579a <=( (not A269)  and  (not A268) );
 a71580a <=( a71579a  and  a71576a );
 a71583a <=( (not A299)  and  A298 );
 a71586a <=( A301  and  A300 );
 a71587a <=( a71586a  and  a71583a );
 a71588a <=( a71587a  and  a71580a );
 a71592a <=( A167  and  (not A169) );
 a71593a <=( A170  and  a71592a );
 a71596a <=( (not A200)  and  (not A166) );
 a71599a <=( A232  and  (not A201) );
 a71600a <=( a71599a  and  a71596a );
 a71601a <=( a71600a  and  a71593a );
 a71604a <=( A265  and  A233 );
 a71607a <=( (not A269)  and  (not A268) );
 a71608a <=( a71607a  and  a71604a );
 a71611a <=( (not A299)  and  A298 );
 a71614a <=( A302  and  A300 );
 a71615a <=( a71614a  and  a71611a );
 a71616a <=( a71615a  and  a71608a );
 a71620a <=( A167  and  (not A169) );
 a71621a <=( A170  and  a71620a );
 a71624a <=( (not A200)  and  (not A166) );
 a71627a <=( (not A233)  and  (not A201) );
 a71628a <=( a71627a  and  a71624a );
 a71629a <=( a71628a  and  a71621a );
 a71632a <=( (not A236)  and  (not A235) );
 a71635a <=( A266  and  A265 );
 a71636a <=( a71635a  and  a71632a );
 a71639a <=( (not A299)  and  A298 );
 a71642a <=( A301  and  A300 );
 a71643a <=( a71642a  and  a71639a );
 a71644a <=( a71643a  and  a71636a );
 a71648a <=( A167  and  (not A169) );
 a71649a <=( A170  and  a71648a );
 a71652a <=( (not A200)  and  (not A166) );
 a71655a <=( (not A233)  and  (not A201) );
 a71656a <=( a71655a  and  a71652a );
 a71657a <=( a71656a  and  a71649a );
 a71660a <=( (not A236)  and  (not A235) );
 a71663a <=( A266  and  A265 );
 a71664a <=( a71663a  and  a71660a );
 a71667a <=( (not A299)  and  A298 );
 a71670a <=( A302  and  A300 );
 a71671a <=( a71670a  and  a71667a );
 a71672a <=( a71671a  and  a71664a );
 a71676a <=( A167  and  (not A169) );
 a71677a <=( A170  and  a71676a );
 a71680a <=( (not A200)  and  (not A166) );
 a71683a <=( (not A233)  and  (not A201) );
 a71684a <=( a71683a  and  a71680a );
 a71685a <=( a71684a  and  a71677a );
 a71688a <=( (not A236)  and  (not A235) );
 a71691a <=( (not A267)  and  (not A266) );
 a71692a <=( a71691a  and  a71688a );
 a71695a <=( (not A299)  and  A298 );
 a71698a <=( A301  and  A300 );
 a71699a <=( a71698a  and  a71695a );
 a71700a <=( a71699a  and  a71692a );
 a71704a <=( A167  and  (not A169) );
 a71705a <=( A170  and  a71704a );
 a71708a <=( (not A200)  and  (not A166) );
 a71711a <=( (not A233)  and  (not A201) );
 a71712a <=( a71711a  and  a71708a );
 a71713a <=( a71712a  and  a71705a );
 a71716a <=( (not A236)  and  (not A235) );
 a71719a <=( (not A267)  and  (not A266) );
 a71720a <=( a71719a  and  a71716a );
 a71723a <=( (not A299)  and  A298 );
 a71726a <=( A302  and  A300 );
 a71727a <=( a71726a  and  a71723a );
 a71728a <=( a71727a  and  a71720a );
 a71732a <=( A167  and  (not A169) );
 a71733a <=( A170  and  a71732a );
 a71736a <=( (not A200)  and  (not A166) );
 a71739a <=( (not A233)  and  (not A201) );
 a71740a <=( a71739a  and  a71736a );
 a71741a <=( a71740a  and  a71733a );
 a71744a <=( (not A236)  and  (not A235) );
 a71747a <=( (not A266)  and  (not A265) );
 a71748a <=( a71747a  and  a71744a );
 a71751a <=( (not A299)  and  A298 );
 a71754a <=( A301  and  A300 );
 a71755a <=( a71754a  and  a71751a );
 a71756a <=( a71755a  and  a71748a );
 a71760a <=( A167  and  (not A169) );
 a71761a <=( A170  and  a71760a );
 a71764a <=( (not A200)  and  (not A166) );
 a71767a <=( (not A233)  and  (not A201) );
 a71768a <=( a71767a  and  a71764a );
 a71769a <=( a71768a  and  a71761a );
 a71772a <=( (not A236)  and  (not A235) );
 a71775a <=( (not A266)  and  (not A265) );
 a71776a <=( a71775a  and  a71772a );
 a71779a <=( (not A299)  and  A298 );
 a71782a <=( A302  and  A300 );
 a71783a <=( a71782a  and  a71779a );
 a71784a <=( a71783a  and  a71776a );
 a71788a <=( A167  and  (not A169) );
 a71789a <=( A170  and  a71788a );
 a71792a <=( (not A200)  and  (not A166) );
 a71795a <=( (not A233)  and  (not A201) );
 a71796a <=( a71795a  and  a71792a );
 a71797a <=( a71796a  and  a71789a );
 a71800a <=( (not A266)  and  (not A234) );
 a71803a <=( (not A269)  and  (not A268) );
 a71804a <=( a71803a  and  a71800a );
 a71807a <=( (not A299)  and  A298 );
 a71810a <=( A301  and  A300 );
 a71811a <=( a71810a  and  a71807a );
 a71812a <=( a71811a  and  a71804a );
 a71816a <=( A167  and  (not A169) );
 a71817a <=( A170  and  a71816a );
 a71820a <=( (not A200)  and  (not A166) );
 a71823a <=( (not A233)  and  (not A201) );
 a71824a <=( a71823a  and  a71820a );
 a71825a <=( a71824a  and  a71817a );
 a71828a <=( (not A266)  and  (not A234) );
 a71831a <=( (not A269)  and  (not A268) );
 a71832a <=( a71831a  and  a71828a );
 a71835a <=( (not A299)  and  A298 );
 a71838a <=( A302  and  A300 );
 a71839a <=( a71838a  and  a71835a );
 a71840a <=( a71839a  and  a71832a );
 a71844a <=( A167  and  (not A169) );
 a71845a <=( A170  and  a71844a );
 a71848a <=( (not A200)  and  (not A166) );
 a71851a <=( (not A232)  and  (not A201) );
 a71852a <=( a71851a  and  a71848a );
 a71853a <=( a71852a  and  a71845a );
 a71856a <=( (not A266)  and  (not A233) );
 a71859a <=( (not A269)  and  (not A268) );
 a71860a <=( a71859a  and  a71856a );
 a71863a <=( (not A299)  and  A298 );
 a71866a <=( A301  and  A300 );
 a71867a <=( a71866a  and  a71863a );
 a71868a <=( a71867a  and  a71860a );
 a71872a <=( A167  and  (not A169) );
 a71873a <=( A170  and  a71872a );
 a71876a <=( (not A200)  and  (not A166) );
 a71879a <=( (not A232)  and  (not A201) );
 a71880a <=( a71879a  and  a71876a );
 a71881a <=( a71880a  and  a71873a );
 a71884a <=( (not A266)  and  (not A233) );
 a71887a <=( (not A269)  and  (not A268) );
 a71888a <=( a71887a  and  a71884a );
 a71891a <=( (not A299)  and  A298 );
 a71894a <=( A302  and  A300 );
 a71895a <=( a71894a  and  a71891a );
 a71896a <=( a71895a  and  a71888a );
 a71900a <=( A167  and  (not A169) );
 a71901a <=( A170  and  a71900a );
 a71904a <=( (not A199)  and  (not A166) );
 a71907a <=( A232  and  (not A200) );
 a71908a <=( a71907a  and  a71904a );
 a71909a <=( a71908a  and  a71901a );
 a71912a <=( A265  and  A233 );
 a71915a <=( (not A269)  and  (not A268) );
 a71916a <=( a71915a  and  a71912a );
 a71919a <=( (not A299)  and  A298 );
 a71922a <=( A301  and  A300 );
 a71923a <=( a71922a  and  a71919a );
 a71924a <=( a71923a  and  a71916a );
 a71928a <=( A167  and  (not A169) );
 a71929a <=( A170  and  a71928a );
 a71932a <=( (not A199)  and  (not A166) );
 a71935a <=( A232  and  (not A200) );
 a71936a <=( a71935a  and  a71932a );
 a71937a <=( a71936a  and  a71929a );
 a71940a <=( A265  and  A233 );
 a71943a <=( (not A269)  and  (not A268) );
 a71944a <=( a71943a  and  a71940a );
 a71947a <=( (not A299)  and  A298 );
 a71950a <=( A302  and  A300 );
 a71951a <=( a71950a  and  a71947a );
 a71952a <=( a71951a  and  a71944a );
 a71956a <=( A167  and  (not A169) );
 a71957a <=( A170  and  a71956a );
 a71960a <=( (not A199)  and  (not A166) );
 a71963a <=( (not A233)  and  (not A200) );
 a71964a <=( a71963a  and  a71960a );
 a71965a <=( a71964a  and  a71957a );
 a71968a <=( (not A236)  and  (not A235) );
 a71971a <=( A266  and  A265 );
 a71972a <=( a71971a  and  a71968a );
 a71975a <=( (not A299)  and  A298 );
 a71978a <=( A301  and  A300 );
 a71979a <=( a71978a  and  a71975a );
 a71980a <=( a71979a  and  a71972a );
 a71984a <=( A167  and  (not A169) );
 a71985a <=( A170  and  a71984a );
 a71988a <=( (not A199)  and  (not A166) );
 a71991a <=( (not A233)  and  (not A200) );
 a71992a <=( a71991a  and  a71988a );
 a71993a <=( a71992a  and  a71985a );
 a71996a <=( (not A236)  and  (not A235) );
 a71999a <=( A266  and  A265 );
 a72000a <=( a71999a  and  a71996a );
 a72003a <=( (not A299)  and  A298 );
 a72006a <=( A302  and  A300 );
 a72007a <=( a72006a  and  a72003a );
 a72008a <=( a72007a  and  a72000a );
 a72012a <=( A167  and  (not A169) );
 a72013a <=( A170  and  a72012a );
 a72016a <=( (not A199)  and  (not A166) );
 a72019a <=( (not A233)  and  (not A200) );
 a72020a <=( a72019a  and  a72016a );
 a72021a <=( a72020a  and  a72013a );
 a72024a <=( (not A236)  and  (not A235) );
 a72027a <=( (not A267)  and  (not A266) );
 a72028a <=( a72027a  and  a72024a );
 a72031a <=( (not A299)  and  A298 );
 a72034a <=( A301  and  A300 );
 a72035a <=( a72034a  and  a72031a );
 a72036a <=( a72035a  and  a72028a );
 a72040a <=( A167  and  (not A169) );
 a72041a <=( A170  and  a72040a );
 a72044a <=( (not A199)  and  (not A166) );
 a72047a <=( (not A233)  and  (not A200) );
 a72048a <=( a72047a  and  a72044a );
 a72049a <=( a72048a  and  a72041a );
 a72052a <=( (not A236)  and  (not A235) );
 a72055a <=( (not A267)  and  (not A266) );
 a72056a <=( a72055a  and  a72052a );
 a72059a <=( (not A299)  and  A298 );
 a72062a <=( A302  and  A300 );
 a72063a <=( a72062a  and  a72059a );
 a72064a <=( a72063a  and  a72056a );
 a72068a <=( A167  and  (not A169) );
 a72069a <=( A170  and  a72068a );
 a72072a <=( (not A199)  and  (not A166) );
 a72075a <=( (not A233)  and  (not A200) );
 a72076a <=( a72075a  and  a72072a );
 a72077a <=( a72076a  and  a72069a );
 a72080a <=( (not A236)  and  (not A235) );
 a72083a <=( (not A266)  and  (not A265) );
 a72084a <=( a72083a  and  a72080a );
 a72087a <=( (not A299)  and  A298 );
 a72090a <=( A301  and  A300 );
 a72091a <=( a72090a  and  a72087a );
 a72092a <=( a72091a  and  a72084a );
 a72096a <=( A167  and  (not A169) );
 a72097a <=( A170  and  a72096a );
 a72100a <=( (not A199)  and  (not A166) );
 a72103a <=( (not A233)  and  (not A200) );
 a72104a <=( a72103a  and  a72100a );
 a72105a <=( a72104a  and  a72097a );
 a72108a <=( (not A236)  and  (not A235) );
 a72111a <=( (not A266)  and  (not A265) );
 a72112a <=( a72111a  and  a72108a );
 a72115a <=( (not A299)  and  A298 );
 a72118a <=( A302  and  A300 );
 a72119a <=( a72118a  and  a72115a );
 a72120a <=( a72119a  and  a72112a );
 a72124a <=( A167  and  (not A169) );
 a72125a <=( A170  and  a72124a );
 a72128a <=( (not A199)  and  (not A166) );
 a72131a <=( (not A233)  and  (not A200) );
 a72132a <=( a72131a  and  a72128a );
 a72133a <=( a72132a  and  a72125a );
 a72136a <=( (not A266)  and  (not A234) );
 a72139a <=( (not A269)  and  (not A268) );
 a72140a <=( a72139a  and  a72136a );
 a72143a <=( (not A299)  and  A298 );
 a72146a <=( A301  and  A300 );
 a72147a <=( a72146a  and  a72143a );
 a72148a <=( a72147a  and  a72140a );
 a72152a <=( A167  and  (not A169) );
 a72153a <=( A170  and  a72152a );
 a72156a <=( (not A199)  and  (not A166) );
 a72159a <=( (not A233)  and  (not A200) );
 a72160a <=( a72159a  and  a72156a );
 a72161a <=( a72160a  and  a72153a );
 a72164a <=( (not A266)  and  (not A234) );
 a72167a <=( (not A269)  and  (not A268) );
 a72168a <=( a72167a  and  a72164a );
 a72171a <=( (not A299)  and  A298 );
 a72174a <=( A302  and  A300 );
 a72175a <=( a72174a  and  a72171a );
 a72176a <=( a72175a  and  a72168a );
 a72180a <=( A167  and  (not A169) );
 a72181a <=( A170  and  a72180a );
 a72184a <=( (not A199)  and  (not A166) );
 a72187a <=( (not A232)  and  (not A200) );
 a72188a <=( a72187a  and  a72184a );
 a72189a <=( a72188a  and  a72181a );
 a72192a <=( (not A266)  and  (not A233) );
 a72195a <=( (not A269)  and  (not A268) );
 a72196a <=( a72195a  and  a72192a );
 a72199a <=( (not A299)  and  A298 );
 a72202a <=( A301  and  A300 );
 a72203a <=( a72202a  and  a72199a );
 a72204a <=( a72203a  and  a72196a );
 a72208a <=( A167  and  (not A169) );
 a72209a <=( A170  and  a72208a );
 a72212a <=( (not A199)  and  (not A166) );
 a72215a <=( (not A232)  and  (not A200) );
 a72216a <=( a72215a  and  a72212a );
 a72217a <=( a72216a  and  a72209a );
 a72220a <=( (not A266)  and  (not A233) );
 a72223a <=( (not A269)  and  (not A268) );
 a72224a <=( a72223a  and  a72220a );
 a72227a <=( (not A299)  and  A298 );
 a72230a <=( A302  and  A300 );
 a72231a <=( a72230a  and  a72227a );
 a72232a <=( a72231a  and  a72224a );
 a72236a <=( (not A167)  and  (not A169) );
 a72237a <=( A170  and  a72236a );
 a72240a <=( A199  and  A166 );
 a72243a <=( A232  and  A200 );
 a72244a <=( a72243a  and  a72240a );
 a72245a <=( a72244a  and  a72237a );
 a72248a <=( A265  and  A233 );
 a72251a <=( (not A269)  and  (not A268) );
 a72252a <=( a72251a  and  a72248a );
 a72255a <=( (not A299)  and  A298 );
 a72258a <=( A301  and  A300 );
 a72259a <=( a72258a  and  a72255a );
 a72260a <=( a72259a  and  a72252a );
 a72264a <=( (not A167)  and  (not A169) );
 a72265a <=( A170  and  a72264a );
 a72268a <=( A199  and  A166 );
 a72271a <=( A232  and  A200 );
 a72272a <=( a72271a  and  a72268a );
 a72273a <=( a72272a  and  a72265a );
 a72276a <=( A265  and  A233 );
 a72279a <=( (not A269)  and  (not A268) );
 a72280a <=( a72279a  and  a72276a );
 a72283a <=( (not A299)  and  A298 );
 a72286a <=( A302  and  A300 );
 a72287a <=( a72286a  and  a72283a );
 a72288a <=( a72287a  and  a72280a );
 a72292a <=( (not A167)  and  (not A169) );
 a72293a <=( A170  and  a72292a );
 a72296a <=( A199  and  A166 );
 a72299a <=( (not A233)  and  A200 );
 a72300a <=( a72299a  and  a72296a );
 a72301a <=( a72300a  and  a72293a );
 a72304a <=( (not A236)  and  (not A235) );
 a72307a <=( A266  and  A265 );
 a72308a <=( a72307a  and  a72304a );
 a72311a <=( (not A299)  and  A298 );
 a72314a <=( A301  and  A300 );
 a72315a <=( a72314a  and  a72311a );
 a72316a <=( a72315a  and  a72308a );
 a72320a <=( (not A167)  and  (not A169) );
 a72321a <=( A170  and  a72320a );
 a72324a <=( A199  and  A166 );
 a72327a <=( (not A233)  and  A200 );
 a72328a <=( a72327a  and  a72324a );
 a72329a <=( a72328a  and  a72321a );
 a72332a <=( (not A236)  and  (not A235) );
 a72335a <=( A266  and  A265 );
 a72336a <=( a72335a  and  a72332a );
 a72339a <=( (not A299)  and  A298 );
 a72342a <=( A302  and  A300 );
 a72343a <=( a72342a  and  a72339a );
 a72344a <=( a72343a  and  a72336a );
 a72348a <=( (not A167)  and  (not A169) );
 a72349a <=( A170  and  a72348a );
 a72352a <=( A199  and  A166 );
 a72355a <=( (not A233)  and  A200 );
 a72356a <=( a72355a  and  a72352a );
 a72357a <=( a72356a  and  a72349a );
 a72360a <=( (not A236)  and  (not A235) );
 a72363a <=( (not A267)  and  (not A266) );
 a72364a <=( a72363a  and  a72360a );
 a72367a <=( (not A299)  and  A298 );
 a72370a <=( A301  and  A300 );
 a72371a <=( a72370a  and  a72367a );
 a72372a <=( a72371a  and  a72364a );
 a72376a <=( (not A167)  and  (not A169) );
 a72377a <=( A170  and  a72376a );
 a72380a <=( A199  and  A166 );
 a72383a <=( (not A233)  and  A200 );
 a72384a <=( a72383a  and  a72380a );
 a72385a <=( a72384a  and  a72377a );
 a72388a <=( (not A236)  and  (not A235) );
 a72391a <=( (not A267)  and  (not A266) );
 a72392a <=( a72391a  and  a72388a );
 a72395a <=( (not A299)  and  A298 );
 a72398a <=( A302  and  A300 );
 a72399a <=( a72398a  and  a72395a );
 a72400a <=( a72399a  and  a72392a );
 a72404a <=( (not A167)  and  (not A169) );
 a72405a <=( A170  and  a72404a );
 a72408a <=( A199  and  A166 );
 a72411a <=( (not A233)  and  A200 );
 a72412a <=( a72411a  and  a72408a );
 a72413a <=( a72412a  and  a72405a );
 a72416a <=( (not A236)  and  (not A235) );
 a72419a <=( (not A266)  and  (not A265) );
 a72420a <=( a72419a  and  a72416a );
 a72423a <=( (not A299)  and  A298 );
 a72426a <=( A301  and  A300 );
 a72427a <=( a72426a  and  a72423a );
 a72428a <=( a72427a  and  a72420a );
 a72432a <=( (not A167)  and  (not A169) );
 a72433a <=( A170  and  a72432a );
 a72436a <=( A199  and  A166 );
 a72439a <=( (not A233)  and  A200 );
 a72440a <=( a72439a  and  a72436a );
 a72441a <=( a72440a  and  a72433a );
 a72444a <=( (not A236)  and  (not A235) );
 a72447a <=( (not A266)  and  (not A265) );
 a72448a <=( a72447a  and  a72444a );
 a72451a <=( (not A299)  and  A298 );
 a72454a <=( A302  and  A300 );
 a72455a <=( a72454a  and  a72451a );
 a72456a <=( a72455a  and  a72448a );
 a72460a <=( (not A167)  and  (not A169) );
 a72461a <=( A170  and  a72460a );
 a72464a <=( A199  and  A166 );
 a72467a <=( (not A233)  and  A200 );
 a72468a <=( a72467a  and  a72464a );
 a72469a <=( a72468a  and  a72461a );
 a72472a <=( (not A266)  and  (not A234) );
 a72475a <=( (not A269)  and  (not A268) );
 a72476a <=( a72475a  and  a72472a );
 a72479a <=( (not A299)  and  A298 );
 a72482a <=( A301  and  A300 );
 a72483a <=( a72482a  and  a72479a );
 a72484a <=( a72483a  and  a72476a );
 a72488a <=( (not A167)  and  (not A169) );
 a72489a <=( A170  and  a72488a );
 a72492a <=( A199  and  A166 );
 a72495a <=( (not A233)  and  A200 );
 a72496a <=( a72495a  and  a72492a );
 a72497a <=( a72496a  and  a72489a );
 a72500a <=( (not A266)  and  (not A234) );
 a72503a <=( (not A269)  and  (not A268) );
 a72504a <=( a72503a  and  a72500a );
 a72507a <=( (not A299)  and  A298 );
 a72510a <=( A302  and  A300 );
 a72511a <=( a72510a  and  a72507a );
 a72512a <=( a72511a  and  a72504a );
 a72516a <=( (not A167)  and  (not A169) );
 a72517a <=( A170  and  a72516a );
 a72520a <=( A199  and  A166 );
 a72523a <=( (not A232)  and  A200 );
 a72524a <=( a72523a  and  a72520a );
 a72525a <=( a72524a  and  a72517a );
 a72528a <=( (not A266)  and  (not A233) );
 a72531a <=( (not A269)  and  (not A268) );
 a72532a <=( a72531a  and  a72528a );
 a72535a <=( (not A299)  and  A298 );
 a72538a <=( A301  and  A300 );
 a72539a <=( a72538a  and  a72535a );
 a72540a <=( a72539a  and  a72532a );
 a72544a <=( (not A167)  and  (not A169) );
 a72545a <=( A170  and  a72544a );
 a72548a <=( A199  and  A166 );
 a72551a <=( (not A232)  and  A200 );
 a72552a <=( a72551a  and  a72548a );
 a72553a <=( a72552a  and  a72545a );
 a72556a <=( (not A266)  and  (not A233) );
 a72559a <=( (not A269)  and  (not A268) );
 a72560a <=( a72559a  and  a72556a );
 a72563a <=( (not A299)  and  A298 );
 a72566a <=( A302  and  A300 );
 a72567a <=( a72566a  and  a72563a );
 a72568a <=( a72567a  and  a72560a );
 a72572a <=( (not A167)  and  (not A169) );
 a72573a <=( A170  and  a72572a );
 a72576a <=( (not A200)  and  A166 );
 a72579a <=( (not A203)  and  (not A202) );
 a72580a <=( a72579a  and  a72576a );
 a72581a <=( a72580a  and  a72573a );
 a72584a <=( A233  and  A232 );
 a72587a <=( (not A267)  and  A265 );
 a72588a <=( a72587a  and  a72584a );
 a72591a <=( (not A299)  and  A298 );
 a72594a <=( A301  and  A300 );
 a72595a <=( a72594a  and  a72591a );
 a72596a <=( a72595a  and  a72588a );
 a72600a <=( (not A167)  and  (not A169) );
 a72601a <=( A170  and  a72600a );
 a72604a <=( (not A200)  and  A166 );
 a72607a <=( (not A203)  and  (not A202) );
 a72608a <=( a72607a  and  a72604a );
 a72609a <=( a72608a  and  a72601a );
 a72612a <=( A233  and  A232 );
 a72615a <=( (not A267)  and  A265 );
 a72616a <=( a72615a  and  a72612a );
 a72619a <=( (not A299)  and  A298 );
 a72622a <=( A302  and  A300 );
 a72623a <=( a72622a  and  a72619a );
 a72624a <=( a72623a  and  a72616a );
 a72628a <=( (not A167)  and  (not A169) );
 a72629a <=( A170  and  a72628a );
 a72632a <=( (not A200)  and  A166 );
 a72635a <=( (not A203)  and  (not A202) );
 a72636a <=( a72635a  and  a72632a );
 a72637a <=( a72636a  and  a72629a );
 a72640a <=( A233  and  A232 );
 a72643a <=( A266  and  A265 );
 a72644a <=( a72643a  and  a72640a );
 a72647a <=( (not A299)  and  A298 );
 a72650a <=( A301  and  A300 );
 a72651a <=( a72650a  and  a72647a );
 a72652a <=( a72651a  and  a72644a );
 a72656a <=( (not A167)  and  (not A169) );
 a72657a <=( A170  and  a72656a );
 a72660a <=( (not A200)  and  A166 );
 a72663a <=( (not A203)  and  (not A202) );
 a72664a <=( a72663a  and  a72660a );
 a72665a <=( a72664a  and  a72657a );
 a72668a <=( A233  and  A232 );
 a72671a <=( A266  and  A265 );
 a72672a <=( a72671a  and  a72668a );
 a72675a <=( (not A299)  and  A298 );
 a72678a <=( A302  and  A300 );
 a72679a <=( a72678a  and  a72675a );
 a72680a <=( a72679a  and  a72672a );
 a72684a <=( (not A167)  and  (not A169) );
 a72685a <=( A170  and  a72684a );
 a72688a <=( (not A200)  and  A166 );
 a72691a <=( (not A203)  and  (not A202) );
 a72692a <=( a72691a  and  a72688a );
 a72693a <=( a72692a  and  a72685a );
 a72696a <=( A233  and  A232 );
 a72699a <=( (not A266)  and  (not A265) );
 a72700a <=( a72699a  and  a72696a );
 a72703a <=( (not A299)  and  A298 );
 a72706a <=( A301  and  A300 );
 a72707a <=( a72706a  and  a72703a );
 a72708a <=( a72707a  and  a72700a );
 a72712a <=( (not A167)  and  (not A169) );
 a72713a <=( A170  and  a72712a );
 a72716a <=( (not A200)  and  A166 );
 a72719a <=( (not A203)  and  (not A202) );
 a72720a <=( a72719a  and  a72716a );
 a72721a <=( a72720a  and  a72713a );
 a72724a <=( A233  and  A232 );
 a72727a <=( (not A266)  and  (not A265) );
 a72728a <=( a72727a  and  a72724a );
 a72731a <=( (not A299)  and  A298 );
 a72734a <=( A302  and  A300 );
 a72735a <=( a72734a  and  a72731a );
 a72736a <=( a72735a  and  a72728a );
 a72740a <=( (not A167)  and  (not A169) );
 a72741a <=( A170  and  a72740a );
 a72744a <=( (not A200)  and  A166 );
 a72747a <=( (not A203)  and  (not A202) );
 a72748a <=( a72747a  and  a72744a );
 a72749a <=( a72748a  and  a72741a );
 a72752a <=( (not A235)  and  (not A233) );
 a72755a <=( (not A266)  and  (not A236) );
 a72756a <=( a72755a  and  a72752a );
 a72759a <=( (not A269)  and  (not A268) );
 a72762a <=( A299  and  (not A298) );
 a72763a <=( a72762a  and  a72759a );
 a72764a <=( a72763a  and  a72756a );
 a72768a <=( (not A167)  and  (not A169) );
 a72769a <=( A170  and  a72768a );
 a72772a <=( (not A200)  and  A166 );
 a72775a <=( (not A203)  and  (not A202) );
 a72776a <=( a72775a  and  a72772a );
 a72777a <=( a72776a  and  a72769a );
 a72780a <=( (not A234)  and  (not A233) );
 a72783a <=( A266  and  A265 );
 a72784a <=( a72783a  and  a72780a );
 a72787a <=( (not A299)  and  A298 );
 a72790a <=( A301  and  A300 );
 a72791a <=( a72790a  and  a72787a );
 a72792a <=( a72791a  and  a72784a );
 a72796a <=( (not A167)  and  (not A169) );
 a72797a <=( A170  and  a72796a );
 a72800a <=( (not A200)  and  A166 );
 a72803a <=( (not A203)  and  (not A202) );
 a72804a <=( a72803a  and  a72800a );
 a72805a <=( a72804a  and  a72797a );
 a72808a <=( (not A234)  and  (not A233) );
 a72811a <=( A266  and  A265 );
 a72812a <=( a72811a  and  a72808a );
 a72815a <=( (not A299)  and  A298 );
 a72818a <=( A302  and  A300 );
 a72819a <=( a72818a  and  a72815a );
 a72820a <=( a72819a  and  a72812a );
 a72824a <=( (not A167)  and  (not A169) );
 a72825a <=( A170  and  a72824a );
 a72828a <=( (not A200)  and  A166 );
 a72831a <=( (not A203)  and  (not A202) );
 a72832a <=( a72831a  and  a72828a );
 a72833a <=( a72832a  and  a72825a );
 a72836a <=( (not A234)  and  (not A233) );
 a72839a <=( (not A267)  and  (not A266) );
 a72840a <=( a72839a  and  a72836a );
 a72843a <=( (not A299)  and  A298 );
 a72846a <=( A301  and  A300 );
 a72847a <=( a72846a  and  a72843a );
 a72848a <=( a72847a  and  a72840a );
 a72852a <=( (not A167)  and  (not A169) );
 a72853a <=( A170  and  a72852a );
 a72856a <=( (not A200)  and  A166 );
 a72859a <=( (not A203)  and  (not A202) );
 a72860a <=( a72859a  and  a72856a );
 a72861a <=( a72860a  and  a72853a );
 a72864a <=( (not A234)  and  (not A233) );
 a72867a <=( (not A267)  and  (not A266) );
 a72868a <=( a72867a  and  a72864a );
 a72871a <=( (not A299)  and  A298 );
 a72874a <=( A302  and  A300 );
 a72875a <=( a72874a  and  a72871a );
 a72876a <=( a72875a  and  a72868a );
 a72880a <=( (not A167)  and  (not A169) );
 a72881a <=( A170  and  a72880a );
 a72884a <=( (not A200)  and  A166 );
 a72887a <=( (not A203)  and  (not A202) );
 a72888a <=( a72887a  and  a72884a );
 a72889a <=( a72888a  and  a72881a );
 a72892a <=( (not A234)  and  (not A233) );
 a72895a <=( (not A266)  and  (not A265) );
 a72896a <=( a72895a  and  a72892a );
 a72899a <=( (not A299)  and  A298 );
 a72902a <=( A301  and  A300 );
 a72903a <=( a72902a  and  a72899a );
 a72904a <=( a72903a  and  a72896a );
 a72908a <=( (not A167)  and  (not A169) );
 a72909a <=( A170  and  a72908a );
 a72912a <=( (not A200)  and  A166 );
 a72915a <=( (not A203)  and  (not A202) );
 a72916a <=( a72915a  and  a72912a );
 a72917a <=( a72916a  and  a72909a );
 a72920a <=( (not A234)  and  (not A233) );
 a72923a <=( (not A266)  and  (not A265) );
 a72924a <=( a72923a  and  a72920a );
 a72927a <=( (not A299)  and  A298 );
 a72930a <=( A302  and  A300 );
 a72931a <=( a72930a  and  a72927a );
 a72932a <=( a72931a  and  a72924a );
 a72936a <=( (not A167)  and  (not A169) );
 a72937a <=( A170  and  a72936a );
 a72940a <=( (not A200)  and  A166 );
 a72943a <=( (not A203)  and  (not A202) );
 a72944a <=( a72943a  and  a72940a );
 a72945a <=( a72944a  and  a72937a );
 a72948a <=( (not A233)  and  A232 );
 a72951a <=( A235  and  A234 );
 a72952a <=( a72951a  and  a72948a );
 a72955a <=( (not A266)  and  A265 );
 a72958a <=( A268  and  A267 );
 a72959a <=( a72958a  and  a72955a );
 a72960a <=( a72959a  and  a72952a );
 a72964a <=( (not A167)  and  (not A169) );
 a72965a <=( A170  and  a72964a );
 a72968a <=( (not A200)  and  A166 );
 a72971a <=( (not A203)  and  (not A202) );
 a72972a <=( a72971a  and  a72968a );
 a72973a <=( a72972a  and  a72965a );
 a72976a <=( (not A233)  and  A232 );
 a72979a <=( A235  and  A234 );
 a72980a <=( a72979a  and  a72976a );
 a72983a <=( (not A266)  and  A265 );
 a72986a <=( A269  and  A267 );
 a72987a <=( a72986a  and  a72983a );
 a72988a <=( a72987a  and  a72980a );
 a72992a <=( (not A167)  and  (not A169) );
 a72993a <=( A170  and  a72992a );
 a72996a <=( (not A200)  and  A166 );
 a72999a <=( (not A203)  and  (not A202) );
 a73000a <=( a72999a  and  a72996a );
 a73001a <=( a73000a  and  a72993a );
 a73004a <=( (not A233)  and  A232 );
 a73007a <=( A236  and  A234 );
 a73008a <=( a73007a  and  a73004a );
 a73011a <=( (not A266)  and  A265 );
 a73014a <=( A268  and  A267 );
 a73015a <=( a73014a  and  a73011a );
 a73016a <=( a73015a  and  a73008a );
 a73020a <=( (not A167)  and  (not A169) );
 a73021a <=( A170  and  a73020a );
 a73024a <=( (not A200)  and  A166 );
 a73027a <=( (not A203)  and  (not A202) );
 a73028a <=( a73027a  and  a73024a );
 a73029a <=( a73028a  and  a73021a );
 a73032a <=( (not A233)  and  A232 );
 a73035a <=( A236  and  A234 );
 a73036a <=( a73035a  and  a73032a );
 a73039a <=( (not A266)  and  A265 );
 a73042a <=( A269  and  A267 );
 a73043a <=( a73042a  and  a73039a );
 a73044a <=( a73043a  and  a73036a );
 a73048a <=( (not A167)  and  (not A169) );
 a73049a <=( A170  and  a73048a );
 a73052a <=( (not A200)  and  A166 );
 a73055a <=( (not A203)  and  (not A202) );
 a73056a <=( a73055a  and  a73052a );
 a73057a <=( a73056a  and  a73049a );
 a73060a <=( (not A233)  and  (not A232) );
 a73063a <=( A266  and  A265 );
 a73064a <=( a73063a  and  a73060a );
 a73067a <=( (not A299)  and  A298 );
 a73070a <=( A301  and  A300 );
 a73071a <=( a73070a  and  a73067a );
 a73072a <=( a73071a  and  a73064a );
 a73076a <=( (not A167)  and  (not A169) );
 a73077a <=( A170  and  a73076a );
 a73080a <=( (not A200)  and  A166 );
 a73083a <=( (not A203)  and  (not A202) );
 a73084a <=( a73083a  and  a73080a );
 a73085a <=( a73084a  and  a73077a );
 a73088a <=( (not A233)  and  (not A232) );
 a73091a <=( A266  and  A265 );
 a73092a <=( a73091a  and  a73088a );
 a73095a <=( (not A299)  and  A298 );
 a73098a <=( A302  and  A300 );
 a73099a <=( a73098a  and  a73095a );
 a73100a <=( a73099a  and  a73092a );
 a73104a <=( (not A167)  and  (not A169) );
 a73105a <=( A170  and  a73104a );
 a73108a <=( (not A200)  and  A166 );
 a73111a <=( (not A203)  and  (not A202) );
 a73112a <=( a73111a  and  a73108a );
 a73113a <=( a73112a  and  a73105a );
 a73116a <=( (not A233)  and  (not A232) );
 a73119a <=( (not A267)  and  (not A266) );
 a73120a <=( a73119a  and  a73116a );
 a73123a <=( (not A299)  and  A298 );
 a73126a <=( A301  and  A300 );
 a73127a <=( a73126a  and  a73123a );
 a73128a <=( a73127a  and  a73120a );
 a73132a <=( (not A167)  and  (not A169) );
 a73133a <=( A170  and  a73132a );
 a73136a <=( (not A200)  and  A166 );
 a73139a <=( (not A203)  and  (not A202) );
 a73140a <=( a73139a  and  a73136a );
 a73141a <=( a73140a  and  a73133a );
 a73144a <=( (not A233)  and  (not A232) );
 a73147a <=( (not A267)  and  (not A266) );
 a73148a <=( a73147a  and  a73144a );
 a73151a <=( (not A299)  and  A298 );
 a73154a <=( A302  and  A300 );
 a73155a <=( a73154a  and  a73151a );
 a73156a <=( a73155a  and  a73148a );
 a73160a <=( (not A167)  and  (not A169) );
 a73161a <=( A170  and  a73160a );
 a73164a <=( (not A200)  and  A166 );
 a73167a <=( (not A203)  and  (not A202) );
 a73168a <=( a73167a  and  a73164a );
 a73169a <=( a73168a  and  a73161a );
 a73172a <=( (not A233)  and  (not A232) );
 a73175a <=( (not A266)  and  (not A265) );
 a73176a <=( a73175a  and  a73172a );
 a73179a <=( (not A299)  and  A298 );
 a73182a <=( A301  and  A300 );
 a73183a <=( a73182a  and  a73179a );
 a73184a <=( a73183a  and  a73176a );
 a73188a <=( (not A167)  and  (not A169) );
 a73189a <=( A170  and  a73188a );
 a73192a <=( (not A200)  and  A166 );
 a73195a <=( (not A203)  and  (not A202) );
 a73196a <=( a73195a  and  a73192a );
 a73197a <=( a73196a  and  a73189a );
 a73200a <=( (not A233)  and  (not A232) );
 a73203a <=( (not A266)  and  (not A265) );
 a73204a <=( a73203a  and  a73200a );
 a73207a <=( (not A299)  and  A298 );
 a73210a <=( A302  and  A300 );
 a73211a <=( a73210a  and  a73207a );
 a73212a <=( a73211a  and  a73204a );
 a73216a <=( (not A167)  and  (not A169) );
 a73217a <=( A170  and  a73216a );
 a73220a <=( (not A200)  and  A166 );
 a73223a <=( A232  and  (not A201) );
 a73224a <=( a73223a  and  a73220a );
 a73225a <=( a73224a  and  a73217a );
 a73228a <=( A265  and  A233 );
 a73231a <=( (not A269)  and  (not A268) );
 a73232a <=( a73231a  and  a73228a );
 a73235a <=( (not A299)  and  A298 );
 a73238a <=( A301  and  A300 );
 a73239a <=( a73238a  and  a73235a );
 a73240a <=( a73239a  and  a73232a );
 a73244a <=( (not A167)  and  (not A169) );
 a73245a <=( A170  and  a73244a );
 a73248a <=( (not A200)  and  A166 );
 a73251a <=( A232  and  (not A201) );
 a73252a <=( a73251a  and  a73248a );
 a73253a <=( a73252a  and  a73245a );
 a73256a <=( A265  and  A233 );
 a73259a <=( (not A269)  and  (not A268) );
 a73260a <=( a73259a  and  a73256a );
 a73263a <=( (not A299)  and  A298 );
 a73266a <=( A302  and  A300 );
 a73267a <=( a73266a  and  a73263a );
 a73268a <=( a73267a  and  a73260a );
 a73272a <=( (not A167)  and  (not A169) );
 a73273a <=( A170  and  a73272a );
 a73276a <=( (not A200)  and  A166 );
 a73279a <=( (not A233)  and  (not A201) );
 a73280a <=( a73279a  and  a73276a );
 a73281a <=( a73280a  and  a73273a );
 a73284a <=( (not A236)  and  (not A235) );
 a73287a <=( A266  and  A265 );
 a73288a <=( a73287a  and  a73284a );
 a73291a <=( (not A299)  and  A298 );
 a73294a <=( A301  and  A300 );
 a73295a <=( a73294a  and  a73291a );
 a73296a <=( a73295a  and  a73288a );
 a73300a <=( (not A167)  and  (not A169) );
 a73301a <=( A170  and  a73300a );
 a73304a <=( (not A200)  and  A166 );
 a73307a <=( (not A233)  and  (not A201) );
 a73308a <=( a73307a  and  a73304a );
 a73309a <=( a73308a  and  a73301a );
 a73312a <=( (not A236)  and  (not A235) );
 a73315a <=( A266  and  A265 );
 a73316a <=( a73315a  and  a73312a );
 a73319a <=( (not A299)  and  A298 );
 a73322a <=( A302  and  A300 );
 a73323a <=( a73322a  and  a73319a );
 a73324a <=( a73323a  and  a73316a );
 a73328a <=( (not A167)  and  (not A169) );
 a73329a <=( A170  and  a73328a );
 a73332a <=( (not A200)  and  A166 );
 a73335a <=( (not A233)  and  (not A201) );
 a73336a <=( a73335a  and  a73332a );
 a73337a <=( a73336a  and  a73329a );
 a73340a <=( (not A236)  and  (not A235) );
 a73343a <=( (not A267)  and  (not A266) );
 a73344a <=( a73343a  and  a73340a );
 a73347a <=( (not A299)  and  A298 );
 a73350a <=( A301  and  A300 );
 a73351a <=( a73350a  and  a73347a );
 a73352a <=( a73351a  and  a73344a );
 a73356a <=( (not A167)  and  (not A169) );
 a73357a <=( A170  and  a73356a );
 a73360a <=( (not A200)  and  A166 );
 a73363a <=( (not A233)  and  (not A201) );
 a73364a <=( a73363a  and  a73360a );
 a73365a <=( a73364a  and  a73357a );
 a73368a <=( (not A236)  and  (not A235) );
 a73371a <=( (not A267)  and  (not A266) );
 a73372a <=( a73371a  and  a73368a );
 a73375a <=( (not A299)  and  A298 );
 a73378a <=( A302  and  A300 );
 a73379a <=( a73378a  and  a73375a );
 a73380a <=( a73379a  and  a73372a );
 a73384a <=( (not A167)  and  (not A169) );
 a73385a <=( A170  and  a73384a );
 a73388a <=( (not A200)  and  A166 );
 a73391a <=( (not A233)  and  (not A201) );
 a73392a <=( a73391a  and  a73388a );
 a73393a <=( a73392a  and  a73385a );
 a73396a <=( (not A236)  and  (not A235) );
 a73399a <=( (not A266)  and  (not A265) );
 a73400a <=( a73399a  and  a73396a );
 a73403a <=( (not A299)  and  A298 );
 a73406a <=( A301  and  A300 );
 a73407a <=( a73406a  and  a73403a );
 a73408a <=( a73407a  and  a73400a );
 a73412a <=( (not A167)  and  (not A169) );
 a73413a <=( A170  and  a73412a );
 a73416a <=( (not A200)  and  A166 );
 a73419a <=( (not A233)  and  (not A201) );
 a73420a <=( a73419a  and  a73416a );
 a73421a <=( a73420a  and  a73413a );
 a73424a <=( (not A236)  and  (not A235) );
 a73427a <=( (not A266)  and  (not A265) );
 a73428a <=( a73427a  and  a73424a );
 a73431a <=( (not A299)  and  A298 );
 a73434a <=( A302  and  A300 );
 a73435a <=( a73434a  and  a73431a );
 a73436a <=( a73435a  and  a73428a );
 a73440a <=( (not A167)  and  (not A169) );
 a73441a <=( A170  and  a73440a );
 a73444a <=( (not A200)  and  A166 );
 a73447a <=( (not A233)  and  (not A201) );
 a73448a <=( a73447a  and  a73444a );
 a73449a <=( a73448a  and  a73441a );
 a73452a <=( (not A266)  and  (not A234) );
 a73455a <=( (not A269)  and  (not A268) );
 a73456a <=( a73455a  and  a73452a );
 a73459a <=( (not A299)  and  A298 );
 a73462a <=( A301  and  A300 );
 a73463a <=( a73462a  and  a73459a );
 a73464a <=( a73463a  and  a73456a );
 a73468a <=( (not A167)  and  (not A169) );
 a73469a <=( A170  and  a73468a );
 a73472a <=( (not A200)  and  A166 );
 a73475a <=( (not A233)  and  (not A201) );
 a73476a <=( a73475a  and  a73472a );
 a73477a <=( a73476a  and  a73469a );
 a73480a <=( (not A266)  and  (not A234) );
 a73483a <=( (not A269)  and  (not A268) );
 a73484a <=( a73483a  and  a73480a );
 a73487a <=( (not A299)  and  A298 );
 a73490a <=( A302  and  A300 );
 a73491a <=( a73490a  and  a73487a );
 a73492a <=( a73491a  and  a73484a );
 a73496a <=( (not A167)  and  (not A169) );
 a73497a <=( A170  and  a73496a );
 a73500a <=( (not A200)  and  A166 );
 a73503a <=( (not A232)  and  (not A201) );
 a73504a <=( a73503a  and  a73500a );
 a73505a <=( a73504a  and  a73497a );
 a73508a <=( (not A266)  and  (not A233) );
 a73511a <=( (not A269)  and  (not A268) );
 a73512a <=( a73511a  and  a73508a );
 a73515a <=( (not A299)  and  A298 );
 a73518a <=( A301  and  A300 );
 a73519a <=( a73518a  and  a73515a );
 a73520a <=( a73519a  and  a73512a );
 a73524a <=( (not A167)  and  (not A169) );
 a73525a <=( A170  and  a73524a );
 a73528a <=( (not A200)  and  A166 );
 a73531a <=( (not A232)  and  (not A201) );
 a73532a <=( a73531a  and  a73528a );
 a73533a <=( a73532a  and  a73525a );
 a73536a <=( (not A266)  and  (not A233) );
 a73539a <=( (not A269)  and  (not A268) );
 a73540a <=( a73539a  and  a73536a );
 a73543a <=( (not A299)  and  A298 );
 a73546a <=( A302  and  A300 );
 a73547a <=( a73546a  and  a73543a );
 a73548a <=( a73547a  and  a73540a );
 a73552a <=( (not A167)  and  (not A169) );
 a73553a <=( A170  and  a73552a );
 a73556a <=( (not A199)  and  A166 );
 a73559a <=( A232  and  (not A200) );
 a73560a <=( a73559a  and  a73556a );
 a73561a <=( a73560a  and  a73553a );
 a73564a <=( A265  and  A233 );
 a73567a <=( (not A269)  and  (not A268) );
 a73568a <=( a73567a  and  a73564a );
 a73571a <=( (not A299)  and  A298 );
 a73574a <=( A301  and  A300 );
 a73575a <=( a73574a  and  a73571a );
 a73576a <=( a73575a  and  a73568a );
 a73580a <=( (not A167)  and  (not A169) );
 a73581a <=( A170  and  a73580a );
 a73584a <=( (not A199)  and  A166 );
 a73587a <=( A232  and  (not A200) );
 a73588a <=( a73587a  and  a73584a );
 a73589a <=( a73588a  and  a73581a );
 a73592a <=( A265  and  A233 );
 a73595a <=( (not A269)  and  (not A268) );
 a73596a <=( a73595a  and  a73592a );
 a73599a <=( (not A299)  and  A298 );
 a73602a <=( A302  and  A300 );
 a73603a <=( a73602a  and  a73599a );
 a73604a <=( a73603a  and  a73596a );
 a73608a <=( (not A167)  and  (not A169) );
 a73609a <=( A170  and  a73608a );
 a73612a <=( (not A199)  and  A166 );
 a73615a <=( (not A233)  and  (not A200) );
 a73616a <=( a73615a  and  a73612a );
 a73617a <=( a73616a  and  a73609a );
 a73620a <=( (not A236)  and  (not A235) );
 a73623a <=( A266  and  A265 );
 a73624a <=( a73623a  and  a73620a );
 a73627a <=( (not A299)  and  A298 );
 a73630a <=( A301  and  A300 );
 a73631a <=( a73630a  and  a73627a );
 a73632a <=( a73631a  and  a73624a );
 a73636a <=( (not A167)  and  (not A169) );
 a73637a <=( A170  and  a73636a );
 a73640a <=( (not A199)  and  A166 );
 a73643a <=( (not A233)  and  (not A200) );
 a73644a <=( a73643a  and  a73640a );
 a73645a <=( a73644a  and  a73637a );
 a73648a <=( (not A236)  and  (not A235) );
 a73651a <=( A266  and  A265 );
 a73652a <=( a73651a  and  a73648a );
 a73655a <=( (not A299)  and  A298 );
 a73658a <=( A302  and  A300 );
 a73659a <=( a73658a  and  a73655a );
 a73660a <=( a73659a  and  a73652a );
 a73664a <=( (not A167)  and  (not A169) );
 a73665a <=( A170  and  a73664a );
 a73668a <=( (not A199)  and  A166 );
 a73671a <=( (not A233)  and  (not A200) );
 a73672a <=( a73671a  and  a73668a );
 a73673a <=( a73672a  and  a73665a );
 a73676a <=( (not A236)  and  (not A235) );
 a73679a <=( (not A267)  and  (not A266) );
 a73680a <=( a73679a  and  a73676a );
 a73683a <=( (not A299)  and  A298 );
 a73686a <=( A301  and  A300 );
 a73687a <=( a73686a  and  a73683a );
 a73688a <=( a73687a  and  a73680a );
 a73692a <=( (not A167)  and  (not A169) );
 a73693a <=( A170  and  a73692a );
 a73696a <=( (not A199)  and  A166 );
 a73699a <=( (not A233)  and  (not A200) );
 a73700a <=( a73699a  and  a73696a );
 a73701a <=( a73700a  and  a73693a );
 a73704a <=( (not A236)  and  (not A235) );
 a73707a <=( (not A267)  and  (not A266) );
 a73708a <=( a73707a  and  a73704a );
 a73711a <=( (not A299)  and  A298 );
 a73714a <=( A302  and  A300 );
 a73715a <=( a73714a  and  a73711a );
 a73716a <=( a73715a  and  a73708a );
 a73720a <=( (not A167)  and  (not A169) );
 a73721a <=( A170  and  a73720a );
 a73724a <=( (not A199)  and  A166 );
 a73727a <=( (not A233)  and  (not A200) );
 a73728a <=( a73727a  and  a73724a );
 a73729a <=( a73728a  and  a73721a );
 a73732a <=( (not A236)  and  (not A235) );
 a73735a <=( (not A266)  and  (not A265) );
 a73736a <=( a73735a  and  a73732a );
 a73739a <=( (not A299)  and  A298 );
 a73742a <=( A301  and  A300 );
 a73743a <=( a73742a  and  a73739a );
 a73744a <=( a73743a  and  a73736a );
 a73748a <=( (not A167)  and  (not A169) );
 a73749a <=( A170  and  a73748a );
 a73752a <=( (not A199)  and  A166 );
 a73755a <=( (not A233)  and  (not A200) );
 a73756a <=( a73755a  and  a73752a );
 a73757a <=( a73756a  and  a73749a );
 a73760a <=( (not A236)  and  (not A235) );
 a73763a <=( (not A266)  and  (not A265) );
 a73764a <=( a73763a  and  a73760a );
 a73767a <=( (not A299)  and  A298 );
 a73770a <=( A302  and  A300 );
 a73771a <=( a73770a  and  a73767a );
 a73772a <=( a73771a  and  a73764a );
 a73776a <=( (not A167)  and  (not A169) );
 a73777a <=( A170  and  a73776a );
 a73780a <=( (not A199)  and  A166 );
 a73783a <=( (not A233)  and  (not A200) );
 a73784a <=( a73783a  and  a73780a );
 a73785a <=( a73784a  and  a73777a );
 a73788a <=( (not A266)  and  (not A234) );
 a73791a <=( (not A269)  and  (not A268) );
 a73792a <=( a73791a  and  a73788a );
 a73795a <=( (not A299)  and  A298 );
 a73798a <=( A301  and  A300 );
 a73799a <=( a73798a  and  a73795a );
 a73800a <=( a73799a  and  a73792a );
 a73804a <=( (not A167)  and  (not A169) );
 a73805a <=( A170  and  a73804a );
 a73808a <=( (not A199)  and  A166 );
 a73811a <=( (not A233)  and  (not A200) );
 a73812a <=( a73811a  and  a73808a );
 a73813a <=( a73812a  and  a73805a );
 a73816a <=( (not A266)  and  (not A234) );
 a73819a <=( (not A269)  and  (not A268) );
 a73820a <=( a73819a  and  a73816a );
 a73823a <=( (not A299)  and  A298 );
 a73826a <=( A302  and  A300 );
 a73827a <=( a73826a  and  a73823a );
 a73828a <=( a73827a  and  a73820a );
 a73832a <=( (not A167)  and  (not A169) );
 a73833a <=( A170  and  a73832a );
 a73836a <=( (not A199)  and  A166 );
 a73839a <=( (not A232)  and  (not A200) );
 a73840a <=( a73839a  and  a73836a );
 a73841a <=( a73840a  and  a73833a );
 a73844a <=( (not A266)  and  (not A233) );
 a73847a <=( (not A269)  and  (not A268) );
 a73848a <=( a73847a  and  a73844a );
 a73851a <=( (not A299)  and  A298 );
 a73854a <=( A301  and  A300 );
 a73855a <=( a73854a  and  a73851a );
 a73856a <=( a73855a  and  a73848a );
 a73860a <=( (not A167)  and  (not A169) );
 a73861a <=( A170  and  a73860a );
 a73864a <=( (not A199)  and  A166 );
 a73867a <=( (not A232)  and  (not A200) );
 a73868a <=( a73867a  and  a73864a );
 a73869a <=( a73868a  and  a73861a );
 a73872a <=( (not A266)  and  (not A233) );
 a73875a <=( (not A269)  and  (not A268) );
 a73876a <=( a73875a  and  a73872a );
 a73879a <=( (not A299)  and  A298 );
 a73882a <=( A302  and  A300 );
 a73883a <=( a73882a  and  a73879a );
 a73884a <=( a73883a  and  a73876a );
 a73888a <=( (not A168)  and  (not A169) );
 a73889a <=( (not A170)  and  a73888a );
 a73892a <=( (not A200)  and  A199 );
 a73895a <=( A202  and  A201 );
 a73896a <=( a73895a  and  a73892a );
 a73897a <=( a73896a  and  a73889a );
 a73900a <=( A233  and  A232 );
 a73903a <=( (not A267)  and  A265 );
 a73904a <=( a73903a  and  a73900a );
 a73907a <=( (not A299)  and  A298 );
 a73910a <=( A301  and  A300 );
 a73911a <=( a73910a  and  a73907a );
 a73912a <=( a73911a  and  a73904a );
 a73916a <=( (not A168)  and  (not A169) );
 a73917a <=( (not A170)  and  a73916a );
 a73920a <=( (not A200)  and  A199 );
 a73923a <=( A202  and  A201 );
 a73924a <=( a73923a  and  a73920a );
 a73925a <=( a73924a  and  a73917a );
 a73928a <=( A233  and  A232 );
 a73931a <=( (not A267)  and  A265 );
 a73932a <=( a73931a  and  a73928a );
 a73935a <=( (not A299)  and  A298 );
 a73938a <=( A302  and  A300 );
 a73939a <=( a73938a  and  a73935a );
 a73940a <=( a73939a  and  a73932a );
 a73944a <=( (not A168)  and  (not A169) );
 a73945a <=( (not A170)  and  a73944a );
 a73948a <=( (not A200)  and  A199 );
 a73951a <=( A202  and  A201 );
 a73952a <=( a73951a  and  a73948a );
 a73953a <=( a73952a  and  a73945a );
 a73956a <=( A233  and  A232 );
 a73959a <=( A266  and  A265 );
 a73960a <=( a73959a  and  a73956a );
 a73963a <=( (not A299)  and  A298 );
 a73966a <=( A301  and  A300 );
 a73967a <=( a73966a  and  a73963a );
 a73968a <=( a73967a  and  a73960a );
 a73972a <=( (not A168)  and  (not A169) );
 a73973a <=( (not A170)  and  a73972a );
 a73976a <=( (not A200)  and  A199 );
 a73979a <=( A202  and  A201 );
 a73980a <=( a73979a  and  a73976a );
 a73981a <=( a73980a  and  a73973a );
 a73984a <=( A233  and  A232 );
 a73987a <=( A266  and  A265 );
 a73988a <=( a73987a  and  a73984a );
 a73991a <=( (not A299)  and  A298 );
 a73994a <=( A302  and  A300 );
 a73995a <=( a73994a  and  a73991a );
 a73996a <=( a73995a  and  a73988a );
 a74000a <=( (not A168)  and  (not A169) );
 a74001a <=( (not A170)  and  a74000a );
 a74004a <=( (not A200)  and  A199 );
 a74007a <=( A202  and  A201 );
 a74008a <=( a74007a  and  a74004a );
 a74009a <=( a74008a  and  a74001a );
 a74012a <=( A233  and  A232 );
 a74015a <=( (not A266)  and  (not A265) );
 a74016a <=( a74015a  and  a74012a );
 a74019a <=( (not A299)  and  A298 );
 a74022a <=( A301  and  A300 );
 a74023a <=( a74022a  and  a74019a );
 a74024a <=( a74023a  and  a74016a );
 a74028a <=( (not A168)  and  (not A169) );
 a74029a <=( (not A170)  and  a74028a );
 a74032a <=( (not A200)  and  A199 );
 a74035a <=( A202  and  A201 );
 a74036a <=( a74035a  and  a74032a );
 a74037a <=( a74036a  and  a74029a );
 a74040a <=( A233  and  A232 );
 a74043a <=( (not A266)  and  (not A265) );
 a74044a <=( a74043a  and  a74040a );
 a74047a <=( (not A299)  and  A298 );
 a74050a <=( A302  and  A300 );
 a74051a <=( a74050a  and  a74047a );
 a74052a <=( a74051a  and  a74044a );
 a74056a <=( (not A168)  and  (not A169) );
 a74057a <=( (not A170)  and  a74056a );
 a74060a <=( (not A200)  and  A199 );
 a74063a <=( A202  and  A201 );
 a74064a <=( a74063a  and  a74060a );
 a74065a <=( a74064a  and  a74057a );
 a74068a <=( (not A235)  and  (not A233) );
 a74071a <=( (not A266)  and  (not A236) );
 a74072a <=( a74071a  and  a74068a );
 a74075a <=( (not A269)  and  (not A268) );
 a74078a <=( A299  and  (not A298) );
 a74079a <=( a74078a  and  a74075a );
 a74080a <=( a74079a  and  a74072a );
 a74084a <=( (not A168)  and  (not A169) );
 a74085a <=( (not A170)  and  a74084a );
 a74088a <=( (not A200)  and  A199 );
 a74091a <=( A202  and  A201 );
 a74092a <=( a74091a  and  a74088a );
 a74093a <=( a74092a  and  a74085a );
 a74096a <=( (not A234)  and  (not A233) );
 a74099a <=( A266  and  A265 );
 a74100a <=( a74099a  and  a74096a );
 a74103a <=( (not A299)  and  A298 );
 a74106a <=( A301  and  A300 );
 a74107a <=( a74106a  and  a74103a );
 a74108a <=( a74107a  and  a74100a );
 a74112a <=( (not A168)  and  (not A169) );
 a74113a <=( (not A170)  and  a74112a );
 a74116a <=( (not A200)  and  A199 );
 a74119a <=( A202  and  A201 );
 a74120a <=( a74119a  and  a74116a );
 a74121a <=( a74120a  and  a74113a );
 a74124a <=( (not A234)  and  (not A233) );
 a74127a <=( A266  and  A265 );
 a74128a <=( a74127a  and  a74124a );
 a74131a <=( (not A299)  and  A298 );
 a74134a <=( A302  and  A300 );
 a74135a <=( a74134a  and  a74131a );
 a74136a <=( a74135a  and  a74128a );
 a74140a <=( (not A168)  and  (not A169) );
 a74141a <=( (not A170)  and  a74140a );
 a74144a <=( (not A200)  and  A199 );
 a74147a <=( A202  and  A201 );
 a74148a <=( a74147a  and  a74144a );
 a74149a <=( a74148a  and  a74141a );
 a74152a <=( (not A234)  and  (not A233) );
 a74155a <=( (not A267)  and  (not A266) );
 a74156a <=( a74155a  and  a74152a );
 a74159a <=( (not A299)  and  A298 );
 a74162a <=( A301  and  A300 );
 a74163a <=( a74162a  and  a74159a );
 a74164a <=( a74163a  and  a74156a );
 a74168a <=( (not A168)  and  (not A169) );
 a74169a <=( (not A170)  and  a74168a );
 a74172a <=( (not A200)  and  A199 );
 a74175a <=( A202  and  A201 );
 a74176a <=( a74175a  and  a74172a );
 a74177a <=( a74176a  and  a74169a );
 a74180a <=( (not A234)  and  (not A233) );
 a74183a <=( (not A267)  and  (not A266) );
 a74184a <=( a74183a  and  a74180a );
 a74187a <=( (not A299)  and  A298 );
 a74190a <=( A302  and  A300 );
 a74191a <=( a74190a  and  a74187a );
 a74192a <=( a74191a  and  a74184a );
 a74196a <=( (not A168)  and  (not A169) );
 a74197a <=( (not A170)  and  a74196a );
 a74200a <=( (not A200)  and  A199 );
 a74203a <=( A202  and  A201 );
 a74204a <=( a74203a  and  a74200a );
 a74205a <=( a74204a  and  a74197a );
 a74208a <=( (not A234)  and  (not A233) );
 a74211a <=( (not A266)  and  (not A265) );
 a74212a <=( a74211a  and  a74208a );
 a74215a <=( (not A299)  and  A298 );
 a74218a <=( A301  and  A300 );
 a74219a <=( a74218a  and  a74215a );
 a74220a <=( a74219a  and  a74212a );
 a74224a <=( (not A168)  and  (not A169) );
 a74225a <=( (not A170)  and  a74224a );
 a74228a <=( (not A200)  and  A199 );
 a74231a <=( A202  and  A201 );
 a74232a <=( a74231a  and  a74228a );
 a74233a <=( a74232a  and  a74225a );
 a74236a <=( (not A234)  and  (not A233) );
 a74239a <=( (not A266)  and  (not A265) );
 a74240a <=( a74239a  and  a74236a );
 a74243a <=( (not A299)  and  A298 );
 a74246a <=( A302  and  A300 );
 a74247a <=( a74246a  and  a74243a );
 a74248a <=( a74247a  and  a74240a );
 a74252a <=( (not A168)  and  (not A169) );
 a74253a <=( (not A170)  and  a74252a );
 a74256a <=( (not A200)  and  A199 );
 a74259a <=( A202  and  A201 );
 a74260a <=( a74259a  and  a74256a );
 a74261a <=( a74260a  and  a74253a );
 a74264a <=( (not A233)  and  A232 );
 a74267a <=( A235  and  A234 );
 a74268a <=( a74267a  and  a74264a );
 a74271a <=( (not A266)  and  A265 );
 a74274a <=( A268  and  A267 );
 a74275a <=( a74274a  and  a74271a );
 a74276a <=( a74275a  and  a74268a );
 a74280a <=( (not A168)  and  (not A169) );
 a74281a <=( (not A170)  and  a74280a );
 a74284a <=( (not A200)  and  A199 );
 a74287a <=( A202  and  A201 );
 a74288a <=( a74287a  and  a74284a );
 a74289a <=( a74288a  and  a74281a );
 a74292a <=( (not A233)  and  A232 );
 a74295a <=( A235  and  A234 );
 a74296a <=( a74295a  and  a74292a );
 a74299a <=( (not A266)  and  A265 );
 a74302a <=( A269  and  A267 );
 a74303a <=( a74302a  and  a74299a );
 a74304a <=( a74303a  and  a74296a );
 a74308a <=( (not A168)  and  (not A169) );
 a74309a <=( (not A170)  and  a74308a );
 a74312a <=( (not A200)  and  A199 );
 a74315a <=( A202  and  A201 );
 a74316a <=( a74315a  and  a74312a );
 a74317a <=( a74316a  and  a74309a );
 a74320a <=( (not A233)  and  A232 );
 a74323a <=( A236  and  A234 );
 a74324a <=( a74323a  and  a74320a );
 a74327a <=( (not A266)  and  A265 );
 a74330a <=( A268  and  A267 );
 a74331a <=( a74330a  and  a74327a );
 a74332a <=( a74331a  and  a74324a );
 a74336a <=( (not A168)  and  (not A169) );
 a74337a <=( (not A170)  and  a74336a );
 a74340a <=( (not A200)  and  A199 );
 a74343a <=( A202  and  A201 );
 a74344a <=( a74343a  and  a74340a );
 a74345a <=( a74344a  and  a74337a );
 a74348a <=( (not A233)  and  A232 );
 a74351a <=( A236  and  A234 );
 a74352a <=( a74351a  and  a74348a );
 a74355a <=( (not A266)  and  A265 );
 a74358a <=( A269  and  A267 );
 a74359a <=( a74358a  and  a74355a );
 a74360a <=( a74359a  and  a74352a );
 a74364a <=( (not A168)  and  (not A169) );
 a74365a <=( (not A170)  and  a74364a );
 a74368a <=( (not A200)  and  A199 );
 a74371a <=( A202  and  A201 );
 a74372a <=( a74371a  and  a74368a );
 a74373a <=( a74372a  and  a74365a );
 a74376a <=( (not A233)  and  (not A232) );
 a74379a <=( A266  and  A265 );
 a74380a <=( a74379a  and  a74376a );
 a74383a <=( (not A299)  and  A298 );
 a74386a <=( A301  and  A300 );
 a74387a <=( a74386a  and  a74383a );
 a74388a <=( a74387a  and  a74380a );
 a74392a <=( (not A168)  and  (not A169) );
 a74393a <=( (not A170)  and  a74392a );
 a74396a <=( (not A200)  and  A199 );
 a74399a <=( A202  and  A201 );
 a74400a <=( a74399a  and  a74396a );
 a74401a <=( a74400a  and  a74393a );
 a74404a <=( (not A233)  and  (not A232) );
 a74407a <=( A266  and  A265 );
 a74408a <=( a74407a  and  a74404a );
 a74411a <=( (not A299)  and  A298 );
 a74414a <=( A302  and  A300 );
 a74415a <=( a74414a  and  a74411a );
 a74416a <=( a74415a  and  a74408a );
 a74420a <=( (not A168)  and  (not A169) );
 a74421a <=( (not A170)  and  a74420a );
 a74424a <=( (not A200)  and  A199 );
 a74427a <=( A202  and  A201 );
 a74428a <=( a74427a  and  a74424a );
 a74429a <=( a74428a  and  a74421a );
 a74432a <=( (not A233)  and  (not A232) );
 a74435a <=( (not A267)  and  (not A266) );
 a74436a <=( a74435a  and  a74432a );
 a74439a <=( (not A299)  and  A298 );
 a74442a <=( A301  and  A300 );
 a74443a <=( a74442a  and  a74439a );
 a74444a <=( a74443a  and  a74436a );
 a74448a <=( (not A168)  and  (not A169) );
 a74449a <=( (not A170)  and  a74448a );
 a74452a <=( (not A200)  and  A199 );
 a74455a <=( A202  and  A201 );
 a74456a <=( a74455a  and  a74452a );
 a74457a <=( a74456a  and  a74449a );
 a74460a <=( (not A233)  and  (not A232) );
 a74463a <=( (not A267)  and  (not A266) );
 a74464a <=( a74463a  and  a74460a );
 a74467a <=( (not A299)  and  A298 );
 a74470a <=( A302  and  A300 );
 a74471a <=( a74470a  and  a74467a );
 a74472a <=( a74471a  and  a74464a );
 a74476a <=( (not A168)  and  (not A169) );
 a74477a <=( (not A170)  and  a74476a );
 a74480a <=( (not A200)  and  A199 );
 a74483a <=( A202  and  A201 );
 a74484a <=( a74483a  and  a74480a );
 a74485a <=( a74484a  and  a74477a );
 a74488a <=( (not A233)  and  (not A232) );
 a74491a <=( (not A266)  and  (not A265) );
 a74492a <=( a74491a  and  a74488a );
 a74495a <=( (not A299)  and  A298 );
 a74498a <=( A301  and  A300 );
 a74499a <=( a74498a  and  a74495a );
 a74500a <=( a74499a  and  a74492a );
 a74504a <=( (not A168)  and  (not A169) );
 a74505a <=( (not A170)  and  a74504a );
 a74508a <=( (not A200)  and  A199 );
 a74511a <=( A202  and  A201 );
 a74512a <=( a74511a  and  a74508a );
 a74513a <=( a74512a  and  a74505a );
 a74516a <=( (not A233)  and  (not A232) );
 a74519a <=( (not A266)  and  (not A265) );
 a74520a <=( a74519a  and  a74516a );
 a74523a <=( (not A299)  and  A298 );
 a74526a <=( A302  and  A300 );
 a74527a <=( a74526a  and  a74523a );
 a74528a <=( a74527a  and  a74520a );
 a74532a <=( (not A168)  and  (not A169) );
 a74533a <=( (not A170)  and  a74532a );
 a74536a <=( (not A200)  and  A199 );
 a74539a <=( A203  and  A201 );
 a74540a <=( a74539a  and  a74536a );
 a74541a <=( a74540a  and  a74533a );
 a74544a <=( A233  and  A232 );
 a74547a <=( (not A267)  and  A265 );
 a74548a <=( a74547a  and  a74544a );
 a74551a <=( (not A299)  and  A298 );
 a74554a <=( A301  and  A300 );
 a74555a <=( a74554a  and  a74551a );
 a74556a <=( a74555a  and  a74548a );
 a74560a <=( (not A168)  and  (not A169) );
 a74561a <=( (not A170)  and  a74560a );
 a74564a <=( (not A200)  and  A199 );
 a74567a <=( A203  and  A201 );
 a74568a <=( a74567a  and  a74564a );
 a74569a <=( a74568a  and  a74561a );
 a74572a <=( A233  and  A232 );
 a74575a <=( (not A267)  and  A265 );
 a74576a <=( a74575a  and  a74572a );
 a74579a <=( (not A299)  and  A298 );
 a74582a <=( A302  and  A300 );
 a74583a <=( a74582a  and  a74579a );
 a74584a <=( a74583a  and  a74576a );
 a74588a <=( (not A168)  and  (not A169) );
 a74589a <=( (not A170)  and  a74588a );
 a74592a <=( (not A200)  and  A199 );
 a74595a <=( A203  and  A201 );
 a74596a <=( a74595a  and  a74592a );
 a74597a <=( a74596a  and  a74589a );
 a74600a <=( A233  and  A232 );
 a74603a <=( A266  and  A265 );
 a74604a <=( a74603a  and  a74600a );
 a74607a <=( (not A299)  and  A298 );
 a74610a <=( A301  and  A300 );
 a74611a <=( a74610a  and  a74607a );
 a74612a <=( a74611a  and  a74604a );
 a74616a <=( (not A168)  and  (not A169) );
 a74617a <=( (not A170)  and  a74616a );
 a74620a <=( (not A200)  and  A199 );
 a74623a <=( A203  and  A201 );
 a74624a <=( a74623a  and  a74620a );
 a74625a <=( a74624a  and  a74617a );
 a74628a <=( A233  and  A232 );
 a74631a <=( A266  and  A265 );
 a74632a <=( a74631a  and  a74628a );
 a74635a <=( (not A299)  and  A298 );
 a74638a <=( A302  and  A300 );
 a74639a <=( a74638a  and  a74635a );
 a74640a <=( a74639a  and  a74632a );
 a74644a <=( (not A168)  and  (not A169) );
 a74645a <=( (not A170)  and  a74644a );
 a74648a <=( (not A200)  and  A199 );
 a74651a <=( A203  and  A201 );
 a74652a <=( a74651a  and  a74648a );
 a74653a <=( a74652a  and  a74645a );
 a74656a <=( A233  and  A232 );
 a74659a <=( (not A266)  and  (not A265) );
 a74660a <=( a74659a  and  a74656a );
 a74663a <=( (not A299)  and  A298 );
 a74666a <=( A301  and  A300 );
 a74667a <=( a74666a  and  a74663a );
 a74668a <=( a74667a  and  a74660a );
 a74672a <=( (not A168)  and  (not A169) );
 a74673a <=( (not A170)  and  a74672a );
 a74676a <=( (not A200)  and  A199 );
 a74679a <=( A203  and  A201 );
 a74680a <=( a74679a  and  a74676a );
 a74681a <=( a74680a  and  a74673a );
 a74684a <=( A233  and  A232 );
 a74687a <=( (not A266)  and  (not A265) );
 a74688a <=( a74687a  and  a74684a );
 a74691a <=( (not A299)  and  A298 );
 a74694a <=( A302  and  A300 );
 a74695a <=( a74694a  and  a74691a );
 a74696a <=( a74695a  and  a74688a );
 a74700a <=( (not A168)  and  (not A169) );
 a74701a <=( (not A170)  and  a74700a );
 a74704a <=( (not A200)  and  A199 );
 a74707a <=( A203  and  A201 );
 a74708a <=( a74707a  and  a74704a );
 a74709a <=( a74708a  and  a74701a );
 a74712a <=( (not A235)  and  (not A233) );
 a74715a <=( (not A266)  and  (not A236) );
 a74716a <=( a74715a  and  a74712a );
 a74719a <=( (not A269)  and  (not A268) );
 a74722a <=( A299  and  (not A298) );
 a74723a <=( a74722a  and  a74719a );
 a74724a <=( a74723a  and  a74716a );
 a74728a <=( (not A168)  and  (not A169) );
 a74729a <=( (not A170)  and  a74728a );
 a74732a <=( (not A200)  and  A199 );
 a74735a <=( A203  and  A201 );
 a74736a <=( a74735a  and  a74732a );
 a74737a <=( a74736a  and  a74729a );
 a74740a <=( (not A234)  and  (not A233) );
 a74743a <=( A266  and  A265 );
 a74744a <=( a74743a  and  a74740a );
 a74747a <=( (not A299)  and  A298 );
 a74750a <=( A301  and  A300 );
 a74751a <=( a74750a  and  a74747a );
 a74752a <=( a74751a  and  a74744a );
 a74756a <=( (not A168)  and  (not A169) );
 a74757a <=( (not A170)  and  a74756a );
 a74760a <=( (not A200)  and  A199 );
 a74763a <=( A203  and  A201 );
 a74764a <=( a74763a  and  a74760a );
 a74765a <=( a74764a  and  a74757a );
 a74768a <=( (not A234)  and  (not A233) );
 a74771a <=( A266  and  A265 );
 a74772a <=( a74771a  and  a74768a );
 a74775a <=( (not A299)  and  A298 );
 a74778a <=( A302  and  A300 );
 a74779a <=( a74778a  and  a74775a );
 a74780a <=( a74779a  and  a74772a );
 a74784a <=( (not A168)  and  (not A169) );
 a74785a <=( (not A170)  and  a74784a );
 a74788a <=( (not A200)  and  A199 );
 a74791a <=( A203  and  A201 );
 a74792a <=( a74791a  and  a74788a );
 a74793a <=( a74792a  and  a74785a );
 a74796a <=( (not A234)  and  (not A233) );
 a74799a <=( (not A267)  and  (not A266) );
 a74800a <=( a74799a  and  a74796a );
 a74803a <=( (not A299)  and  A298 );
 a74806a <=( A301  and  A300 );
 a74807a <=( a74806a  and  a74803a );
 a74808a <=( a74807a  and  a74800a );
 a74812a <=( (not A168)  and  (not A169) );
 a74813a <=( (not A170)  and  a74812a );
 a74816a <=( (not A200)  and  A199 );
 a74819a <=( A203  and  A201 );
 a74820a <=( a74819a  and  a74816a );
 a74821a <=( a74820a  and  a74813a );
 a74824a <=( (not A234)  and  (not A233) );
 a74827a <=( (not A267)  and  (not A266) );
 a74828a <=( a74827a  and  a74824a );
 a74831a <=( (not A299)  and  A298 );
 a74834a <=( A302  and  A300 );
 a74835a <=( a74834a  and  a74831a );
 a74836a <=( a74835a  and  a74828a );
 a74840a <=( (not A168)  and  (not A169) );
 a74841a <=( (not A170)  and  a74840a );
 a74844a <=( (not A200)  and  A199 );
 a74847a <=( A203  and  A201 );
 a74848a <=( a74847a  and  a74844a );
 a74849a <=( a74848a  and  a74841a );
 a74852a <=( (not A234)  and  (not A233) );
 a74855a <=( (not A266)  and  (not A265) );
 a74856a <=( a74855a  and  a74852a );
 a74859a <=( (not A299)  and  A298 );
 a74862a <=( A301  and  A300 );
 a74863a <=( a74862a  and  a74859a );
 a74864a <=( a74863a  and  a74856a );
 a74868a <=( (not A168)  and  (not A169) );
 a74869a <=( (not A170)  and  a74868a );
 a74872a <=( (not A200)  and  A199 );
 a74875a <=( A203  and  A201 );
 a74876a <=( a74875a  and  a74872a );
 a74877a <=( a74876a  and  a74869a );
 a74880a <=( (not A234)  and  (not A233) );
 a74883a <=( (not A266)  and  (not A265) );
 a74884a <=( a74883a  and  a74880a );
 a74887a <=( (not A299)  and  A298 );
 a74890a <=( A302  and  A300 );
 a74891a <=( a74890a  and  a74887a );
 a74892a <=( a74891a  and  a74884a );
 a74896a <=( (not A168)  and  (not A169) );
 a74897a <=( (not A170)  and  a74896a );
 a74900a <=( (not A200)  and  A199 );
 a74903a <=( A203  and  A201 );
 a74904a <=( a74903a  and  a74900a );
 a74905a <=( a74904a  and  a74897a );
 a74908a <=( (not A233)  and  A232 );
 a74911a <=( A235  and  A234 );
 a74912a <=( a74911a  and  a74908a );
 a74915a <=( (not A266)  and  A265 );
 a74918a <=( A268  and  A267 );
 a74919a <=( a74918a  and  a74915a );
 a74920a <=( a74919a  and  a74912a );
 a74924a <=( (not A168)  and  (not A169) );
 a74925a <=( (not A170)  and  a74924a );
 a74928a <=( (not A200)  and  A199 );
 a74931a <=( A203  and  A201 );
 a74932a <=( a74931a  and  a74928a );
 a74933a <=( a74932a  and  a74925a );
 a74936a <=( (not A233)  and  A232 );
 a74939a <=( A235  and  A234 );
 a74940a <=( a74939a  and  a74936a );
 a74943a <=( (not A266)  and  A265 );
 a74946a <=( A269  and  A267 );
 a74947a <=( a74946a  and  a74943a );
 a74948a <=( a74947a  and  a74940a );
 a74952a <=( (not A168)  and  (not A169) );
 a74953a <=( (not A170)  and  a74952a );
 a74956a <=( (not A200)  and  A199 );
 a74959a <=( A203  and  A201 );
 a74960a <=( a74959a  and  a74956a );
 a74961a <=( a74960a  and  a74953a );
 a74964a <=( (not A233)  and  A232 );
 a74967a <=( A236  and  A234 );
 a74968a <=( a74967a  and  a74964a );
 a74971a <=( (not A266)  and  A265 );
 a74974a <=( A268  and  A267 );
 a74975a <=( a74974a  and  a74971a );
 a74976a <=( a74975a  and  a74968a );
 a74980a <=( (not A168)  and  (not A169) );
 a74981a <=( (not A170)  and  a74980a );
 a74984a <=( (not A200)  and  A199 );
 a74987a <=( A203  and  A201 );
 a74988a <=( a74987a  and  a74984a );
 a74989a <=( a74988a  and  a74981a );
 a74992a <=( (not A233)  and  A232 );
 a74995a <=( A236  and  A234 );
 a74996a <=( a74995a  and  a74992a );
 a74999a <=( (not A266)  and  A265 );
 a75002a <=( A269  and  A267 );
 a75003a <=( a75002a  and  a74999a );
 a75004a <=( a75003a  and  a74996a );
 a75008a <=( (not A168)  and  (not A169) );
 a75009a <=( (not A170)  and  a75008a );
 a75012a <=( (not A200)  and  A199 );
 a75015a <=( A203  and  A201 );
 a75016a <=( a75015a  and  a75012a );
 a75017a <=( a75016a  and  a75009a );
 a75020a <=( (not A233)  and  (not A232) );
 a75023a <=( A266  and  A265 );
 a75024a <=( a75023a  and  a75020a );
 a75027a <=( (not A299)  and  A298 );
 a75030a <=( A301  and  A300 );
 a75031a <=( a75030a  and  a75027a );
 a75032a <=( a75031a  and  a75024a );
 a75036a <=( (not A168)  and  (not A169) );
 a75037a <=( (not A170)  and  a75036a );
 a75040a <=( (not A200)  and  A199 );
 a75043a <=( A203  and  A201 );
 a75044a <=( a75043a  and  a75040a );
 a75045a <=( a75044a  and  a75037a );
 a75048a <=( (not A233)  and  (not A232) );
 a75051a <=( A266  and  A265 );
 a75052a <=( a75051a  and  a75048a );
 a75055a <=( (not A299)  and  A298 );
 a75058a <=( A302  and  A300 );
 a75059a <=( a75058a  and  a75055a );
 a75060a <=( a75059a  and  a75052a );
 a75064a <=( (not A168)  and  (not A169) );
 a75065a <=( (not A170)  and  a75064a );
 a75068a <=( (not A200)  and  A199 );
 a75071a <=( A203  and  A201 );
 a75072a <=( a75071a  and  a75068a );
 a75073a <=( a75072a  and  a75065a );
 a75076a <=( (not A233)  and  (not A232) );
 a75079a <=( (not A267)  and  (not A266) );
 a75080a <=( a75079a  and  a75076a );
 a75083a <=( (not A299)  and  A298 );
 a75086a <=( A301  and  A300 );
 a75087a <=( a75086a  and  a75083a );
 a75088a <=( a75087a  and  a75080a );
 a75092a <=( (not A168)  and  (not A169) );
 a75093a <=( (not A170)  and  a75092a );
 a75096a <=( (not A200)  and  A199 );
 a75099a <=( A203  and  A201 );
 a75100a <=( a75099a  and  a75096a );
 a75101a <=( a75100a  and  a75093a );
 a75104a <=( (not A233)  and  (not A232) );
 a75107a <=( (not A267)  and  (not A266) );
 a75108a <=( a75107a  and  a75104a );
 a75111a <=( (not A299)  and  A298 );
 a75114a <=( A302  and  A300 );
 a75115a <=( a75114a  and  a75111a );
 a75116a <=( a75115a  and  a75108a );
 a75120a <=( (not A168)  and  (not A169) );
 a75121a <=( (not A170)  and  a75120a );
 a75124a <=( (not A200)  and  A199 );
 a75127a <=( A203  and  A201 );
 a75128a <=( a75127a  and  a75124a );
 a75129a <=( a75128a  and  a75121a );
 a75132a <=( (not A233)  and  (not A232) );
 a75135a <=( (not A266)  and  (not A265) );
 a75136a <=( a75135a  and  a75132a );
 a75139a <=( (not A299)  and  A298 );
 a75142a <=( A301  and  A300 );
 a75143a <=( a75142a  and  a75139a );
 a75144a <=( a75143a  and  a75136a );
 a75148a <=( (not A168)  and  (not A169) );
 a75149a <=( (not A170)  and  a75148a );
 a75152a <=( (not A200)  and  A199 );
 a75155a <=( A203  and  A201 );
 a75156a <=( a75155a  and  a75152a );
 a75157a <=( a75156a  and  a75149a );
 a75160a <=( (not A233)  and  (not A232) );
 a75163a <=( (not A266)  and  (not A265) );
 a75164a <=( a75163a  and  a75160a );
 a75167a <=( (not A299)  and  A298 );
 a75170a <=( A302  and  A300 );
 a75171a <=( a75170a  and  a75167a );
 a75172a <=( a75171a  and  a75164a );
 a75175a <=( (not A167)  and  A170 );
 a75178a <=( A199  and  (not A166) );
 a75179a <=( a75178a  and  a75175a );
 a75182a <=( A201  and  (not A200) );
 a75185a <=( A232  and  A202 );
 a75186a <=( a75185a  and  a75182a );
 a75187a <=( a75186a  and  a75179a );
 a75190a <=( A265  and  A233 );
 a75193a <=( (not A269)  and  (not A268) );
 a75194a <=( a75193a  and  a75190a );
 a75197a <=( (not A299)  and  A298 );
 a75200a <=( A301  and  A300 );
 a75201a <=( a75200a  and  a75197a );
 a75202a <=( a75201a  and  a75194a );
 a75205a <=( (not A167)  and  A170 );
 a75208a <=( A199  and  (not A166) );
 a75209a <=( a75208a  and  a75205a );
 a75212a <=( A201  and  (not A200) );
 a75215a <=( A232  and  A202 );
 a75216a <=( a75215a  and  a75212a );
 a75217a <=( a75216a  and  a75209a );
 a75220a <=( A265  and  A233 );
 a75223a <=( (not A269)  and  (not A268) );
 a75224a <=( a75223a  and  a75220a );
 a75227a <=( (not A299)  and  A298 );
 a75230a <=( A302  and  A300 );
 a75231a <=( a75230a  and  a75227a );
 a75232a <=( a75231a  and  a75224a );
 a75235a <=( (not A167)  and  A170 );
 a75238a <=( A199  and  (not A166) );
 a75239a <=( a75238a  and  a75235a );
 a75242a <=( A201  and  (not A200) );
 a75245a <=( (not A233)  and  A202 );
 a75246a <=( a75245a  and  a75242a );
 a75247a <=( a75246a  and  a75239a );
 a75250a <=( (not A236)  and  (not A235) );
 a75253a <=( A266  and  A265 );
 a75254a <=( a75253a  and  a75250a );
 a75257a <=( (not A299)  and  A298 );
 a75260a <=( A301  and  A300 );
 a75261a <=( a75260a  and  a75257a );
 a75262a <=( a75261a  and  a75254a );
 a75265a <=( (not A167)  and  A170 );
 a75268a <=( A199  and  (not A166) );
 a75269a <=( a75268a  and  a75265a );
 a75272a <=( A201  and  (not A200) );
 a75275a <=( (not A233)  and  A202 );
 a75276a <=( a75275a  and  a75272a );
 a75277a <=( a75276a  and  a75269a );
 a75280a <=( (not A236)  and  (not A235) );
 a75283a <=( A266  and  A265 );
 a75284a <=( a75283a  and  a75280a );
 a75287a <=( (not A299)  and  A298 );
 a75290a <=( A302  and  A300 );
 a75291a <=( a75290a  and  a75287a );
 a75292a <=( a75291a  and  a75284a );
 a75295a <=( (not A167)  and  A170 );
 a75298a <=( A199  and  (not A166) );
 a75299a <=( a75298a  and  a75295a );
 a75302a <=( A201  and  (not A200) );
 a75305a <=( (not A233)  and  A202 );
 a75306a <=( a75305a  and  a75302a );
 a75307a <=( a75306a  and  a75299a );
 a75310a <=( (not A236)  and  (not A235) );
 a75313a <=( (not A267)  and  (not A266) );
 a75314a <=( a75313a  and  a75310a );
 a75317a <=( (not A299)  and  A298 );
 a75320a <=( A301  and  A300 );
 a75321a <=( a75320a  and  a75317a );
 a75322a <=( a75321a  and  a75314a );
 a75325a <=( (not A167)  and  A170 );
 a75328a <=( A199  and  (not A166) );
 a75329a <=( a75328a  and  a75325a );
 a75332a <=( A201  and  (not A200) );
 a75335a <=( (not A233)  and  A202 );
 a75336a <=( a75335a  and  a75332a );
 a75337a <=( a75336a  and  a75329a );
 a75340a <=( (not A236)  and  (not A235) );
 a75343a <=( (not A267)  and  (not A266) );
 a75344a <=( a75343a  and  a75340a );
 a75347a <=( (not A299)  and  A298 );
 a75350a <=( A302  and  A300 );
 a75351a <=( a75350a  and  a75347a );
 a75352a <=( a75351a  and  a75344a );
 a75355a <=( (not A167)  and  A170 );
 a75358a <=( A199  and  (not A166) );
 a75359a <=( a75358a  and  a75355a );
 a75362a <=( A201  and  (not A200) );
 a75365a <=( (not A233)  and  A202 );
 a75366a <=( a75365a  and  a75362a );
 a75367a <=( a75366a  and  a75359a );
 a75370a <=( (not A236)  and  (not A235) );
 a75373a <=( (not A266)  and  (not A265) );
 a75374a <=( a75373a  and  a75370a );
 a75377a <=( (not A299)  and  A298 );
 a75380a <=( A301  and  A300 );
 a75381a <=( a75380a  and  a75377a );
 a75382a <=( a75381a  and  a75374a );
 a75385a <=( (not A167)  and  A170 );
 a75388a <=( A199  and  (not A166) );
 a75389a <=( a75388a  and  a75385a );
 a75392a <=( A201  and  (not A200) );
 a75395a <=( (not A233)  and  A202 );
 a75396a <=( a75395a  and  a75392a );
 a75397a <=( a75396a  and  a75389a );
 a75400a <=( (not A236)  and  (not A235) );
 a75403a <=( (not A266)  and  (not A265) );
 a75404a <=( a75403a  and  a75400a );
 a75407a <=( (not A299)  and  A298 );
 a75410a <=( A302  and  A300 );
 a75411a <=( a75410a  and  a75407a );
 a75412a <=( a75411a  and  a75404a );
 a75415a <=( (not A167)  and  A170 );
 a75418a <=( A199  and  (not A166) );
 a75419a <=( a75418a  and  a75415a );
 a75422a <=( A201  and  (not A200) );
 a75425a <=( (not A233)  and  A202 );
 a75426a <=( a75425a  and  a75422a );
 a75427a <=( a75426a  and  a75419a );
 a75430a <=( (not A266)  and  (not A234) );
 a75433a <=( (not A269)  and  (not A268) );
 a75434a <=( a75433a  and  a75430a );
 a75437a <=( (not A299)  and  A298 );
 a75440a <=( A301  and  A300 );
 a75441a <=( a75440a  and  a75437a );
 a75442a <=( a75441a  and  a75434a );
 a75445a <=( (not A167)  and  A170 );
 a75448a <=( A199  and  (not A166) );
 a75449a <=( a75448a  and  a75445a );
 a75452a <=( A201  and  (not A200) );
 a75455a <=( (not A233)  and  A202 );
 a75456a <=( a75455a  and  a75452a );
 a75457a <=( a75456a  and  a75449a );
 a75460a <=( (not A266)  and  (not A234) );
 a75463a <=( (not A269)  and  (not A268) );
 a75464a <=( a75463a  and  a75460a );
 a75467a <=( (not A299)  and  A298 );
 a75470a <=( A302  and  A300 );
 a75471a <=( a75470a  and  a75467a );
 a75472a <=( a75471a  and  a75464a );
 a75475a <=( (not A167)  and  A170 );
 a75478a <=( A199  and  (not A166) );
 a75479a <=( a75478a  and  a75475a );
 a75482a <=( A201  and  (not A200) );
 a75485a <=( (not A232)  and  A202 );
 a75486a <=( a75485a  and  a75482a );
 a75487a <=( a75486a  and  a75479a );
 a75490a <=( (not A266)  and  (not A233) );
 a75493a <=( (not A269)  and  (not A268) );
 a75494a <=( a75493a  and  a75490a );
 a75497a <=( (not A299)  and  A298 );
 a75500a <=( A301  and  A300 );
 a75501a <=( a75500a  and  a75497a );
 a75502a <=( a75501a  and  a75494a );
 a75505a <=( (not A167)  and  A170 );
 a75508a <=( A199  and  (not A166) );
 a75509a <=( a75508a  and  a75505a );
 a75512a <=( A201  and  (not A200) );
 a75515a <=( (not A232)  and  A202 );
 a75516a <=( a75515a  and  a75512a );
 a75517a <=( a75516a  and  a75509a );
 a75520a <=( (not A266)  and  (not A233) );
 a75523a <=( (not A269)  and  (not A268) );
 a75524a <=( a75523a  and  a75520a );
 a75527a <=( (not A299)  and  A298 );
 a75530a <=( A302  and  A300 );
 a75531a <=( a75530a  and  a75527a );
 a75532a <=( a75531a  and  a75524a );
 a75535a <=( (not A167)  and  A170 );
 a75538a <=( A199  and  (not A166) );
 a75539a <=( a75538a  and  a75535a );
 a75542a <=( A201  and  (not A200) );
 a75545a <=( A232  and  A203 );
 a75546a <=( a75545a  and  a75542a );
 a75547a <=( a75546a  and  a75539a );
 a75550a <=( A265  and  A233 );
 a75553a <=( (not A269)  and  (not A268) );
 a75554a <=( a75553a  and  a75550a );
 a75557a <=( (not A299)  and  A298 );
 a75560a <=( A301  and  A300 );
 a75561a <=( a75560a  and  a75557a );
 a75562a <=( a75561a  and  a75554a );
 a75565a <=( (not A167)  and  A170 );
 a75568a <=( A199  and  (not A166) );
 a75569a <=( a75568a  and  a75565a );
 a75572a <=( A201  and  (not A200) );
 a75575a <=( A232  and  A203 );
 a75576a <=( a75575a  and  a75572a );
 a75577a <=( a75576a  and  a75569a );
 a75580a <=( A265  and  A233 );
 a75583a <=( (not A269)  and  (not A268) );
 a75584a <=( a75583a  and  a75580a );
 a75587a <=( (not A299)  and  A298 );
 a75590a <=( A302  and  A300 );
 a75591a <=( a75590a  and  a75587a );
 a75592a <=( a75591a  and  a75584a );
 a75595a <=( (not A167)  and  A170 );
 a75598a <=( A199  and  (not A166) );
 a75599a <=( a75598a  and  a75595a );
 a75602a <=( A201  and  (not A200) );
 a75605a <=( (not A233)  and  A203 );
 a75606a <=( a75605a  and  a75602a );
 a75607a <=( a75606a  and  a75599a );
 a75610a <=( (not A236)  and  (not A235) );
 a75613a <=( A266  and  A265 );
 a75614a <=( a75613a  and  a75610a );
 a75617a <=( (not A299)  and  A298 );
 a75620a <=( A301  and  A300 );
 a75621a <=( a75620a  and  a75617a );
 a75622a <=( a75621a  and  a75614a );
 a75625a <=( (not A167)  and  A170 );
 a75628a <=( A199  and  (not A166) );
 a75629a <=( a75628a  and  a75625a );
 a75632a <=( A201  and  (not A200) );
 a75635a <=( (not A233)  and  A203 );
 a75636a <=( a75635a  and  a75632a );
 a75637a <=( a75636a  and  a75629a );
 a75640a <=( (not A236)  and  (not A235) );
 a75643a <=( A266  and  A265 );
 a75644a <=( a75643a  and  a75640a );
 a75647a <=( (not A299)  and  A298 );
 a75650a <=( A302  and  A300 );
 a75651a <=( a75650a  and  a75647a );
 a75652a <=( a75651a  and  a75644a );
 a75655a <=( (not A167)  and  A170 );
 a75658a <=( A199  and  (not A166) );
 a75659a <=( a75658a  and  a75655a );
 a75662a <=( A201  and  (not A200) );
 a75665a <=( (not A233)  and  A203 );
 a75666a <=( a75665a  and  a75662a );
 a75667a <=( a75666a  and  a75659a );
 a75670a <=( (not A236)  and  (not A235) );
 a75673a <=( (not A267)  and  (not A266) );
 a75674a <=( a75673a  and  a75670a );
 a75677a <=( (not A299)  and  A298 );
 a75680a <=( A301  and  A300 );
 a75681a <=( a75680a  and  a75677a );
 a75682a <=( a75681a  and  a75674a );
 a75685a <=( (not A167)  and  A170 );
 a75688a <=( A199  and  (not A166) );
 a75689a <=( a75688a  and  a75685a );
 a75692a <=( A201  and  (not A200) );
 a75695a <=( (not A233)  and  A203 );
 a75696a <=( a75695a  and  a75692a );
 a75697a <=( a75696a  and  a75689a );
 a75700a <=( (not A236)  and  (not A235) );
 a75703a <=( (not A267)  and  (not A266) );
 a75704a <=( a75703a  and  a75700a );
 a75707a <=( (not A299)  and  A298 );
 a75710a <=( A302  and  A300 );
 a75711a <=( a75710a  and  a75707a );
 a75712a <=( a75711a  and  a75704a );
 a75715a <=( (not A167)  and  A170 );
 a75718a <=( A199  and  (not A166) );
 a75719a <=( a75718a  and  a75715a );
 a75722a <=( A201  and  (not A200) );
 a75725a <=( (not A233)  and  A203 );
 a75726a <=( a75725a  and  a75722a );
 a75727a <=( a75726a  and  a75719a );
 a75730a <=( (not A236)  and  (not A235) );
 a75733a <=( (not A266)  and  (not A265) );
 a75734a <=( a75733a  and  a75730a );
 a75737a <=( (not A299)  and  A298 );
 a75740a <=( A301  and  A300 );
 a75741a <=( a75740a  and  a75737a );
 a75742a <=( a75741a  and  a75734a );
 a75745a <=( (not A167)  and  A170 );
 a75748a <=( A199  and  (not A166) );
 a75749a <=( a75748a  and  a75745a );
 a75752a <=( A201  and  (not A200) );
 a75755a <=( (not A233)  and  A203 );
 a75756a <=( a75755a  and  a75752a );
 a75757a <=( a75756a  and  a75749a );
 a75760a <=( (not A236)  and  (not A235) );
 a75763a <=( (not A266)  and  (not A265) );
 a75764a <=( a75763a  and  a75760a );
 a75767a <=( (not A299)  and  A298 );
 a75770a <=( A302  and  A300 );
 a75771a <=( a75770a  and  a75767a );
 a75772a <=( a75771a  and  a75764a );
 a75775a <=( (not A167)  and  A170 );
 a75778a <=( A199  and  (not A166) );
 a75779a <=( a75778a  and  a75775a );
 a75782a <=( A201  and  (not A200) );
 a75785a <=( (not A233)  and  A203 );
 a75786a <=( a75785a  and  a75782a );
 a75787a <=( a75786a  and  a75779a );
 a75790a <=( (not A266)  and  (not A234) );
 a75793a <=( (not A269)  and  (not A268) );
 a75794a <=( a75793a  and  a75790a );
 a75797a <=( (not A299)  and  A298 );
 a75800a <=( A301  and  A300 );
 a75801a <=( a75800a  and  a75797a );
 a75802a <=( a75801a  and  a75794a );
 a75805a <=( (not A167)  and  A170 );
 a75808a <=( A199  and  (not A166) );
 a75809a <=( a75808a  and  a75805a );
 a75812a <=( A201  and  (not A200) );
 a75815a <=( (not A233)  and  A203 );
 a75816a <=( a75815a  and  a75812a );
 a75817a <=( a75816a  and  a75809a );
 a75820a <=( (not A266)  and  (not A234) );
 a75823a <=( (not A269)  and  (not A268) );
 a75824a <=( a75823a  and  a75820a );
 a75827a <=( (not A299)  and  A298 );
 a75830a <=( A302  and  A300 );
 a75831a <=( a75830a  and  a75827a );
 a75832a <=( a75831a  and  a75824a );
 a75835a <=( (not A167)  and  A170 );
 a75838a <=( A199  and  (not A166) );
 a75839a <=( a75838a  and  a75835a );
 a75842a <=( A201  and  (not A200) );
 a75845a <=( (not A232)  and  A203 );
 a75846a <=( a75845a  and  a75842a );
 a75847a <=( a75846a  and  a75839a );
 a75850a <=( (not A266)  and  (not A233) );
 a75853a <=( (not A269)  and  (not A268) );
 a75854a <=( a75853a  and  a75850a );
 a75857a <=( (not A299)  and  A298 );
 a75860a <=( A301  and  A300 );
 a75861a <=( a75860a  and  a75857a );
 a75862a <=( a75861a  and  a75854a );
 a75865a <=( (not A167)  and  A170 );
 a75868a <=( A199  and  (not A166) );
 a75869a <=( a75868a  and  a75865a );
 a75872a <=( A201  and  (not A200) );
 a75875a <=( (not A232)  and  A203 );
 a75876a <=( a75875a  and  a75872a );
 a75877a <=( a75876a  and  a75869a );
 a75880a <=( (not A266)  and  (not A233) );
 a75883a <=( (not A269)  and  (not A268) );
 a75884a <=( a75883a  and  a75880a );
 a75887a <=( (not A299)  and  A298 );
 a75890a <=( A302  and  A300 );
 a75891a <=( a75890a  and  a75887a );
 a75892a <=( a75891a  and  a75884a );
 a75895a <=( (not A168)  and  A170 );
 a75898a <=( A166  and  A167 );
 a75899a <=( a75898a  and  a75895a );
 a75902a <=( A200  and  (not A199) );
 a75905a <=( (not A235)  and  (not A233) );
 a75906a <=( a75905a  and  a75902a );
 a75907a <=( a75906a  and  a75899a );
 a75910a <=( (not A266)  and  (not A236) );
 a75913a <=( (not A269)  and  (not A268) );
 a75914a <=( a75913a  and  a75910a );
 a75917a <=( (not A299)  and  A298 );
 a75920a <=( A301  and  A300 );
 a75921a <=( a75920a  and  a75917a );
 a75922a <=( a75921a  and  a75914a );
 a75925a <=( (not A168)  and  A170 );
 a75928a <=( A166  and  A167 );
 a75929a <=( a75928a  and  a75925a );
 a75932a <=( A200  and  (not A199) );
 a75935a <=( (not A235)  and  (not A233) );
 a75936a <=( a75935a  and  a75932a );
 a75937a <=( a75936a  and  a75929a );
 a75940a <=( (not A266)  and  (not A236) );
 a75943a <=( (not A269)  and  (not A268) );
 a75944a <=( a75943a  and  a75940a );
 a75947a <=( (not A299)  and  A298 );
 a75950a <=( A302  and  A300 );
 a75951a <=( a75950a  and  a75947a );
 a75952a <=( a75951a  and  a75944a );
 a75955a <=( (not A168)  and  (not A170) );
 a75958a <=( (not A166)  and  A167 );
 a75959a <=( a75958a  and  a75955a );
 a75962a <=( A200  and  (not A199) );
 a75965a <=( (not A235)  and  (not A233) );
 a75966a <=( a75965a  and  a75962a );
 a75967a <=( a75966a  and  a75959a );
 a75970a <=( (not A266)  and  (not A236) );
 a75973a <=( (not A269)  and  (not A268) );
 a75974a <=( a75973a  and  a75970a );
 a75977a <=( (not A299)  and  A298 );
 a75980a <=( A301  and  A300 );
 a75981a <=( a75980a  and  a75977a );
 a75982a <=( a75981a  and  a75974a );
 a75985a <=( (not A168)  and  (not A170) );
 a75988a <=( (not A166)  and  A167 );
 a75989a <=( a75988a  and  a75985a );
 a75992a <=( A200  and  (not A199) );
 a75995a <=( (not A235)  and  (not A233) );
 a75996a <=( a75995a  and  a75992a );
 a75997a <=( a75996a  and  a75989a );
 a76000a <=( (not A266)  and  (not A236) );
 a76003a <=( (not A269)  and  (not A268) );
 a76004a <=( a76003a  and  a76000a );
 a76007a <=( (not A299)  and  A298 );
 a76010a <=( A302  and  A300 );
 a76011a <=( a76010a  and  a76007a );
 a76012a <=( a76011a  and  a76004a );
 a76015a <=( (not A168)  and  (not A170) );
 a76018a <=( A166  and  (not A167) );
 a76019a <=( a76018a  and  a76015a );
 a76022a <=( A200  and  (not A199) );
 a76025a <=( (not A235)  and  (not A233) );
 a76026a <=( a76025a  and  a76022a );
 a76027a <=( a76026a  and  a76019a );
 a76030a <=( (not A266)  and  (not A236) );
 a76033a <=( (not A269)  and  (not A268) );
 a76034a <=( a76033a  and  a76030a );
 a76037a <=( (not A299)  and  A298 );
 a76040a <=( A301  and  A300 );
 a76041a <=( a76040a  and  a76037a );
 a76042a <=( a76041a  and  a76034a );
 a76045a <=( (not A168)  and  (not A170) );
 a76048a <=( A166  and  (not A167) );
 a76049a <=( a76048a  and  a76045a );
 a76052a <=( A200  and  (not A199) );
 a76055a <=( (not A235)  and  (not A233) );
 a76056a <=( a76055a  and  a76052a );
 a76057a <=( a76056a  and  a76049a );
 a76060a <=( (not A266)  and  (not A236) );
 a76063a <=( (not A269)  and  (not A268) );
 a76064a <=( a76063a  and  a76060a );
 a76067a <=( (not A299)  and  A298 );
 a76070a <=( A302  and  A300 );
 a76071a <=( a76070a  and  a76067a );
 a76072a <=( a76071a  and  a76064a );
 a76075a <=( (not A168)  and  A169 );
 a76078a <=( (not A166)  and  A167 );
 a76079a <=( a76078a  and  a76075a );
 a76082a <=( A200  and  (not A199) );
 a76085a <=( (not A235)  and  (not A233) );
 a76086a <=( a76085a  and  a76082a );
 a76087a <=( a76086a  and  a76079a );
 a76090a <=( (not A266)  and  (not A236) );
 a76093a <=( (not A269)  and  (not A268) );
 a76094a <=( a76093a  and  a76090a );
 a76097a <=( (not A299)  and  A298 );
 a76100a <=( A301  and  A300 );
 a76101a <=( a76100a  and  a76097a );
 a76102a <=( a76101a  and  a76094a );
 a76105a <=( (not A168)  and  A169 );
 a76108a <=( (not A166)  and  A167 );
 a76109a <=( a76108a  and  a76105a );
 a76112a <=( A200  and  (not A199) );
 a76115a <=( (not A235)  and  (not A233) );
 a76116a <=( a76115a  and  a76112a );
 a76117a <=( a76116a  and  a76109a );
 a76120a <=( (not A266)  and  (not A236) );
 a76123a <=( (not A269)  and  (not A268) );
 a76124a <=( a76123a  and  a76120a );
 a76127a <=( (not A299)  and  A298 );
 a76130a <=( A302  and  A300 );
 a76131a <=( a76130a  and  a76127a );
 a76132a <=( a76131a  and  a76124a );
 a76135a <=( (not A168)  and  A169 );
 a76138a <=( (not A166)  and  A167 );
 a76139a <=( a76138a  and  a76135a );
 a76142a <=( (not A200)  and  A199 );
 a76145a <=( A202  and  A201 );
 a76146a <=( a76145a  and  a76142a );
 a76147a <=( a76146a  and  a76139a );
 a76150a <=( A233  and  A232 );
 a76153a <=( (not A267)  and  A265 );
 a76154a <=( a76153a  and  a76150a );
 a76157a <=( (not A299)  and  A298 );
 a76160a <=( A301  and  A300 );
 a76161a <=( a76160a  and  a76157a );
 a76162a <=( a76161a  and  a76154a );
 a76165a <=( (not A168)  and  A169 );
 a76168a <=( (not A166)  and  A167 );
 a76169a <=( a76168a  and  a76165a );
 a76172a <=( (not A200)  and  A199 );
 a76175a <=( A202  and  A201 );
 a76176a <=( a76175a  and  a76172a );
 a76177a <=( a76176a  and  a76169a );
 a76180a <=( A233  and  A232 );
 a76183a <=( (not A267)  and  A265 );
 a76184a <=( a76183a  and  a76180a );
 a76187a <=( (not A299)  and  A298 );
 a76190a <=( A302  and  A300 );
 a76191a <=( a76190a  and  a76187a );
 a76192a <=( a76191a  and  a76184a );
 a76195a <=( (not A168)  and  A169 );
 a76198a <=( (not A166)  and  A167 );
 a76199a <=( a76198a  and  a76195a );
 a76202a <=( (not A200)  and  A199 );
 a76205a <=( A202  and  A201 );
 a76206a <=( a76205a  and  a76202a );
 a76207a <=( a76206a  and  a76199a );
 a76210a <=( A233  and  A232 );
 a76213a <=( A266  and  A265 );
 a76214a <=( a76213a  and  a76210a );
 a76217a <=( (not A299)  and  A298 );
 a76220a <=( A301  and  A300 );
 a76221a <=( a76220a  and  a76217a );
 a76222a <=( a76221a  and  a76214a );
 a76225a <=( (not A168)  and  A169 );
 a76228a <=( (not A166)  and  A167 );
 a76229a <=( a76228a  and  a76225a );
 a76232a <=( (not A200)  and  A199 );
 a76235a <=( A202  and  A201 );
 a76236a <=( a76235a  and  a76232a );
 a76237a <=( a76236a  and  a76229a );
 a76240a <=( A233  and  A232 );
 a76243a <=( A266  and  A265 );
 a76244a <=( a76243a  and  a76240a );
 a76247a <=( (not A299)  and  A298 );
 a76250a <=( A302  and  A300 );
 a76251a <=( a76250a  and  a76247a );
 a76252a <=( a76251a  and  a76244a );
 a76255a <=( (not A168)  and  A169 );
 a76258a <=( (not A166)  and  A167 );
 a76259a <=( a76258a  and  a76255a );
 a76262a <=( (not A200)  and  A199 );
 a76265a <=( A202  and  A201 );
 a76266a <=( a76265a  and  a76262a );
 a76267a <=( a76266a  and  a76259a );
 a76270a <=( A233  and  A232 );
 a76273a <=( (not A266)  and  (not A265) );
 a76274a <=( a76273a  and  a76270a );
 a76277a <=( (not A299)  and  A298 );
 a76280a <=( A301  and  A300 );
 a76281a <=( a76280a  and  a76277a );
 a76282a <=( a76281a  and  a76274a );
 a76285a <=( (not A168)  and  A169 );
 a76288a <=( (not A166)  and  A167 );
 a76289a <=( a76288a  and  a76285a );
 a76292a <=( (not A200)  and  A199 );
 a76295a <=( A202  and  A201 );
 a76296a <=( a76295a  and  a76292a );
 a76297a <=( a76296a  and  a76289a );
 a76300a <=( A233  and  A232 );
 a76303a <=( (not A266)  and  (not A265) );
 a76304a <=( a76303a  and  a76300a );
 a76307a <=( (not A299)  and  A298 );
 a76310a <=( A302  and  A300 );
 a76311a <=( a76310a  and  a76307a );
 a76312a <=( a76311a  and  a76304a );
 a76315a <=( (not A168)  and  A169 );
 a76318a <=( (not A166)  and  A167 );
 a76319a <=( a76318a  and  a76315a );
 a76322a <=( (not A200)  and  A199 );
 a76325a <=( A202  and  A201 );
 a76326a <=( a76325a  and  a76322a );
 a76327a <=( a76326a  and  a76319a );
 a76330a <=( (not A235)  and  (not A233) );
 a76333a <=( (not A266)  and  (not A236) );
 a76334a <=( a76333a  and  a76330a );
 a76337a <=( (not A269)  and  (not A268) );
 a76340a <=( A299  and  (not A298) );
 a76341a <=( a76340a  and  a76337a );
 a76342a <=( a76341a  and  a76334a );
 a76345a <=( (not A168)  and  A169 );
 a76348a <=( (not A166)  and  A167 );
 a76349a <=( a76348a  and  a76345a );
 a76352a <=( (not A200)  and  A199 );
 a76355a <=( A202  and  A201 );
 a76356a <=( a76355a  and  a76352a );
 a76357a <=( a76356a  and  a76349a );
 a76360a <=( (not A234)  and  (not A233) );
 a76363a <=( A266  and  A265 );
 a76364a <=( a76363a  and  a76360a );
 a76367a <=( (not A299)  and  A298 );
 a76370a <=( A301  and  A300 );
 a76371a <=( a76370a  and  a76367a );
 a76372a <=( a76371a  and  a76364a );
 a76375a <=( (not A168)  and  A169 );
 a76378a <=( (not A166)  and  A167 );
 a76379a <=( a76378a  and  a76375a );
 a76382a <=( (not A200)  and  A199 );
 a76385a <=( A202  and  A201 );
 a76386a <=( a76385a  and  a76382a );
 a76387a <=( a76386a  and  a76379a );
 a76390a <=( (not A234)  and  (not A233) );
 a76393a <=( A266  and  A265 );
 a76394a <=( a76393a  and  a76390a );
 a76397a <=( (not A299)  and  A298 );
 a76400a <=( A302  and  A300 );
 a76401a <=( a76400a  and  a76397a );
 a76402a <=( a76401a  and  a76394a );
 a76405a <=( (not A168)  and  A169 );
 a76408a <=( (not A166)  and  A167 );
 a76409a <=( a76408a  and  a76405a );
 a76412a <=( (not A200)  and  A199 );
 a76415a <=( A202  and  A201 );
 a76416a <=( a76415a  and  a76412a );
 a76417a <=( a76416a  and  a76409a );
 a76420a <=( (not A234)  and  (not A233) );
 a76423a <=( (not A267)  and  (not A266) );
 a76424a <=( a76423a  and  a76420a );
 a76427a <=( (not A299)  and  A298 );
 a76430a <=( A301  and  A300 );
 a76431a <=( a76430a  and  a76427a );
 a76432a <=( a76431a  and  a76424a );
 a76435a <=( (not A168)  and  A169 );
 a76438a <=( (not A166)  and  A167 );
 a76439a <=( a76438a  and  a76435a );
 a76442a <=( (not A200)  and  A199 );
 a76445a <=( A202  and  A201 );
 a76446a <=( a76445a  and  a76442a );
 a76447a <=( a76446a  and  a76439a );
 a76450a <=( (not A234)  and  (not A233) );
 a76453a <=( (not A267)  and  (not A266) );
 a76454a <=( a76453a  and  a76450a );
 a76457a <=( (not A299)  and  A298 );
 a76460a <=( A302  and  A300 );
 a76461a <=( a76460a  and  a76457a );
 a76462a <=( a76461a  and  a76454a );
 a76465a <=( (not A168)  and  A169 );
 a76468a <=( (not A166)  and  A167 );
 a76469a <=( a76468a  and  a76465a );
 a76472a <=( (not A200)  and  A199 );
 a76475a <=( A202  and  A201 );
 a76476a <=( a76475a  and  a76472a );
 a76477a <=( a76476a  and  a76469a );
 a76480a <=( (not A234)  and  (not A233) );
 a76483a <=( (not A266)  and  (not A265) );
 a76484a <=( a76483a  and  a76480a );
 a76487a <=( (not A299)  and  A298 );
 a76490a <=( A301  and  A300 );
 a76491a <=( a76490a  and  a76487a );
 a76492a <=( a76491a  and  a76484a );
 a76495a <=( (not A168)  and  A169 );
 a76498a <=( (not A166)  and  A167 );
 a76499a <=( a76498a  and  a76495a );
 a76502a <=( (not A200)  and  A199 );
 a76505a <=( A202  and  A201 );
 a76506a <=( a76505a  and  a76502a );
 a76507a <=( a76506a  and  a76499a );
 a76510a <=( (not A234)  and  (not A233) );
 a76513a <=( (not A266)  and  (not A265) );
 a76514a <=( a76513a  and  a76510a );
 a76517a <=( (not A299)  and  A298 );
 a76520a <=( A302  and  A300 );
 a76521a <=( a76520a  and  a76517a );
 a76522a <=( a76521a  and  a76514a );
 a76525a <=( (not A168)  and  A169 );
 a76528a <=( (not A166)  and  A167 );
 a76529a <=( a76528a  and  a76525a );
 a76532a <=( (not A200)  and  A199 );
 a76535a <=( A202  and  A201 );
 a76536a <=( a76535a  and  a76532a );
 a76537a <=( a76536a  and  a76529a );
 a76540a <=( (not A233)  and  A232 );
 a76543a <=( A235  and  A234 );
 a76544a <=( a76543a  and  a76540a );
 a76547a <=( (not A266)  and  A265 );
 a76550a <=( A268  and  A267 );
 a76551a <=( a76550a  and  a76547a );
 a76552a <=( a76551a  and  a76544a );
 a76555a <=( (not A168)  and  A169 );
 a76558a <=( (not A166)  and  A167 );
 a76559a <=( a76558a  and  a76555a );
 a76562a <=( (not A200)  and  A199 );
 a76565a <=( A202  and  A201 );
 a76566a <=( a76565a  and  a76562a );
 a76567a <=( a76566a  and  a76559a );
 a76570a <=( (not A233)  and  A232 );
 a76573a <=( A235  and  A234 );
 a76574a <=( a76573a  and  a76570a );
 a76577a <=( (not A266)  and  A265 );
 a76580a <=( A269  and  A267 );
 a76581a <=( a76580a  and  a76577a );
 a76582a <=( a76581a  and  a76574a );
 a76585a <=( (not A168)  and  A169 );
 a76588a <=( (not A166)  and  A167 );
 a76589a <=( a76588a  and  a76585a );
 a76592a <=( (not A200)  and  A199 );
 a76595a <=( A202  and  A201 );
 a76596a <=( a76595a  and  a76592a );
 a76597a <=( a76596a  and  a76589a );
 a76600a <=( (not A233)  and  A232 );
 a76603a <=( A236  and  A234 );
 a76604a <=( a76603a  and  a76600a );
 a76607a <=( (not A266)  and  A265 );
 a76610a <=( A268  and  A267 );
 a76611a <=( a76610a  and  a76607a );
 a76612a <=( a76611a  and  a76604a );
 a76615a <=( (not A168)  and  A169 );
 a76618a <=( (not A166)  and  A167 );
 a76619a <=( a76618a  and  a76615a );
 a76622a <=( (not A200)  and  A199 );
 a76625a <=( A202  and  A201 );
 a76626a <=( a76625a  and  a76622a );
 a76627a <=( a76626a  and  a76619a );
 a76630a <=( (not A233)  and  A232 );
 a76633a <=( A236  and  A234 );
 a76634a <=( a76633a  and  a76630a );
 a76637a <=( (not A266)  and  A265 );
 a76640a <=( A269  and  A267 );
 a76641a <=( a76640a  and  a76637a );
 a76642a <=( a76641a  and  a76634a );
 a76645a <=( (not A168)  and  A169 );
 a76648a <=( (not A166)  and  A167 );
 a76649a <=( a76648a  and  a76645a );
 a76652a <=( (not A200)  and  A199 );
 a76655a <=( A202  and  A201 );
 a76656a <=( a76655a  and  a76652a );
 a76657a <=( a76656a  and  a76649a );
 a76660a <=( (not A233)  and  (not A232) );
 a76663a <=( A266  and  A265 );
 a76664a <=( a76663a  and  a76660a );
 a76667a <=( (not A299)  and  A298 );
 a76670a <=( A301  and  A300 );
 a76671a <=( a76670a  and  a76667a );
 a76672a <=( a76671a  and  a76664a );
 a76675a <=( (not A168)  and  A169 );
 a76678a <=( (not A166)  and  A167 );
 a76679a <=( a76678a  and  a76675a );
 a76682a <=( (not A200)  and  A199 );
 a76685a <=( A202  and  A201 );
 a76686a <=( a76685a  and  a76682a );
 a76687a <=( a76686a  and  a76679a );
 a76690a <=( (not A233)  and  (not A232) );
 a76693a <=( A266  and  A265 );
 a76694a <=( a76693a  and  a76690a );
 a76697a <=( (not A299)  and  A298 );
 a76700a <=( A302  and  A300 );
 a76701a <=( a76700a  and  a76697a );
 a76702a <=( a76701a  and  a76694a );
 a76705a <=( (not A168)  and  A169 );
 a76708a <=( (not A166)  and  A167 );
 a76709a <=( a76708a  and  a76705a );
 a76712a <=( (not A200)  and  A199 );
 a76715a <=( A202  and  A201 );
 a76716a <=( a76715a  and  a76712a );
 a76717a <=( a76716a  and  a76709a );
 a76720a <=( (not A233)  and  (not A232) );
 a76723a <=( (not A267)  and  (not A266) );
 a76724a <=( a76723a  and  a76720a );
 a76727a <=( (not A299)  and  A298 );
 a76730a <=( A301  and  A300 );
 a76731a <=( a76730a  and  a76727a );
 a76732a <=( a76731a  and  a76724a );
 a76735a <=( (not A168)  and  A169 );
 a76738a <=( (not A166)  and  A167 );
 a76739a <=( a76738a  and  a76735a );
 a76742a <=( (not A200)  and  A199 );
 a76745a <=( A202  and  A201 );
 a76746a <=( a76745a  and  a76742a );
 a76747a <=( a76746a  and  a76739a );
 a76750a <=( (not A233)  and  (not A232) );
 a76753a <=( (not A267)  and  (not A266) );
 a76754a <=( a76753a  and  a76750a );
 a76757a <=( (not A299)  and  A298 );
 a76760a <=( A302  and  A300 );
 a76761a <=( a76760a  and  a76757a );
 a76762a <=( a76761a  and  a76754a );
 a76765a <=( (not A168)  and  A169 );
 a76768a <=( (not A166)  and  A167 );
 a76769a <=( a76768a  and  a76765a );
 a76772a <=( (not A200)  and  A199 );
 a76775a <=( A202  and  A201 );
 a76776a <=( a76775a  and  a76772a );
 a76777a <=( a76776a  and  a76769a );
 a76780a <=( (not A233)  and  (not A232) );
 a76783a <=( (not A266)  and  (not A265) );
 a76784a <=( a76783a  and  a76780a );
 a76787a <=( (not A299)  and  A298 );
 a76790a <=( A301  and  A300 );
 a76791a <=( a76790a  and  a76787a );
 a76792a <=( a76791a  and  a76784a );
 a76795a <=( (not A168)  and  A169 );
 a76798a <=( (not A166)  and  A167 );
 a76799a <=( a76798a  and  a76795a );
 a76802a <=( (not A200)  and  A199 );
 a76805a <=( A202  and  A201 );
 a76806a <=( a76805a  and  a76802a );
 a76807a <=( a76806a  and  a76799a );
 a76810a <=( (not A233)  and  (not A232) );
 a76813a <=( (not A266)  and  (not A265) );
 a76814a <=( a76813a  and  a76810a );
 a76817a <=( (not A299)  and  A298 );
 a76820a <=( A302  and  A300 );
 a76821a <=( a76820a  and  a76817a );
 a76822a <=( a76821a  and  a76814a );
 a76825a <=( (not A168)  and  A169 );
 a76828a <=( (not A166)  and  A167 );
 a76829a <=( a76828a  and  a76825a );
 a76832a <=( (not A200)  and  A199 );
 a76835a <=( A203  and  A201 );
 a76836a <=( a76835a  and  a76832a );
 a76837a <=( a76836a  and  a76829a );
 a76840a <=( A233  and  A232 );
 a76843a <=( (not A267)  and  A265 );
 a76844a <=( a76843a  and  a76840a );
 a76847a <=( (not A299)  and  A298 );
 a76850a <=( A301  and  A300 );
 a76851a <=( a76850a  and  a76847a );
 a76852a <=( a76851a  and  a76844a );
 a76855a <=( (not A168)  and  A169 );
 a76858a <=( (not A166)  and  A167 );
 a76859a <=( a76858a  and  a76855a );
 a76862a <=( (not A200)  and  A199 );
 a76865a <=( A203  and  A201 );
 a76866a <=( a76865a  and  a76862a );
 a76867a <=( a76866a  and  a76859a );
 a76870a <=( A233  and  A232 );
 a76873a <=( (not A267)  and  A265 );
 a76874a <=( a76873a  and  a76870a );
 a76877a <=( (not A299)  and  A298 );
 a76880a <=( A302  and  A300 );
 a76881a <=( a76880a  and  a76877a );
 a76882a <=( a76881a  and  a76874a );
 a76885a <=( (not A168)  and  A169 );
 a76888a <=( (not A166)  and  A167 );
 a76889a <=( a76888a  and  a76885a );
 a76892a <=( (not A200)  and  A199 );
 a76895a <=( A203  and  A201 );
 a76896a <=( a76895a  and  a76892a );
 a76897a <=( a76896a  and  a76889a );
 a76900a <=( A233  and  A232 );
 a76903a <=( A266  and  A265 );
 a76904a <=( a76903a  and  a76900a );
 a76907a <=( (not A299)  and  A298 );
 a76910a <=( A301  and  A300 );
 a76911a <=( a76910a  and  a76907a );
 a76912a <=( a76911a  and  a76904a );
 a76915a <=( (not A168)  and  A169 );
 a76918a <=( (not A166)  and  A167 );
 a76919a <=( a76918a  and  a76915a );
 a76922a <=( (not A200)  and  A199 );
 a76925a <=( A203  and  A201 );
 a76926a <=( a76925a  and  a76922a );
 a76927a <=( a76926a  and  a76919a );
 a76930a <=( A233  and  A232 );
 a76933a <=( A266  and  A265 );
 a76934a <=( a76933a  and  a76930a );
 a76937a <=( (not A299)  and  A298 );
 a76940a <=( A302  and  A300 );
 a76941a <=( a76940a  and  a76937a );
 a76942a <=( a76941a  and  a76934a );
 a76945a <=( (not A168)  and  A169 );
 a76948a <=( (not A166)  and  A167 );
 a76949a <=( a76948a  and  a76945a );
 a76952a <=( (not A200)  and  A199 );
 a76955a <=( A203  and  A201 );
 a76956a <=( a76955a  and  a76952a );
 a76957a <=( a76956a  and  a76949a );
 a76960a <=( A233  and  A232 );
 a76963a <=( (not A266)  and  (not A265) );
 a76964a <=( a76963a  and  a76960a );
 a76967a <=( (not A299)  and  A298 );
 a76970a <=( A301  and  A300 );
 a76971a <=( a76970a  and  a76967a );
 a76972a <=( a76971a  and  a76964a );
 a76975a <=( (not A168)  and  A169 );
 a76978a <=( (not A166)  and  A167 );
 a76979a <=( a76978a  and  a76975a );
 a76982a <=( (not A200)  and  A199 );
 a76985a <=( A203  and  A201 );
 a76986a <=( a76985a  and  a76982a );
 a76987a <=( a76986a  and  a76979a );
 a76990a <=( A233  and  A232 );
 a76993a <=( (not A266)  and  (not A265) );
 a76994a <=( a76993a  and  a76990a );
 a76997a <=( (not A299)  and  A298 );
 a77000a <=( A302  and  A300 );
 a77001a <=( a77000a  and  a76997a );
 a77002a <=( a77001a  and  a76994a );
 a77005a <=( (not A168)  and  A169 );
 a77008a <=( (not A166)  and  A167 );
 a77009a <=( a77008a  and  a77005a );
 a77012a <=( (not A200)  and  A199 );
 a77015a <=( A203  and  A201 );
 a77016a <=( a77015a  and  a77012a );
 a77017a <=( a77016a  and  a77009a );
 a77020a <=( (not A235)  and  (not A233) );
 a77023a <=( (not A266)  and  (not A236) );
 a77024a <=( a77023a  and  a77020a );
 a77027a <=( (not A269)  and  (not A268) );
 a77030a <=( A299  and  (not A298) );
 a77031a <=( a77030a  and  a77027a );
 a77032a <=( a77031a  and  a77024a );
 a77035a <=( (not A168)  and  A169 );
 a77038a <=( (not A166)  and  A167 );
 a77039a <=( a77038a  and  a77035a );
 a77042a <=( (not A200)  and  A199 );
 a77045a <=( A203  and  A201 );
 a77046a <=( a77045a  and  a77042a );
 a77047a <=( a77046a  and  a77039a );
 a77050a <=( (not A234)  and  (not A233) );
 a77053a <=( A266  and  A265 );
 a77054a <=( a77053a  and  a77050a );
 a77057a <=( (not A299)  and  A298 );
 a77060a <=( A301  and  A300 );
 a77061a <=( a77060a  and  a77057a );
 a77062a <=( a77061a  and  a77054a );
 a77065a <=( (not A168)  and  A169 );
 a77068a <=( (not A166)  and  A167 );
 a77069a <=( a77068a  and  a77065a );
 a77072a <=( (not A200)  and  A199 );
 a77075a <=( A203  and  A201 );
 a77076a <=( a77075a  and  a77072a );
 a77077a <=( a77076a  and  a77069a );
 a77080a <=( (not A234)  and  (not A233) );
 a77083a <=( A266  and  A265 );
 a77084a <=( a77083a  and  a77080a );
 a77087a <=( (not A299)  and  A298 );
 a77090a <=( A302  and  A300 );
 a77091a <=( a77090a  and  a77087a );
 a77092a <=( a77091a  and  a77084a );
 a77095a <=( (not A168)  and  A169 );
 a77098a <=( (not A166)  and  A167 );
 a77099a <=( a77098a  and  a77095a );
 a77102a <=( (not A200)  and  A199 );
 a77105a <=( A203  and  A201 );
 a77106a <=( a77105a  and  a77102a );
 a77107a <=( a77106a  and  a77099a );
 a77110a <=( (not A234)  and  (not A233) );
 a77113a <=( (not A267)  and  (not A266) );
 a77114a <=( a77113a  and  a77110a );
 a77117a <=( (not A299)  and  A298 );
 a77120a <=( A301  and  A300 );
 a77121a <=( a77120a  and  a77117a );
 a77122a <=( a77121a  and  a77114a );
 a77125a <=( (not A168)  and  A169 );
 a77128a <=( (not A166)  and  A167 );
 a77129a <=( a77128a  and  a77125a );
 a77132a <=( (not A200)  and  A199 );
 a77135a <=( A203  and  A201 );
 a77136a <=( a77135a  and  a77132a );
 a77137a <=( a77136a  and  a77129a );
 a77140a <=( (not A234)  and  (not A233) );
 a77143a <=( (not A267)  and  (not A266) );
 a77144a <=( a77143a  and  a77140a );
 a77147a <=( (not A299)  and  A298 );
 a77150a <=( A302  and  A300 );
 a77151a <=( a77150a  and  a77147a );
 a77152a <=( a77151a  and  a77144a );
 a77155a <=( (not A168)  and  A169 );
 a77158a <=( (not A166)  and  A167 );
 a77159a <=( a77158a  and  a77155a );
 a77162a <=( (not A200)  and  A199 );
 a77165a <=( A203  and  A201 );
 a77166a <=( a77165a  and  a77162a );
 a77167a <=( a77166a  and  a77159a );
 a77170a <=( (not A234)  and  (not A233) );
 a77173a <=( (not A266)  and  (not A265) );
 a77174a <=( a77173a  and  a77170a );
 a77177a <=( (not A299)  and  A298 );
 a77180a <=( A301  and  A300 );
 a77181a <=( a77180a  and  a77177a );
 a77182a <=( a77181a  and  a77174a );
 a77185a <=( (not A168)  and  A169 );
 a77188a <=( (not A166)  and  A167 );
 a77189a <=( a77188a  and  a77185a );
 a77192a <=( (not A200)  and  A199 );
 a77195a <=( A203  and  A201 );
 a77196a <=( a77195a  and  a77192a );
 a77197a <=( a77196a  and  a77189a );
 a77200a <=( (not A234)  and  (not A233) );
 a77203a <=( (not A266)  and  (not A265) );
 a77204a <=( a77203a  and  a77200a );
 a77207a <=( (not A299)  and  A298 );
 a77210a <=( A302  and  A300 );
 a77211a <=( a77210a  and  a77207a );
 a77212a <=( a77211a  and  a77204a );
 a77215a <=( (not A168)  and  A169 );
 a77218a <=( (not A166)  and  A167 );
 a77219a <=( a77218a  and  a77215a );
 a77222a <=( (not A200)  and  A199 );
 a77225a <=( A203  and  A201 );
 a77226a <=( a77225a  and  a77222a );
 a77227a <=( a77226a  and  a77219a );
 a77230a <=( (not A233)  and  A232 );
 a77233a <=( A235  and  A234 );
 a77234a <=( a77233a  and  a77230a );
 a77237a <=( (not A266)  and  A265 );
 a77240a <=( A268  and  A267 );
 a77241a <=( a77240a  and  a77237a );
 a77242a <=( a77241a  and  a77234a );
 a77245a <=( (not A168)  and  A169 );
 a77248a <=( (not A166)  and  A167 );
 a77249a <=( a77248a  and  a77245a );
 a77252a <=( (not A200)  and  A199 );
 a77255a <=( A203  and  A201 );
 a77256a <=( a77255a  and  a77252a );
 a77257a <=( a77256a  and  a77249a );
 a77260a <=( (not A233)  and  A232 );
 a77263a <=( A235  and  A234 );
 a77264a <=( a77263a  and  a77260a );
 a77267a <=( (not A266)  and  A265 );
 a77270a <=( A269  and  A267 );
 a77271a <=( a77270a  and  a77267a );
 a77272a <=( a77271a  and  a77264a );
 a77275a <=( (not A168)  and  A169 );
 a77278a <=( (not A166)  and  A167 );
 a77279a <=( a77278a  and  a77275a );
 a77282a <=( (not A200)  and  A199 );
 a77285a <=( A203  and  A201 );
 a77286a <=( a77285a  and  a77282a );
 a77287a <=( a77286a  and  a77279a );
 a77290a <=( (not A233)  and  A232 );
 a77293a <=( A236  and  A234 );
 a77294a <=( a77293a  and  a77290a );
 a77297a <=( (not A266)  and  A265 );
 a77300a <=( A268  and  A267 );
 a77301a <=( a77300a  and  a77297a );
 a77302a <=( a77301a  and  a77294a );
 a77305a <=( (not A168)  and  A169 );
 a77308a <=( (not A166)  and  A167 );
 a77309a <=( a77308a  and  a77305a );
 a77312a <=( (not A200)  and  A199 );
 a77315a <=( A203  and  A201 );
 a77316a <=( a77315a  and  a77312a );
 a77317a <=( a77316a  and  a77309a );
 a77320a <=( (not A233)  and  A232 );
 a77323a <=( A236  and  A234 );
 a77324a <=( a77323a  and  a77320a );
 a77327a <=( (not A266)  and  A265 );
 a77330a <=( A269  and  A267 );
 a77331a <=( a77330a  and  a77327a );
 a77332a <=( a77331a  and  a77324a );
 a77335a <=( (not A168)  and  A169 );
 a77338a <=( (not A166)  and  A167 );
 a77339a <=( a77338a  and  a77335a );
 a77342a <=( (not A200)  and  A199 );
 a77345a <=( A203  and  A201 );
 a77346a <=( a77345a  and  a77342a );
 a77347a <=( a77346a  and  a77339a );
 a77350a <=( (not A233)  and  (not A232) );
 a77353a <=( A266  and  A265 );
 a77354a <=( a77353a  and  a77350a );
 a77357a <=( (not A299)  and  A298 );
 a77360a <=( A301  and  A300 );
 a77361a <=( a77360a  and  a77357a );
 a77362a <=( a77361a  and  a77354a );
 a77365a <=( (not A168)  and  A169 );
 a77368a <=( (not A166)  and  A167 );
 a77369a <=( a77368a  and  a77365a );
 a77372a <=( (not A200)  and  A199 );
 a77375a <=( A203  and  A201 );
 a77376a <=( a77375a  and  a77372a );
 a77377a <=( a77376a  and  a77369a );
 a77380a <=( (not A233)  and  (not A232) );
 a77383a <=( A266  and  A265 );
 a77384a <=( a77383a  and  a77380a );
 a77387a <=( (not A299)  and  A298 );
 a77390a <=( A302  and  A300 );
 a77391a <=( a77390a  and  a77387a );
 a77392a <=( a77391a  and  a77384a );
 a77395a <=( (not A168)  and  A169 );
 a77398a <=( (not A166)  and  A167 );
 a77399a <=( a77398a  and  a77395a );
 a77402a <=( (not A200)  and  A199 );
 a77405a <=( A203  and  A201 );
 a77406a <=( a77405a  and  a77402a );
 a77407a <=( a77406a  and  a77399a );
 a77410a <=( (not A233)  and  (not A232) );
 a77413a <=( (not A267)  and  (not A266) );
 a77414a <=( a77413a  and  a77410a );
 a77417a <=( (not A299)  and  A298 );
 a77420a <=( A301  and  A300 );
 a77421a <=( a77420a  and  a77417a );
 a77422a <=( a77421a  and  a77414a );
 a77425a <=( (not A168)  and  A169 );
 a77428a <=( (not A166)  and  A167 );
 a77429a <=( a77428a  and  a77425a );
 a77432a <=( (not A200)  and  A199 );
 a77435a <=( A203  and  A201 );
 a77436a <=( a77435a  and  a77432a );
 a77437a <=( a77436a  and  a77429a );
 a77440a <=( (not A233)  and  (not A232) );
 a77443a <=( (not A267)  and  (not A266) );
 a77444a <=( a77443a  and  a77440a );
 a77447a <=( (not A299)  and  A298 );
 a77450a <=( A302  and  A300 );
 a77451a <=( a77450a  and  a77447a );
 a77452a <=( a77451a  and  a77444a );
 a77455a <=( (not A168)  and  A169 );
 a77458a <=( (not A166)  and  A167 );
 a77459a <=( a77458a  and  a77455a );
 a77462a <=( (not A200)  and  A199 );
 a77465a <=( A203  and  A201 );
 a77466a <=( a77465a  and  a77462a );
 a77467a <=( a77466a  and  a77459a );
 a77470a <=( (not A233)  and  (not A232) );
 a77473a <=( (not A266)  and  (not A265) );
 a77474a <=( a77473a  and  a77470a );
 a77477a <=( (not A299)  and  A298 );
 a77480a <=( A301  and  A300 );
 a77481a <=( a77480a  and  a77477a );
 a77482a <=( a77481a  and  a77474a );
 a77485a <=( (not A168)  and  A169 );
 a77488a <=( (not A166)  and  A167 );
 a77489a <=( a77488a  and  a77485a );
 a77492a <=( (not A200)  and  A199 );
 a77495a <=( A203  and  A201 );
 a77496a <=( a77495a  and  a77492a );
 a77497a <=( a77496a  and  a77489a );
 a77500a <=( (not A233)  and  (not A232) );
 a77503a <=( (not A266)  and  (not A265) );
 a77504a <=( a77503a  and  a77500a );
 a77507a <=( (not A299)  and  A298 );
 a77510a <=( A302  and  A300 );
 a77511a <=( a77510a  and  a77507a );
 a77512a <=( a77511a  and  a77504a );
 a77515a <=( (not A168)  and  A169 );
 a77518a <=( A166  and  (not A167) );
 a77519a <=( a77518a  and  a77515a );
 a77522a <=( A200  and  (not A199) );
 a77525a <=( (not A235)  and  (not A233) );
 a77526a <=( a77525a  and  a77522a );
 a77527a <=( a77526a  and  a77519a );
 a77530a <=( (not A266)  and  (not A236) );
 a77533a <=( (not A269)  and  (not A268) );
 a77534a <=( a77533a  and  a77530a );
 a77537a <=( (not A299)  and  A298 );
 a77540a <=( A301  and  A300 );
 a77541a <=( a77540a  and  a77537a );
 a77542a <=( a77541a  and  a77534a );
 a77545a <=( (not A168)  and  A169 );
 a77548a <=( A166  and  (not A167) );
 a77549a <=( a77548a  and  a77545a );
 a77552a <=( A200  and  (not A199) );
 a77555a <=( (not A235)  and  (not A233) );
 a77556a <=( a77555a  and  a77552a );
 a77557a <=( a77556a  and  a77549a );
 a77560a <=( (not A266)  and  (not A236) );
 a77563a <=( (not A269)  and  (not A268) );
 a77564a <=( a77563a  and  a77560a );
 a77567a <=( (not A299)  and  A298 );
 a77570a <=( A302  and  A300 );
 a77571a <=( a77570a  and  a77567a );
 a77572a <=( a77571a  and  a77564a );
 a77575a <=( (not A168)  and  A169 );
 a77578a <=( A166  and  (not A167) );
 a77579a <=( a77578a  and  a77575a );
 a77582a <=( (not A200)  and  A199 );
 a77585a <=( A202  and  A201 );
 a77586a <=( a77585a  and  a77582a );
 a77587a <=( a77586a  and  a77579a );
 a77590a <=( A233  and  A232 );
 a77593a <=( (not A267)  and  A265 );
 a77594a <=( a77593a  and  a77590a );
 a77597a <=( (not A299)  and  A298 );
 a77600a <=( A301  and  A300 );
 a77601a <=( a77600a  and  a77597a );
 a77602a <=( a77601a  and  a77594a );
 a77605a <=( (not A168)  and  A169 );
 a77608a <=( A166  and  (not A167) );
 a77609a <=( a77608a  and  a77605a );
 a77612a <=( (not A200)  and  A199 );
 a77615a <=( A202  and  A201 );
 a77616a <=( a77615a  and  a77612a );
 a77617a <=( a77616a  and  a77609a );
 a77620a <=( A233  and  A232 );
 a77623a <=( (not A267)  and  A265 );
 a77624a <=( a77623a  and  a77620a );
 a77627a <=( (not A299)  and  A298 );
 a77630a <=( A302  and  A300 );
 a77631a <=( a77630a  and  a77627a );
 a77632a <=( a77631a  and  a77624a );
 a77635a <=( (not A168)  and  A169 );
 a77638a <=( A166  and  (not A167) );
 a77639a <=( a77638a  and  a77635a );
 a77642a <=( (not A200)  and  A199 );
 a77645a <=( A202  and  A201 );
 a77646a <=( a77645a  and  a77642a );
 a77647a <=( a77646a  and  a77639a );
 a77650a <=( A233  and  A232 );
 a77653a <=( A266  and  A265 );
 a77654a <=( a77653a  and  a77650a );
 a77657a <=( (not A299)  and  A298 );
 a77660a <=( A301  and  A300 );
 a77661a <=( a77660a  and  a77657a );
 a77662a <=( a77661a  and  a77654a );
 a77665a <=( (not A168)  and  A169 );
 a77668a <=( A166  and  (not A167) );
 a77669a <=( a77668a  and  a77665a );
 a77672a <=( (not A200)  and  A199 );
 a77675a <=( A202  and  A201 );
 a77676a <=( a77675a  and  a77672a );
 a77677a <=( a77676a  and  a77669a );
 a77680a <=( A233  and  A232 );
 a77683a <=( A266  and  A265 );
 a77684a <=( a77683a  and  a77680a );
 a77687a <=( (not A299)  and  A298 );
 a77690a <=( A302  and  A300 );
 a77691a <=( a77690a  and  a77687a );
 a77692a <=( a77691a  and  a77684a );
 a77695a <=( (not A168)  and  A169 );
 a77698a <=( A166  and  (not A167) );
 a77699a <=( a77698a  and  a77695a );
 a77702a <=( (not A200)  and  A199 );
 a77705a <=( A202  and  A201 );
 a77706a <=( a77705a  and  a77702a );
 a77707a <=( a77706a  and  a77699a );
 a77710a <=( A233  and  A232 );
 a77713a <=( (not A266)  and  (not A265) );
 a77714a <=( a77713a  and  a77710a );
 a77717a <=( (not A299)  and  A298 );
 a77720a <=( A301  and  A300 );
 a77721a <=( a77720a  and  a77717a );
 a77722a <=( a77721a  and  a77714a );
 a77725a <=( (not A168)  and  A169 );
 a77728a <=( A166  and  (not A167) );
 a77729a <=( a77728a  and  a77725a );
 a77732a <=( (not A200)  and  A199 );
 a77735a <=( A202  and  A201 );
 a77736a <=( a77735a  and  a77732a );
 a77737a <=( a77736a  and  a77729a );
 a77740a <=( A233  and  A232 );
 a77743a <=( (not A266)  and  (not A265) );
 a77744a <=( a77743a  and  a77740a );
 a77747a <=( (not A299)  and  A298 );
 a77750a <=( A302  and  A300 );
 a77751a <=( a77750a  and  a77747a );
 a77752a <=( a77751a  and  a77744a );
 a77755a <=( (not A168)  and  A169 );
 a77758a <=( A166  and  (not A167) );
 a77759a <=( a77758a  and  a77755a );
 a77762a <=( (not A200)  and  A199 );
 a77765a <=( A202  and  A201 );
 a77766a <=( a77765a  and  a77762a );
 a77767a <=( a77766a  and  a77759a );
 a77770a <=( (not A235)  and  (not A233) );
 a77773a <=( (not A266)  and  (not A236) );
 a77774a <=( a77773a  and  a77770a );
 a77777a <=( (not A269)  and  (not A268) );
 a77780a <=( A299  and  (not A298) );
 a77781a <=( a77780a  and  a77777a );
 a77782a <=( a77781a  and  a77774a );
 a77785a <=( (not A168)  and  A169 );
 a77788a <=( A166  and  (not A167) );
 a77789a <=( a77788a  and  a77785a );
 a77792a <=( (not A200)  and  A199 );
 a77795a <=( A202  and  A201 );
 a77796a <=( a77795a  and  a77792a );
 a77797a <=( a77796a  and  a77789a );
 a77800a <=( (not A234)  and  (not A233) );
 a77803a <=( A266  and  A265 );
 a77804a <=( a77803a  and  a77800a );
 a77807a <=( (not A299)  and  A298 );
 a77810a <=( A301  and  A300 );
 a77811a <=( a77810a  and  a77807a );
 a77812a <=( a77811a  and  a77804a );
 a77815a <=( (not A168)  and  A169 );
 a77818a <=( A166  and  (not A167) );
 a77819a <=( a77818a  and  a77815a );
 a77822a <=( (not A200)  and  A199 );
 a77825a <=( A202  and  A201 );
 a77826a <=( a77825a  and  a77822a );
 a77827a <=( a77826a  and  a77819a );
 a77830a <=( (not A234)  and  (not A233) );
 a77833a <=( A266  and  A265 );
 a77834a <=( a77833a  and  a77830a );
 a77837a <=( (not A299)  and  A298 );
 a77840a <=( A302  and  A300 );
 a77841a <=( a77840a  and  a77837a );
 a77842a <=( a77841a  and  a77834a );
 a77845a <=( (not A168)  and  A169 );
 a77848a <=( A166  and  (not A167) );
 a77849a <=( a77848a  and  a77845a );
 a77852a <=( (not A200)  and  A199 );
 a77855a <=( A202  and  A201 );
 a77856a <=( a77855a  and  a77852a );
 a77857a <=( a77856a  and  a77849a );
 a77860a <=( (not A234)  and  (not A233) );
 a77863a <=( (not A267)  and  (not A266) );
 a77864a <=( a77863a  and  a77860a );
 a77867a <=( (not A299)  and  A298 );
 a77870a <=( A301  and  A300 );
 a77871a <=( a77870a  and  a77867a );
 a77872a <=( a77871a  and  a77864a );
 a77875a <=( (not A168)  and  A169 );
 a77878a <=( A166  and  (not A167) );
 a77879a <=( a77878a  and  a77875a );
 a77882a <=( (not A200)  and  A199 );
 a77885a <=( A202  and  A201 );
 a77886a <=( a77885a  and  a77882a );
 a77887a <=( a77886a  and  a77879a );
 a77890a <=( (not A234)  and  (not A233) );
 a77893a <=( (not A267)  and  (not A266) );
 a77894a <=( a77893a  and  a77890a );
 a77897a <=( (not A299)  and  A298 );
 a77900a <=( A302  and  A300 );
 a77901a <=( a77900a  and  a77897a );
 a77902a <=( a77901a  and  a77894a );
 a77905a <=( (not A168)  and  A169 );
 a77908a <=( A166  and  (not A167) );
 a77909a <=( a77908a  and  a77905a );
 a77912a <=( (not A200)  and  A199 );
 a77915a <=( A202  and  A201 );
 a77916a <=( a77915a  and  a77912a );
 a77917a <=( a77916a  and  a77909a );
 a77920a <=( (not A234)  and  (not A233) );
 a77923a <=( (not A266)  and  (not A265) );
 a77924a <=( a77923a  and  a77920a );
 a77927a <=( (not A299)  and  A298 );
 a77930a <=( A301  and  A300 );
 a77931a <=( a77930a  and  a77927a );
 a77932a <=( a77931a  and  a77924a );
 a77935a <=( (not A168)  and  A169 );
 a77938a <=( A166  and  (not A167) );
 a77939a <=( a77938a  and  a77935a );
 a77942a <=( (not A200)  and  A199 );
 a77945a <=( A202  and  A201 );
 a77946a <=( a77945a  and  a77942a );
 a77947a <=( a77946a  and  a77939a );
 a77950a <=( (not A234)  and  (not A233) );
 a77953a <=( (not A266)  and  (not A265) );
 a77954a <=( a77953a  and  a77950a );
 a77957a <=( (not A299)  and  A298 );
 a77960a <=( A302  and  A300 );
 a77961a <=( a77960a  and  a77957a );
 a77962a <=( a77961a  and  a77954a );
 a77965a <=( (not A168)  and  A169 );
 a77968a <=( A166  and  (not A167) );
 a77969a <=( a77968a  and  a77965a );
 a77972a <=( (not A200)  and  A199 );
 a77975a <=( A202  and  A201 );
 a77976a <=( a77975a  and  a77972a );
 a77977a <=( a77976a  and  a77969a );
 a77980a <=( (not A233)  and  A232 );
 a77983a <=( A235  and  A234 );
 a77984a <=( a77983a  and  a77980a );
 a77987a <=( (not A266)  and  A265 );
 a77990a <=( A268  and  A267 );
 a77991a <=( a77990a  and  a77987a );
 a77992a <=( a77991a  and  a77984a );
 a77995a <=( (not A168)  and  A169 );
 a77998a <=( A166  and  (not A167) );
 a77999a <=( a77998a  and  a77995a );
 a78002a <=( (not A200)  and  A199 );
 a78005a <=( A202  and  A201 );
 a78006a <=( a78005a  and  a78002a );
 a78007a <=( a78006a  and  a77999a );
 a78010a <=( (not A233)  and  A232 );
 a78013a <=( A235  and  A234 );
 a78014a <=( a78013a  and  a78010a );
 a78017a <=( (not A266)  and  A265 );
 a78020a <=( A269  and  A267 );
 a78021a <=( a78020a  and  a78017a );
 a78022a <=( a78021a  and  a78014a );
 a78025a <=( (not A168)  and  A169 );
 a78028a <=( A166  and  (not A167) );
 a78029a <=( a78028a  and  a78025a );
 a78032a <=( (not A200)  and  A199 );
 a78035a <=( A202  and  A201 );
 a78036a <=( a78035a  and  a78032a );
 a78037a <=( a78036a  and  a78029a );
 a78040a <=( (not A233)  and  A232 );
 a78043a <=( A236  and  A234 );
 a78044a <=( a78043a  and  a78040a );
 a78047a <=( (not A266)  and  A265 );
 a78050a <=( A268  and  A267 );
 a78051a <=( a78050a  and  a78047a );
 a78052a <=( a78051a  and  a78044a );
 a78055a <=( (not A168)  and  A169 );
 a78058a <=( A166  and  (not A167) );
 a78059a <=( a78058a  and  a78055a );
 a78062a <=( (not A200)  and  A199 );
 a78065a <=( A202  and  A201 );
 a78066a <=( a78065a  and  a78062a );
 a78067a <=( a78066a  and  a78059a );
 a78070a <=( (not A233)  and  A232 );
 a78073a <=( A236  and  A234 );
 a78074a <=( a78073a  and  a78070a );
 a78077a <=( (not A266)  and  A265 );
 a78080a <=( A269  and  A267 );
 a78081a <=( a78080a  and  a78077a );
 a78082a <=( a78081a  and  a78074a );
 a78085a <=( (not A168)  and  A169 );
 a78088a <=( A166  and  (not A167) );
 a78089a <=( a78088a  and  a78085a );
 a78092a <=( (not A200)  and  A199 );
 a78095a <=( A202  and  A201 );
 a78096a <=( a78095a  and  a78092a );
 a78097a <=( a78096a  and  a78089a );
 a78100a <=( (not A233)  and  (not A232) );
 a78103a <=( A266  and  A265 );
 a78104a <=( a78103a  and  a78100a );
 a78107a <=( (not A299)  and  A298 );
 a78110a <=( A301  and  A300 );
 a78111a <=( a78110a  and  a78107a );
 a78112a <=( a78111a  and  a78104a );
 a78115a <=( (not A168)  and  A169 );
 a78118a <=( A166  and  (not A167) );
 a78119a <=( a78118a  and  a78115a );
 a78122a <=( (not A200)  and  A199 );
 a78125a <=( A202  and  A201 );
 a78126a <=( a78125a  and  a78122a );
 a78127a <=( a78126a  and  a78119a );
 a78130a <=( (not A233)  and  (not A232) );
 a78133a <=( A266  and  A265 );
 a78134a <=( a78133a  and  a78130a );
 a78137a <=( (not A299)  and  A298 );
 a78140a <=( A302  and  A300 );
 a78141a <=( a78140a  and  a78137a );
 a78142a <=( a78141a  and  a78134a );
 a78145a <=( (not A168)  and  A169 );
 a78148a <=( A166  and  (not A167) );
 a78149a <=( a78148a  and  a78145a );
 a78152a <=( (not A200)  and  A199 );
 a78155a <=( A202  and  A201 );
 a78156a <=( a78155a  and  a78152a );
 a78157a <=( a78156a  and  a78149a );
 a78160a <=( (not A233)  and  (not A232) );
 a78163a <=( (not A267)  and  (not A266) );
 a78164a <=( a78163a  and  a78160a );
 a78167a <=( (not A299)  and  A298 );
 a78170a <=( A301  and  A300 );
 a78171a <=( a78170a  and  a78167a );
 a78172a <=( a78171a  and  a78164a );
 a78175a <=( (not A168)  and  A169 );
 a78178a <=( A166  and  (not A167) );
 a78179a <=( a78178a  and  a78175a );
 a78182a <=( (not A200)  and  A199 );
 a78185a <=( A202  and  A201 );
 a78186a <=( a78185a  and  a78182a );
 a78187a <=( a78186a  and  a78179a );
 a78190a <=( (not A233)  and  (not A232) );
 a78193a <=( (not A267)  and  (not A266) );
 a78194a <=( a78193a  and  a78190a );
 a78197a <=( (not A299)  and  A298 );
 a78200a <=( A302  and  A300 );
 a78201a <=( a78200a  and  a78197a );
 a78202a <=( a78201a  and  a78194a );
 a78205a <=( (not A168)  and  A169 );
 a78208a <=( A166  and  (not A167) );
 a78209a <=( a78208a  and  a78205a );
 a78212a <=( (not A200)  and  A199 );
 a78215a <=( A202  and  A201 );
 a78216a <=( a78215a  and  a78212a );
 a78217a <=( a78216a  and  a78209a );
 a78220a <=( (not A233)  and  (not A232) );
 a78223a <=( (not A266)  and  (not A265) );
 a78224a <=( a78223a  and  a78220a );
 a78227a <=( (not A299)  and  A298 );
 a78230a <=( A301  and  A300 );
 a78231a <=( a78230a  and  a78227a );
 a78232a <=( a78231a  and  a78224a );
 a78235a <=( (not A168)  and  A169 );
 a78238a <=( A166  and  (not A167) );
 a78239a <=( a78238a  and  a78235a );
 a78242a <=( (not A200)  and  A199 );
 a78245a <=( A202  and  A201 );
 a78246a <=( a78245a  and  a78242a );
 a78247a <=( a78246a  and  a78239a );
 a78250a <=( (not A233)  and  (not A232) );
 a78253a <=( (not A266)  and  (not A265) );
 a78254a <=( a78253a  and  a78250a );
 a78257a <=( (not A299)  and  A298 );
 a78260a <=( A302  and  A300 );
 a78261a <=( a78260a  and  a78257a );
 a78262a <=( a78261a  and  a78254a );
 a78265a <=( (not A168)  and  A169 );
 a78268a <=( A166  and  (not A167) );
 a78269a <=( a78268a  and  a78265a );
 a78272a <=( (not A200)  and  A199 );
 a78275a <=( A203  and  A201 );
 a78276a <=( a78275a  and  a78272a );
 a78277a <=( a78276a  and  a78269a );
 a78280a <=( A233  and  A232 );
 a78283a <=( (not A267)  and  A265 );
 a78284a <=( a78283a  and  a78280a );
 a78287a <=( (not A299)  and  A298 );
 a78290a <=( A301  and  A300 );
 a78291a <=( a78290a  and  a78287a );
 a78292a <=( a78291a  and  a78284a );
 a78295a <=( (not A168)  and  A169 );
 a78298a <=( A166  and  (not A167) );
 a78299a <=( a78298a  and  a78295a );
 a78302a <=( (not A200)  and  A199 );
 a78305a <=( A203  and  A201 );
 a78306a <=( a78305a  and  a78302a );
 a78307a <=( a78306a  and  a78299a );
 a78310a <=( A233  and  A232 );
 a78313a <=( (not A267)  and  A265 );
 a78314a <=( a78313a  and  a78310a );
 a78317a <=( (not A299)  and  A298 );
 a78320a <=( A302  and  A300 );
 a78321a <=( a78320a  and  a78317a );
 a78322a <=( a78321a  and  a78314a );
 a78325a <=( (not A168)  and  A169 );
 a78328a <=( A166  and  (not A167) );
 a78329a <=( a78328a  and  a78325a );
 a78332a <=( (not A200)  and  A199 );
 a78335a <=( A203  and  A201 );
 a78336a <=( a78335a  and  a78332a );
 a78337a <=( a78336a  and  a78329a );
 a78340a <=( A233  and  A232 );
 a78343a <=( A266  and  A265 );
 a78344a <=( a78343a  and  a78340a );
 a78347a <=( (not A299)  and  A298 );
 a78350a <=( A301  and  A300 );
 a78351a <=( a78350a  and  a78347a );
 a78352a <=( a78351a  and  a78344a );
 a78355a <=( (not A168)  and  A169 );
 a78358a <=( A166  and  (not A167) );
 a78359a <=( a78358a  and  a78355a );
 a78362a <=( (not A200)  and  A199 );
 a78365a <=( A203  and  A201 );
 a78366a <=( a78365a  and  a78362a );
 a78367a <=( a78366a  and  a78359a );
 a78370a <=( A233  and  A232 );
 a78373a <=( A266  and  A265 );
 a78374a <=( a78373a  and  a78370a );
 a78377a <=( (not A299)  and  A298 );
 a78380a <=( A302  and  A300 );
 a78381a <=( a78380a  and  a78377a );
 a78382a <=( a78381a  and  a78374a );
 a78385a <=( (not A168)  and  A169 );
 a78388a <=( A166  and  (not A167) );
 a78389a <=( a78388a  and  a78385a );
 a78392a <=( (not A200)  and  A199 );
 a78395a <=( A203  and  A201 );
 a78396a <=( a78395a  and  a78392a );
 a78397a <=( a78396a  and  a78389a );
 a78400a <=( A233  and  A232 );
 a78403a <=( (not A266)  and  (not A265) );
 a78404a <=( a78403a  and  a78400a );
 a78407a <=( (not A299)  and  A298 );
 a78410a <=( A301  and  A300 );
 a78411a <=( a78410a  and  a78407a );
 a78412a <=( a78411a  and  a78404a );
 a78415a <=( (not A168)  and  A169 );
 a78418a <=( A166  and  (not A167) );
 a78419a <=( a78418a  and  a78415a );
 a78422a <=( (not A200)  and  A199 );
 a78425a <=( A203  and  A201 );
 a78426a <=( a78425a  and  a78422a );
 a78427a <=( a78426a  and  a78419a );
 a78430a <=( A233  and  A232 );
 a78433a <=( (not A266)  and  (not A265) );
 a78434a <=( a78433a  and  a78430a );
 a78437a <=( (not A299)  and  A298 );
 a78440a <=( A302  and  A300 );
 a78441a <=( a78440a  and  a78437a );
 a78442a <=( a78441a  and  a78434a );
 a78445a <=( (not A168)  and  A169 );
 a78448a <=( A166  and  (not A167) );
 a78449a <=( a78448a  and  a78445a );
 a78452a <=( (not A200)  and  A199 );
 a78455a <=( A203  and  A201 );
 a78456a <=( a78455a  and  a78452a );
 a78457a <=( a78456a  and  a78449a );
 a78460a <=( (not A235)  and  (not A233) );
 a78463a <=( (not A266)  and  (not A236) );
 a78464a <=( a78463a  and  a78460a );
 a78467a <=( (not A269)  and  (not A268) );
 a78470a <=( A299  and  (not A298) );
 a78471a <=( a78470a  and  a78467a );
 a78472a <=( a78471a  and  a78464a );
 a78475a <=( (not A168)  and  A169 );
 a78478a <=( A166  and  (not A167) );
 a78479a <=( a78478a  and  a78475a );
 a78482a <=( (not A200)  and  A199 );
 a78485a <=( A203  and  A201 );
 a78486a <=( a78485a  and  a78482a );
 a78487a <=( a78486a  and  a78479a );
 a78490a <=( (not A234)  and  (not A233) );
 a78493a <=( A266  and  A265 );
 a78494a <=( a78493a  and  a78490a );
 a78497a <=( (not A299)  and  A298 );
 a78500a <=( A301  and  A300 );
 a78501a <=( a78500a  and  a78497a );
 a78502a <=( a78501a  and  a78494a );
 a78505a <=( (not A168)  and  A169 );
 a78508a <=( A166  and  (not A167) );
 a78509a <=( a78508a  and  a78505a );
 a78512a <=( (not A200)  and  A199 );
 a78515a <=( A203  and  A201 );
 a78516a <=( a78515a  and  a78512a );
 a78517a <=( a78516a  and  a78509a );
 a78520a <=( (not A234)  and  (not A233) );
 a78523a <=( A266  and  A265 );
 a78524a <=( a78523a  and  a78520a );
 a78527a <=( (not A299)  and  A298 );
 a78530a <=( A302  and  A300 );
 a78531a <=( a78530a  and  a78527a );
 a78532a <=( a78531a  and  a78524a );
 a78535a <=( (not A168)  and  A169 );
 a78538a <=( A166  and  (not A167) );
 a78539a <=( a78538a  and  a78535a );
 a78542a <=( (not A200)  and  A199 );
 a78545a <=( A203  and  A201 );
 a78546a <=( a78545a  and  a78542a );
 a78547a <=( a78546a  and  a78539a );
 a78550a <=( (not A234)  and  (not A233) );
 a78553a <=( (not A267)  and  (not A266) );
 a78554a <=( a78553a  and  a78550a );
 a78557a <=( (not A299)  and  A298 );
 a78560a <=( A301  and  A300 );
 a78561a <=( a78560a  and  a78557a );
 a78562a <=( a78561a  and  a78554a );
 a78565a <=( (not A168)  and  A169 );
 a78568a <=( A166  and  (not A167) );
 a78569a <=( a78568a  and  a78565a );
 a78572a <=( (not A200)  and  A199 );
 a78575a <=( A203  and  A201 );
 a78576a <=( a78575a  and  a78572a );
 a78577a <=( a78576a  and  a78569a );
 a78580a <=( (not A234)  and  (not A233) );
 a78583a <=( (not A267)  and  (not A266) );
 a78584a <=( a78583a  and  a78580a );
 a78587a <=( (not A299)  and  A298 );
 a78590a <=( A302  and  A300 );
 a78591a <=( a78590a  and  a78587a );
 a78592a <=( a78591a  and  a78584a );
 a78595a <=( (not A168)  and  A169 );
 a78598a <=( A166  and  (not A167) );
 a78599a <=( a78598a  and  a78595a );
 a78602a <=( (not A200)  and  A199 );
 a78605a <=( A203  and  A201 );
 a78606a <=( a78605a  and  a78602a );
 a78607a <=( a78606a  and  a78599a );
 a78610a <=( (not A234)  and  (not A233) );
 a78613a <=( (not A266)  and  (not A265) );
 a78614a <=( a78613a  and  a78610a );
 a78617a <=( (not A299)  and  A298 );
 a78620a <=( A301  and  A300 );
 a78621a <=( a78620a  and  a78617a );
 a78622a <=( a78621a  and  a78614a );
 a78625a <=( (not A168)  and  A169 );
 a78628a <=( A166  and  (not A167) );
 a78629a <=( a78628a  and  a78625a );
 a78632a <=( (not A200)  and  A199 );
 a78635a <=( A203  and  A201 );
 a78636a <=( a78635a  and  a78632a );
 a78637a <=( a78636a  and  a78629a );
 a78640a <=( (not A234)  and  (not A233) );
 a78643a <=( (not A266)  and  (not A265) );
 a78644a <=( a78643a  and  a78640a );
 a78647a <=( (not A299)  and  A298 );
 a78650a <=( A302  and  A300 );
 a78651a <=( a78650a  and  a78647a );
 a78652a <=( a78651a  and  a78644a );
 a78655a <=( (not A168)  and  A169 );
 a78658a <=( A166  and  (not A167) );
 a78659a <=( a78658a  and  a78655a );
 a78662a <=( (not A200)  and  A199 );
 a78665a <=( A203  and  A201 );
 a78666a <=( a78665a  and  a78662a );
 a78667a <=( a78666a  and  a78659a );
 a78670a <=( (not A233)  and  A232 );
 a78673a <=( A235  and  A234 );
 a78674a <=( a78673a  and  a78670a );
 a78677a <=( (not A266)  and  A265 );
 a78680a <=( A268  and  A267 );
 a78681a <=( a78680a  and  a78677a );
 a78682a <=( a78681a  and  a78674a );
 a78685a <=( (not A168)  and  A169 );
 a78688a <=( A166  and  (not A167) );
 a78689a <=( a78688a  and  a78685a );
 a78692a <=( (not A200)  and  A199 );
 a78695a <=( A203  and  A201 );
 a78696a <=( a78695a  and  a78692a );
 a78697a <=( a78696a  and  a78689a );
 a78700a <=( (not A233)  and  A232 );
 a78703a <=( A235  and  A234 );
 a78704a <=( a78703a  and  a78700a );
 a78707a <=( (not A266)  and  A265 );
 a78710a <=( A269  and  A267 );
 a78711a <=( a78710a  and  a78707a );
 a78712a <=( a78711a  and  a78704a );
 a78715a <=( (not A168)  and  A169 );
 a78718a <=( A166  and  (not A167) );
 a78719a <=( a78718a  and  a78715a );
 a78722a <=( (not A200)  and  A199 );
 a78725a <=( A203  and  A201 );
 a78726a <=( a78725a  and  a78722a );
 a78727a <=( a78726a  and  a78719a );
 a78730a <=( (not A233)  and  A232 );
 a78733a <=( A236  and  A234 );
 a78734a <=( a78733a  and  a78730a );
 a78737a <=( (not A266)  and  A265 );
 a78740a <=( A268  and  A267 );
 a78741a <=( a78740a  and  a78737a );
 a78742a <=( a78741a  and  a78734a );
 a78745a <=( (not A168)  and  A169 );
 a78748a <=( A166  and  (not A167) );
 a78749a <=( a78748a  and  a78745a );
 a78752a <=( (not A200)  and  A199 );
 a78755a <=( A203  and  A201 );
 a78756a <=( a78755a  and  a78752a );
 a78757a <=( a78756a  and  a78749a );
 a78760a <=( (not A233)  and  A232 );
 a78763a <=( A236  and  A234 );
 a78764a <=( a78763a  and  a78760a );
 a78767a <=( (not A266)  and  A265 );
 a78770a <=( A269  and  A267 );
 a78771a <=( a78770a  and  a78767a );
 a78772a <=( a78771a  and  a78764a );
 a78775a <=( (not A168)  and  A169 );
 a78778a <=( A166  and  (not A167) );
 a78779a <=( a78778a  and  a78775a );
 a78782a <=( (not A200)  and  A199 );
 a78785a <=( A203  and  A201 );
 a78786a <=( a78785a  and  a78782a );
 a78787a <=( a78786a  and  a78779a );
 a78790a <=( (not A233)  and  (not A232) );
 a78793a <=( A266  and  A265 );
 a78794a <=( a78793a  and  a78790a );
 a78797a <=( (not A299)  and  A298 );
 a78800a <=( A301  and  A300 );
 a78801a <=( a78800a  and  a78797a );
 a78802a <=( a78801a  and  a78794a );
 a78805a <=( (not A168)  and  A169 );
 a78808a <=( A166  and  (not A167) );
 a78809a <=( a78808a  and  a78805a );
 a78812a <=( (not A200)  and  A199 );
 a78815a <=( A203  and  A201 );
 a78816a <=( a78815a  and  a78812a );
 a78817a <=( a78816a  and  a78809a );
 a78820a <=( (not A233)  and  (not A232) );
 a78823a <=( A266  and  A265 );
 a78824a <=( a78823a  and  a78820a );
 a78827a <=( (not A299)  and  A298 );
 a78830a <=( A302  and  A300 );
 a78831a <=( a78830a  and  a78827a );
 a78832a <=( a78831a  and  a78824a );
 a78835a <=( (not A168)  and  A169 );
 a78838a <=( A166  and  (not A167) );
 a78839a <=( a78838a  and  a78835a );
 a78842a <=( (not A200)  and  A199 );
 a78845a <=( A203  and  A201 );
 a78846a <=( a78845a  and  a78842a );
 a78847a <=( a78846a  and  a78839a );
 a78850a <=( (not A233)  and  (not A232) );
 a78853a <=( (not A267)  and  (not A266) );
 a78854a <=( a78853a  and  a78850a );
 a78857a <=( (not A299)  and  A298 );
 a78860a <=( A301  and  A300 );
 a78861a <=( a78860a  and  a78857a );
 a78862a <=( a78861a  and  a78854a );
 a78865a <=( (not A168)  and  A169 );
 a78868a <=( A166  and  (not A167) );
 a78869a <=( a78868a  and  a78865a );
 a78872a <=( (not A200)  and  A199 );
 a78875a <=( A203  and  A201 );
 a78876a <=( a78875a  and  a78872a );
 a78877a <=( a78876a  and  a78869a );
 a78880a <=( (not A233)  and  (not A232) );
 a78883a <=( (not A267)  and  (not A266) );
 a78884a <=( a78883a  and  a78880a );
 a78887a <=( (not A299)  and  A298 );
 a78890a <=( A302  and  A300 );
 a78891a <=( a78890a  and  a78887a );
 a78892a <=( a78891a  and  a78884a );
 a78895a <=( (not A168)  and  A169 );
 a78898a <=( A166  and  (not A167) );
 a78899a <=( a78898a  and  a78895a );
 a78902a <=( (not A200)  and  A199 );
 a78905a <=( A203  and  A201 );
 a78906a <=( a78905a  and  a78902a );
 a78907a <=( a78906a  and  a78899a );
 a78910a <=( (not A233)  and  (not A232) );
 a78913a <=( (not A266)  and  (not A265) );
 a78914a <=( a78913a  and  a78910a );
 a78917a <=( (not A299)  and  A298 );
 a78920a <=( A301  and  A300 );
 a78921a <=( a78920a  and  a78917a );
 a78922a <=( a78921a  and  a78914a );
 a78925a <=( (not A168)  and  A169 );
 a78928a <=( A166  and  (not A167) );
 a78929a <=( a78928a  and  a78925a );
 a78932a <=( (not A200)  and  A199 );
 a78935a <=( A203  and  A201 );
 a78936a <=( a78935a  and  a78932a );
 a78937a <=( a78936a  and  a78929a );
 a78940a <=( (not A233)  and  (not A232) );
 a78943a <=( (not A266)  and  (not A265) );
 a78944a <=( a78943a  and  a78940a );
 a78947a <=( (not A299)  and  A298 );
 a78950a <=( A302  and  A300 );
 a78951a <=( a78950a  and  a78947a );
 a78952a <=( a78951a  and  a78944a );
 a78955a <=( A169  and  A170 );
 a78958a <=( A199  and  (not A168) );
 a78959a <=( a78958a  and  a78955a );
 a78962a <=( A201  and  (not A200) );
 a78965a <=( A232  and  A202 );
 a78966a <=( a78965a  and  a78962a );
 a78967a <=( a78966a  and  a78959a );
 a78970a <=( A265  and  A233 );
 a78973a <=( (not A269)  and  (not A268) );
 a78974a <=( a78973a  and  a78970a );
 a78977a <=( (not A299)  and  A298 );
 a78980a <=( A301  and  A300 );
 a78981a <=( a78980a  and  a78977a );
 a78982a <=( a78981a  and  a78974a );
 a78985a <=( A169  and  A170 );
 a78988a <=( A199  and  (not A168) );
 a78989a <=( a78988a  and  a78985a );
 a78992a <=( A201  and  (not A200) );
 a78995a <=( A232  and  A202 );
 a78996a <=( a78995a  and  a78992a );
 a78997a <=( a78996a  and  a78989a );
 a79000a <=( A265  and  A233 );
 a79003a <=( (not A269)  and  (not A268) );
 a79004a <=( a79003a  and  a79000a );
 a79007a <=( (not A299)  and  A298 );
 a79010a <=( A302  and  A300 );
 a79011a <=( a79010a  and  a79007a );
 a79012a <=( a79011a  and  a79004a );
 a79015a <=( A169  and  A170 );
 a79018a <=( A199  and  (not A168) );
 a79019a <=( a79018a  and  a79015a );
 a79022a <=( A201  and  (not A200) );
 a79025a <=( (not A233)  and  A202 );
 a79026a <=( a79025a  and  a79022a );
 a79027a <=( a79026a  and  a79019a );
 a79030a <=( (not A236)  and  (not A235) );
 a79033a <=( A266  and  A265 );
 a79034a <=( a79033a  and  a79030a );
 a79037a <=( (not A299)  and  A298 );
 a79040a <=( A301  and  A300 );
 a79041a <=( a79040a  and  a79037a );
 a79042a <=( a79041a  and  a79034a );
 a79045a <=( A169  and  A170 );
 a79048a <=( A199  and  (not A168) );
 a79049a <=( a79048a  and  a79045a );
 a79052a <=( A201  and  (not A200) );
 a79055a <=( (not A233)  and  A202 );
 a79056a <=( a79055a  and  a79052a );
 a79057a <=( a79056a  and  a79049a );
 a79060a <=( (not A236)  and  (not A235) );
 a79063a <=( A266  and  A265 );
 a79064a <=( a79063a  and  a79060a );
 a79067a <=( (not A299)  and  A298 );
 a79070a <=( A302  and  A300 );
 a79071a <=( a79070a  and  a79067a );
 a79072a <=( a79071a  and  a79064a );
 a79075a <=( A169  and  A170 );
 a79078a <=( A199  and  (not A168) );
 a79079a <=( a79078a  and  a79075a );
 a79082a <=( A201  and  (not A200) );
 a79085a <=( (not A233)  and  A202 );
 a79086a <=( a79085a  and  a79082a );
 a79087a <=( a79086a  and  a79079a );
 a79090a <=( (not A236)  and  (not A235) );
 a79093a <=( (not A267)  and  (not A266) );
 a79094a <=( a79093a  and  a79090a );
 a79097a <=( (not A299)  and  A298 );
 a79100a <=( A301  and  A300 );
 a79101a <=( a79100a  and  a79097a );
 a79102a <=( a79101a  and  a79094a );
 a79105a <=( A169  and  A170 );
 a79108a <=( A199  and  (not A168) );
 a79109a <=( a79108a  and  a79105a );
 a79112a <=( A201  and  (not A200) );
 a79115a <=( (not A233)  and  A202 );
 a79116a <=( a79115a  and  a79112a );
 a79117a <=( a79116a  and  a79109a );
 a79120a <=( (not A236)  and  (not A235) );
 a79123a <=( (not A267)  and  (not A266) );
 a79124a <=( a79123a  and  a79120a );
 a79127a <=( (not A299)  and  A298 );
 a79130a <=( A302  and  A300 );
 a79131a <=( a79130a  and  a79127a );
 a79132a <=( a79131a  and  a79124a );
 a79135a <=( A169  and  A170 );
 a79138a <=( A199  and  (not A168) );
 a79139a <=( a79138a  and  a79135a );
 a79142a <=( A201  and  (not A200) );
 a79145a <=( (not A233)  and  A202 );
 a79146a <=( a79145a  and  a79142a );
 a79147a <=( a79146a  and  a79139a );
 a79150a <=( (not A236)  and  (not A235) );
 a79153a <=( (not A266)  and  (not A265) );
 a79154a <=( a79153a  and  a79150a );
 a79157a <=( (not A299)  and  A298 );
 a79160a <=( A301  and  A300 );
 a79161a <=( a79160a  and  a79157a );
 a79162a <=( a79161a  and  a79154a );
 a79165a <=( A169  and  A170 );
 a79168a <=( A199  and  (not A168) );
 a79169a <=( a79168a  and  a79165a );
 a79172a <=( A201  and  (not A200) );
 a79175a <=( (not A233)  and  A202 );
 a79176a <=( a79175a  and  a79172a );
 a79177a <=( a79176a  and  a79169a );
 a79180a <=( (not A236)  and  (not A235) );
 a79183a <=( (not A266)  and  (not A265) );
 a79184a <=( a79183a  and  a79180a );
 a79187a <=( (not A299)  and  A298 );
 a79190a <=( A302  and  A300 );
 a79191a <=( a79190a  and  a79187a );
 a79192a <=( a79191a  and  a79184a );
 a79195a <=( A169  and  A170 );
 a79198a <=( A199  and  (not A168) );
 a79199a <=( a79198a  and  a79195a );
 a79202a <=( A201  and  (not A200) );
 a79205a <=( A232  and  A203 );
 a79206a <=( a79205a  and  a79202a );
 a79207a <=( a79206a  and  a79199a );
 a79210a <=( A265  and  A233 );
 a79213a <=( (not A269)  and  (not A268) );
 a79214a <=( a79213a  and  a79210a );
 a79217a <=( (not A299)  and  A298 );
 a79220a <=( A301  and  A300 );
 a79221a <=( a79220a  and  a79217a );
 a79222a <=( a79221a  and  a79214a );
 a79225a <=( A169  and  A170 );
 a79228a <=( A199  and  (not A168) );
 a79229a <=( a79228a  and  a79225a );
 a79232a <=( A201  and  (not A200) );
 a79235a <=( A232  and  A203 );
 a79236a <=( a79235a  and  a79232a );
 a79237a <=( a79236a  and  a79229a );
 a79240a <=( A265  and  A233 );
 a79243a <=( (not A269)  and  (not A268) );
 a79244a <=( a79243a  and  a79240a );
 a79247a <=( (not A299)  and  A298 );
 a79250a <=( A302  and  A300 );
 a79251a <=( a79250a  and  a79247a );
 a79252a <=( a79251a  and  a79244a );
 a79255a <=( A169  and  A170 );
 a79258a <=( A199  and  (not A168) );
 a79259a <=( a79258a  and  a79255a );
 a79262a <=( A201  and  (not A200) );
 a79265a <=( (not A233)  and  A203 );
 a79266a <=( a79265a  and  a79262a );
 a79267a <=( a79266a  and  a79259a );
 a79270a <=( (not A236)  and  (not A235) );
 a79273a <=( A266  and  A265 );
 a79274a <=( a79273a  and  a79270a );
 a79277a <=( (not A299)  and  A298 );
 a79280a <=( A301  and  A300 );
 a79281a <=( a79280a  and  a79277a );
 a79282a <=( a79281a  and  a79274a );
 a79285a <=( A169  and  A170 );
 a79288a <=( A199  and  (not A168) );
 a79289a <=( a79288a  and  a79285a );
 a79292a <=( A201  and  (not A200) );
 a79295a <=( (not A233)  and  A203 );
 a79296a <=( a79295a  and  a79292a );
 a79297a <=( a79296a  and  a79289a );
 a79300a <=( (not A236)  and  (not A235) );
 a79303a <=( A266  and  A265 );
 a79304a <=( a79303a  and  a79300a );
 a79307a <=( (not A299)  and  A298 );
 a79310a <=( A302  and  A300 );
 a79311a <=( a79310a  and  a79307a );
 a79312a <=( a79311a  and  a79304a );
 a79315a <=( A169  and  A170 );
 a79318a <=( A199  and  (not A168) );
 a79319a <=( a79318a  and  a79315a );
 a79322a <=( A201  and  (not A200) );
 a79325a <=( (not A233)  and  A203 );
 a79326a <=( a79325a  and  a79322a );
 a79327a <=( a79326a  and  a79319a );
 a79330a <=( (not A236)  and  (not A235) );
 a79333a <=( (not A267)  and  (not A266) );
 a79334a <=( a79333a  and  a79330a );
 a79337a <=( (not A299)  and  A298 );
 a79340a <=( A301  and  A300 );
 a79341a <=( a79340a  and  a79337a );
 a79342a <=( a79341a  and  a79334a );
 a79345a <=( A169  and  A170 );
 a79348a <=( A199  and  (not A168) );
 a79349a <=( a79348a  and  a79345a );
 a79352a <=( A201  and  (not A200) );
 a79355a <=( (not A233)  and  A203 );
 a79356a <=( a79355a  and  a79352a );
 a79357a <=( a79356a  and  a79349a );
 a79360a <=( (not A236)  and  (not A235) );
 a79363a <=( (not A267)  and  (not A266) );
 a79364a <=( a79363a  and  a79360a );
 a79367a <=( (not A299)  and  A298 );
 a79370a <=( A302  and  A300 );
 a79371a <=( a79370a  and  a79367a );
 a79372a <=( a79371a  and  a79364a );
 a79375a <=( A169  and  A170 );
 a79378a <=( A199  and  (not A168) );
 a79379a <=( a79378a  and  a79375a );
 a79382a <=( A201  and  (not A200) );
 a79385a <=( (not A233)  and  A203 );
 a79386a <=( a79385a  and  a79382a );
 a79387a <=( a79386a  and  a79379a );
 a79390a <=( (not A236)  and  (not A235) );
 a79393a <=( (not A266)  and  (not A265) );
 a79394a <=( a79393a  and  a79390a );
 a79397a <=( (not A299)  and  A298 );
 a79400a <=( A301  and  A300 );
 a79401a <=( a79400a  and  a79397a );
 a79402a <=( a79401a  and  a79394a );
 a79405a <=( A169  and  A170 );
 a79408a <=( A199  and  (not A168) );
 a79409a <=( a79408a  and  a79405a );
 a79412a <=( A201  and  (not A200) );
 a79415a <=( (not A233)  and  A203 );
 a79416a <=( a79415a  and  a79412a );
 a79417a <=( a79416a  and  a79409a );
 a79420a <=( (not A236)  and  (not A235) );
 a79423a <=( (not A266)  and  (not A265) );
 a79424a <=( a79423a  and  a79420a );
 a79427a <=( (not A299)  and  A298 );
 a79430a <=( A302  and  A300 );
 a79431a <=( a79430a  and  a79427a );
 a79432a <=( a79431a  and  a79424a );
 a79435a <=( A169  and  A170 );
 a79438a <=( A166  and  (not A168) );
 a79439a <=( a79438a  and  a79435a );
 a79442a <=( (not A200)  and  A199 );
 a79445a <=( A202  and  A201 );
 a79446a <=( a79445a  and  a79442a );
 a79447a <=( a79446a  and  a79439a );
 a79450a <=( (not A234)  and  (not A233) );
 a79453a <=( (not A267)  and  (not A266) );
 a79454a <=( a79453a  and  a79450a );
 a79457a <=( (not A299)  and  A298 );
 a79460a <=( A301  and  A300 );
 a79461a <=( a79460a  and  a79457a );
 a79462a <=( a79461a  and  a79454a );
 a79465a <=( A169  and  A170 );
 a79468a <=( A166  and  (not A168) );
 a79469a <=( a79468a  and  a79465a );
 a79472a <=( (not A200)  and  A199 );
 a79475a <=( A202  and  A201 );
 a79476a <=( a79475a  and  a79472a );
 a79477a <=( a79476a  and  a79469a );
 a79480a <=( (not A234)  and  (not A233) );
 a79483a <=( (not A267)  and  (not A266) );
 a79484a <=( a79483a  and  a79480a );
 a79487a <=( (not A299)  and  A298 );
 a79490a <=( A302  and  A300 );
 a79491a <=( a79490a  and  a79487a );
 a79492a <=( a79491a  and  a79484a );
 a79495a <=( A169  and  A170 );
 a79498a <=( A166  and  (not A168) );
 a79499a <=( a79498a  and  a79495a );
 a79502a <=( (not A200)  and  A199 );
 a79505a <=( A202  and  A201 );
 a79506a <=( a79505a  and  a79502a );
 a79507a <=( a79506a  and  a79499a );
 a79510a <=( (not A234)  and  (not A233) );
 a79513a <=( (not A266)  and  (not A265) );
 a79514a <=( a79513a  and  a79510a );
 a79517a <=( (not A299)  and  A298 );
 a79520a <=( A301  and  A300 );
 a79521a <=( a79520a  and  a79517a );
 a79522a <=( a79521a  and  a79514a );
 a79525a <=( A169  and  A170 );
 a79528a <=( A166  and  (not A168) );
 a79529a <=( a79528a  and  a79525a );
 a79532a <=( (not A200)  and  A199 );
 a79535a <=( A202  and  A201 );
 a79536a <=( a79535a  and  a79532a );
 a79537a <=( a79536a  and  a79529a );
 a79540a <=( (not A234)  and  (not A233) );
 a79543a <=( (not A266)  and  (not A265) );
 a79544a <=( a79543a  and  a79540a );
 a79547a <=( (not A299)  and  A298 );
 a79550a <=( A302  and  A300 );
 a79551a <=( a79550a  and  a79547a );
 a79552a <=( a79551a  and  a79544a );
 a79555a <=( A169  and  A170 );
 a79558a <=( A166  and  (not A168) );
 a79559a <=( a79558a  and  a79555a );
 a79562a <=( (not A200)  and  A199 );
 a79565a <=( A202  and  A201 );
 a79566a <=( a79565a  and  a79562a );
 a79567a <=( a79566a  and  a79559a );
 a79570a <=( (not A233)  and  (not A232) );
 a79573a <=( (not A267)  and  (not A266) );
 a79574a <=( a79573a  and  a79570a );
 a79577a <=( (not A299)  and  A298 );
 a79580a <=( A301  and  A300 );
 a79581a <=( a79580a  and  a79577a );
 a79582a <=( a79581a  and  a79574a );
 a79585a <=( A169  and  A170 );
 a79588a <=( A166  and  (not A168) );
 a79589a <=( a79588a  and  a79585a );
 a79592a <=( (not A200)  and  A199 );
 a79595a <=( A202  and  A201 );
 a79596a <=( a79595a  and  a79592a );
 a79597a <=( a79596a  and  a79589a );
 a79600a <=( (not A233)  and  (not A232) );
 a79603a <=( (not A267)  and  (not A266) );
 a79604a <=( a79603a  and  a79600a );
 a79607a <=( (not A299)  and  A298 );
 a79610a <=( A302  and  A300 );
 a79611a <=( a79610a  and  a79607a );
 a79612a <=( a79611a  and  a79604a );
 a79615a <=( A169  and  A170 );
 a79618a <=( A166  and  (not A168) );
 a79619a <=( a79618a  and  a79615a );
 a79622a <=( (not A200)  and  A199 );
 a79625a <=( A202  and  A201 );
 a79626a <=( a79625a  and  a79622a );
 a79627a <=( a79626a  and  a79619a );
 a79630a <=( (not A233)  and  (not A232) );
 a79633a <=( (not A266)  and  (not A265) );
 a79634a <=( a79633a  and  a79630a );
 a79637a <=( (not A299)  and  A298 );
 a79640a <=( A301  and  A300 );
 a79641a <=( a79640a  and  a79637a );
 a79642a <=( a79641a  and  a79634a );
 a79645a <=( A169  and  A170 );
 a79648a <=( A166  and  (not A168) );
 a79649a <=( a79648a  and  a79645a );
 a79652a <=( (not A200)  and  A199 );
 a79655a <=( A202  and  A201 );
 a79656a <=( a79655a  and  a79652a );
 a79657a <=( a79656a  and  a79649a );
 a79660a <=( (not A233)  and  (not A232) );
 a79663a <=( (not A266)  and  (not A265) );
 a79664a <=( a79663a  and  a79660a );
 a79667a <=( (not A299)  and  A298 );
 a79670a <=( A302  and  A300 );
 a79671a <=( a79670a  and  a79667a );
 a79672a <=( a79671a  and  a79664a );
 a79675a <=( A169  and  A170 );
 a79678a <=( A166  and  (not A168) );
 a79679a <=( a79678a  and  a79675a );
 a79682a <=( (not A200)  and  A199 );
 a79685a <=( A203  and  A201 );
 a79686a <=( a79685a  and  a79682a );
 a79687a <=( a79686a  and  a79679a );
 a79690a <=( (not A234)  and  (not A233) );
 a79693a <=( (not A267)  and  (not A266) );
 a79694a <=( a79693a  and  a79690a );
 a79697a <=( (not A299)  and  A298 );
 a79700a <=( A301  and  A300 );
 a79701a <=( a79700a  and  a79697a );
 a79702a <=( a79701a  and  a79694a );
 a79705a <=( A169  and  A170 );
 a79708a <=( A166  and  (not A168) );
 a79709a <=( a79708a  and  a79705a );
 a79712a <=( (not A200)  and  A199 );
 a79715a <=( A203  and  A201 );
 a79716a <=( a79715a  and  a79712a );
 a79717a <=( a79716a  and  a79709a );
 a79720a <=( (not A234)  and  (not A233) );
 a79723a <=( (not A267)  and  (not A266) );
 a79724a <=( a79723a  and  a79720a );
 a79727a <=( (not A299)  and  A298 );
 a79730a <=( A302  and  A300 );
 a79731a <=( a79730a  and  a79727a );
 a79732a <=( a79731a  and  a79724a );
 a79735a <=( A169  and  A170 );
 a79738a <=( A166  and  (not A168) );
 a79739a <=( a79738a  and  a79735a );
 a79742a <=( (not A200)  and  A199 );
 a79745a <=( A203  and  A201 );
 a79746a <=( a79745a  and  a79742a );
 a79747a <=( a79746a  and  a79739a );
 a79750a <=( (not A234)  and  (not A233) );
 a79753a <=( (not A266)  and  (not A265) );
 a79754a <=( a79753a  and  a79750a );
 a79757a <=( (not A299)  and  A298 );
 a79760a <=( A301  and  A300 );
 a79761a <=( a79760a  and  a79757a );
 a79762a <=( a79761a  and  a79754a );
 a79765a <=( A169  and  A170 );
 a79768a <=( A166  and  (not A168) );
 a79769a <=( a79768a  and  a79765a );
 a79772a <=( (not A200)  and  A199 );
 a79775a <=( A203  and  A201 );
 a79776a <=( a79775a  and  a79772a );
 a79777a <=( a79776a  and  a79769a );
 a79780a <=( (not A234)  and  (not A233) );
 a79783a <=( (not A266)  and  (not A265) );
 a79784a <=( a79783a  and  a79780a );
 a79787a <=( (not A299)  and  A298 );
 a79790a <=( A302  and  A300 );
 a79791a <=( a79790a  and  a79787a );
 a79792a <=( a79791a  and  a79784a );
 a79795a <=( A169  and  A170 );
 a79798a <=( A166  and  (not A168) );
 a79799a <=( a79798a  and  a79795a );
 a79802a <=( (not A200)  and  A199 );
 a79805a <=( A203  and  A201 );
 a79806a <=( a79805a  and  a79802a );
 a79807a <=( a79806a  and  a79799a );
 a79810a <=( (not A233)  and  (not A232) );
 a79813a <=( (not A267)  and  (not A266) );
 a79814a <=( a79813a  and  a79810a );
 a79817a <=( (not A299)  and  A298 );
 a79820a <=( A301  and  A300 );
 a79821a <=( a79820a  and  a79817a );
 a79822a <=( a79821a  and  a79814a );
 a79825a <=( A169  and  A170 );
 a79828a <=( A166  and  (not A168) );
 a79829a <=( a79828a  and  a79825a );
 a79832a <=( (not A200)  and  A199 );
 a79835a <=( A203  and  A201 );
 a79836a <=( a79835a  and  a79832a );
 a79837a <=( a79836a  and  a79829a );
 a79840a <=( (not A233)  and  (not A232) );
 a79843a <=( (not A267)  and  (not A266) );
 a79844a <=( a79843a  and  a79840a );
 a79847a <=( (not A299)  and  A298 );
 a79850a <=( A302  and  A300 );
 a79851a <=( a79850a  and  a79847a );
 a79852a <=( a79851a  and  a79844a );
 a79855a <=( A169  and  A170 );
 a79858a <=( A166  and  (not A168) );
 a79859a <=( a79858a  and  a79855a );
 a79862a <=( (not A200)  and  A199 );
 a79865a <=( A203  and  A201 );
 a79866a <=( a79865a  and  a79862a );
 a79867a <=( a79866a  and  a79859a );
 a79870a <=( (not A233)  and  (not A232) );
 a79873a <=( (not A266)  and  (not A265) );
 a79874a <=( a79873a  and  a79870a );
 a79877a <=( (not A299)  and  A298 );
 a79880a <=( A301  and  A300 );
 a79881a <=( a79880a  and  a79877a );
 a79882a <=( a79881a  and  a79874a );
 a79885a <=( A169  and  A170 );
 a79888a <=( A166  and  (not A168) );
 a79889a <=( a79888a  and  a79885a );
 a79892a <=( (not A200)  and  A199 );
 a79895a <=( A203  and  A201 );
 a79896a <=( a79895a  and  a79892a );
 a79897a <=( a79896a  and  a79889a );
 a79900a <=( (not A233)  and  (not A232) );
 a79903a <=( (not A266)  and  (not A265) );
 a79904a <=( a79903a  and  a79900a );
 a79907a <=( (not A299)  and  A298 );
 a79910a <=( A302  and  A300 );
 a79911a <=( a79910a  and  a79907a );
 a79912a <=( a79911a  and  a79904a );
 a79915a <=( A169  and  (not A170) );
 a79918a <=( A166  and  A167 );
 a79919a <=( a79918a  and  a79915a );
 a79922a <=( A200  and  A199 );
 a79925a <=( (not A235)  and  (not A233) );
 a79926a <=( a79925a  and  a79922a );
 a79927a <=( a79926a  and  a79919a );
 a79930a <=( (not A266)  and  (not A236) );
 a79933a <=( (not A269)  and  (not A268) );
 a79934a <=( a79933a  and  a79930a );
 a79937a <=( (not A299)  and  A298 );
 a79940a <=( A301  and  A300 );
 a79941a <=( a79940a  and  a79937a );
 a79942a <=( a79941a  and  a79934a );
 a79945a <=( A169  and  (not A170) );
 a79948a <=( A166  and  A167 );
 a79949a <=( a79948a  and  a79945a );
 a79952a <=( A200  and  A199 );
 a79955a <=( (not A235)  and  (not A233) );
 a79956a <=( a79955a  and  a79952a );
 a79957a <=( a79956a  and  a79949a );
 a79960a <=( (not A266)  and  (not A236) );
 a79963a <=( (not A269)  and  (not A268) );
 a79964a <=( a79963a  and  a79960a );
 a79967a <=( (not A299)  and  A298 );
 a79970a <=( A302  and  A300 );
 a79971a <=( a79970a  and  a79967a );
 a79972a <=( a79971a  and  a79964a );
 a79975a <=( A169  and  (not A170) );
 a79978a <=( A166  and  A167 );
 a79979a <=( a79978a  and  a79975a );
 a79982a <=( (not A202)  and  (not A200) );
 a79985a <=( A232  and  (not A203) );
 a79986a <=( a79985a  and  a79982a );
 a79987a <=( a79986a  and  a79979a );
 a79990a <=( A265  and  A233 );
 a79993a <=( (not A269)  and  (not A268) );
 a79994a <=( a79993a  and  a79990a );
 a79997a <=( (not A299)  and  A298 );
 a80000a <=( A301  and  A300 );
 a80001a <=( a80000a  and  a79997a );
 a80002a <=( a80001a  and  a79994a );
 a80005a <=( A169  and  (not A170) );
 a80008a <=( A166  and  A167 );
 a80009a <=( a80008a  and  a80005a );
 a80012a <=( (not A202)  and  (not A200) );
 a80015a <=( A232  and  (not A203) );
 a80016a <=( a80015a  and  a80012a );
 a80017a <=( a80016a  and  a80009a );
 a80020a <=( A265  and  A233 );
 a80023a <=( (not A269)  and  (not A268) );
 a80024a <=( a80023a  and  a80020a );
 a80027a <=( (not A299)  and  A298 );
 a80030a <=( A302  and  A300 );
 a80031a <=( a80030a  and  a80027a );
 a80032a <=( a80031a  and  a80024a );
 a80035a <=( A169  and  (not A170) );
 a80038a <=( A166  and  A167 );
 a80039a <=( a80038a  and  a80035a );
 a80042a <=( (not A202)  and  (not A200) );
 a80045a <=( (not A233)  and  (not A203) );
 a80046a <=( a80045a  and  a80042a );
 a80047a <=( a80046a  and  a80039a );
 a80050a <=( (not A236)  and  (not A235) );
 a80053a <=( A266  and  A265 );
 a80054a <=( a80053a  and  a80050a );
 a80057a <=( (not A299)  and  A298 );
 a80060a <=( A301  and  A300 );
 a80061a <=( a80060a  and  a80057a );
 a80062a <=( a80061a  and  a80054a );
 a80065a <=( A169  and  (not A170) );
 a80068a <=( A166  and  A167 );
 a80069a <=( a80068a  and  a80065a );
 a80072a <=( (not A202)  and  (not A200) );
 a80075a <=( (not A233)  and  (not A203) );
 a80076a <=( a80075a  and  a80072a );
 a80077a <=( a80076a  and  a80069a );
 a80080a <=( (not A236)  and  (not A235) );
 a80083a <=( A266  and  A265 );
 a80084a <=( a80083a  and  a80080a );
 a80087a <=( (not A299)  and  A298 );
 a80090a <=( A302  and  A300 );
 a80091a <=( a80090a  and  a80087a );
 a80092a <=( a80091a  and  a80084a );
 a80095a <=( A169  and  (not A170) );
 a80098a <=( A166  and  A167 );
 a80099a <=( a80098a  and  a80095a );
 a80102a <=( (not A202)  and  (not A200) );
 a80105a <=( (not A233)  and  (not A203) );
 a80106a <=( a80105a  and  a80102a );
 a80107a <=( a80106a  and  a80099a );
 a80110a <=( (not A236)  and  (not A235) );
 a80113a <=( (not A267)  and  (not A266) );
 a80114a <=( a80113a  and  a80110a );
 a80117a <=( (not A299)  and  A298 );
 a80120a <=( A301  and  A300 );
 a80121a <=( a80120a  and  a80117a );
 a80122a <=( a80121a  and  a80114a );
 a80125a <=( A169  and  (not A170) );
 a80128a <=( A166  and  A167 );
 a80129a <=( a80128a  and  a80125a );
 a80132a <=( (not A202)  and  (not A200) );
 a80135a <=( (not A233)  and  (not A203) );
 a80136a <=( a80135a  and  a80132a );
 a80137a <=( a80136a  and  a80129a );
 a80140a <=( (not A236)  and  (not A235) );
 a80143a <=( (not A267)  and  (not A266) );
 a80144a <=( a80143a  and  a80140a );
 a80147a <=( (not A299)  and  A298 );
 a80150a <=( A302  and  A300 );
 a80151a <=( a80150a  and  a80147a );
 a80152a <=( a80151a  and  a80144a );
 a80155a <=( A169  and  (not A170) );
 a80158a <=( A166  and  A167 );
 a80159a <=( a80158a  and  a80155a );
 a80162a <=( (not A202)  and  (not A200) );
 a80165a <=( (not A233)  and  (not A203) );
 a80166a <=( a80165a  and  a80162a );
 a80167a <=( a80166a  and  a80159a );
 a80170a <=( (not A236)  and  (not A235) );
 a80173a <=( (not A266)  and  (not A265) );
 a80174a <=( a80173a  and  a80170a );
 a80177a <=( (not A299)  and  A298 );
 a80180a <=( A301  and  A300 );
 a80181a <=( a80180a  and  a80177a );
 a80182a <=( a80181a  and  a80174a );
 a80185a <=( A169  and  (not A170) );
 a80188a <=( A166  and  A167 );
 a80189a <=( a80188a  and  a80185a );
 a80192a <=( (not A202)  and  (not A200) );
 a80195a <=( (not A233)  and  (not A203) );
 a80196a <=( a80195a  and  a80192a );
 a80197a <=( a80196a  and  a80189a );
 a80200a <=( (not A236)  and  (not A235) );
 a80203a <=( (not A266)  and  (not A265) );
 a80204a <=( a80203a  and  a80200a );
 a80207a <=( (not A299)  and  A298 );
 a80210a <=( A302  and  A300 );
 a80211a <=( a80210a  and  a80207a );
 a80212a <=( a80211a  and  a80204a );
 a80215a <=( A169  and  (not A170) );
 a80218a <=( A166  and  A167 );
 a80219a <=( a80218a  and  a80215a );
 a80222a <=( (not A202)  and  (not A200) );
 a80225a <=( (not A233)  and  (not A203) );
 a80226a <=( a80225a  and  a80222a );
 a80227a <=( a80226a  and  a80219a );
 a80230a <=( (not A266)  and  (not A234) );
 a80233a <=( (not A269)  and  (not A268) );
 a80234a <=( a80233a  and  a80230a );
 a80237a <=( (not A299)  and  A298 );
 a80240a <=( A301  and  A300 );
 a80241a <=( a80240a  and  a80237a );
 a80242a <=( a80241a  and  a80234a );
 a80245a <=( A169  and  (not A170) );
 a80248a <=( A166  and  A167 );
 a80249a <=( a80248a  and  a80245a );
 a80252a <=( (not A202)  and  (not A200) );
 a80255a <=( (not A233)  and  (not A203) );
 a80256a <=( a80255a  and  a80252a );
 a80257a <=( a80256a  and  a80249a );
 a80260a <=( (not A266)  and  (not A234) );
 a80263a <=( (not A269)  and  (not A268) );
 a80264a <=( a80263a  and  a80260a );
 a80267a <=( (not A299)  and  A298 );
 a80270a <=( A302  and  A300 );
 a80271a <=( a80270a  and  a80267a );
 a80272a <=( a80271a  and  a80264a );
 a80275a <=( A169  and  (not A170) );
 a80278a <=( A166  and  A167 );
 a80279a <=( a80278a  and  a80275a );
 a80282a <=( (not A202)  and  (not A200) );
 a80285a <=( (not A232)  and  (not A203) );
 a80286a <=( a80285a  and  a80282a );
 a80287a <=( a80286a  and  a80279a );
 a80290a <=( (not A266)  and  (not A233) );
 a80293a <=( (not A269)  and  (not A268) );
 a80294a <=( a80293a  and  a80290a );
 a80297a <=( (not A299)  and  A298 );
 a80300a <=( A301  and  A300 );
 a80301a <=( a80300a  and  a80297a );
 a80302a <=( a80301a  and  a80294a );
 a80305a <=( A169  and  (not A170) );
 a80308a <=( A166  and  A167 );
 a80309a <=( a80308a  and  a80305a );
 a80312a <=( (not A202)  and  (not A200) );
 a80315a <=( (not A232)  and  (not A203) );
 a80316a <=( a80315a  and  a80312a );
 a80317a <=( a80316a  and  a80309a );
 a80320a <=( (not A266)  and  (not A233) );
 a80323a <=( (not A269)  and  (not A268) );
 a80324a <=( a80323a  and  a80320a );
 a80327a <=( (not A299)  and  A298 );
 a80330a <=( A302  and  A300 );
 a80331a <=( a80330a  and  a80327a );
 a80332a <=( a80331a  and  a80324a );
 a80335a <=( A169  and  (not A170) );
 a80338a <=( A166  and  A167 );
 a80339a <=( a80338a  and  a80335a );
 a80342a <=( (not A201)  and  (not A200) );
 a80345a <=( (not A235)  and  (not A233) );
 a80346a <=( a80345a  and  a80342a );
 a80347a <=( a80346a  and  a80339a );
 a80350a <=( (not A266)  and  (not A236) );
 a80353a <=( (not A269)  and  (not A268) );
 a80354a <=( a80353a  and  a80350a );
 a80357a <=( (not A299)  and  A298 );
 a80360a <=( A301  and  A300 );
 a80361a <=( a80360a  and  a80357a );
 a80362a <=( a80361a  and  a80354a );
 a80365a <=( A169  and  (not A170) );
 a80368a <=( A166  and  A167 );
 a80369a <=( a80368a  and  a80365a );
 a80372a <=( (not A201)  and  (not A200) );
 a80375a <=( (not A235)  and  (not A233) );
 a80376a <=( a80375a  and  a80372a );
 a80377a <=( a80376a  and  a80369a );
 a80380a <=( (not A266)  and  (not A236) );
 a80383a <=( (not A269)  and  (not A268) );
 a80384a <=( a80383a  and  a80380a );
 a80387a <=( (not A299)  and  A298 );
 a80390a <=( A302  and  A300 );
 a80391a <=( a80390a  and  a80387a );
 a80392a <=( a80391a  and  a80384a );
 a80395a <=( A169  and  (not A170) );
 a80398a <=( A166  and  A167 );
 a80399a <=( a80398a  and  a80395a );
 a80402a <=( (not A200)  and  (not A199) );
 a80405a <=( (not A235)  and  (not A233) );
 a80406a <=( a80405a  and  a80402a );
 a80407a <=( a80406a  and  a80399a );
 a80410a <=( (not A266)  and  (not A236) );
 a80413a <=( (not A269)  and  (not A268) );
 a80414a <=( a80413a  and  a80410a );
 a80417a <=( (not A299)  and  A298 );
 a80420a <=( A301  and  A300 );
 a80421a <=( a80420a  and  a80417a );
 a80422a <=( a80421a  and  a80414a );
 a80425a <=( A169  and  (not A170) );
 a80428a <=( A166  and  A167 );
 a80429a <=( a80428a  and  a80425a );
 a80432a <=( (not A200)  and  (not A199) );
 a80435a <=( (not A235)  and  (not A233) );
 a80436a <=( a80435a  and  a80432a );
 a80437a <=( a80436a  and  a80429a );
 a80440a <=( (not A266)  and  (not A236) );
 a80443a <=( (not A269)  and  (not A268) );
 a80444a <=( a80443a  and  a80440a );
 a80447a <=( (not A299)  and  A298 );
 a80450a <=( A302  and  A300 );
 a80451a <=( a80450a  and  a80447a );
 a80452a <=( a80451a  and  a80444a );
 a80455a <=( A169  and  (not A170) );
 a80458a <=( (not A166)  and  (not A167) );
 a80459a <=( a80458a  and  a80455a );
 a80462a <=( A200  and  A199 );
 a80465a <=( (not A235)  and  (not A233) );
 a80466a <=( a80465a  and  a80462a );
 a80467a <=( a80466a  and  a80459a );
 a80470a <=( (not A266)  and  (not A236) );
 a80473a <=( (not A269)  and  (not A268) );
 a80474a <=( a80473a  and  a80470a );
 a80477a <=( (not A299)  and  A298 );
 a80480a <=( A301  and  A300 );
 a80481a <=( a80480a  and  a80477a );
 a80482a <=( a80481a  and  a80474a );
 a80485a <=( A169  and  (not A170) );
 a80488a <=( (not A166)  and  (not A167) );
 a80489a <=( a80488a  and  a80485a );
 a80492a <=( A200  and  A199 );
 a80495a <=( (not A235)  and  (not A233) );
 a80496a <=( a80495a  and  a80492a );
 a80497a <=( a80496a  and  a80489a );
 a80500a <=( (not A266)  and  (not A236) );
 a80503a <=( (not A269)  and  (not A268) );
 a80504a <=( a80503a  and  a80500a );
 a80507a <=( (not A299)  and  A298 );
 a80510a <=( A302  and  A300 );
 a80511a <=( a80510a  and  a80507a );
 a80512a <=( a80511a  and  a80504a );
 a80515a <=( A169  and  (not A170) );
 a80518a <=( (not A166)  and  (not A167) );
 a80519a <=( a80518a  and  a80515a );
 a80522a <=( (not A202)  and  (not A200) );
 a80525a <=( A232  and  (not A203) );
 a80526a <=( a80525a  and  a80522a );
 a80527a <=( a80526a  and  a80519a );
 a80530a <=( A265  and  A233 );
 a80533a <=( (not A269)  and  (not A268) );
 a80534a <=( a80533a  and  a80530a );
 a80537a <=( (not A299)  and  A298 );
 a80540a <=( A301  and  A300 );
 a80541a <=( a80540a  and  a80537a );
 a80542a <=( a80541a  and  a80534a );
 a80545a <=( A169  and  (not A170) );
 a80548a <=( (not A166)  and  (not A167) );
 a80549a <=( a80548a  and  a80545a );
 a80552a <=( (not A202)  and  (not A200) );
 a80555a <=( A232  and  (not A203) );
 a80556a <=( a80555a  and  a80552a );
 a80557a <=( a80556a  and  a80549a );
 a80560a <=( A265  and  A233 );
 a80563a <=( (not A269)  and  (not A268) );
 a80564a <=( a80563a  and  a80560a );
 a80567a <=( (not A299)  and  A298 );
 a80570a <=( A302  and  A300 );
 a80571a <=( a80570a  and  a80567a );
 a80572a <=( a80571a  and  a80564a );
 a80575a <=( A169  and  (not A170) );
 a80578a <=( (not A166)  and  (not A167) );
 a80579a <=( a80578a  and  a80575a );
 a80582a <=( (not A202)  and  (not A200) );
 a80585a <=( (not A233)  and  (not A203) );
 a80586a <=( a80585a  and  a80582a );
 a80587a <=( a80586a  and  a80579a );
 a80590a <=( (not A236)  and  (not A235) );
 a80593a <=( A266  and  A265 );
 a80594a <=( a80593a  and  a80590a );
 a80597a <=( (not A299)  and  A298 );
 a80600a <=( A301  and  A300 );
 a80601a <=( a80600a  and  a80597a );
 a80602a <=( a80601a  and  a80594a );
 a80605a <=( A169  and  (not A170) );
 a80608a <=( (not A166)  and  (not A167) );
 a80609a <=( a80608a  and  a80605a );
 a80612a <=( (not A202)  and  (not A200) );
 a80615a <=( (not A233)  and  (not A203) );
 a80616a <=( a80615a  and  a80612a );
 a80617a <=( a80616a  and  a80609a );
 a80620a <=( (not A236)  and  (not A235) );
 a80623a <=( A266  and  A265 );
 a80624a <=( a80623a  and  a80620a );
 a80627a <=( (not A299)  and  A298 );
 a80630a <=( A302  and  A300 );
 a80631a <=( a80630a  and  a80627a );
 a80632a <=( a80631a  and  a80624a );
 a80635a <=( A169  and  (not A170) );
 a80638a <=( (not A166)  and  (not A167) );
 a80639a <=( a80638a  and  a80635a );
 a80642a <=( (not A202)  and  (not A200) );
 a80645a <=( (not A233)  and  (not A203) );
 a80646a <=( a80645a  and  a80642a );
 a80647a <=( a80646a  and  a80639a );
 a80650a <=( (not A236)  and  (not A235) );
 a80653a <=( (not A267)  and  (not A266) );
 a80654a <=( a80653a  and  a80650a );
 a80657a <=( (not A299)  and  A298 );
 a80660a <=( A301  and  A300 );
 a80661a <=( a80660a  and  a80657a );
 a80662a <=( a80661a  and  a80654a );
 a80665a <=( A169  and  (not A170) );
 a80668a <=( (not A166)  and  (not A167) );
 a80669a <=( a80668a  and  a80665a );
 a80672a <=( (not A202)  and  (not A200) );
 a80675a <=( (not A233)  and  (not A203) );
 a80676a <=( a80675a  and  a80672a );
 a80677a <=( a80676a  and  a80669a );
 a80680a <=( (not A236)  and  (not A235) );
 a80683a <=( (not A267)  and  (not A266) );
 a80684a <=( a80683a  and  a80680a );
 a80687a <=( (not A299)  and  A298 );
 a80690a <=( A302  and  A300 );
 a80691a <=( a80690a  and  a80687a );
 a80692a <=( a80691a  and  a80684a );
 a80695a <=( A169  and  (not A170) );
 a80698a <=( (not A166)  and  (not A167) );
 a80699a <=( a80698a  and  a80695a );
 a80702a <=( (not A202)  and  (not A200) );
 a80705a <=( (not A233)  and  (not A203) );
 a80706a <=( a80705a  and  a80702a );
 a80707a <=( a80706a  and  a80699a );
 a80710a <=( (not A236)  and  (not A235) );
 a80713a <=( (not A266)  and  (not A265) );
 a80714a <=( a80713a  and  a80710a );
 a80717a <=( (not A299)  and  A298 );
 a80720a <=( A301  and  A300 );
 a80721a <=( a80720a  and  a80717a );
 a80722a <=( a80721a  and  a80714a );
 a80725a <=( A169  and  (not A170) );
 a80728a <=( (not A166)  and  (not A167) );
 a80729a <=( a80728a  and  a80725a );
 a80732a <=( (not A202)  and  (not A200) );
 a80735a <=( (not A233)  and  (not A203) );
 a80736a <=( a80735a  and  a80732a );
 a80737a <=( a80736a  and  a80729a );
 a80740a <=( (not A236)  and  (not A235) );
 a80743a <=( (not A266)  and  (not A265) );
 a80744a <=( a80743a  and  a80740a );
 a80747a <=( (not A299)  and  A298 );
 a80750a <=( A302  and  A300 );
 a80751a <=( a80750a  and  a80747a );
 a80752a <=( a80751a  and  a80744a );
 a80755a <=( A169  and  (not A170) );
 a80758a <=( (not A166)  and  (not A167) );
 a80759a <=( a80758a  and  a80755a );
 a80762a <=( (not A202)  and  (not A200) );
 a80765a <=( (not A233)  and  (not A203) );
 a80766a <=( a80765a  and  a80762a );
 a80767a <=( a80766a  and  a80759a );
 a80770a <=( (not A266)  and  (not A234) );
 a80773a <=( (not A269)  and  (not A268) );
 a80774a <=( a80773a  and  a80770a );
 a80777a <=( (not A299)  and  A298 );
 a80780a <=( A301  and  A300 );
 a80781a <=( a80780a  and  a80777a );
 a80782a <=( a80781a  and  a80774a );
 a80785a <=( A169  and  (not A170) );
 a80788a <=( (not A166)  and  (not A167) );
 a80789a <=( a80788a  and  a80785a );
 a80792a <=( (not A202)  and  (not A200) );
 a80795a <=( (not A233)  and  (not A203) );
 a80796a <=( a80795a  and  a80792a );
 a80797a <=( a80796a  and  a80789a );
 a80800a <=( (not A266)  and  (not A234) );
 a80803a <=( (not A269)  and  (not A268) );
 a80804a <=( a80803a  and  a80800a );
 a80807a <=( (not A299)  and  A298 );
 a80810a <=( A302  and  A300 );
 a80811a <=( a80810a  and  a80807a );
 a80812a <=( a80811a  and  a80804a );
 a80815a <=( A169  and  (not A170) );
 a80818a <=( (not A166)  and  (not A167) );
 a80819a <=( a80818a  and  a80815a );
 a80822a <=( (not A202)  and  (not A200) );
 a80825a <=( (not A232)  and  (not A203) );
 a80826a <=( a80825a  and  a80822a );
 a80827a <=( a80826a  and  a80819a );
 a80830a <=( (not A266)  and  (not A233) );
 a80833a <=( (not A269)  and  (not A268) );
 a80834a <=( a80833a  and  a80830a );
 a80837a <=( (not A299)  and  A298 );
 a80840a <=( A301  and  A300 );
 a80841a <=( a80840a  and  a80837a );
 a80842a <=( a80841a  and  a80834a );
 a80845a <=( A169  and  (not A170) );
 a80848a <=( (not A166)  and  (not A167) );
 a80849a <=( a80848a  and  a80845a );
 a80852a <=( (not A202)  and  (not A200) );
 a80855a <=( (not A232)  and  (not A203) );
 a80856a <=( a80855a  and  a80852a );
 a80857a <=( a80856a  and  a80849a );
 a80860a <=( (not A266)  and  (not A233) );
 a80863a <=( (not A269)  and  (not A268) );
 a80864a <=( a80863a  and  a80860a );
 a80867a <=( (not A299)  and  A298 );
 a80870a <=( A302  and  A300 );
 a80871a <=( a80870a  and  a80867a );
 a80872a <=( a80871a  and  a80864a );
 a80875a <=( A169  and  (not A170) );
 a80878a <=( (not A166)  and  (not A167) );
 a80879a <=( a80878a  and  a80875a );
 a80882a <=( (not A201)  and  (not A200) );
 a80885a <=( (not A235)  and  (not A233) );
 a80886a <=( a80885a  and  a80882a );
 a80887a <=( a80886a  and  a80879a );
 a80890a <=( (not A266)  and  (not A236) );
 a80893a <=( (not A269)  and  (not A268) );
 a80894a <=( a80893a  and  a80890a );
 a80897a <=( (not A299)  and  A298 );
 a80900a <=( A301  and  A300 );
 a80901a <=( a80900a  and  a80897a );
 a80902a <=( a80901a  and  a80894a );
 a80905a <=( A169  and  (not A170) );
 a80908a <=( (not A166)  and  (not A167) );
 a80909a <=( a80908a  and  a80905a );
 a80912a <=( (not A201)  and  (not A200) );
 a80915a <=( (not A235)  and  (not A233) );
 a80916a <=( a80915a  and  a80912a );
 a80917a <=( a80916a  and  a80909a );
 a80920a <=( (not A266)  and  (not A236) );
 a80923a <=( (not A269)  and  (not A268) );
 a80924a <=( a80923a  and  a80920a );
 a80927a <=( (not A299)  and  A298 );
 a80930a <=( A302  and  A300 );
 a80931a <=( a80930a  and  a80927a );
 a80932a <=( a80931a  and  a80924a );
 a80935a <=( A169  and  (not A170) );
 a80938a <=( (not A166)  and  (not A167) );
 a80939a <=( a80938a  and  a80935a );
 a80942a <=( (not A200)  and  (not A199) );
 a80945a <=( (not A235)  and  (not A233) );
 a80946a <=( a80945a  and  a80942a );
 a80947a <=( a80946a  and  a80939a );
 a80950a <=( (not A266)  and  (not A236) );
 a80953a <=( (not A269)  and  (not A268) );
 a80954a <=( a80953a  and  a80950a );
 a80957a <=( (not A299)  and  A298 );
 a80960a <=( A301  and  A300 );
 a80961a <=( a80960a  and  a80957a );
 a80962a <=( a80961a  and  a80954a );
 a80965a <=( A169  and  (not A170) );
 a80968a <=( (not A166)  and  (not A167) );
 a80969a <=( a80968a  and  a80965a );
 a80972a <=( (not A200)  and  (not A199) );
 a80975a <=( (not A235)  and  (not A233) );
 a80976a <=( a80975a  and  a80972a );
 a80977a <=( a80976a  and  a80969a );
 a80980a <=( (not A266)  and  (not A236) );
 a80983a <=( (not A269)  and  (not A268) );
 a80984a <=( a80983a  and  a80980a );
 a80987a <=( (not A299)  and  A298 );
 a80990a <=( A302  and  A300 );
 a80991a <=( a80990a  and  a80987a );
 a80992a <=( a80991a  and  a80984a );
 a80995a <=( (not A167)  and  (not A169) );
 a80998a <=( A199  and  (not A166) );
 a80999a <=( a80998a  and  a80995a );
 a81002a <=( A201  and  (not A200) );
 a81005a <=( A232  and  A202 );
 a81006a <=( a81005a  and  a81002a );
 a81007a <=( a81006a  and  a80999a );
 a81010a <=( A265  and  A233 );
 a81013a <=( (not A269)  and  (not A268) );
 a81014a <=( a81013a  and  a81010a );
 a81017a <=( (not A299)  and  A298 );
 a81020a <=( A301  and  A300 );
 a81021a <=( a81020a  and  a81017a );
 a81022a <=( a81021a  and  a81014a );
 a81025a <=( (not A167)  and  (not A169) );
 a81028a <=( A199  and  (not A166) );
 a81029a <=( a81028a  and  a81025a );
 a81032a <=( A201  and  (not A200) );
 a81035a <=( A232  and  A202 );
 a81036a <=( a81035a  and  a81032a );
 a81037a <=( a81036a  and  a81029a );
 a81040a <=( A265  and  A233 );
 a81043a <=( (not A269)  and  (not A268) );
 a81044a <=( a81043a  and  a81040a );
 a81047a <=( (not A299)  and  A298 );
 a81050a <=( A302  and  A300 );
 a81051a <=( a81050a  and  a81047a );
 a81052a <=( a81051a  and  a81044a );
 a81055a <=( (not A167)  and  (not A169) );
 a81058a <=( A199  and  (not A166) );
 a81059a <=( a81058a  and  a81055a );
 a81062a <=( A201  and  (not A200) );
 a81065a <=( (not A233)  and  A202 );
 a81066a <=( a81065a  and  a81062a );
 a81067a <=( a81066a  and  a81059a );
 a81070a <=( (not A236)  and  (not A235) );
 a81073a <=( A266  and  A265 );
 a81074a <=( a81073a  and  a81070a );
 a81077a <=( (not A299)  and  A298 );
 a81080a <=( A301  and  A300 );
 a81081a <=( a81080a  and  a81077a );
 a81082a <=( a81081a  and  a81074a );
 a81085a <=( (not A167)  and  (not A169) );
 a81088a <=( A199  and  (not A166) );
 a81089a <=( a81088a  and  a81085a );
 a81092a <=( A201  and  (not A200) );
 a81095a <=( (not A233)  and  A202 );
 a81096a <=( a81095a  and  a81092a );
 a81097a <=( a81096a  and  a81089a );
 a81100a <=( (not A236)  and  (not A235) );
 a81103a <=( A266  and  A265 );
 a81104a <=( a81103a  and  a81100a );
 a81107a <=( (not A299)  and  A298 );
 a81110a <=( A302  and  A300 );
 a81111a <=( a81110a  and  a81107a );
 a81112a <=( a81111a  and  a81104a );
 a81115a <=( (not A167)  and  (not A169) );
 a81118a <=( A199  and  (not A166) );
 a81119a <=( a81118a  and  a81115a );
 a81122a <=( A201  and  (not A200) );
 a81125a <=( (not A233)  and  A202 );
 a81126a <=( a81125a  and  a81122a );
 a81127a <=( a81126a  and  a81119a );
 a81130a <=( (not A236)  and  (not A235) );
 a81133a <=( (not A267)  and  (not A266) );
 a81134a <=( a81133a  and  a81130a );
 a81137a <=( (not A299)  and  A298 );
 a81140a <=( A301  and  A300 );
 a81141a <=( a81140a  and  a81137a );
 a81142a <=( a81141a  and  a81134a );
 a81145a <=( (not A167)  and  (not A169) );
 a81148a <=( A199  and  (not A166) );
 a81149a <=( a81148a  and  a81145a );
 a81152a <=( A201  and  (not A200) );
 a81155a <=( (not A233)  and  A202 );
 a81156a <=( a81155a  and  a81152a );
 a81157a <=( a81156a  and  a81149a );
 a81160a <=( (not A236)  and  (not A235) );
 a81163a <=( (not A267)  and  (not A266) );
 a81164a <=( a81163a  and  a81160a );
 a81167a <=( (not A299)  and  A298 );
 a81170a <=( A302  and  A300 );
 a81171a <=( a81170a  and  a81167a );
 a81172a <=( a81171a  and  a81164a );
 a81175a <=( (not A167)  and  (not A169) );
 a81178a <=( A199  and  (not A166) );
 a81179a <=( a81178a  and  a81175a );
 a81182a <=( A201  and  (not A200) );
 a81185a <=( (not A233)  and  A202 );
 a81186a <=( a81185a  and  a81182a );
 a81187a <=( a81186a  and  a81179a );
 a81190a <=( (not A236)  and  (not A235) );
 a81193a <=( (not A266)  and  (not A265) );
 a81194a <=( a81193a  and  a81190a );
 a81197a <=( (not A299)  and  A298 );
 a81200a <=( A301  and  A300 );
 a81201a <=( a81200a  and  a81197a );
 a81202a <=( a81201a  and  a81194a );
 a81205a <=( (not A167)  and  (not A169) );
 a81208a <=( A199  and  (not A166) );
 a81209a <=( a81208a  and  a81205a );
 a81212a <=( A201  and  (not A200) );
 a81215a <=( (not A233)  and  A202 );
 a81216a <=( a81215a  and  a81212a );
 a81217a <=( a81216a  and  a81209a );
 a81220a <=( (not A236)  and  (not A235) );
 a81223a <=( (not A266)  and  (not A265) );
 a81224a <=( a81223a  and  a81220a );
 a81227a <=( (not A299)  and  A298 );
 a81230a <=( A302  and  A300 );
 a81231a <=( a81230a  and  a81227a );
 a81232a <=( a81231a  and  a81224a );
 a81235a <=( (not A167)  and  (not A169) );
 a81238a <=( A199  and  (not A166) );
 a81239a <=( a81238a  and  a81235a );
 a81242a <=( A201  and  (not A200) );
 a81245a <=( (not A233)  and  A202 );
 a81246a <=( a81245a  and  a81242a );
 a81247a <=( a81246a  and  a81239a );
 a81250a <=( (not A266)  and  (not A234) );
 a81253a <=( (not A269)  and  (not A268) );
 a81254a <=( a81253a  and  a81250a );
 a81257a <=( (not A299)  and  A298 );
 a81260a <=( A301  and  A300 );
 a81261a <=( a81260a  and  a81257a );
 a81262a <=( a81261a  and  a81254a );
 a81265a <=( (not A167)  and  (not A169) );
 a81268a <=( A199  and  (not A166) );
 a81269a <=( a81268a  and  a81265a );
 a81272a <=( A201  and  (not A200) );
 a81275a <=( (not A233)  and  A202 );
 a81276a <=( a81275a  and  a81272a );
 a81277a <=( a81276a  and  a81269a );
 a81280a <=( (not A266)  and  (not A234) );
 a81283a <=( (not A269)  and  (not A268) );
 a81284a <=( a81283a  and  a81280a );
 a81287a <=( (not A299)  and  A298 );
 a81290a <=( A302  and  A300 );
 a81291a <=( a81290a  and  a81287a );
 a81292a <=( a81291a  and  a81284a );
 a81295a <=( (not A167)  and  (not A169) );
 a81298a <=( A199  and  (not A166) );
 a81299a <=( a81298a  and  a81295a );
 a81302a <=( A201  and  (not A200) );
 a81305a <=( (not A232)  and  A202 );
 a81306a <=( a81305a  and  a81302a );
 a81307a <=( a81306a  and  a81299a );
 a81310a <=( (not A266)  and  (not A233) );
 a81313a <=( (not A269)  and  (not A268) );
 a81314a <=( a81313a  and  a81310a );
 a81317a <=( (not A299)  and  A298 );
 a81320a <=( A301  and  A300 );
 a81321a <=( a81320a  and  a81317a );
 a81322a <=( a81321a  and  a81314a );
 a81325a <=( (not A167)  and  (not A169) );
 a81328a <=( A199  and  (not A166) );
 a81329a <=( a81328a  and  a81325a );
 a81332a <=( A201  and  (not A200) );
 a81335a <=( (not A232)  and  A202 );
 a81336a <=( a81335a  and  a81332a );
 a81337a <=( a81336a  and  a81329a );
 a81340a <=( (not A266)  and  (not A233) );
 a81343a <=( (not A269)  and  (not A268) );
 a81344a <=( a81343a  and  a81340a );
 a81347a <=( (not A299)  and  A298 );
 a81350a <=( A302  and  A300 );
 a81351a <=( a81350a  and  a81347a );
 a81352a <=( a81351a  and  a81344a );
 a81355a <=( (not A167)  and  (not A169) );
 a81358a <=( A199  and  (not A166) );
 a81359a <=( a81358a  and  a81355a );
 a81362a <=( A201  and  (not A200) );
 a81365a <=( A232  and  A203 );
 a81366a <=( a81365a  and  a81362a );
 a81367a <=( a81366a  and  a81359a );
 a81370a <=( A265  and  A233 );
 a81373a <=( (not A269)  and  (not A268) );
 a81374a <=( a81373a  and  a81370a );
 a81377a <=( (not A299)  and  A298 );
 a81380a <=( A301  and  A300 );
 a81381a <=( a81380a  and  a81377a );
 a81382a <=( a81381a  and  a81374a );
 a81385a <=( (not A167)  and  (not A169) );
 a81388a <=( A199  and  (not A166) );
 a81389a <=( a81388a  and  a81385a );
 a81392a <=( A201  and  (not A200) );
 a81395a <=( A232  and  A203 );
 a81396a <=( a81395a  and  a81392a );
 a81397a <=( a81396a  and  a81389a );
 a81400a <=( A265  and  A233 );
 a81403a <=( (not A269)  and  (not A268) );
 a81404a <=( a81403a  and  a81400a );
 a81407a <=( (not A299)  and  A298 );
 a81410a <=( A302  and  A300 );
 a81411a <=( a81410a  and  a81407a );
 a81412a <=( a81411a  and  a81404a );
 a81415a <=( (not A167)  and  (not A169) );
 a81418a <=( A199  and  (not A166) );
 a81419a <=( a81418a  and  a81415a );
 a81422a <=( A201  and  (not A200) );
 a81425a <=( (not A233)  and  A203 );
 a81426a <=( a81425a  and  a81422a );
 a81427a <=( a81426a  and  a81419a );
 a81430a <=( (not A236)  and  (not A235) );
 a81433a <=( A266  and  A265 );
 a81434a <=( a81433a  and  a81430a );
 a81437a <=( (not A299)  and  A298 );
 a81440a <=( A301  and  A300 );
 a81441a <=( a81440a  and  a81437a );
 a81442a <=( a81441a  and  a81434a );
 a81445a <=( (not A167)  and  (not A169) );
 a81448a <=( A199  and  (not A166) );
 a81449a <=( a81448a  and  a81445a );
 a81452a <=( A201  and  (not A200) );
 a81455a <=( (not A233)  and  A203 );
 a81456a <=( a81455a  and  a81452a );
 a81457a <=( a81456a  and  a81449a );
 a81460a <=( (not A236)  and  (not A235) );
 a81463a <=( A266  and  A265 );
 a81464a <=( a81463a  and  a81460a );
 a81467a <=( (not A299)  and  A298 );
 a81470a <=( A302  and  A300 );
 a81471a <=( a81470a  and  a81467a );
 a81472a <=( a81471a  and  a81464a );
 a81475a <=( (not A167)  and  (not A169) );
 a81478a <=( A199  and  (not A166) );
 a81479a <=( a81478a  and  a81475a );
 a81482a <=( A201  and  (not A200) );
 a81485a <=( (not A233)  and  A203 );
 a81486a <=( a81485a  and  a81482a );
 a81487a <=( a81486a  and  a81479a );
 a81490a <=( (not A236)  and  (not A235) );
 a81493a <=( (not A267)  and  (not A266) );
 a81494a <=( a81493a  and  a81490a );
 a81497a <=( (not A299)  and  A298 );
 a81500a <=( A301  and  A300 );
 a81501a <=( a81500a  and  a81497a );
 a81502a <=( a81501a  and  a81494a );
 a81505a <=( (not A167)  and  (not A169) );
 a81508a <=( A199  and  (not A166) );
 a81509a <=( a81508a  and  a81505a );
 a81512a <=( A201  and  (not A200) );
 a81515a <=( (not A233)  and  A203 );
 a81516a <=( a81515a  and  a81512a );
 a81517a <=( a81516a  and  a81509a );
 a81520a <=( (not A236)  and  (not A235) );
 a81523a <=( (not A267)  and  (not A266) );
 a81524a <=( a81523a  and  a81520a );
 a81527a <=( (not A299)  and  A298 );
 a81530a <=( A302  and  A300 );
 a81531a <=( a81530a  and  a81527a );
 a81532a <=( a81531a  and  a81524a );
 a81535a <=( (not A167)  and  (not A169) );
 a81538a <=( A199  and  (not A166) );
 a81539a <=( a81538a  and  a81535a );
 a81542a <=( A201  and  (not A200) );
 a81545a <=( (not A233)  and  A203 );
 a81546a <=( a81545a  and  a81542a );
 a81547a <=( a81546a  and  a81539a );
 a81550a <=( (not A236)  and  (not A235) );
 a81553a <=( (not A266)  and  (not A265) );
 a81554a <=( a81553a  and  a81550a );
 a81557a <=( (not A299)  and  A298 );
 a81560a <=( A301  and  A300 );
 a81561a <=( a81560a  and  a81557a );
 a81562a <=( a81561a  and  a81554a );
 a81565a <=( (not A167)  and  (not A169) );
 a81568a <=( A199  and  (not A166) );
 a81569a <=( a81568a  and  a81565a );
 a81572a <=( A201  and  (not A200) );
 a81575a <=( (not A233)  and  A203 );
 a81576a <=( a81575a  and  a81572a );
 a81577a <=( a81576a  and  a81569a );
 a81580a <=( (not A236)  and  (not A235) );
 a81583a <=( (not A266)  and  (not A265) );
 a81584a <=( a81583a  and  a81580a );
 a81587a <=( (not A299)  and  A298 );
 a81590a <=( A302  and  A300 );
 a81591a <=( a81590a  and  a81587a );
 a81592a <=( a81591a  and  a81584a );
 a81595a <=( (not A167)  and  (not A169) );
 a81598a <=( A199  and  (not A166) );
 a81599a <=( a81598a  and  a81595a );
 a81602a <=( A201  and  (not A200) );
 a81605a <=( (not A233)  and  A203 );
 a81606a <=( a81605a  and  a81602a );
 a81607a <=( a81606a  and  a81599a );
 a81610a <=( (not A266)  and  (not A234) );
 a81613a <=( (not A269)  and  (not A268) );
 a81614a <=( a81613a  and  a81610a );
 a81617a <=( (not A299)  and  A298 );
 a81620a <=( A301  and  A300 );
 a81621a <=( a81620a  and  a81617a );
 a81622a <=( a81621a  and  a81614a );
 a81625a <=( (not A167)  and  (not A169) );
 a81628a <=( A199  and  (not A166) );
 a81629a <=( a81628a  and  a81625a );
 a81632a <=( A201  and  (not A200) );
 a81635a <=( (not A233)  and  A203 );
 a81636a <=( a81635a  and  a81632a );
 a81637a <=( a81636a  and  a81629a );
 a81640a <=( (not A266)  and  (not A234) );
 a81643a <=( (not A269)  and  (not A268) );
 a81644a <=( a81643a  and  a81640a );
 a81647a <=( (not A299)  and  A298 );
 a81650a <=( A302  and  A300 );
 a81651a <=( a81650a  and  a81647a );
 a81652a <=( a81651a  and  a81644a );
 a81655a <=( (not A167)  and  (not A169) );
 a81658a <=( A199  and  (not A166) );
 a81659a <=( a81658a  and  a81655a );
 a81662a <=( A201  and  (not A200) );
 a81665a <=( (not A232)  and  A203 );
 a81666a <=( a81665a  and  a81662a );
 a81667a <=( a81666a  and  a81659a );
 a81670a <=( (not A266)  and  (not A233) );
 a81673a <=( (not A269)  and  (not A268) );
 a81674a <=( a81673a  and  a81670a );
 a81677a <=( (not A299)  and  A298 );
 a81680a <=( A301  and  A300 );
 a81681a <=( a81680a  and  a81677a );
 a81682a <=( a81681a  and  a81674a );
 a81685a <=( (not A167)  and  (not A169) );
 a81688a <=( A199  and  (not A166) );
 a81689a <=( a81688a  and  a81685a );
 a81692a <=( A201  and  (not A200) );
 a81695a <=( (not A232)  and  A203 );
 a81696a <=( a81695a  and  a81692a );
 a81697a <=( a81696a  and  a81689a );
 a81700a <=( (not A266)  and  (not A233) );
 a81703a <=( (not A269)  and  (not A268) );
 a81704a <=( a81703a  and  a81700a );
 a81707a <=( (not A299)  and  A298 );
 a81710a <=( A302  and  A300 );
 a81711a <=( a81710a  and  a81707a );
 a81712a <=( a81711a  and  a81704a );
 a81715a <=( (not A168)  and  (not A169) );
 a81718a <=( A166  and  A167 );
 a81719a <=( a81718a  and  a81715a );
 a81722a <=( A200  and  (not A199) );
 a81725a <=( (not A235)  and  (not A233) );
 a81726a <=( a81725a  and  a81722a );
 a81727a <=( a81726a  and  a81719a );
 a81730a <=( (not A266)  and  (not A236) );
 a81733a <=( (not A269)  and  (not A268) );
 a81734a <=( a81733a  and  a81730a );
 a81737a <=( (not A299)  and  A298 );
 a81740a <=( A301  and  A300 );
 a81741a <=( a81740a  and  a81737a );
 a81742a <=( a81741a  and  a81734a );
 a81745a <=( (not A168)  and  (not A169) );
 a81748a <=( A166  and  A167 );
 a81749a <=( a81748a  and  a81745a );
 a81752a <=( A200  and  (not A199) );
 a81755a <=( (not A235)  and  (not A233) );
 a81756a <=( a81755a  and  a81752a );
 a81757a <=( a81756a  and  a81749a );
 a81760a <=( (not A266)  and  (not A236) );
 a81763a <=( (not A269)  and  (not A268) );
 a81764a <=( a81763a  and  a81760a );
 a81767a <=( (not A299)  and  A298 );
 a81770a <=( A302  and  A300 );
 a81771a <=( a81770a  and  a81767a );
 a81772a <=( a81771a  and  a81764a );
 a81775a <=( (not A168)  and  (not A169) );
 a81778a <=( A166  and  A167 );
 a81779a <=( a81778a  and  a81775a );
 a81782a <=( (not A200)  and  A199 );
 a81785a <=( A202  and  A201 );
 a81786a <=( a81785a  and  a81782a );
 a81787a <=( a81786a  and  a81779a );
 a81790a <=( A233  and  A232 );
 a81793a <=( (not A267)  and  A265 );
 a81794a <=( a81793a  and  a81790a );
 a81797a <=( (not A299)  and  A298 );
 a81800a <=( A301  and  A300 );
 a81801a <=( a81800a  and  a81797a );
 a81802a <=( a81801a  and  a81794a );
 a81805a <=( (not A168)  and  (not A169) );
 a81808a <=( A166  and  A167 );
 a81809a <=( a81808a  and  a81805a );
 a81812a <=( (not A200)  and  A199 );
 a81815a <=( A202  and  A201 );
 a81816a <=( a81815a  and  a81812a );
 a81817a <=( a81816a  and  a81809a );
 a81820a <=( A233  and  A232 );
 a81823a <=( (not A267)  and  A265 );
 a81824a <=( a81823a  and  a81820a );
 a81827a <=( (not A299)  and  A298 );
 a81830a <=( A302  and  A300 );
 a81831a <=( a81830a  and  a81827a );
 a81832a <=( a81831a  and  a81824a );
 a81835a <=( (not A168)  and  (not A169) );
 a81838a <=( A166  and  A167 );
 a81839a <=( a81838a  and  a81835a );
 a81842a <=( (not A200)  and  A199 );
 a81845a <=( A202  and  A201 );
 a81846a <=( a81845a  and  a81842a );
 a81847a <=( a81846a  and  a81839a );
 a81850a <=( A233  and  A232 );
 a81853a <=( A266  and  A265 );
 a81854a <=( a81853a  and  a81850a );
 a81857a <=( (not A299)  and  A298 );
 a81860a <=( A301  and  A300 );
 a81861a <=( a81860a  and  a81857a );
 a81862a <=( a81861a  and  a81854a );
 a81865a <=( (not A168)  and  (not A169) );
 a81868a <=( A166  and  A167 );
 a81869a <=( a81868a  and  a81865a );
 a81872a <=( (not A200)  and  A199 );
 a81875a <=( A202  and  A201 );
 a81876a <=( a81875a  and  a81872a );
 a81877a <=( a81876a  and  a81869a );
 a81880a <=( A233  and  A232 );
 a81883a <=( A266  and  A265 );
 a81884a <=( a81883a  and  a81880a );
 a81887a <=( (not A299)  and  A298 );
 a81890a <=( A302  and  A300 );
 a81891a <=( a81890a  and  a81887a );
 a81892a <=( a81891a  and  a81884a );
 a81895a <=( (not A168)  and  (not A169) );
 a81898a <=( A166  and  A167 );
 a81899a <=( a81898a  and  a81895a );
 a81902a <=( (not A200)  and  A199 );
 a81905a <=( A202  and  A201 );
 a81906a <=( a81905a  and  a81902a );
 a81907a <=( a81906a  and  a81899a );
 a81910a <=( A233  and  A232 );
 a81913a <=( (not A266)  and  (not A265) );
 a81914a <=( a81913a  and  a81910a );
 a81917a <=( (not A299)  and  A298 );
 a81920a <=( A301  and  A300 );
 a81921a <=( a81920a  and  a81917a );
 a81922a <=( a81921a  and  a81914a );
 a81925a <=( (not A168)  and  (not A169) );
 a81928a <=( A166  and  A167 );
 a81929a <=( a81928a  and  a81925a );
 a81932a <=( (not A200)  and  A199 );
 a81935a <=( A202  and  A201 );
 a81936a <=( a81935a  and  a81932a );
 a81937a <=( a81936a  and  a81929a );
 a81940a <=( A233  and  A232 );
 a81943a <=( (not A266)  and  (not A265) );
 a81944a <=( a81943a  and  a81940a );
 a81947a <=( (not A299)  and  A298 );
 a81950a <=( A302  and  A300 );
 a81951a <=( a81950a  and  a81947a );
 a81952a <=( a81951a  and  a81944a );
 a81955a <=( (not A168)  and  (not A169) );
 a81958a <=( A166  and  A167 );
 a81959a <=( a81958a  and  a81955a );
 a81962a <=( (not A200)  and  A199 );
 a81965a <=( A202  and  A201 );
 a81966a <=( a81965a  and  a81962a );
 a81967a <=( a81966a  and  a81959a );
 a81970a <=( (not A235)  and  (not A233) );
 a81973a <=( (not A266)  and  (not A236) );
 a81974a <=( a81973a  and  a81970a );
 a81977a <=( (not A269)  and  (not A268) );
 a81980a <=( A299  and  (not A298) );
 a81981a <=( a81980a  and  a81977a );
 a81982a <=( a81981a  and  a81974a );
 a81985a <=( (not A168)  and  (not A169) );
 a81988a <=( A166  and  A167 );
 a81989a <=( a81988a  and  a81985a );
 a81992a <=( (not A200)  and  A199 );
 a81995a <=( A202  and  A201 );
 a81996a <=( a81995a  and  a81992a );
 a81997a <=( a81996a  and  a81989a );
 a82000a <=( (not A234)  and  (not A233) );
 a82003a <=( A266  and  A265 );
 a82004a <=( a82003a  and  a82000a );
 a82007a <=( (not A299)  and  A298 );
 a82010a <=( A301  and  A300 );
 a82011a <=( a82010a  and  a82007a );
 a82012a <=( a82011a  and  a82004a );
 a82015a <=( (not A168)  and  (not A169) );
 a82018a <=( A166  and  A167 );
 a82019a <=( a82018a  and  a82015a );
 a82022a <=( (not A200)  and  A199 );
 a82025a <=( A202  and  A201 );
 a82026a <=( a82025a  and  a82022a );
 a82027a <=( a82026a  and  a82019a );
 a82030a <=( (not A234)  and  (not A233) );
 a82033a <=( A266  and  A265 );
 a82034a <=( a82033a  and  a82030a );
 a82037a <=( (not A299)  and  A298 );
 a82040a <=( A302  and  A300 );
 a82041a <=( a82040a  and  a82037a );
 a82042a <=( a82041a  and  a82034a );
 a82045a <=( (not A168)  and  (not A169) );
 a82048a <=( A166  and  A167 );
 a82049a <=( a82048a  and  a82045a );
 a82052a <=( (not A200)  and  A199 );
 a82055a <=( A202  and  A201 );
 a82056a <=( a82055a  and  a82052a );
 a82057a <=( a82056a  and  a82049a );
 a82060a <=( (not A234)  and  (not A233) );
 a82063a <=( (not A267)  and  (not A266) );
 a82064a <=( a82063a  and  a82060a );
 a82067a <=( (not A299)  and  A298 );
 a82070a <=( A301  and  A300 );
 a82071a <=( a82070a  and  a82067a );
 a82072a <=( a82071a  and  a82064a );
 a82075a <=( (not A168)  and  (not A169) );
 a82078a <=( A166  and  A167 );
 a82079a <=( a82078a  and  a82075a );
 a82082a <=( (not A200)  and  A199 );
 a82085a <=( A202  and  A201 );
 a82086a <=( a82085a  and  a82082a );
 a82087a <=( a82086a  and  a82079a );
 a82090a <=( (not A234)  and  (not A233) );
 a82093a <=( (not A267)  and  (not A266) );
 a82094a <=( a82093a  and  a82090a );
 a82097a <=( (not A299)  and  A298 );
 a82100a <=( A302  and  A300 );
 a82101a <=( a82100a  and  a82097a );
 a82102a <=( a82101a  and  a82094a );
 a82105a <=( (not A168)  and  (not A169) );
 a82108a <=( A166  and  A167 );
 a82109a <=( a82108a  and  a82105a );
 a82112a <=( (not A200)  and  A199 );
 a82115a <=( A202  and  A201 );
 a82116a <=( a82115a  and  a82112a );
 a82117a <=( a82116a  and  a82109a );
 a82120a <=( (not A234)  and  (not A233) );
 a82123a <=( (not A266)  and  (not A265) );
 a82124a <=( a82123a  and  a82120a );
 a82127a <=( (not A299)  and  A298 );
 a82130a <=( A301  and  A300 );
 a82131a <=( a82130a  and  a82127a );
 a82132a <=( a82131a  and  a82124a );
 a82135a <=( (not A168)  and  (not A169) );
 a82138a <=( A166  and  A167 );
 a82139a <=( a82138a  and  a82135a );
 a82142a <=( (not A200)  and  A199 );
 a82145a <=( A202  and  A201 );
 a82146a <=( a82145a  and  a82142a );
 a82147a <=( a82146a  and  a82139a );
 a82150a <=( (not A234)  and  (not A233) );
 a82153a <=( (not A266)  and  (not A265) );
 a82154a <=( a82153a  and  a82150a );
 a82157a <=( (not A299)  and  A298 );
 a82160a <=( A302  and  A300 );
 a82161a <=( a82160a  and  a82157a );
 a82162a <=( a82161a  and  a82154a );
 a82165a <=( (not A168)  and  (not A169) );
 a82168a <=( A166  and  A167 );
 a82169a <=( a82168a  and  a82165a );
 a82172a <=( (not A200)  and  A199 );
 a82175a <=( A202  and  A201 );
 a82176a <=( a82175a  and  a82172a );
 a82177a <=( a82176a  and  a82169a );
 a82180a <=( (not A233)  and  A232 );
 a82183a <=( A235  and  A234 );
 a82184a <=( a82183a  and  a82180a );
 a82187a <=( (not A266)  and  A265 );
 a82190a <=( A268  and  A267 );
 a82191a <=( a82190a  and  a82187a );
 a82192a <=( a82191a  and  a82184a );
 a82195a <=( (not A168)  and  (not A169) );
 a82198a <=( A166  and  A167 );
 a82199a <=( a82198a  and  a82195a );
 a82202a <=( (not A200)  and  A199 );
 a82205a <=( A202  and  A201 );
 a82206a <=( a82205a  and  a82202a );
 a82207a <=( a82206a  and  a82199a );
 a82210a <=( (not A233)  and  A232 );
 a82213a <=( A235  and  A234 );
 a82214a <=( a82213a  and  a82210a );
 a82217a <=( (not A266)  and  A265 );
 a82220a <=( A269  and  A267 );
 a82221a <=( a82220a  and  a82217a );
 a82222a <=( a82221a  and  a82214a );
 a82225a <=( (not A168)  and  (not A169) );
 a82228a <=( A166  and  A167 );
 a82229a <=( a82228a  and  a82225a );
 a82232a <=( (not A200)  and  A199 );
 a82235a <=( A202  and  A201 );
 a82236a <=( a82235a  and  a82232a );
 a82237a <=( a82236a  and  a82229a );
 a82240a <=( (not A233)  and  A232 );
 a82243a <=( A236  and  A234 );
 a82244a <=( a82243a  and  a82240a );
 a82247a <=( (not A266)  and  A265 );
 a82250a <=( A268  and  A267 );
 a82251a <=( a82250a  and  a82247a );
 a82252a <=( a82251a  and  a82244a );
 a82255a <=( (not A168)  and  (not A169) );
 a82258a <=( A166  and  A167 );
 a82259a <=( a82258a  and  a82255a );
 a82262a <=( (not A200)  and  A199 );
 a82265a <=( A202  and  A201 );
 a82266a <=( a82265a  and  a82262a );
 a82267a <=( a82266a  and  a82259a );
 a82270a <=( (not A233)  and  A232 );
 a82273a <=( A236  and  A234 );
 a82274a <=( a82273a  and  a82270a );
 a82277a <=( (not A266)  and  A265 );
 a82280a <=( A269  and  A267 );
 a82281a <=( a82280a  and  a82277a );
 a82282a <=( a82281a  and  a82274a );
 a82285a <=( (not A168)  and  (not A169) );
 a82288a <=( A166  and  A167 );
 a82289a <=( a82288a  and  a82285a );
 a82292a <=( (not A200)  and  A199 );
 a82295a <=( A202  and  A201 );
 a82296a <=( a82295a  and  a82292a );
 a82297a <=( a82296a  and  a82289a );
 a82300a <=( (not A233)  and  (not A232) );
 a82303a <=( A266  and  A265 );
 a82304a <=( a82303a  and  a82300a );
 a82307a <=( (not A299)  and  A298 );
 a82310a <=( A301  and  A300 );
 a82311a <=( a82310a  and  a82307a );
 a82312a <=( a82311a  and  a82304a );
 a82315a <=( (not A168)  and  (not A169) );
 a82318a <=( A166  and  A167 );
 a82319a <=( a82318a  and  a82315a );
 a82322a <=( (not A200)  and  A199 );
 a82325a <=( A202  and  A201 );
 a82326a <=( a82325a  and  a82322a );
 a82327a <=( a82326a  and  a82319a );
 a82330a <=( (not A233)  and  (not A232) );
 a82333a <=( A266  and  A265 );
 a82334a <=( a82333a  and  a82330a );
 a82337a <=( (not A299)  and  A298 );
 a82340a <=( A302  and  A300 );
 a82341a <=( a82340a  and  a82337a );
 a82342a <=( a82341a  and  a82334a );
 a82345a <=( (not A168)  and  (not A169) );
 a82348a <=( A166  and  A167 );
 a82349a <=( a82348a  and  a82345a );
 a82352a <=( (not A200)  and  A199 );
 a82355a <=( A202  and  A201 );
 a82356a <=( a82355a  and  a82352a );
 a82357a <=( a82356a  and  a82349a );
 a82360a <=( (not A233)  and  (not A232) );
 a82363a <=( (not A267)  and  (not A266) );
 a82364a <=( a82363a  and  a82360a );
 a82367a <=( (not A299)  and  A298 );
 a82370a <=( A301  and  A300 );
 a82371a <=( a82370a  and  a82367a );
 a82372a <=( a82371a  and  a82364a );
 a82375a <=( (not A168)  and  (not A169) );
 a82378a <=( A166  and  A167 );
 a82379a <=( a82378a  and  a82375a );
 a82382a <=( (not A200)  and  A199 );
 a82385a <=( A202  and  A201 );
 a82386a <=( a82385a  and  a82382a );
 a82387a <=( a82386a  and  a82379a );
 a82390a <=( (not A233)  and  (not A232) );
 a82393a <=( (not A267)  and  (not A266) );
 a82394a <=( a82393a  and  a82390a );
 a82397a <=( (not A299)  and  A298 );
 a82400a <=( A302  and  A300 );
 a82401a <=( a82400a  and  a82397a );
 a82402a <=( a82401a  and  a82394a );
 a82405a <=( (not A168)  and  (not A169) );
 a82408a <=( A166  and  A167 );
 a82409a <=( a82408a  and  a82405a );
 a82412a <=( (not A200)  and  A199 );
 a82415a <=( A202  and  A201 );
 a82416a <=( a82415a  and  a82412a );
 a82417a <=( a82416a  and  a82409a );
 a82420a <=( (not A233)  and  (not A232) );
 a82423a <=( (not A266)  and  (not A265) );
 a82424a <=( a82423a  and  a82420a );
 a82427a <=( (not A299)  and  A298 );
 a82430a <=( A301  and  A300 );
 a82431a <=( a82430a  and  a82427a );
 a82432a <=( a82431a  and  a82424a );
 a82435a <=( (not A168)  and  (not A169) );
 a82438a <=( A166  and  A167 );
 a82439a <=( a82438a  and  a82435a );
 a82442a <=( (not A200)  and  A199 );
 a82445a <=( A202  and  A201 );
 a82446a <=( a82445a  and  a82442a );
 a82447a <=( a82446a  and  a82439a );
 a82450a <=( (not A233)  and  (not A232) );
 a82453a <=( (not A266)  and  (not A265) );
 a82454a <=( a82453a  and  a82450a );
 a82457a <=( (not A299)  and  A298 );
 a82460a <=( A302  and  A300 );
 a82461a <=( a82460a  and  a82457a );
 a82462a <=( a82461a  and  a82454a );
 a82465a <=( (not A168)  and  (not A169) );
 a82468a <=( A166  and  A167 );
 a82469a <=( a82468a  and  a82465a );
 a82472a <=( (not A200)  and  A199 );
 a82475a <=( A203  and  A201 );
 a82476a <=( a82475a  and  a82472a );
 a82477a <=( a82476a  and  a82469a );
 a82480a <=( A233  and  A232 );
 a82483a <=( (not A267)  and  A265 );
 a82484a <=( a82483a  and  a82480a );
 a82487a <=( (not A299)  and  A298 );
 a82490a <=( A301  and  A300 );
 a82491a <=( a82490a  and  a82487a );
 a82492a <=( a82491a  and  a82484a );
 a82495a <=( (not A168)  and  (not A169) );
 a82498a <=( A166  and  A167 );
 a82499a <=( a82498a  and  a82495a );
 a82502a <=( (not A200)  and  A199 );
 a82505a <=( A203  and  A201 );
 a82506a <=( a82505a  and  a82502a );
 a82507a <=( a82506a  and  a82499a );
 a82510a <=( A233  and  A232 );
 a82513a <=( (not A267)  and  A265 );
 a82514a <=( a82513a  and  a82510a );
 a82517a <=( (not A299)  and  A298 );
 a82520a <=( A302  and  A300 );
 a82521a <=( a82520a  and  a82517a );
 a82522a <=( a82521a  and  a82514a );
 a82525a <=( (not A168)  and  (not A169) );
 a82528a <=( A166  and  A167 );
 a82529a <=( a82528a  and  a82525a );
 a82532a <=( (not A200)  and  A199 );
 a82535a <=( A203  and  A201 );
 a82536a <=( a82535a  and  a82532a );
 a82537a <=( a82536a  and  a82529a );
 a82540a <=( A233  and  A232 );
 a82543a <=( A266  and  A265 );
 a82544a <=( a82543a  and  a82540a );
 a82547a <=( (not A299)  and  A298 );
 a82550a <=( A301  and  A300 );
 a82551a <=( a82550a  and  a82547a );
 a82552a <=( a82551a  and  a82544a );
 a82555a <=( (not A168)  and  (not A169) );
 a82558a <=( A166  and  A167 );
 a82559a <=( a82558a  and  a82555a );
 a82562a <=( (not A200)  and  A199 );
 a82565a <=( A203  and  A201 );
 a82566a <=( a82565a  and  a82562a );
 a82567a <=( a82566a  and  a82559a );
 a82570a <=( A233  and  A232 );
 a82573a <=( A266  and  A265 );
 a82574a <=( a82573a  and  a82570a );
 a82577a <=( (not A299)  and  A298 );
 a82580a <=( A302  and  A300 );
 a82581a <=( a82580a  and  a82577a );
 a82582a <=( a82581a  and  a82574a );
 a82585a <=( (not A168)  and  (not A169) );
 a82588a <=( A166  and  A167 );
 a82589a <=( a82588a  and  a82585a );
 a82592a <=( (not A200)  and  A199 );
 a82595a <=( A203  and  A201 );
 a82596a <=( a82595a  and  a82592a );
 a82597a <=( a82596a  and  a82589a );
 a82600a <=( A233  and  A232 );
 a82603a <=( (not A266)  and  (not A265) );
 a82604a <=( a82603a  and  a82600a );
 a82607a <=( (not A299)  and  A298 );
 a82610a <=( A301  and  A300 );
 a82611a <=( a82610a  and  a82607a );
 a82612a <=( a82611a  and  a82604a );
 a82615a <=( (not A168)  and  (not A169) );
 a82618a <=( A166  and  A167 );
 a82619a <=( a82618a  and  a82615a );
 a82622a <=( (not A200)  and  A199 );
 a82625a <=( A203  and  A201 );
 a82626a <=( a82625a  and  a82622a );
 a82627a <=( a82626a  and  a82619a );
 a82630a <=( A233  and  A232 );
 a82633a <=( (not A266)  and  (not A265) );
 a82634a <=( a82633a  and  a82630a );
 a82637a <=( (not A299)  and  A298 );
 a82640a <=( A302  and  A300 );
 a82641a <=( a82640a  and  a82637a );
 a82642a <=( a82641a  and  a82634a );
 a82645a <=( (not A168)  and  (not A169) );
 a82648a <=( A166  and  A167 );
 a82649a <=( a82648a  and  a82645a );
 a82652a <=( (not A200)  and  A199 );
 a82655a <=( A203  and  A201 );
 a82656a <=( a82655a  and  a82652a );
 a82657a <=( a82656a  and  a82649a );
 a82660a <=( (not A235)  and  (not A233) );
 a82663a <=( (not A266)  and  (not A236) );
 a82664a <=( a82663a  and  a82660a );
 a82667a <=( (not A269)  and  (not A268) );
 a82670a <=( A299  and  (not A298) );
 a82671a <=( a82670a  and  a82667a );
 a82672a <=( a82671a  and  a82664a );
 a82675a <=( (not A168)  and  (not A169) );
 a82678a <=( A166  and  A167 );
 a82679a <=( a82678a  and  a82675a );
 a82682a <=( (not A200)  and  A199 );
 a82685a <=( A203  and  A201 );
 a82686a <=( a82685a  and  a82682a );
 a82687a <=( a82686a  and  a82679a );
 a82690a <=( (not A234)  and  (not A233) );
 a82693a <=( A266  and  A265 );
 a82694a <=( a82693a  and  a82690a );
 a82697a <=( (not A299)  and  A298 );
 a82700a <=( A301  and  A300 );
 a82701a <=( a82700a  and  a82697a );
 a82702a <=( a82701a  and  a82694a );
 a82705a <=( (not A168)  and  (not A169) );
 a82708a <=( A166  and  A167 );
 a82709a <=( a82708a  and  a82705a );
 a82712a <=( (not A200)  and  A199 );
 a82715a <=( A203  and  A201 );
 a82716a <=( a82715a  and  a82712a );
 a82717a <=( a82716a  and  a82709a );
 a82720a <=( (not A234)  and  (not A233) );
 a82723a <=( A266  and  A265 );
 a82724a <=( a82723a  and  a82720a );
 a82727a <=( (not A299)  and  A298 );
 a82730a <=( A302  and  A300 );
 a82731a <=( a82730a  and  a82727a );
 a82732a <=( a82731a  and  a82724a );
 a82735a <=( (not A168)  and  (not A169) );
 a82738a <=( A166  and  A167 );
 a82739a <=( a82738a  and  a82735a );
 a82742a <=( (not A200)  and  A199 );
 a82745a <=( A203  and  A201 );
 a82746a <=( a82745a  and  a82742a );
 a82747a <=( a82746a  and  a82739a );
 a82750a <=( (not A234)  and  (not A233) );
 a82753a <=( (not A267)  and  (not A266) );
 a82754a <=( a82753a  and  a82750a );
 a82757a <=( (not A299)  and  A298 );
 a82760a <=( A301  and  A300 );
 a82761a <=( a82760a  and  a82757a );
 a82762a <=( a82761a  and  a82754a );
 a82765a <=( (not A168)  and  (not A169) );
 a82768a <=( A166  and  A167 );
 a82769a <=( a82768a  and  a82765a );
 a82772a <=( (not A200)  and  A199 );
 a82775a <=( A203  and  A201 );
 a82776a <=( a82775a  and  a82772a );
 a82777a <=( a82776a  and  a82769a );
 a82780a <=( (not A234)  and  (not A233) );
 a82783a <=( (not A267)  and  (not A266) );
 a82784a <=( a82783a  and  a82780a );
 a82787a <=( (not A299)  and  A298 );
 a82790a <=( A302  and  A300 );
 a82791a <=( a82790a  and  a82787a );
 a82792a <=( a82791a  and  a82784a );
 a82795a <=( (not A168)  and  (not A169) );
 a82798a <=( A166  and  A167 );
 a82799a <=( a82798a  and  a82795a );
 a82802a <=( (not A200)  and  A199 );
 a82805a <=( A203  and  A201 );
 a82806a <=( a82805a  and  a82802a );
 a82807a <=( a82806a  and  a82799a );
 a82810a <=( (not A234)  and  (not A233) );
 a82813a <=( (not A266)  and  (not A265) );
 a82814a <=( a82813a  and  a82810a );
 a82817a <=( (not A299)  and  A298 );
 a82820a <=( A301  and  A300 );
 a82821a <=( a82820a  and  a82817a );
 a82822a <=( a82821a  and  a82814a );
 a82825a <=( (not A168)  and  (not A169) );
 a82828a <=( A166  and  A167 );
 a82829a <=( a82828a  and  a82825a );
 a82832a <=( (not A200)  and  A199 );
 a82835a <=( A203  and  A201 );
 a82836a <=( a82835a  and  a82832a );
 a82837a <=( a82836a  and  a82829a );
 a82840a <=( (not A234)  and  (not A233) );
 a82843a <=( (not A266)  and  (not A265) );
 a82844a <=( a82843a  and  a82840a );
 a82847a <=( (not A299)  and  A298 );
 a82850a <=( A302  and  A300 );
 a82851a <=( a82850a  and  a82847a );
 a82852a <=( a82851a  and  a82844a );
 a82855a <=( (not A168)  and  (not A169) );
 a82858a <=( A166  and  A167 );
 a82859a <=( a82858a  and  a82855a );
 a82862a <=( (not A200)  and  A199 );
 a82865a <=( A203  and  A201 );
 a82866a <=( a82865a  and  a82862a );
 a82867a <=( a82866a  and  a82859a );
 a82870a <=( (not A233)  and  A232 );
 a82873a <=( A235  and  A234 );
 a82874a <=( a82873a  and  a82870a );
 a82877a <=( (not A266)  and  A265 );
 a82880a <=( A268  and  A267 );
 a82881a <=( a82880a  and  a82877a );
 a82882a <=( a82881a  and  a82874a );
 a82885a <=( (not A168)  and  (not A169) );
 a82888a <=( A166  and  A167 );
 a82889a <=( a82888a  and  a82885a );
 a82892a <=( (not A200)  and  A199 );
 a82895a <=( A203  and  A201 );
 a82896a <=( a82895a  and  a82892a );
 a82897a <=( a82896a  and  a82889a );
 a82900a <=( (not A233)  and  A232 );
 a82903a <=( A235  and  A234 );
 a82904a <=( a82903a  and  a82900a );
 a82907a <=( (not A266)  and  A265 );
 a82910a <=( A269  and  A267 );
 a82911a <=( a82910a  and  a82907a );
 a82912a <=( a82911a  and  a82904a );
 a82915a <=( (not A168)  and  (not A169) );
 a82918a <=( A166  and  A167 );
 a82919a <=( a82918a  and  a82915a );
 a82922a <=( (not A200)  and  A199 );
 a82925a <=( A203  and  A201 );
 a82926a <=( a82925a  and  a82922a );
 a82927a <=( a82926a  and  a82919a );
 a82930a <=( (not A233)  and  A232 );
 a82933a <=( A236  and  A234 );
 a82934a <=( a82933a  and  a82930a );
 a82937a <=( (not A266)  and  A265 );
 a82940a <=( A268  and  A267 );
 a82941a <=( a82940a  and  a82937a );
 a82942a <=( a82941a  and  a82934a );
 a82945a <=( (not A168)  and  (not A169) );
 a82948a <=( A166  and  A167 );
 a82949a <=( a82948a  and  a82945a );
 a82952a <=( (not A200)  and  A199 );
 a82955a <=( A203  and  A201 );
 a82956a <=( a82955a  and  a82952a );
 a82957a <=( a82956a  and  a82949a );
 a82960a <=( (not A233)  and  A232 );
 a82963a <=( A236  and  A234 );
 a82964a <=( a82963a  and  a82960a );
 a82967a <=( (not A266)  and  A265 );
 a82970a <=( A269  and  A267 );
 a82971a <=( a82970a  and  a82967a );
 a82972a <=( a82971a  and  a82964a );
 a82975a <=( (not A168)  and  (not A169) );
 a82978a <=( A166  and  A167 );
 a82979a <=( a82978a  and  a82975a );
 a82982a <=( (not A200)  and  A199 );
 a82985a <=( A203  and  A201 );
 a82986a <=( a82985a  and  a82982a );
 a82987a <=( a82986a  and  a82979a );
 a82990a <=( (not A233)  and  (not A232) );
 a82993a <=( A266  and  A265 );
 a82994a <=( a82993a  and  a82990a );
 a82997a <=( (not A299)  and  A298 );
 a83000a <=( A301  and  A300 );
 a83001a <=( a83000a  and  a82997a );
 a83002a <=( a83001a  and  a82994a );
 a83005a <=( (not A168)  and  (not A169) );
 a83008a <=( A166  and  A167 );
 a83009a <=( a83008a  and  a83005a );
 a83012a <=( (not A200)  and  A199 );
 a83015a <=( A203  and  A201 );
 a83016a <=( a83015a  and  a83012a );
 a83017a <=( a83016a  and  a83009a );
 a83020a <=( (not A233)  and  (not A232) );
 a83023a <=( A266  and  A265 );
 a83024a <=( a83023a  and  a83020a );
 a83027a <=( (not A299)  and  A298 );
 a83030a <=( A302  and  A300 );
 a83031a <=( a83030a  and  a83027a );
 a83032a <=( a83031a  and  a83024a );
 a83035a <=( (not A168)  and  (not A169) );
 a83038a <=( A166  and  A167 );
 a83039a <=( a83038a  and  a83035a );
 a83042a <=( (not A200)  and  A199 );
 a83045a <=( A203  and  A201 );
 a83046a <=( a83045a  and  a83042a );
 a83047a <=( a83046a  and  a83039a );
 a83050a <=( (not A233)  and  (not A232) );
 a83053a <=( (not A267)  and  (not A266) );
 a83054a <=( a83053a  and  a83050a );
 a83057a <=( (not A299)  and  A298 );
 a83060a <=( A301  and  A300 );
 a83061a <=( a83060a  and  a83057a );
 a83062a <=( a83061a  and  a83054a );
 a83065a <=( (not A168)  and  (not A169) );
 a83068a <=( A166  and  A167 );
 a83069a <=( a83068a  and  a83065a );
 a83072a <=( (not A200)  and  A199 );
 a83075a <=( A203  and  A201 );
 a83076a <=( a83075a  and  a83072a );
 a83077a <=( a83076a  and  a83069a );
 a83080a <=( (not A233)  and  (not A232) );
 a83083a <=( (not A267)  and  (not A266) );
 a83084a <=( a83083a  and  a83080a );
 a83087a <=( (not A299)  and  A298 );
 a83090a <=( A302  and  A300 );
 a83091a <=( a83090a  and  a83087a );
 a83092a <=( a83091a  and  a83084a );
 a83095a <=( (not A168)  and  (not A169) );
 a83098a <=( A166  and  A167 );
 a83099a <=( a83098a  and  a83095a );
 a83102a <=( (not A200)  and  A199 );
 a83105a <=( A203  and  A201 );
 a83106a <=( a83105a  and  a83102a );
 a83107a <=( a83106a  and  a83099a );
 a83110a <=( (not A233)  and  (not A232) );
 a83113a <=( (not A266)  and  (not A265) );
 a83114a <=( a83113a  and  a83110a );
 a83117a <=( (not A299)  and  A298 );
 a83120a <=( A301  and  A300 );
 a83121a <=( a83120a  and  a83117a );
 a83122a <=( a83121a  and  a83114a );
 a83125a <=( (not A168)  and  (not A169) );
 a83128a <=( A166  and  A167 );
 a83129a <=( a83128a  and  a83125a );
 a83132a <=( (not A200)  and  A199 );
 a83135a <=( A203  and  A201 );
 a83136a <=( a83135a  and  a83132a );
 a83137a <=( a83136a  and  a83129a );
 a83140a <=( (not A233)  and  (not A232) );
 a83143a <=( (not A266)  and  (not A265) );
 a83144a <=( a83143a  and  a83140a );
 a83147a <=( (not A299)  and  A298 );
 a83150a <=( A302  and  A300 );
 a83151a <=( a83150a  and  a83147a );
 a83152a <=( a83151a  and  a83144a );
 a83155a <=( (not A169)  and  A170 );
 a83158a <=( (not A166)  and  A167 );
 a83159a <=( a83158a  and  a83155a );
 a83162a <=( A200  and  A199 );
 a83165a <=( (not A235)  and  (not A233) );
 a83166a <=( a83165a  and  a83162a );
 a83167a <=( a83166a  and  a83159a );
 a83170a <=( (not A266)  and  (not A236) );
 a83173a <=( (not A269)  and  (not A268) );
 a83174a <=( a83173a  and  a83170a );
 a83177a <=( (not A299)  and  A298 );
 a83180a <=( A301  and  A300 );
 a83181a <=( a83180a  and  a83177a );
 a83182a <=( a83181a  and  a83174a );
 a83185a <=( (not A169)  and  A170 );
 a83188a <=( (not A166)  and  A167 );
 a83189a <=( a83188a  and  a83185a );
 a83192a <=( A200  and  A199 );
 a83195a <=( (not A235)  and  (not A233) );
 a83196a <=( a83195a  and  a83192a );
 a83197a <=( a83196a  and  a83189a );
 a83200a <=( (not A266)  and  (not A236) );
 a83203a <=( (not A269)  and  (not A268) );
 a83204a <=( a83203a  and  a83200a );
 a83207a <=( (not A299)  and  A298 );
 a83210a <=( A302  and  A300 );
 a83211a <=( a83210a  and  a83207a );
 a83212a <=( a83211a  and  a83204a );
 a83215a <=( (not A169)  and  A170 );
 a83218a <=( (not A166)  and  A167 );
 a83219a <=( a83218a  and  a83215a );
 a83222a <=( (not A202)  and  (not A200) );
 a83225a <=( A232  and  (not A203) );
 a83226a <=( a83225a  and  a83222a );
 a83227a <=( a83226a  and  a83219a );
 a83230a <=( A265  and  A233 );
 a83233a <=( (not A269)  and  (not A268) );
 a83234a <=( a83233a  and  a83230a );
 a83237a <=( (not A299)  and  A298 );
 a83240a <=( A301  and  A300 );
 a83241a <=( a83240a  and  a83237a );
 a83242a <=( a83241a  and  a83234a );
 a83245a <=( (not A169)  and  A170 );
 a83248a <=( (not A166)  and  A167 );
 a83249a <=( a83248a  and  a83245a );
 a83252a <=( (not A202)  and  (not A200) );
 a83255a <=( A232  and  (not A203) );
 a83256a <=( a83255a  and  a83252a );
 a83257a <=( a83256a  and  a83249a );
 a83260a <=( A265  and  A233 );
 a83263a <=( (not A269)  and  (not A268) );
 a83264a <=( a83263a  and  a83260a );
 a83267a <=( (not A299)  and  A298 );
 a83270a <=( A302  and  A300 );
 a83271a <=( a83270a  and  a83267a );
 a83272a <=( a83271a  and  a83264a );
 a83275a <=( (not A169)  and  A170 );
 a83278a <=( (not A166)  and  A167 );
 a83279a <=( a83278a  and  a83275a );
 a83282a <=( (not A202)  and  (not A200) );
 a83285a <=( (not A233)  and  (not A203) );
 a83286a <=( a83285a  and  a83282a );
 a83287a <=( a83286a  and  a83279a );
 a83290a <=( (not A236)  and  (not A235) );
 a83293a <=( A266  and  A265 );
 a83294a <=( a83293a  and  a83290a );
 a83297a <=( (not A299)  and  A298 );
 a83300a <=( A301  and  A300 );
 a83301a <=( a83300a  and  a83297a );
 a83302a <=( a83301a  and  a83294a );
 a83305a <=( (not A169)  and  A170 );
 a83308a <=( (not A166)  and  A167 );
 a83309a <=( a83308a  and  a83305a );
 a83312a <=( (not A202)  and  (not A200) );
 a83315a <=( (not A233)  and  (not A203) );
 a83316a <=( a83315a  and  a83312a );
 a83317a <=( a83316a  and  a83309a );
 a83320a <=( (not A236)  and  (not A235) );
 a83323a <=( A266  and  A265 );
 a83324a <=( a83323a  and  a83320a );
 a83327a <=( (not A299)  and  A298 );
 a83330a <=( A302  and  A300 );
 a83331a <=( a83330a  and  a83327a );
 a83332a <=( a83331a  and  a83324a );
 a83335a <=( (not A169)  and  A170 );
 a83338a <=( (not A166)  and  A167 );
 a83339a <=( a83338a  and  a83335a );
 a83342a <=( (not A202)  and  (not A200) );
 a83345a <=( (not A233)  and  (not A203) );
 a83346a <=( a83345a  and  a83342a );
 a83347a <=( a83346a  and  a83339a );
 a83350a <=( (not A236)  and  (not A235) );
 a83353a <=( (not A267)  and  (not A266) );
 a83354a <=( a83353a  and  a83350a );
 a83357a <=( (not A299)  and  A298 );
 a83360a <=( A301  and  A300 );
 a83361a <=( a83360a  and  a83357a );
 a83362a <=( a83361a  and  a83354a );
 a83365a <=( (not A169)  and  A170 );
 a83368a <=( (not A166)  and  A167 );
 a83369a <=( a83368a  and  a83365a );
 a83372a <=( (not A202)  and  (not A200) );
 a83375a <=( (not A233)  and  (not A203) );
 a83376a <=( a83375a  and  a83372a );
 a83377a <=( a83376a  and  a83369a );
 a83380a <=( (not A236)  and  (not A235) );
 a83383a <=( (not A267)  and  (not A266) );
 a83384a <=( a83383a  and  a83380a );
 a83387a <=( (not A299)  and  A298 );
 a83390a <=( A302  and  A300 );
 a83391a <=( a83390a  and  a83387a );
 a83392a <=( a83391a  and  a83384a );
 a83395a <=( (not A169)  and  A170 );
 a83398a <=( (not A166)  and  A167 );
 a83399a <=( a83398a  and  a83395a );
 a83402a <=( (not A202)  and  (not A200) );
 a83405a <=( (not A233)  and  (not A203) );
 a83406a <=( a83405a  and  a83402a );
 a83407a <=( a83406a  and  a83399a );
 a83410a <=( (not A236)  and  (not A235) );
 a83413a <=( (not A266)  and  (not A265) );
 a83414a <=( a83413a  and  a83410a );
 a83417a <=( (not A299)  and  A298 );
 a83420a <=( A301  and  A300 );
 a83421a <=( a83420a  and  a83417a );
 a83422a <=( a83421a  and  a83414a );
 a83425a <=( (not A169)  and  A170 );
 a83428a <=( (not A166)  and  A167 );
 a83429a <=( a83428a  and  a83425a );
 a83432a <=( (not A202)  and  (not A200) );
 a83435a <=( (not A233)  and  (not A203) );
 a83436a <=( a83435a  and  a83432a );
 a83437a <=( a83436a  and  a83429a );
 a83440a <=( (not A236)  and  (not A235) );
 a83443a <=( (not A266)  and  (not A265) );
 a83444a <=( a83443a  and  a83440a );
 a83447a <=( (not A299)  and  A298 );
 a83450a <=( A302  and  A300 );
 a83451a <=( a83450a  and  a83447a );
 a83452a <=( a83451a  and  a83444a );
 a83455a <=( (not A169)  and  A170 );
 a83458a <=( (not A166)  and  A167 );
 a83459a <=( a83458a  and  a83455a );
 a83462a <=( (not A202)  and  (not A200) );
 a83465a <=( (not A233)  and  (not A203) );
 a83466a <=( a83465a  and  a83462a );
 a83467a <=( a83466a  and  a83459a );
 a83470a <=( (not A266)  and  (not A234) );
 a83473a <=( (not A269)  and  (not A268) );
 a83474a <=( a83473a  and  a83470a );
 a83477a <=( (not A299)  and  A298 );
 a83480a <=( A301  and  A300 );
 a83481a <=( a83480a  and  a83477a );
 a83482a <=( a83481a  and  a83474a );
 a83485a <=( (not A169)  and  A170 );
 a83488a <=( (not A166)  and  A167 );
 a83489a <=( a83488a  and  a83485a );
 a83492a <=( (not A202)  and  (not A200) );
 a83495a <=( (not A233)  and  (not A203) );
 a83496a <=( a83495a  and  a83492a );
 a83497a <=( a83496a  and  a83489a );
 a83500a <=( (not A266)  and  (not A234) );
 a83503a <=( (not A269)  and  (not A268) );
 a83504a <=( a83503a  and  a83500a );
 a83507a <=( (not A299)  and  A298 );
 a83510a <=( A302  and  A300 );
 a83511a <=( a83510a  and  a83507a );
 a83512a <=( a83511a  and  a83504a );
 a83515a <=( (not A169)  and  A170 );
 a83518a <=( (not A166)  and  A167 );
 a83519a <=( a83518a  and  a83515a );
 a83522a <=( (not A202)  and  (not A200) );
 a83525a <=( (not A232)  and  (not A203) );
 a83526a <=( a83525a  and  a83522a );
 a83527a <=( a83526a  and  a83519a );
 a83530a <=( (not A266)  and  (not A233) );
 a83533a <=( (not A269)  and  (not A268) );
 a83534a <=( a83533a  and  a83530a );
 a83537a <=( (not A299)  and  A298 );
 a83540a <=( A301  and  A300 );
 a83541a <=( a83540a  and  a83537a );
 a83542a <=( a83541a  and  a83534a );
 a83545a <=( (not A169)  and  A170 );
 a83548a <=( (not A166)  and  A167 );
 a83549a <=( a83548a  and  a83545a );
 a83552a <=( (not A202)  and  (not A200) );
 a83555a <=( (not A232)  and  (not A203) );
 a83556a <=( a83555a  and  a83552a );
 a83557a <=( a83556a  and  a83549a );
 a83560a <=( (not A266)  and  (not A233) );
 a83563a <=( (not A269)  and  (not A268) );
 a83564a <=( a83563a  and  a83560a );
 a83567a <=( (not A299)  and  A298 );
 a83570a <=( A302  and  A300 );
 a83571a <=( a83570a  and  a83567a );
 a83572a <=( a83571a  and  a83564a );
 a83575a <=( (not A169)  and  A170 );
 a83578a <=( (not A166)  and  A167 );
 a83579a <=( a83578a  and  a83575a );
 a83582a <=( (not A201)  and  (not A200) );
 a83585a <=( (not A235)  and  (not A233) );
 a83586a <=( a83585a  and  a83582a );
 a83587a <=( a83586a  and  a83579a );
 a83590a <=( (not A266)  and  (not A236) );
 a83593a <=( (not A269)  and  (not A268) );
 a83594a <=( a83593a  and  a83590a );
 a83597a <=( (not A299)  and  A298 );
 a83600a <=( A301  and  A300 );
 a83601a <=( a83600a  and  a83597a );
 a83602a <=( a83601a  and  a83594a );
 a83605a <=( (not A169)  and  A170 );
 a83608a <=( (not A166)  and  A167 );
 a83609a <=( a83608a  and  a83605a );
 a83612a <=( (not A201)  and  (not A200) );
 a83615a <=( (not A235)  and  (not A233) );
 a83616a <=( a83615a  and  a83612a );
 a83617a <=( a83616a  and  a83609a );
 a83620a <=( (not A266)  and  (not A236) );
 a83623a <=( (not A269)  and  (not A268) );
 a83624a <=( a83623a  and  a83620a );
 a83627a <=( (not A299)  and  A298 );
 a83630a <=( A302  and  A300 );
 a83631a <=( a83630a  and  a83627a );
 a83632a <=( a83631a  and  a83624a );
 a83635a <=( (not A169)  and  A170 );
 a83638a <=( (not A166)  and  A167 );
 a83639a <=( a83638a  and  a83635a );
 a83642a <=( (not A200)  and  (not A199) );
 a83645a <=( (not A235)  and  (not A233) );
 a83646a <=( a83645a  and  a83642a );
 a83647a <=( a83646a  and  a83639a );
 a83650a <=( (not A266)  and  (not A236) );
 a83653a <=( (not A269)  and  (not A268) );
 a83654a <=( a83653a  and  a83650a );
 a83657a <=( (not A299)  and  A298 );
 a83660a <=( A301  and  A300 );
 a83661a <=( a83660a  and  a83657a );
 a83662a <=( a83661a  and  a83654a );
 a83665a <=( (not A169)  and  A170 );
 a83668a <=( (not A166)  and  A167 );
 a83669a <=( a83668a  and  a83665a );
 a83672a <=( (not A200)  and  (not A199) );
 a83675a <=( (not A235)  and  (not A233) );
 a83676a <=( a83675a  and  a83672a );
 a83677a <=( a83676a  and  a83669a );
 a83680a <=( (not A266)  and  (not A236) );
 a83683a <=( (not A269)  and  (not A268) );
 a83684a <=( a83683a  and  a83680a );
 a83687a <=( (not A299)  and  A298 );
 a83690a <=( A302  and  A300 );
 a83691a <=( a83690a  and  a83687a );
 a83692a <=( a83691a  and  a83684a );
 a83695a <=( (not A169)  and  A170 );
 a83698a <=( A166  and  (not A167) );
 a83699a <=( a83698a  and  a83695a );
 a83702a <=( A200  and  A199 );
 a83705a <=( (not A235)  and  (not A233) );
 a83706a <=( a83705a  and  a83702a );
 a83707a <=( a83706a  and  a83699a );
 a83710a <=( (not A266)  and  (not A236) );
 a83713a <=( (not A269)  and  (not A268) );
 a83714a <=( a83713a  and  a83710a );
 a83717a <=( (not A299)  and  A298 );
 a83720a <=( A301  and  A300 );
 a83721a <=( a83720a  and  a83717a );
 a83722a <=( a83721a  and  a83714a );
 a83725a <=( (not A169)  and  A170 );
 a83728a <=( A166  and  (not A167) );
 a83729a <=( a83728a  and  a83725a );
 a83732a <=( A200  and  A199 );
 a83735a <=( (not A235)  and  (not A233) );
 a83736a <=( a83735a  and  a83732a );
 a83737a <=( a83736a  and  a83729a );
 a83740a <=( (not A266)  and  (not A236) );
 a83743a <=( (not A269)  and  (not A268) );
 a83744a <=( a83743a  and  a83740a );
 a83747a <=( (not A299)  and  A298 );
 a83750a <=( A302  and  A300 );
 a83751a <=( a83750a  and  a83747a );
 a83752a <=( a83751a  and  a83744a );
 a83755a <=( (not A169)  and  A170 );
 a83758a <=( A166  and  (not A167) );
 a83759a <=( a83758a  and  a83755a );
 a83762a <=( (not A202)  and  (not A200) );
 a83765a <=( A232  and  (not A203) );
 a83766a <=( a83765a  and  a83762a );
 a83767a <=( a83766a  and  a83759a );
 a83770a <=( A265  and  A233 );
 a83773a <=( (not A269)  and  (not A268) );
 a83774a <=( a83773a  and  a83770a );
 a83777a <=( (not A299)  and  A298 );
 a83780a <=( A301  and  A300 );
 a83781a <=( a83780a  and  a83777a );
 a83782a <=( a83781a  and  a83774a );
 a83785a <=( (not A169)  and  A170 );
 a83788a <=( A166  and  (not A167) );
 a83789a <=( a83788a  and  a83785a );
 a83792a <=( (not A202)  and  (not A200) );
 a83795a <=( A232  and  (not A203) );
 a83796a <=( a83795a  and  a83792a );
 a83797a <=( a83796a  and  a83789a );
 a83800a <=( A265  and  A233 );
 a83803a <=( (not A269)  and  (not A268) );
 a83804a <=( a83803a  and  a83800a );
 a83807a <=( (not A299)  and  A298 );
 a83810a <=( A302  and  A300 );
 a83811a <=( a83810a  and  a83807a );
 a83812a <=( a83811a  and  a83804a );
 a83815a <=( (not A169)  and  A170 );
 a83818a <=( A166  and  (not A167) );
 a83819a <=( a83818a  and  a83815a );
 a83822a <=( (not A202)  and  (not A200) );
 a83825a <=( (not A233)  and  (not A203) );
 a83826a <=( a83825a  and  a83822a );
 a83827a <=( a83826a  and  a83819a );
 a83830a <=( (not A236)  and  (not A235) );
 a83833a <=( A266  and  A265 );
 a83834a <=( a83833a  and  a83830a );
 a83837a <=( (not A299)  and  A298 );
 a83840a <=( A301  and  A300 );
 a83841a <=( a83840a  and  a83837a );
 a83842a <=( a83841a  and  a83834a );
 a83845a <=( (not A169)  and  A170 );
 a83848a <=( A166  and  (not A167) );
 a83849a <=( a83848a  and  a83845a );
 a83852a <=( (not A202)  and  (not A200) );
 a83855a <=( (not A233)  and  (not A203) );
 a83856a <=( a83855a  and  a83852a );
 a83857a <=( a83856a  and  a83849a );
 a83860a <=( (not A236)  and  (not A235) );
 a83863a <=( A266  and  A265 );
 a83864a <=( a83863a  and  a83860a );
 a83867a <=( (not A299)  and  A298 );
 a83870a <=( A302  and  A300 );
 a83871a <=( a83870a  and  a83867a );
 a83872a <=( a83871a  and  a83864a );
 a83875a <=( (not A169)  and  A170 );
 a83878a <=( A166  and  (not A167) );
 a83879a <=( a83878a  and  a83875a );
 a83882a <=( (not A202)  and  (not A200) );
 a83885a <=( (not A233)  and  (not A203) );
 a83886a <=( a83885a  and  a83882a );
 a83887a <=( a83886a  and  a83879a );
 a83890a <=( (not A236)  and  (not A235) );
 a83893a <=( (not A267)  and  (not A266) );
 a83894a <=( a83893a  and  a83890a );
 a83897a <=( (not A299)  and  A298 );
 a83900a <=( A301  and  A300 );
 a83901a <=( a83900a  and  a83897a );
 a83902a <=( a83901a  and  a83894a );
 a83905a <=( (not A169)  and  A170 );
 a83908a <=( A166  and  (not A167) );
 a83909a <=( a83908a  and  a83905a );
 a83912a <=( (not A202)  and  (not A200) );
 a83915a <=( (not A233)  and  (not A203) );
 a83916a <=( a83915a  and  a83912a );
 a83917a <=( a83916a  and  a83909a );
 a83920a <=( (not A236)  and  (not A235) );
 a83923a <=( (not A267)  and  (not A266) );
 a83924a <=( a83923a  and  a83920a );
 a83927a <=( (not A299)  and  A298 );
 a83930a <=( A302  and  A300 );
 a83931a <=( a83930a  and  a83927a );
 a83932a <=( a83931a  and  a83924a );
 a83935a <=( (not A169)  and  A170 );
 a83938a <=( A166  and  (not A167) );
 a83939a <=( a83938a  and  a83935a );
 a83942a <=( (not A202)  and  (not A200) );
 a83945a <=( (not A233)  and  (not A203) );
 a83946a <=( a83945a  and  a83942a );
 a83947a <=( a83946a  and  a83939a );
 a83950a <=( (not A236)  and  (not A235) );
 a83953a <=( (not A266)  and  (not A265) );
 a83954a <=( a83953a  and  a83950a );
 a83957a <=( (not A299)  and  A298 );
 a83960a <=( A301  and  A300 );
 a83961a <=( a83960a  and  a83957a );
 a83962a <=( a83961a  and  a83954a );
 a83965a <=( (not A169)  and  A170 );
 a83968a <=( A166  and  (not A167) );
 a83969a <=( a83968a  and  a83965a );
 a83972a <=( (not A202)  and  (not A200) );
 a83975a <=( (not A233)  and  (not A203) );
 a83976a <=( a83975a  and  a83972a );
 a83977a <=( a83976a  and  a83969a );
 a83980a <=( (not A236)  and  (not A235) );
 a83983a <=( (not A266)  and  (not A265) );
 a83984a <=( a83983a  and  a83980a );
 a83987a <=( (not A299)  and  A298 );
 a83990a <=( A302  and  A300 );
 a83991a <=( a83990a  and  a83987a );
 a83992a <=( a83991a  and  a83984a );
 a83995a <=( (not A169)  and  A170 );
 a83998a <=( A166  and  (not A167) );
 a83999a <=( a83998a  and  a83995a );
 a84002a <=( (not A202)  and  (not A200) );
 a84005a <=( (not A233)  and  (not A203) );
 a84006a <=( a84005a  and  a84002a );
 a84007a <=( a84006a  and  a83999a );
 a84010a <=( (not A266)  and  (not A234) );
 a84013a <=( (not A269)  and  (not A268) );
 a84014a <=( a84013a  and  a84010a );
 a84017a <=( (not A299)  and  A298 );
 a84020a <=( A301  and  A300 );
 a84021a <=( a84020a  and  a84017a );
 a84022a <=( a84021a  and  a84014a );
 a84025a <=( (not A169)  and  A170 );
 a84028a <=( A166  and  (not A167) );
 a84029a <=( a84028a  and  a84025a );
 a84032a <=( (not A202)  and  (not A200) );
 a84035a <=( (not A233)  and  (not A203) );
 a84036a <=( a84035a  and  a84032a );
 a84037a <=( a84036a  and  a84029a );
 a84040a <=( (not A266)  and  (not A234) );
 a84043a <=( (not A269)  and  (not A268) );
 a84044a <=( a84043a  and  a84040a );
 a84047a <=( (not A299)  and  A298 );
 a84050a <=( A302  and  A300 );
 a84051a <=( a84050a  and  a84047a );
 a84052a <=( a84051a  and  a84044a );
 a84055a <=( (not A169)  and  A170 );
 a84058a <=( A166  and  (not A167) );
 a84059a <=( a84058a  and  a84055a );
 a84062a <=( (not A202)  and  (not A200) );
 a84065a <=( (not A232)  and  (not A203) );
 a84066a <=( a84065a  and  a84062a );
 a84067a <=( a84066a  and  a84059a );
 a84070a <=( (not A266)  and  (not A233) );
 a84073a <=( (not A269)  and  (not A268) );
 a84074a <=( a84073a  and  a84070a );
 a84077a <=( (not A299)  and  A298 );
 a84080a <=( A301  and  A300 );
 a84081a <=( a84080a  and  a84077a );
 a84082a <=( a84081a  and  a84074a );
 a84085a <=( (not A169)  and  A170 );
 a84088a <=( A166  and  (not A167) );
 a84089a <=( a84088a  and  a84085a );
 a84092a <=( (not A202)  and  (not A200) );
 a84095a <=( (not A232)  and  (not A203) );
 a84096a <=( a84095a  and  a84092a );
 a84097a <=( a84096a  and  a84089a );
 a84100a <=( (not A266)  and  (not A233) );
 a84103a <=( (not A269)  and  (not A268) );
 a84104a <=( a84103a  and  a84100a );
 a84107a <=( (not A299)  and  A298 );
 a84110a <=( A302  and  A300 );
 a84111a <=( a84110a  and  a84107a );
 a84112a <=( a84111a  and  a84104a );
 a84115a <=( (not A169)  and  A170 );
 a84118a <=( A166  and  (not A167) );
 a84119a <=( a84118a  and  a84115a );
 a84122a <=( (not A201)  and  (not A200) );
 a84125a <=( (not A235)  and  (not A233) );
 a84126a <=( a84125a  and  a84122a );
 a84127a <=( a84126a  and  a84119a );
 a84130a <=( (not A266)  and  (not A236) );
 a84133a <=( (not A269)  and  (not A268) );
 a84134a <=( a84133a  and  a84130a );
 a84137a <=( (not A299)  and  A298 );
 a84140a <=( A301  and  A300 );
 a84141a <=( a84140a  and  a84137a );
 a84142a <=( a84141a  and  a84134a );
 a84145a <=( (not A169)  and  A170 );
 a84148a <=( A166  and  (not A167) );
 a84149a <=( a84148a  and  a84145a );
 a84152a <=( (not A201)  and  (not A200) );
 a84155a <=( (not A235)  and  (not A233) );
 a84156a <=( a84155a  and  a84152a );
 a84157a <=( a84156a  and  a84149a );
 a84160a <=( (not A266)  and  (not A236) );
 a84163a <=( (not A269)  and  (not A268) );
 a84164a <=( a84163a  and  a84160a );
 a84167a <=( (not A299)  and  A298 );
 a84170a <=( A302  and  A300 );
 a84171a <=( a84170a  and  a84167a );
 a84172a <=( a84171a  and  a84164a );
 a84175a <=( (not A169)  and  A170 );
 a84178a <=( A166  and  (not A167) );
 a84179a <=( a84178a  and  a84175a );
 a84182a <=( (not A200)  and  (not A199) );
 a84185a <=( (not A235)  and  (not A233) );
 a84186a <=( a84185a  and  a84182a );
 a84187a <=( a84186a  and  a84179a );
 a84190a <=( (not A266)  and  (not A236) );
 a84193a <=( (not A269)  and  (not A268) );
 a84194a <=( a84193a  and  a84190a );
 a84197a <=( (not A299)  and  A298 );
 a84200a <=( A301  and  A300 );
 a84201a <=( a84200a  and  a84197a );
 a84202a <=( a84201a  and  a84194a );
 a84205a <=( (not A169)  and  A170 );
 a84208a <=( A166  and  (not A167) );
 a84209a <=( a84208a  and  a84205a );
 a84212a <=( (not A200)  and  (not A199) );
 a84215a <=( (not A235)  and  (not A233) );
 a84216a <=( a84215a  and  a84212a );
 a84217a <=( a84216a  and  a84209a );
 a84220a <=( (not A266)  and  (not A236) );
 a84223a <=( (not A269)  and  (not A268) );
 a84224a <=( a84223a  and  a84220a );
 a84227a <=( (not A299)  and  A298 );
 a84230a <=( A302  and  A300 );
 a84231a <=( a84230a  and  a84227a );
 a84232a <=( a84231a  and  a84224a );
 a84235a <=( (not A169)  and  (not A170) );
 a84238a <=( A199  and  (not A168) );
 a84239a <=( a84238a  and  a84235a );
 a84242a <=( A201  and  (not A200) );
 a84245a <=( A232  and  A202 );
 a84246a <=( a84245a  and  a84242a );
 a84247a <=( a84246a  and  a84239a );
 a84250a <=( A265  and  A233 );
 a84253a <=( (not A269)  and  (not A268) );
 a84254a <=( a84253a  and  a84250a );
 a84257a <=( (not A299)  and  A298 );
 a84260a <=( A301  and  A300 );
 a84261a <=( a84260a  and  a84257a );
 a84262a <=( a84261a  and  a84254a );
 a84265a <=( (not A169)  and  (not A170) );
 a84268a <=( A199  and  (not A168) );
 a84269a <=( a84268a  and  a84265a );
 a84272a <=( A201  and  (not A200) );
 a84275a <=( A232  and  A202 );
 a84276a <=( a84275a  and  a84272a );
 a84277a <=( a84276a  and  a84269a );
 a84280a <=( A265  and  A233 );
 a84283a <=( (not A269)  and  (not A268) );
 a84284a <=( a84283a  and  a84280a );
 a84287a <=( (not A299)  and  A298 );
 a84290a <=( A302  and  A300 );
 a84291a <=( a84290a  and  a84287a );
 a84292a <=( a84291a  and  a84284a );
 a84295a <=( (not A169)  and  (not A170) );
 a84298a <=( A199  and  (not A168) );
 a84299a <=( a84298a  and  a84295a );
 a84302a <=( A201  and  (not A200) );
 a84305a <=( (not A233)  and  A202 );
 a84306a <=( a84305a  and  a84302a );
 a84307a <=( a84306a  and  a84299a );
 a84310a <=( (not A236)  and  (not A235) );
 a84313a <=( A266  and  A265 );
 a84314a <=( a84313a  and  a84310a );
 a84317a <=( (not A299)  and  A298 );
 a84320a <=( A301  and  A300 );
 a84321a <=( a84320a  and  a84317a );
 a84322a <=( a84321a  and  a84314a );
 a84325a <=( (not A169)  and  (not A170) );
 a84328a <=( A199  and  (not A168) );
 a84329a <=( a84328a  and  a84325a );
 a84332a <=( A201  and  (not A200) );
 a84335a <=( (not A233)  and  A202 );
 a84336a <=( a84335a  and  a84332a );
 a84337a <=( a84336a  and  a84329a );
 a84340a <=( (not A236)  and  (not A235) );
 a84343a <=( A266  and  A265 );
 a84344a <=( a84343a  and  a84340a );
 a84347a <=( (not A299)  and  A298 );
 a84350a <=( A302  and  A300 );
 a84351a <=( a84350a  and  a84347a );
 a84352a <=( a84351a  and  a84344a );
 a84355a <=( (not A169)  and  (not A170) );
 a84358a <=( A199  and  (not A168) );
 a84359a <=( a84358a  and  a84355a );
 a84362a <=( A201  and  (not A200) );
 a84365a <=( (not A233)  and  A202 );
 a84366a <=( a84365a  and  a84362a );
 a84367a <=( a84366a  and  a84359a );
 a84370a <=( (not A236)  and  (not A235) );
 a84373a <=( (not A267)  and  (not A266) );
 a84374a <=( a84373a  and  a84370a );
 a84377a <=( (not A299)  and  A298 );
 a84380a <=( A301  and  A300 );
 a84381a <=( a84380a  and  a84377a );
 a84382a <=( a84381a  and  a84374a );
 a84385a <=( (not A169)  and  (not A170) );
 a84388a <=( A199  and  (not A168) );
 a84389a <=( a84388a  and  a84385a );
 a84392a <=( A201  and  (not A200) );
 a84395a <=( (not A233)  and  A202 );
 a84396a <=( a84395a  and  a84392a );
 a84397a <=( a84396a  and  a84389a );
 a84400a <=( (not A236)  and  (not A235) );
 a84403a <=( (not A267)  and  (not A266) );
 a84404a <=( a84403a  and  a84400a );
 a84407a <=( (not A299)  and  A298 );
 a84410a <=( A302  and  A300 );
 a84411a <=( a84410a  and  a84407a );
 a84412a <=( a84411a  and  a84404a );
 a84415a <=( (not A169)  and  (not A170) );
 a84418a <=( A199  and  (not A168) );
 a84419a <=( a84418a  and  a84415a );
 a84422a <=( A201  and  (not A200) );
 a84425a <=( (not A233)  and  A202 );
 a84426a <=( a84425a  and  a84422a );
 a84427a <=( a84426a  and  a84419a );
 a84430a <=( (not A236)  and  (not A235) );
 a84433a <=( (not A266)  and  (not A265) );
 a84434a <=( a84433a  and  a84430a );
 a84437a <=( (not A299)  and  A298 );
 a84440a <=( A301  and  A300 );
 a84441a <=( a84440a  and  a84437a );
 a84442a <=( a84441a  and  a84434a );
 a84445a <=( (not A169)  and  (not A170) );
 a84448a <=( A199  and  (not A168) );
 a84449a <=( a84448a  and  a84445a );
 a84452a <=( A201  and  (not A200) );
 a84455a <=( (not A233)  and  A202 );
 a84456a <=( a84455a  and  a84452a );
 a84457a <=( a84456a  and  a84449a );
 a84460a <=( (not A236)  and  (not A235) );
 a84463a <=( (not A266)  and  (not A265) );
 a84464a <=( a84463a  and  a84460a );
 a84467a <=( (not A299)  and  A298 );
 a84470a <=( A302  and  A300 );
 a84471a <=( a84470a  and  a84467a );
 a84472a <=( a84471a  and  a84464a );
 a84475a <=( (not A169)  and  (not A170) );
 a84478a <=( A199  and  (not A168) );
 a84479a <=( a84478a  and  a84475a );
 a84482a <=( A201  and  (not A200) );
 a84485a <=( (not A233)  and  A202 );
 a84486a <=( a84485a  and  a84482a );
 a84487a <=( a84486a  and  a84479a );
 a84490a <=( (not A266)  and  (not A234) );
 a84493a <=( (not A269)  and  (not A268) );
 a84494a <=( a84493a  and  a84490a );
 a84497a <=( (not A299)  and  A298 );
 a84500a <=( A301  and  A300 );
 a84501a <=( a84500a  and  a84497a );
 a84502a <=( a84501a  and  a84494a );
 a84505a <=( (not A169)  and  (not A170) );
 a84508a <=( A199  and  (not A168) );
 a84509a <=( a84508a  and  a84505a );
 a84512a <=( A201  and  (not A200) );
 a84515a <=( (not A233)  and  A202 );
 a84516a <=( a84515a  and  a84512a );
 a84517a <=( a84516a  and  a84509a );
 a84520a <=( (not A266)  and  (not A234) );
 a84523a <=( (not A269)  and  (not A268) );
 a84524a <=( a84523a  and  a84520a );
 a84527a <=( (not A299)  and  A298 );
 a84530a <=( A302  and  A300 );
 a84531a <=( a84530a  and  a84527a );
 a84532a <=( a84531a  and  a84524a );
 a84535a <=( (not A169)  and  (not A170) );
 a84538a <=( A199  and  (not A168) );
 a84539a <=( a84538a  and  a84535a );
 a84542a <=( A201  and  (not A200) );
 a84545a <=( (not A232)  and  A202 );
 a84546a <=( a84545a  and  a84542a );
 a84547a <=( a84546a  and  a84539a );
 a84550a <=( (not A266)  and  (not A233) );
 a84553a <=( (not A269)  and  (not A268) );
 a84554a <=( a84553a  and  a84550a );
 a84557a <=( (not A299)  and  A298 );
 a84560a <=( A301  and  A300 );
 a84561a <=( a84560a  and  a84557a );
 a84562a <=( a84561a  and  a84554a );
 a84565a <=( (not A169)  and  (not A170) );
 a84568a <=( A199  and  (not A168) );
 a84569a <=( a84568a  and  a84565a );
 a84572a <=( A201  and  (not A200) );
 a84575a <=( (not A232)  and  A202 );
 a84576a <=( a84575a  and  a84572a );
 a84577a <=( a84576a  and  a84569a );
 a84580a <=( (not A266)  and  (not A233) );
 a84583a <=( (not A269)  and  (not A268) );
 a84584a <=( a84583a  and  a84580a );
 a84587a <=( (not A299)  and  A298 );
 a84590a <=( A302  and  A300 );
 a84591a <=( a84590a  and  a84587a );
 a84592a <=( a84591a  and  a84584a );
 a84595a <=( (not A169)  and  (not A170) );
 a84598a <=( A199  and  (not A168) );
 a84599a <=( a84598a  and  a84595a );
 a84602a <=( A201  and  (not A200) );
 a84605a <=( A232  and  A203 );
 a84606a <=( a84605a  and  a84602a );
 a84607a <=( a84606a  and  a84599a );
 a84610a <=( A265  and  A233 );
 a84613a <=( (not A269)  and  (not A268) );
 a84614a <=( a84613a  and  a84610a );
 a84617a <=( (not A299)  and  A298 );
 a84620a <=( A301  and  A300 );
 a84621a <=( a84620a  and  a84617a );
 a84622a <=( a84621a  and  a84614a );
 a84625a <=( (not A169)  and  (not A170) );
 a84628a <=( A199  and  (not A168) );
 a84629a <=( a84628a  and  a84625a );
 a84632a <=( A201  and  (not A200) );
 a84635a <=( A232  and  A203 );
 a84636a <=( a84635a  and  a84632a );
 a84637a <=( a84636a  and  a84629a );
 a84640a <=( A265  and  A233 );
 a84643a <=( (not A269)  and  (not A268) );
 a84644a <=( a84643a  and  a84640a );
 a84647a <=( (not A299)  and  A298 );
 a84650a <=( A302  and  A300 );
 a84651a <=( a84650a  and  a84647a );
 a84652a <=( a84651a  and  a84644a );
 a84655a <=( (not A169)  and  (not A170) );
 a84658a <=( A199  and  (not A168) );
 a84659a <=( a84658a  and  a84655a );
 a84662a <=( A201  and  (not A200) );
 a84665a <=( (not A233)  and  A203 );
 a84666a <=( a84665a  and  a84662a );
 a84667a <=( a84666a  and  a84659a );
 a84670a <=( (not A236)  and  (not A235) );
 a84673a <=( A266  and  A265 );
 a84674a <=( a84673a  and  a84670a );
 a84677a <=( (not A299)  and  A298 );
 a84680a <=( A301  and  A300 );
 a84681a <=( a84680a  and  a84677a );
 a84682a <=( a84681a  and  a84674a );
 a84685a <=( (not A169)  and  (not A170) );
 a84688a <=( A199  and  (not A168) );
 a84689a <=( a84688a  and  a84685a );
 a84692a <=( A201  and  (not A200) );
 a84695a <=( (not A233)  and  A203 );
 a84696a <=( a84695a  and  a84692a );
 a84697a <=( a84696a  and  a84689a );
 a84700a <=( (not A236)  and  (not A235) );
 a84703a <=( A266  and  A265 );
 a84704a <=( a84703a  and  a84700a );
 a84707a <=( (not A299)  and  A298 );
 a84710a <=( A302  and  A300 );
 a84711a <=( a84710a  and  a84707a );
 a84712a <=( a84711a  and  a84704a );
 a84715a <=( (not A169)  and  (not A170) );
 a84718a <=( A199  and  (not A168) );
 a84719a <=( a84718a  and  a84715a );
 a84722a <=( A201  and  (not A200) );
 a84725a <=( (not A233)  and  A203 );
 a84726a <=( a84725a  and  a84722a );
 a84727a <=( a84726a  and  a84719a );
 a84730a <=( (not A236)  and  (not A235) );
 a84733a <=( (not A267)  and  (not A266) );
 a84734a <=( a84733a  and  a84730a );
 a84737a <=( (not A299)  and  A298 );
 a84740a <=( A301  and  A300 );
 a84741a <=( a84740a  and  a84737a );
 a84742a <=( a84741a  and  a84734a );
 a84745a <=( (not A169)  and  (not A170) );
 a84748a <=( A199  and  (not A168) );
 a84749a <=( a84748a  and  a84745a );
 a84752a <=( A201  and  (not A200) );
 a84755a <=( (not A233)  and  A203 );
 a84756a <=( a84755a  and  a84752a );
 a84757a <=( a84756a  and  a84749a );
 a84760a <=( (not A236)  and  (not A235) );
 a84763a <=( (not A267)  and  (not A266) );
 a84764a <=( a84763a  and  a84760a );
 a84767a <=( (not A299)  and  A298 );
 a84770a <=( A302  and  A300 );
 a84771a <=( a84770a  and  a84767a );
 a84772a <=( a84771a  and  a84764a );
 a84775a <=( (not A169)  and  (not A170) );
 a84778a <=( A199  and  (not A168) );
 a84779a <=( a84778a  and  a84775a );
 a84782a <=( A201  and  (not A200) );
 a84785a <=( (not A233)  and  A203 );
 a84786a <=( a84785a  and  a84782a );
 a84787a <=( a84786a  and  a84779a );
 a84790a <=( (not A236)  and  (not A235) );
 a84793a <=( (not A266)  and  (not A265) );
 a84794a <=( a84793a  and  a84790a );
 a84797a <=( (not A299)  and  A298 );
 a84800a <=( A301  and  A300 );
 a84801a <=( a84800a  and  a84797a );
 a84802a <=( a84801a  and  a84794a );
 a84805a <=( (not A169)  and  (not A170) );
 a84808a <=( A199  and  (not A168) );
 a84809a <=( a84808a  and  a84805a );
 a84812a <=( A201  and  (not A200) );
 a84815a <=( (not A233)  and  A203 );
 a84816a <=( a84815a  and  a84812a );
 a84817a <=( a84816a  and  a84809a );
 a84820a <=( (not A236)  and  (not A235) );
 a84823a <=( (not A266)  and  (not A265) );
 a84824a <=( a84823a  and  a84820a );
 a84827a <=( (not A299)  and  A298 );
 a84830a <=( A302  and  A300 );
 a84831a <=( a84830a  and  a84827a );
 a84832a <=( a84831a  and  a84824a );
 a84835a <=( (not A169)  and  (not A170) );
 a84838a <=( A199  and  (not A168) );
 a84839a <=( a84838a  and  a84835a );
 a84842a <=( A201  and  (not A200) );
 a84845a <=( (not A233)  and  A203 );
 a84846a <=( a84845a  and  a84842a );
 a84847a <=( a84846a  and  a84839a );
 a84850a <=( (not A266)  and  (not A234) );
 a84853a <=( (not A269)  and  (not A268) );
 a84854a <=( a84853a  and  a84850a );
 a84857a <=( (not A299)  and  A298 );
 a84860a <=( A301  and  A300 );
 a84861a <=( a84860a  and  a84857a );
 a84862a <=( a84861a  and  a84854a );
 a84865a <=( (not A169)  and  (not A170) );
 a84868a <=( A199  and  (not A168) );
 a84869a <=( a84868a  and  a84865a );
 a84872a <=( A201  and  (not A200) );
 a84875a <=( (not A233)  and  A203 );
 a84876a <=( a84875a  and  a84872a );
 a84877a <=( a84876a  and  a84869a );
 a84880a <=( (not A266)  and  (not A234) );
 a84883a <=( (not A269)  and  (not A268) );
 a84884a <=( a84883a  and  a84880a );
 a84887a <=( (not A299)  and  A298 );
 a84890a <=( A302  and  A300 );
 a84891a <=( a84890a  and  a84887a );
 a84892a <=( a84891a  and  a84884a );
 a84895a <=( (not A169)  and  (not A170) );
 a84898a <=( A199  and  (not A168) );
 a84899a <=( a84898a  and  a84895a );
 a84902a <=( A201  and  (not A200) );
 a84905a <=( (not A232)  and  A203 );
 a84906a <=( a84905a  and  a84902a );
 a84907a <=( a84906a  and  a84899a );
 a84910a <=( (not A266)  and  (not A233) );
 a84913a <=( (not A269)  and  (not A268) );
 a84914a <=( a84913a  and  a84910a );
 a84917a <=( (not A299)  and  A298 );
 a84920a <=( A301  and  A300 );
 a84921a <=( a84920a  and  a84917a );
 a84922a <=( a84921a  and  a84914a );
 a84925a <=( (not A169)  and  (not A170) );
 a84928a <=( A199  and  (not A168) );
 a84929a <=( a84928a  and  a84925a );
 a84932a <=( A201  and  (not A200) );
 a84935a <=( (not A232)  and  A203 );
 a84936a <=( a84935a  and  a84932a );
 a84937a <=( a84936a  and  a84929a );
 a84940a <=( (not A266)  and  (not A233) );
 a84943a <=( (not A269)  and  (not A268) );
 a84944a <=( a84943a  and  a84940a );
 a84947a <=( (not A299)  and  A298 );
 a84950a <=( A302  and  A300 );
 a84951a <=( a84950a  and  a84947a );
 a84952a <=( a84951a  and  a84944a );
 a84955a <=( (not A167)  and  A170 );
 a84958a <=( A199  and  (not A166) );
 a84959a <=( a84958a  and  a84955a );
 a84962a <=( A201  and  (not A200) );
 a84965a <=( (not A233)  and  A202 );
 a84966a <=( a84965a  and  a84962a );
 a84967a <=( a84966a  and  a84959a );
 a84970a <=( (not A236)  and  (not A235) );
 a84973a <=( (not A268)  and  (not A266) );
 a84974a <=( a84973a  and  a84970a );
 a84977a <=( A298  and  (not A269) );
 a84981a <=( A301  and  A300 );
 a84982a <=( (not A299)  and  a84981a );
 a84983a <=( a84982a  and  a84977a );
 a84984a <=( a84983a  and  a84974a );
 a84987a <=( (not A167)  and  A170 );
 a84990a <=( A199  and  (not A166) );
 a84991a <=( a84990a  and  a84987a );
 a84994a <=( A201  and  (not A200) );
 a84997a <=( (not A233)  and  A202 );
 a84998a <=( a84997a  and  a84994a );
 a84999a <=( a84998a  and  a84991a );
 a85002a <=( (not A236)  and  (not A235) );
 a85005a <=( (not A268)  and  (not A266) );
 a85006a <=( a85005a  and  a85002a );
 a85009a <=( A298  and  (not A269) );
 a85013a <=( A302  and  A300 );
 a85014a <=( (not A299)  and  a85013a );
 a85015a <=( a85014a  and  a85009a );
 a85016a <=( a85015a  and  a85006a );
 a85019a <=( (not A167)  and  A170 );
 a85022a <=( A199  and  (not A166) );
 a85023a <=( a85022a  and  a85019a );
 a85026a <=( A201  and  (not A200) );
 a85029a <=( (not A233)  and  A203 );
 a85030a <=( a85029a  and  a85026a );
 a85031a <=( a85030a  and  a85023a );
 a85034a <=( (not A236)  and  (not A235) );
 a85037a <=( (not A268)  and  (not A266) );
 a85038a <=( a85037a  and  a85034a );
 a85041a <=( A298  and  (not A269) );
 a85045a <=( A301  and  A300 );
 a85046a <=( (not A299)  and  a85045a );
 a85047a <=( a85046a  and  a85041a );
 a85048a <=( a85047a  and  a85038a );
 a85051a <=( (not A167)  and  A170 );
 a85054a <=( A199  and  (not A166) );
 a85055a <=( a85054a  and  a85051a );
 a85058a <=( A201  and  (not A200) );
 a85061a <=( (not A233)  and  A203 );
 a85062a <=( a85061a  and  a85058a );
 a85063a <=( a85062a  and  a85055a );
 a85066a <=( (not A236)  and  (not A235) );
 a85069a <=( (not A268)  and  (not A266) );
 a85070a <=( a85069a  and  a85066a );
 a85073a <=( A298  and  (not A269) );
 a85077a <=( A302  and  A300 );
 a85078a <=( (not A299)  and  a85077a );
 a85079a <=( a85078a  and  a85073a );
 a85080a <=( a85079a  and  a85070a );
 a85083a <=( (not A168)  and  A169 );
 a85086a <=( (not A166)  and  A167 );
 a85087a <=( a85086a  and  a85083a );
 a85090a <=( (not A200)  and  A199 );
 a85093a <=( A202  and  A201 );
 a85094a <=( a85093a  and  a85090a );
 a85095a <=( a85094a  and  a85087a );
 a85098a <=( A233  and  A232 );
 a85101a <=( (not A268)  and  A265 );
 a85102a <=( a85101a  and  a85098a );
 a85105a <=( A298  and  (not A269) );
 a85109a <=( A301  and  A300 );
 a85110a <=( (not A299)  and  a85109a );
 a85111a <=( a85110a  and  a85105a );
 a85112a <=( a85111a  and  a85102a );
 a85115a <=( (not A168)  and  A169 );
 a85118a <=( (not A166)  and  A167 );
 a85119a <=( a85118a  and  a85115a );
 a85122a <=( (not A200)  and  A199 );
 a85125a <=( A202  and  A201 );
 a85126a <=( a85125a  and  a85122a );
 a85127a <=( a85126a  and  a85119a );
 a85130a <=( A233  and  A232 );
 a85133a <=( (not A268)  and  A265 );
 a85134a <=( a85133a  and  a85130a );
 a85137a <=( A298  and  (not A269) );
 a85141a <=( A302  and  A300 );
 a85142a <=( (not A299)  and  a85141a );
 a85143a <=( a85142a  and  a85137a );
 a85144a <=( a85143a  and  a85134a );
 a85147a <=( (not A168)  and  A169 );
 a85150a <=( (not A166)  and  A167 );
 a85151a <=( a85150a  and  a85147a );
 a85154a <=( (not A200)  and  A199 );
 a85157a <=( A202  and  A201 );
 a85158a <=( a85157a  and  a85154a );
 a85159a <=( a85158a  and  a85151a );
 a85162a <=( (not A235)  and  (not A233) );
 a85165a <=( A265  and  (not A236) );
 a85166a <=( a85165a  and  a85162a );
 a85169a <=( A298  and  A266 );
 a85173a <=( A301  and  A300 );
 a85174a <=( (not A299)  and  a85173a );
 a85175a <=( a85174a  and  a85169a );
 a85176a <=( a85175a  and  a85166a );
 a85179a <=( (not A168)  and  A169 );
 a85182a <=( (not A166)  and  A167 );
 a85183a <=( a85182a  and  a85179a );
 a85186a <=( (not A200)  and  A199 );
 a85189a <=( A202  and  A201 );
 a85190a <=( a85189a  and  a85186a );
 a85191a <=( a85190a  and  a85183a );
 a85194a <=( (not A235)  and  (not A233) );
 a85197a <=( A265  and  (not A236) );
 a85198a <=( a85197a  and  a85194a );
 a85201a <=( A298  and  A266 );
 a85205a <=( A302  and  A300 );
 a85206a <=( (not A299)  and  a85205a );
 a85207a <=( a85206a  and  a85201a );
 a85208a <=( a85207a  and  a85198a );
 a85211a <=( (not A168)  and  A169 );
 a85214a <=( (not A166)  and  A167 );
 a85215a <=( a85214a  and  a85211a );
 a85218a <=( (not A200)  and  A199 );
 a85221a <=( A202  and  A201 );
 a85222a <=( a85221a  and  a85218a );
 a85223a <=( a85222a  and  a85215a );
 a85226a <=( (not A235)  and  (not A233) );
 a85229a <=( (not A266)  and  (not A236) );
 a85230a <=( a85229a  and  a85226a );
 a85233a <=( A298  and  (not A267) );
 a85237a <=( A301  and  A300 );
 a85238a <=( (not A299)  and  a85237a );
 a85239a <=( a85238a  and  a85233a );
 a85240a <=( a85239a  and  a85230a );
 a85243a <=( (not A168)  and  A169 );
 a85246a <=( (not A166)  and  A167 );
 a85247a <=( a85246a  and  a85243a );
 a85250a <=( (not A200)  and  A199 );
 a85253a <=( A202  and  A201 );
 a85254a <=( a85253a  and  a85250a );
 a85255a <=( a85254a  and  a85247a );
 a85258a <=( (not A235)  and  (not A233) );
 a85261a <=( (not A266)  and  (not A236) );
 a85262a <=( a85261a  and  a85258a );
 a85265a <=( A298  and  (not A267) );
 a85269a <=( A302  and  A300 );
 a85270a <=( (not A299)  and  a85269a );
 a85271a <=( a85270a  and  a85265a );
 a85272a <=( a85271a  and  a85262a );
 a85275a <=( (not A168)  and  A169 );
 a85278a <=( (not A166)  and  A167 );
 a85279a <=( a85278a  and  a85275a );
 a85282a <=( (not A200)  and  A199 );
 a85285a <=( A202  and  A201 );
 a85286a <=( a85285a  and  a85282a );
 a85287a <=( a85286a  and  a85279a );
 a85290a <=( (not A235)  and  (not A233) );
 a85293a <=( (not A265)  and  (not A236) );
 a85294a <=( a85293a  and  a85290a );
 a85297a <=( A298  and  (not A266) );
 a85301a <=( A301  and  A300 );
 a85302a <=( (not A299)  and  a85301a );
 a85303a <=( a85302a  and  a85297a );
 a85304a <=( a85303a  and  a85294a );
 a85307a <=( (not A168)  and  A169 );
 a85310a <=( (not A166)  and  A167 );
 a85311a <=( a85310a  and  a85307a );
 a85314a <=( (not A200)  and  A199 );
 a85317a <=( A202  and  A201 );
 a85318a <=( a85317a  and  a85314a );
 a85319a <=( a85318a  and  a85311a );
 a85322a <=( (not A235)  and  (not A233) );
 a85325a <=( (not A265)  and  (not A236) );
 a85326a <=( a85325a  and  a85322a );
 a85329a <=( A298  and  (not A266) );
 a85333a <=( A302  and  A300 );
 a85334a <=( (not A299)  and  a85333a );
 a85335a <=( a85334a  and  a85329a );
 a85336a <=( a85335a  and  a85326a );
 a85339a <=( (not A168)  and  A169 );
 a85342a <=( (not A166)  and  A167 );
 a85343a <=( a85342a  and  a85339a );
 a85346a <=( (not A200)  and  A199 );
 a85349a <=( A202  and  A201 );
 a85350a <=( a85349a  and  a85346a );
 a85351a <=( a85350a  and  a85343a );
 a85354a <=( (not A234)  and  (not A233) );
 a85357a <=( (not A268)  and  (not A266) );
 a85358a <=( a85357a  and  a85354a );
 a85361a <=( A298  and  (not A269) );
 a85365a <=( A301  and  A300 );
 a85366a <=( (not A299)  and  a85365a );
 a85367a <=( a85366a  and  a85361a );
 a85368a <=( a85367a  and  a85358a );
 a85371a <=( (not A168)  and  A169 );
 a85374a <=( (not A166)  and  A167 );
 a85375a <=( a85374a  and  a85371a );
 a85378a <=( (not A200)  and  A199 );
 a85381a <=( A202  and  A201 );
 a85382a <=( a85381a  and  a85378a );
 a85383a <=( a85382a  and  a85375a );
 a85386a <=( (not A234)  and  (not A233) );
 a85389a <=( (not A268)  and  (not A266) );
 a85390a <=( a85389a  and  a85386a );
 a85393a <=( A298  and  (not A269) );
 a85397a <=( A302  and  A300 );
 a85398a <=( (not A299)  and  a85397a );
 a85399a <=( a85398a  and  a85393a );
 a85400a <=( a85399a  and  a85390a );
 a85403a <=( (not A168)  and  A169 );
 a85406a <=( (not A166)  and  A167 );
 a85407a <=( a85406a  and  a85403a );
 a85410a <=( (not A200)  and  A199 );
 a85413a <=( A202  and  A201 );
 a85414a <=( a85413a  and  a85410a );
 a85415a <=( a85414a  and  a85407a );
 a85418a <=( (not A233)  and  (not A232) );
 a85421a <=( (not A268)  and  (not A266) );
 a85422a <=( a85421a  and  a85418a );
 a85425a <=( A298  and  (not A269) );
 a85429a <=( A301  and  A300 );
 a85430a <=( (not A299)  and  a85429a );
 a85431a <=( a85430a  and  a85425a );
 a85432a <=( a85431a  and  a85422a );
 a85435a <=( (not A168)  and  A169 );
 a85438a <=( (not A166)  and  A167 );
 a85439a <=( a85438a  and  a85435a );
 a85442a <=( (not A200)  and  A199 );
 a85445a <=( A202  and  A201 );
 a85446a <=( a85445a  and  a85442a );
 a85447a <=( a85446a  and  a85439a );
 a85450a <=( (not A233)  and  (not A232) );
 a85453a <=( (not A268)  and  (not A266) );
 a85454a <=( a85453a  and  a85450a );
 a85457a <=( A298  and  (not A269) );
 a85461a <=( A302  and  A300 );
 a85462a <=( (not A299)  and  a85461a );
 a85463a <=( a85462a  and  a85457a );
 a85464a <=( a85463a  and  a85454a );
 a85467a <=( (not A168)  and  A169 );
 a85470a <=( (not A166)  and  A167 );
 a85471a <=( a85470a  and  a85467a );
 a85474a <=( (not A200)  and  A199 );
 a85477a <=( A203  and  A201 );
 a85478a <=( a85477a  and  a85474a );
 a85479a <=( a85478a  and  a85471a );
 a85482a <=( A233  and  A232 );
 a85485a <=( (not A268)  and  A265 );
 a85486a <=( a85485a  and  a85482a );
 a85489a <=( A298  and  (not A269) );
 a85493a <=( A301  and  A300 );
 a85494a <=( (not A299)  and  a85493a );
 a85495a <=( a85494a  and  a85489a );
 a85496a <=( a85495a  and  a85486a );
 a85499a <=( (not A168)  and  A169 );
 a85502a <=( (not A166)  and  A167 );
 a85503a <=( a85502a  and  a85499a );
 a85506a <=( (not A200)  and  A199 );
 a85509a <=( A203  and  A201 );
 a85510a <=( a85509a  and  a85506a );
 a85511a <=( a85510a  and  a85503a );
 a85514a <=( A233  and  A232 );
 a85517a <=( (not A268)  and  A265 );
 a85518a <=( a85517a  and  a85514a );
 a85521a <=( A298  and  (not A269) );
 a85525a <=( A302  and  A300 );
 a85526a <=( (not A299)  and  a85525a );
 a85527a <=( a85526a  and  a85521a );
 a85528a <=( a85527a  and  a85518a );
 a85531a <=( (not A168)  and  A169 );
 a85534a <=( (not A166)  and  A167 );
 a85535a <=( a85534a  and  a85531a );
 a85538a <=( (not A200)  and  A199 );
 a85541a <=( A203  and  A201 );
 a85542a <=( a85541a  and  a85538a );
 a85543a <=( a85542a  and  a85535a );
 a85546a <=( (not A235)  and  (not A233) );
 a85549a <=( A265  and  (not A236) );
 a85550a <=( a85549a  and  a85546a );
 a85553a <=( A298  and  A266 );
 a85557a <=( A301  and  A300 );
 a85558a <=( (not A299)  and  a85557a );
 a85559a <=( a85558a  and  a85553a );
 a85560a <=( a85559a  and  a85550a );
 a85563a <=( (not A168)  and  A169 );
 a85566a <=( (not A166)  and  A167 );
 a85567a <=( a85566a  and  a85563a );
 a85570a <=( (not A200)  and  A199 );
 a85573a <=( A203  and  A201 );
 a85574a <=( a85573a  and  a85570a );
 a85575a <=( a85574a  and  a85567a );
 a85578a <=( (not A235)  and  (not A233) );
 a85581a <=( A265  and  (not A236) );
 a85582a <=( a85581a  and  a85578a );
 a85585a <=( A298  and  A266 );
 a85589a <=( A302  and  A300 );
 a85590a <=( (not A299)  and  a85589a );
 a85591a <=( a85590a  and  a85585a );
 a85592a <=( a85591a  and  a85582a );
 a85595a <=( (not A168)  and  A169 );
 a85598a <=( (not A166)  and  A167 );
 a85599a <=( a85598a  and  a85595a );
 a85602a <=( (not A200)  and  A199 );
 a85605a <=( A203  and  A201 );
 a85606a <=( a85605a  and  a85602a );
 a85607a <=( a85606a  and  a85599a );
 a85610a <=( (not A235)  and  (not A233) );
 a85613a <=( (not A266)  and  (not A236) );
 a85614a <=( a85613a  and  a85610a );
 a85617a <=( A298  and  (not A267) );
 a85621a <=( A301  and  A300 );
 a85622a <=( (not A299)  and  a85621a );
 a85623a <=( a85622a  and  a85617a );
 a85624a <=( a85623a  and  a85614a );
 a85627a <=( (not A168)  and  A169 );
 a85630a <=( (not A166)  and  A167 );
 a85631a <=( a85630a  and  a85627a );
 a85634a <=( (not A200)  and  A199 );
 a85637a <=( A203  and  A201 );
 a85638a <=( a85637a  and  a85634a );
 a85639a <=( a85638a  and  a85631a );
 a85642a <=( (not A235)  and  (not A233) );
 a85645a <=( (not A266)  and  (not A236) );
 a85646a <=( a85645a  and  a85642a );
 a85649a <=( A298  and  (not A267) );
 a85653a <=( A302  and  A300 );
 a85654a <=( (not A299)  and  a85653a );
 a85655a <=( a85654a  and  a85649a );
 a85656a <=( a85655a  and  a85646a );
 a85659a <=( (not A168)  and  A169 );
 a85662a <=( (not A166)  and  A167 );
 a85663a <=( a85662a  and  a85659a );
 a85666a <=( (not A200)  and  A199 );
 a85669a <=( A203  and  A201 );
 a85670a <=( a85669a  and  a85666a );
 a85671a <=( a85670a  and  a85663a );
 a85674a <=( (not A235)  and  (not A233) );
 a85677a <=( (not A265)  and  (not A236) );
 a85678a <=( a85677a  and  a85674a );
 a85681a <=( A298  and  (not A266) );
 a85685a <=( A301  and  A300 );
 a85686a <=( (not A299)  and  a85685a );
 a85687a <=( a85686a  and  a85681a );
 a85688a <=( a85687a  and  a85678a );
 a85691a <=( (not A168)  and  A169 );
 a85694a <=( (not A166)  and  A167 );
 a85695a <=( a85694a  and  a85691a );
 a85698a <=( (not A200)  and  A199 );
 a85701a <=( A203  and  A201 );
 a85702a <=( a85701a  and  a85698a );
 a85703a <=( a85702a  and  a85695a );
 a85706a <=( (not A235)  and  (not A233) );
 a85709a <=( (not A265)  and  (not A236) );
 a85710a <=( a85709a  and  a85706a );
 a85713a <=( A298  and  (not A266) );
 a85717a <=( A302  and  A300 );
 a85718a <=( (not A299)  and  a85717a );
 a85719a <=( a85718a  and  a85713a );
 a85720a <=( a85719a  and  a85710a );
 a85723a <=( (not A168)  and  A169 );
 a85726a <=( (not A166)  and  A167 );
 a85727a <=( a85726a  and  a85723a );
 a85730a <=( (not A200)  and  A199 );
 a85733a <=( A203  and  A201 );
 a85734a <=( a85733a  and  a85730a );
 a85735a <=( a85734a  and  a85727a );
 a85738a <=( (not A234)  and  (not A233) );
 a85741a <=( (not A268)  and  (not A266) );
 a85742a <=( a85741a  and  a85738a );
 a85745a <=( A298  and  (not A269) );
 a85749a <=( A301  and  A300 );
 a85750a <=( (not A299)  and  a85749a );
 a85751a <=( a85750a  and  a85745a );
 a85752a <=( a85751a  and  a85742a );
 a85755a <=( (not A168)  and  A169 );
 a85758a <=( (not A166)  and  A167 );
 a85759a <=( a85758a  and  a85755a );
 a85762a <=( (not A200)  and  A199 );
 a85765a <=( A203  and  A201 );
 a85766a <=( a85765a  and  a85762a );
 a85767a <=( a85766a  and  a85759a );
 a85770a <=( (not A234)  and  (not A233) );
 a85773a <=( (not A268)  and  (not A266) );
 a85774a <=( a85773a  and  a85770a );
 a85777a <=( A298  and  (not A269) );
 a85781a <=( A302  and  A300 );
 a85782a <=( (not A299)  and  a85781a );
 a85783a <=( a85782a  and  a85777a );
 a85784a <=( a85783a  and  a85774a );
 a85787a <=( (not A168)  and  A169 );
 a85790a <=( (not A166)  and  A167 );
 a85791a <=( a85790a  and  a85787a );
 a85794a <=( (not A200)  and  A199 );
 a85797a <=( A203  and  A201 );
 a85798a <=( a85797a  and  a85794a );
 a85799a <=( a85798a  and  a85791a );
 a85802a <=( (not A233)  and  (not A232) );
 a85805a <=( (not A268)  and  (not A266) );
 a85806a <=( a85805a  and  a85802a );
 a85809a <=( A298  and  (not A269) );
 a85813a <=( A301  and  A300 );
 a85814a <=( (not A299)  and  a85813a );
 a85815a <=( a85814a  and  a85809a );
 a85816a <=( a85815a  and  a85806a );
 a85819a <=( (not A168)  and  A169 );
 a85822a <=( (not A166)  and  A167 );
 a85823a <=( a85822a  and  a85819a );
 a85826a <=( (not A200)  and  A199 );
 a85829a <=( A203  and  A201 );
 a85830a <=( a85829a  and  a85826a );
 a85831a <=( a85830a  and  a85823a );
 a85834a <=( (not A233)  and  (not A232) );
 a85837a <=( (not A268)  and  (not A266) );
 a85838a <=( a85837a  and  a85834a );
 a85841a <=( A298  and  (not A269) );
 a85845a <=( A302  and  A300 );
 a85846a <=( (not A299)  and  a85845a );
 a85847a <=( a85846a  and  a85841a );
 a85848a <=( a85847a  and  a85838a );
 a85851a <=( (not A168)  and  A169 );
 a85854a <=( A166  and  (not A167) );
 a85855a <=( a85854a  and  a85851a );
 a85858a <=( (not A200)  and  A199 );
 a85861a <=( A202  and  A201 );
 a85862a <=( a85861a  and  a85858a );
 a85863a <=( a85862a  and  a85855a );
 a85866a <=( A233  and  A232 );
 a85869a <=( (not A268)  and  A265 );
 a85870a <=( a85869a  and  a85866a );
 a85873a <=( A298  and  (not A269) );
 a85877a <=( A301  and  A300 );
 a85878a <=( (not A299)  and  a85877a );
 a85879a <=( a85878a  and  a85873a );
 a85880a <=( a85879a  and  a85870a );
 a85883a <=( (not A168)  and  A169 );
 a85886a <=( A166  and  (not A167) );
 a85887a <=( a85886a  and  a85883a );
 a85890a <=( (not A200)  and  A199 );
 a85893a <=( A202  and  A201 );
 a85894a <=( a85893a  and  a85890a );
 a85895a <=( a85894a  and  a85887a );
 a85898a <=( A233  and  A232 );
 a85901a <=( (not A268)  and  A265 );
 a85902a <=( a85901a  and  a85898a );
 a85905a <=( A298  and  (not A269) );
 a85909a <=( A302  and  A300 );
 a85910a <=( (not A299)  and  a85909a );
 a85911a <=( a85910a  and  a85905a );
 a85912a <=( a85911a  and  a85902a );
 a85915a <=( (not A168)  and  A169 );
 a85918a <=( A166  and  (not A167) );
 a85919a <=( a85918a  and  a85915a );
 a85922a <=( (not A200)  and  A199 );
 a85925a <=( A202  and  A201 );
 a85926a <=( a85925a  and  a85922a );
 a85927a <=( a85926a  and  a85919a );
 a85930a <=( (not A235)  and  (not A233) );
 a85933a <=( A265  and  (not A236) );
 a85934a <=( a85933a  and  a85930a );
 a85937a <=( A298  and  A266 );
 a85941a <=( A301  and  A300 );
 a85942a <=( (not A299)  and  a85941a );
 a85943a <=( a85942a  and  a85937a );
 a85944a <=( a85943a  and  a85934a );
 a85947a <=( (not A168)  and  A169 );
 a85950a <=( A166  and  (not A167) );
 a85951a <=( a85950a  and  a85947a );
 a85954a <=( (not A200)  and  A199 );
 a85957a <=( A202  and  A201 );
 a85958a <=( a85957a  and  a85954a );
 a85959a <=( a85958a  and  a85951a );
 a85962a <=( (not A235)  and  (not A233) );
 a85965a <=( A265  and  (not A236) );
 a85966a <=( a85965a  and  a85962a );
 a85969a <=( A298  and  A266 );
 a85973a <=( A302  and  A300 );
 a85974a <=( (not A299)  and  a85973a );
 a85975a <=( a85974a  and  a85969a );
 a85976a <=( a85975a  and  a85966a );
 a85979a <=( (not A168)  and  A169 );
 a85982a <=( A166  and  (not A167) );
 a85983a <=( a85982a  and  a85979a );
 a85986a <=( (not A200)  and  A199 );
 a85989a <=( A202  and  A201 );
 a85990a <=( a85989a  and  a85986a );
 a85991a <=( a85990a  and  a85983a );
 a85994a <=( (not A235)  and  (not A233) );
 a85997a <=( (not A266)  and  (not A236) );
 a85998a <=( a85997a  and  a85994a );
 a86001a <=( A298  and  (not A267) );
 a86005a <=( A301  and  A300 );
 a86006a <=( (not A299)  and  a86005a );
 a86007a <=( a86006a  and  a86001a );
 a86008a <=( a86007a  and  a85998a );
 a86011a <=( (not A168)  and  A169 );
 a86014a <=( A166  and  (not A167) );
 a86015a <=( a86014a  and  a86011a );
 a86018a <=( (not A200)  and  A199 );
 a86021a <=( A202  and  A201 );
 a86022a <=( a86021a  and  a86018a );
 a86023a <=( a86022a  and  a86015a );
 a86026a <=( (not A235)  and  (not A233) );
 a86029a <=( (not A266)  and  (not A236) );
 a86030a <=( a86029a  and  a86026a );
 a86033a <=( A298  and  (not A267) );
 a86037a <=( A302  and  A300 );
 a86038a <=( (not A299)  and  a86037a );
 a86039a <=( a86038a  and  a86033a );
 a86040a <=( a86039a  and  a86030a );
 a86043a <=( (not A168)  and  A169 );
 a86046a <=( A166  and  (not A167) );
 a86047a <=( a86046a  and  a86043a );
 a86050a <=( (not A200)  and  A199 );
 a86053a <=( A202  and  A201 );
 a86054a <=( a86053a  and  a86050a );
 a86055a <=( a86054a  and  a86047a );
 a86058a <=( (not A235)  and  (not A233) );
 a86061a <=( (not A265)  and  (not A236) );
 a86062a <=( a86061a  and  a86058a );
 a86065a <=( A298  and  (not A266) );
 a86069a <=( A301  and  A300 );
 a86070a <=( (not A299)  and  a86069a );
 a86071a <=( a86070a  and  a86065a );
 a86072a <=( a86071a  and  a86062a );
 a86075a <=( (not A168)  and  A169 );
 a86078a <=( A166  and  (not A167) );
 a86079a <=( a86078a  and  a86075a );
 a86082a <=( (not A200)  and  A199 );
 a86085a <=( A202  and  A201 );
 a86086a <=( a86085a  and  a86082a );
 a86087a <=( a86086a  and  a86079a );
 a86090a <=( (not A235)  and  (not A233) );
 a86093a <=( (not A265)  and  (not A236) );
 a86094a <=( a86093a  and  a86090a );
 a86097a <=( A298  and  (not A266) );
 a86101a <=( A302  and  A300 );
 a86102a <=( (not A299)  and  a86101a );
 a86103a <=( a86102a  and  a86097a );
 a86104a <=( a86103a  and  a86094a );
 a86107a <=( (not A168)  and  A169 );
 a86110a <=( A166  and  (not A167) );
 a86111a <=( a86110a  and  a86107a );
 a86114a <=( (not A200)  and  A199 );
 a86117a <=( A202  and  A201 );
 a86118a <=( a86117a  and  a86114a );
 a86119a <=( a86118a  and  a86111a );
 a86122a <=( (not A234)  and  (not A233) );
 a86125a <=( (not A268)  and  (not A266) );
 a86126a <=( a86125a  and  a86122a );
 a86129a <=( A298  and  (not A269) );
 a86133a <=( A301  and  A300 );
 a86134a <=( (not A299)  and  a86133a );
 a86135a <=( a86134a  and  a86129a );
 a86136a <=( a86135a  and  a86126a );
 a86139a <=( (not A168)  and  A169 );
 a86142a <=( A166  and  (not A167) );
 a86143a <=( a86142a  and  a86139a );
 a86146a <=( (not A200)  and  A199 );
 a86149a <=( A202  and  A201 );
 a86150a <=( a86149a  and  a86146a );
 a86151a <=( a86150a  and  a86143a );
 a86154a <=( (not A234)  and  (not A233) );
 a86157a <=( (not A268)  and  (not A266) );
 a86158a <=( a86157a  and  a86154a );
 a86161a <=( A298  and  (not A269) );
 a86165a <=( A302  and  A300 );
 a86166a <=( (not A299)  and  a86165a );
 a86167a <=( a86166a  and  a86161a );
 a86168a <=( a86167a  and  a86158a );
 a86171a <=( (not A168)  and  A169 );
 a86174a <=( A166  and  (not A167) );
 a86175a <=( a86174a  and  a86171a );
 a86178a <=( (not A200)  and  A199 );
 a86181a <=( A202  and  A201 );
 a86182a <=( a86181a  and  a86178a );
 a86183a <=( a86182a  and  a86175a );
 a86186a <=( (not A233)  and  (not A232) );
 a86189a <=( (not A268)  and  (not A266) );
 a86190a <=( a86189a  and  a86186a );
 a86193a <=( A298  and  (not A269) );
 a86197a <=( A301  and  A300 );
 a86198a <=( (not A299)  and  a86197a );
 a86199a <=( a86198a  and  a86193a );
 a86200a <=( a86199a  and  a86190a );
 a86203a <=( (not A168)  and  A169 );
 a86206a <=( A166  and  (not A167) );
 a86207a <=( a86206a  and  a86203a );
 a86210a <=( (not A200)  and  A199 );
 a86213a <=( A202  and  A201 );
 a86214a <=( a86213a  and  a86210a );
 a86215a <=( a86214a  and  a86207a );
 a86218a <=( (not A233)  and  (not A232) );
 a86221a <=( (not A268)  and  (not A266) );
 a86222a <=( a86221a  and  a86218a );
 a86225a <=( A298  and  (not A269) );
 a86229a <=( A302  and  A300 );
 a86230a <=( (not A299)  and  a86229a );
 a86231a <=( a86230a  and  a86225a );
 a86232a <=( a86231a  and  a86222a );
 a86235a <=( (not A168)  and  A169 );
 a86238a <=( A166  and  (not A167) );
 a86239a <=( a86238a  and  a86235a );
 a86242a <=( (not A200)  and  A199 );
 a86245a <=( A203  and  A201 );
 a86246a <=( a86245a  and  a86242a );
 a86247a <=( a86246a  and  a86239a );
 a86250a <=( A233  and  A232 );
 a86253a <=( (not A268)  and  A265 );
 a86254a <=( a86253a  and  a86250a );
 a86257a <=( A298  and  (not A269) );
 a86261a <=( A301  and  A300 );
 a86262a <=( (not A299)  and  a86261a );
 a86263a <=( a86262a  and  a86257a );
 a86264a <=( a86263a  and  a86254a );
 a86267a <=( (not A168)  and  A169 );
 a86270a <=( A166  and  (not A167) );
 a86271a <=( a86270a  and  a86267a );
 a86274a <=( (not A200)  and  A199 );
 a86277a <=( A203  and  A201 );
 a86278a <=( a86277a  and  a86274a );
 a86279a <=( a86278a  and  a86271a );
 a86282a <=( A233  and  A232 );
 a86285a <=( (not A268)  and  A265 );
 a86286a <=( a86285a  and  a86282a );
 a86289a <=( A298  and  (not A269) );
 a86293a <=( A302  and  A300 );
 a86294a <=( (not A299)  and  a86293a );
 a86295a <=( a86294a  and  a86289a );
 a86296a <=( a86295a  and  a86286a );
 a86299a <=( (not A168)  and  A169 );
 a86302a <=( A166  and  (not A167) );
 a86303a <=( a86302a  and  a86299a );
 a86306a <=( (not A200)  and  A199 );
 a86309a <=( A203  and  A201 );
 a86310a <=( a86309a  and  a86306a );
 a86311a <=( a86310a  and  a86303a );
 a86314a <=( (not A235)  and  (not A233) );
 a86317a <=( A265  and  (not A236) );
 a86318a <=( a86317a  and  a86314a );
 a86321a <=( A298  and  A266 );
 a86325a <=( A301  and  A300 );
 a86326a <=( (not A299)  and  a86325a );
 a86327a <=( a86326a  and  a86321a );
 a86328a <=( a86327a  and  a86318a );
 a86331a <=( (not A168)  and  A169 );
 a86334a <=( A166  and  (not A167) );
 a86335a <=( a86334a  and  a86331a );
 a86338a <=( (not A200)  and  A199 );
 a86341a <=( A203  and  A201 );
 a86342a <=( a86341a  and  a86338a );
 a86343a <=( a86342a  and  a86335a );
 a86346a <=( (not A235)  and  (not A233) );
 a86349a <=( A265  and  (not A236) );
 a86350a <=( a86349a  and  a86346a );
 a86353a <=( A298  and  A266 );
 a86357a <=( A302  and  A300 );
 a86358a <=( (not A299)  and  a86357a );
 a86359a <=( a86358a  and  a86353a );
 a86360a <=( a86359a  and  a86350a );
 a86363a <=( (not A168)  and  A169 );
 a86366a <=( A166  and  (not A167) );
 a86367a <=( a86366a  and  a86363a );
 a86370a <=( (not A200)  and  A199 );
 a86373a <=( A203  and  A201 );
 a86374a <=( a86373a  and  a86370a );
 a86375a <=( a86374a  and  a86367a );
 a86378a <=( (not A235)  and  (not A233) );
 a86381a <=( (not A266)  and  (not A236) );
 a86382a <=( a86381a  and  a86378a );
 a86385a <=( A298  and  (not A267) );
 a86389a <=( A301  and  A300 );
 a86390a <=( (not A299)  and  a86389a );
 a86391a <=( a86390a  and  a86385a );
 a86392a <=( a86391a  and  a86382a );
 a86395a <=( (not A168)  and  A169 );
 a86398a <=( A166  and  (not A167) );
 a86399a <=( a86398a  and  a86395a );
 a86402a <=( (not A200)  and  A199 );
 a86405a <=( A203  and  A201 );
 a86406a <=( a86405a  and  a86402a );
 a86407a <=( a86406a  and  a86399a );
 a86410a <=( (not A235)  and  (not A233) );
 a86413a <=( (not A266)  and  (not A236) );
 a86414a <=( a86413a  and  a86410a );
 a86417a <=( A298  and  (not A267) );
 a86421a <=( A302  and  A300 );
 a86422a <=( (not A299)  and  a86421a );
 a86423a <=( a86422a  and  a86417a );
 a86424a <=( a86423a  and  a86414a );
 a86427a <=( (not A168)  and  A169 );
 a86430a <=( A166  and  (not A167) );
 a86431a <=( a86430a  and  a86427a );
 a86434a <=( (not A200)  and  A199 );
 a86437a <=( A203  and  A201 );
 a86438a <=( a86437a  and  a86434a );
 a86439a <=( a86438a  and  a86431a );
 a86442a <=( (not A235)  and  (not A233) );
 a86445a <=( (not A265)  and  (not A236) );
 a86446a <=( a86445a  and  a86442a );
 a86449a <=( A298  and  (not A266) );
 a86453a <=( A301  and  A300 );
 a86454a <=( (not A299)  and  a86453a );
 a86455a <=( a86454a  and  a86449a );
 a86456a <=( a86455a  and  a86446a );
 a86459a <=( (not A168)  and  A169 );
 a86462a <=( A166  and  (not A167) );
 a86463a <=( a86462a  and  a86459a );
 a86466a <=( (not A200)  and  A199 );
 a86469a <=( A203  and  A201 );
 a86470a <=( a86469a  and  a86466a );
 a86471a <=( a86470a  and  a86463a );
 a86474a <=( (not A235)  and  (not A233) );
 a86477a <=( (not A265)  and  (not A236) );
 a86478a <=( a86477a  and  a86474a );
 a86481a <=( A298  and  (not A266) );
 a86485a <=( A302  and  A300 );
 a86486a <=( (not A299)  and  a86485a );
 a86487a <=( a86486a  and  a86481a );
 a86488a <=( a86487a  and  a86478a );
 a86491a <=( (not A168)  and  A169 );
 a86494a <=( A166  and  (not A167) );
 a86495a <=( a86494a  and  a86491a );
 a86498a <=( (not A200)  and  A199 );
 a86501a <=( A203  and  A201 );
 a86502a <=( a86501a  and  a86498a );
 a86503a <=( a86502a  and  a86495a );
 a86506a <=( (not A234)  and  (not A233) );
 a86509a <=( (not A268)  and  (not A266) );
 a86510a <=( a86509a  and  a86506a );
 a86513a <=( A298  and  (not A269) );
 a86517a <=( A301  and  A300 );
 a86518a <=( (not A299)  and  a86517a );
 a86519a <=( a86518a  and  a86513a );
 a86520a <=( a86519a  and  a86510a );
 a86523a <=( (not A168)  and  A169 );
 a86526a <=( A166  and  (not A167) );
 a86527a <=( a86526a  and  a86523a );
 a86530a <=( (not A200)  and  A199 );
 a86533a <=( A203  and  A201 );
 a86534a <=( a86533a  and  a86530a );
 a86535a <=( a86534a  and  a86527a );
 a86538a <=( (not A234)  and  (not A233) );
 a86541a <=( (not A268)  and  (not A266) );
 a86542a <=( a86541a  and  a86538a );
 a86545a <=( A298  and  (not A269) );
 a86549a <=( A302  and  A300 );
 a86550a <=( (not A299)  and  a86549a );
 a86551a <=( a86550a  and  a86545a );
 a86552a <=( a86551a  and  a86542a );
 a86555a <=( (not A168)  and  A169 );
 a86558a <=( A166  and  (not A167) );
 a86559a <=( a86558a  and  a86555a );
 a86562a <=( (not A200)  and  A199 );
 a86565a <=( A203  and  A201 );
 a86566a <=( a86565a  and  a86562a );
 a86567a <=( a86566a  and  a86559a );
 a86570a <=( (not A233)  and  (not A232) );
 a86573a <=( (not A268)  and  (not A266) );
 a86574a <=( a86573a  and  a86570a );
 a86577a <=( A298  and  (not A269) );
 a86581a <=( A301  and  A300 );
 a86582a <=( (not A299)  and  a86581a );
 a86583a <=( a86582a  and  a86577a );
 a86584a <=( a86583a  and  a86574a );
 a86587a <=( (not A168)  and  A169 );
 a86590a <=( A166  and  (not A167) );
 a86591a <=( a86590a  and  a86587a );
 a86594a <=( (not A200)  and  A199 );
 a86597a <=( A203  and  A201 );
 a86598a <=( a86597a  and  a86594a );
 a86599a <=( a86598a  and  a86591a );
 a86602a <=( (not A233)  and  (not A232) );
 a86605a <=( (not A268)  and  (not A266) );
 a86606a <=( a86605a  and  a86602a );
 a86609a <=( A298  and  (not A269) );
 a86613a <=( A302  and  A300 );
 a86614a <=( (not A299)  and  a86613a );
 a86615a <=( a86614a  and  a86609a );
 a86616a <=( a86615a  and  a86606a );
 a86619a <=( A169  and  A170 );
 a86622a <=( A199  and  (not A168) );
 a86623a <=( a86622a  and  a86619a );
 a86626a <=( A201  and  (not A200) );
 a86629a <=( (not A233)  and  A202 );
 a86630a <=( a86629a  and  a86626a );
 a86631a <=( a86630a  and  a86623a );
 a86634a <=( (not A236)  and  (not A235) );
 a86637a <=( (not A268)  and  (not A266) );
 a86638a <=( a86637a  and  a86634a );
 a86641a <=( A298  and  (not A269) );
 a86645a <=( A301  and  A300 );
 a86646a <=( (not A299)  and  a86645a );
 a86647a <=( a86646a  and  a86641a );
 a86648a <=( a86647a  and  a86638a );
 a86651a <=( A169  and  A170 );
 a86654a <=( A199  and  (not A168) );
 a86655a <=( a86654a  and  a86651a );
 a86658a <=( A201  and  (not A200) );
 a86661a <=( (not A233)  and  A202 );
 a86662a <=( a86661a  and  a86658a );
 a86663a <=( a86662a  and  a86655a );
 a86666a <=( (not A236)  and  (not A235) );
 a86669a <=( (not A268)  and  (not A266) );
 a86670a <=( a86669a  and  a86666a );
 a86673a <=( A298  and  (not A269) );
 a86677a <=( A302  and  A300 );
 a86678a <=( (not A299)  and  a86677a );
 a86679a <=( a86678a  and  a86673a );
 a86680a <=( a86679a  and  a86670a );
 a86683a <=( A169  and  A170 );
 a86686a <=( A199  and  (not A168) );
 a86687a <=( a86686a  and  a86683a );
 a86690a <=( A201  and  (not A200) );
 a86693a <=( (not A233)  and  A203 );
 a86694a <=( a86693a  and  a86690a );
 a86695a <=( a86694a  and  a86687a );
 a86698a <=( (not A236)  and  (not A235) );
 a86701a <=( (not A268)  and  (not A266) );
 a86702a <=( a86701a  and  a86698a );
 a86705a <=( A298  and  (not A269) );
 a86709a <=( A301  and  A300 );
 a86710a <=( (not A299)  and  a86709a );
 a86711a <=( a86710a  and  a86705a );
 a86712a <=( a86711a  and  a86702a );
 a86715a <=( A169  and  A170 );
 a86718a <=( A199  and  (not A168) );
 a86719a <=( a86718a  and  a86715a );
 a86722a <=( A201  and  (not A200) );
 a86725a <=( (not A233)  and  A203 );
 a86726a <=( a86725a  and  a86722a );
 a86727a <=( a86726a  and  a86719a );
 a86730a <=( (not A236)  and  (not A235) );
 a86733a <=( (not A268)  and  (not A266) );
 a86734a <=( a86733a  and  a86730a );
 a86737a <=( A298  and  (not A269) );
 a86741a <=( A302  and  A300 );
 a86742a <=( (not A299)  and  a86741a );
 a86743a <=( a86742a  and  a86737a );
 a86744a <=( a86743a  and  a86734a );
 a86747a <=( A169  and  A170 );
 a86750a <=( A166  and  (not A168) );
 a86751a <=( a86750a  and  a86747a );
 a86754a <=( (not A200)  and  A199 );
 a86757a <=( A202  and  A201 );
 a86758a <=( a86757a  and  a86754a );
 a86759a <=( a86758a  and  a86751a );
 a86762a <=( (not A234)  and  (not A233) );
 a86765a <=( (not A268)  and  (not A266) );
 a86766a <=( a86765a  and  a86762a );
 a86769a <=( A298  and  (not A269) );
 a86773a <=( A301  and  A300 );
 a86774a <=( (not A299)  and  a86773a );
 a86775a <=( a86774a  and  a86769a );
 a86776a <=( a86775a  and  a86766a );
 a86779a <=( A169  and  A170 );
 a86782a <=( A166  and  (not A168) );
 a86783a <=( a86782a  and  a86779a );
 a86786a <=( (not A200)  and  A199 );
 a86789a <=( A202  and  A201 );
 a86790a <=( a86789a  and  a86786a );
 a86791a <=( a86790a  and  a86783a );
 a86794a <=( (not A234)  and  (not A233) );
 a86797a <=( (not A268)  and  (not A266) );
 a86798a <=( a86797a  and  a86794a );
 a86801a <=( A298  and  (not A269) );
 a86805a <=( A302  and  A300 );
 a86806a <=( (not A299)  and  a86805a );
 a86807a <=( a86806a  and  a86801a );
 a86808a <=( a86807a  and  a86798a );
 a86811a <=( A169  and  A170 );
 a86814a <=( A166  and  (not A168) );
 a86815a <=( a86814a  and  a86811a );
 a86818a <=( (not A200)  and  A199 );
 a86821a <=( A202  and  A201 );
 a86822a <=( a86821a  and  a86818a );
 a86823a <=( a86822a  and  a86815a );
 a86826a <=( (not A233)  and  (not A232) );
 a86829a <=( (not A268)  and  (not A266) );
 a86830a <=( a86829a  and  a86826a );
 a86833a <=( A298  and  (not A269) );
 a86837a <=( A301  and  A300 );
 a86838a <=( (not A299)  and  a86837a );
 a86839a <=( a86838a  and  a86833a );
 a86840a <=( a86839a  and  a86830a );
 a86843a <=( A169  and  A170 );
 a86846a <=( A166  and  (not A168) );
 a86847a <=( a86846a  and  a86843a );
 a86850a <=( (not A200)  and  A199 );
 a86853a <=( A202  and  A201 );
 a86854a <=( a86853a  and  a86850a );
 a86855a <=( a86854a  and  a86847a );
 a86858a <=( (not A233)  and  (not A232) );
 a86861a <=( (not A268)  and  (not A266) );
 a86862a <=( a86861a  and  a86858a );
 a86865a <=( A298  and  (not A269) );
 a86869a <=( A302  and  A300 );
 a86870a <=( (not A299)  and  a86869a );
 a86871a <=( a86870a  and  a86865a );
 a86872a <=( a86871a  and  a86862a );
 a86875a <=( A169  and  A170 );
 a86878a <=( A166  and  (not A168) );
 a86879a <=( a86878a  and  a86875a );
 a86882a <=( (not A200)  and  A199 );
 a86885a <=( A203  and  A201 );
 a86886a <=( a86885a  and  a86882a );
 a86887a <=( a86886a  and  a86879a );
 a86890a <=( (not A234)  and  (not A233) );
 a86893a <=( (not A268)  and  (not A266) );
 a86894a <=( a86893a  and  a86890a );
 a86897a <=( A298  and  (not A269) );
 a86901a <=( A301  and  A300 );
 a86902a <=( (not A299)  and  a86901a );
 a86903a <=( a86902a  and  a86897a );
 a86904a <=( a86903a  and  a86894a );
 a86907a <=( A169  and  A170 );
 a86910a <=( A166  and  (not A168) );
 a86911a <=( a86910a  and  a86907a );
 a86914a <=( (not A200)  and  A199 );
 a86917a <=( A203  and  A201 );
 a86918a <=( a86917a  and  a86914a );
 a86919a <=( a86918a  and  a86911a );
 a86922a <=( (not A234)  and  (not A233) );
 a86925a <=( (not A268)  and  (not A266) );
 a86926a <=( a86925a  and  a86922a );
 a86929a <=( A298  and  (not A269) );
 a86933a <=( A302  and  A300 );
 a86934a <=( (not A299)  and  a86933a );
 a86935a <=( a86934a  and  a86929a );
 a86936a <=( a86935a  and  a86926a );
 a86939a <=( A169  and  A170 );
 a86942a <=( A166  and  (not A168) );
 a86943a <=( a86942a  and  a86939a );
 a86946a <=( (not A200)  and  A199 );
 a86949a <=( A203  and  A201 );
 a86950a <=( a86949a  and  a86946a );
 a86951a <=( a86950a  and  a86943a );
 a86954a <=( (not A233)  and  (not A232) );
 a86957a <=( (not A268)  and  (not A266) );
 a86958a <=( a86957a  and  a86954a );
 a86961a <=( A298  and  (not A269) );
 a86965a <=( A301  and  A300 );
 a86966a <=( (not A299)  and  a86965a );
 a86967a <=( a86966a  and  a86961a );
 a86968a <=( a86967a  and  a86958a );
 a86971a <=( A169  and  A170 );
 a86974a <=( A166  and  (not A168) );
 a86975a <=( a86974a  and  a86971a );
 a86978a <=( (not A200)  and  A199 );
 a86981a <=( A203  and  A201 );
 a86982a <=( a86981a  and  a86978a );
 a86983a <=( a86982a  and  a86975a );
 a86986a <=( (not A233)  and  (not A232) );
 a86989a <=( (not A268)  and  (not A266) );
 a86990a <=( a86989a  and  a86986a );
 a86993a <=( A298  and  (not A269) );
 a86997a <=( A302  and  A300 );
 a86998a <=( (not A299)  and  a86997a );
 a86999a <=( a86998a  and  a86993a );
 a87000a <=( a86999a  and  a86990a );
 a87003a <=( A169  and  (not A170) );
 a87006a <=( A166  and  A167 );
 a87007a <=( a87006a  and  a87003a );
 a87010a <=( (not A202)  and  (not A200) );
 a87013a <=( (not A233)  and  (not A203) );
 a87014a <=( a87013a  and  a87010a );
 a87015a <=( a87014a  and  a87007a );
 a87018a <=( (not A236)  and  (not A235) );
 a87021a <=( (not A268)  and  (not A266) );
 a87022a <=( a87021a  and  a87018a );
 a87025a <=( A298  and  (not A269) );
 a87029a <=( A301  and  A300 );
 a87030a <=( (not A299)  and  a87029a );
 a87031a <=( a87030a  and  a87025a );
 a87032a <=( a87031a  and  a87022a );
 a87035a <=( A169  and  (not A170) );
 a87038a <=( A166  and  A167 );
 a87039a <=( a87038a  and  a87035a );
 a87042a <=( (not A202)  and  (not A200) );
 a87045a <=( (not A233)  and  (not A203) );
 a87046a <=( a87045a  and  a87042a );
 a87047a <=( a87046a  and  a87039a );
 a87050a <=( (not A236)  and  (not A235) );
 a87053a <=( (not A268)  and  (not A266) );
 a87054a <=( a87053a  and  a87050a );
 a87057a <=( A298  and  (not A269) );
 a87061a <=( A302  and  A300 );
 a87062a <=( (not A299)  and  a87061a );
 a87063a <=( a87062a  and  a87057a );
 a87064a <=( a87063a  and  a87054a );
 a87067a <=( A169  and  (not A170) );
 a87070a <=( (not A166)  and  (not A167) );
 a87071a <=( a87070a  and  a87067a );
 a87074a <=( (not A202)  and  (not A200) );
 a87077a <=( (not A233)  and  (not A203) );
 a87078a <=( a87077a  and  a87074a );
 a87079a <=( a87078a  and  a87071a );
 a87082a <=( (not A236)  and  (not A235) );
 a87085a <=( (not A268)  and  (not A266) );
 a87086a <=( a87085a  and  a87082a );
 a87089a <=( A298  and  (not A269) );
 a87093a <=( A301  and  A300 );
 a87094a <=( (not A299)  and  a87093a );
 a87095a <=( a87094a  and  a87089a );
 a87096a <=( a87095a  and  a87086a );
 a87099a <=( A169  and  (not A170) );
 a87102a <=( (not A166)  and  (not A167) );
 a87103a <=( a87102a  and  a87099a );
 a87106a <=( (not A202)  and  (not A200) );
 a87109a <=( (not A233)  and  (not A203) );
 a87110a <=( a87109a  and  a87106a );
 a87111a <=( a87110a  and  a87103a );
 a87114a <=( (not A236)  and  (not A235) );
 a87117a <=( (not A268)  and  (not A266) );
 a87118a <=( a87117a  and  a87114a );
 a87121a <=( A298  and  (not A269) );
 a87125a <=( A302  and  A300 );
 a87126a <=( (not A299)  and  a87125a );
 a87127a <=( a87126a  and  a87121a );
 a87128a <=( a87127a  and  a87118a );
 a87131a <=( (not A167)  and  (not A169) );
 a87134a <=( A199  and  (not A166) );
 a87135a <=( a87134a  and  a87131a );
 a87138a <=( A201  and  (not A200) );
 a87141a <=( (not A233)  and  A202 );
 a87142a <=( a87141a  and  a87138a );
 a87143a <=( a87142a  and  a87135a );
 a87146a <=( (not A236)  and  (not A235) );
 a87149a <=( (not A268)  and  (not A266) );
 a87150a <=( a87149a  and  a87146a );
 a87153a <=( A298  and  (not A269) );
 a87157a <=( A301  and  A300 );
 a87158a <=( (not A299)  and  a87157a );
 a87159a <=( a87158a  and  a87153a );
 a87160a <=( a87159a  and  a87150a );
 a87163a <=( (not A167)  and  (not A169) );
 a87166a <=( A199  and  (not A166) );
 a87167a <=( a87166a  and  a87163a );
 a87170a <=( A201  and  (not A200) );
 a87173a <=( (not A233)  and  A202 );
 a87174a <=( a87173a  and  a87170a );
 a87175a <=( a87174a  and  a87167a );
 a87178a <=( (not A236)  and  (not A235) );
 a87181a <=( (not A268)  and  (not A266) );
 a87182a <=( a87181a  and  a87178a );
 a87185a <=( A298  and  (not A269) );
 a87189a <=( A302  and  A300 );
 a87190a <=( (not A299)  and  a87189a );
 a87191a <=( a87190a  and  a87185a );
 a87192a <=( a87191a  and  a87182a );
 a87195a <=( (not A167)  and  (not A169) );
 a87198a <=( A199  and  (not A166) );
 a87199a <=( a87198a  and  a87195a );
 a87202a <=( A201  and  (not A200) );
 a87205a <=( (not A233)  and  A203 );
 a87206a <=( a87205a  and  a87202a );
 a87207a <=( a87206a  and  a87199a );
 a87210a <=( (not A236)  and  (not A235) );
 a87213a <=( (not A268)  and  (not A266) );
 a87214a <=( a87213a  and  a87210a );
 a87217a <=( A298  and  (not A269) );
 a87221a <=( A301  and  A300 );
 a87222a <=( (not A299)  and  a87221a );
 a87223a <=( a87222a  and  a87217a );
 a87224a <=( a87223a  and  a87214a );
 a87227a <=( (not A167)  and  (not A169) );
 a87230a <=( A199  and  (not A166) );
 a87231a <=( a87230a  and  a87227a );
 a87234a <=( A201  and  (not A200) );
 a87237a <=( (not A233)  and  A203 );
 a87238a <=( a87237a  and  a87234a );
 a87239a <=( a87238a  and  a87231a );
 a87242a <=( (not A236)  and  (not A235) );
 a87245a <=( (not A268)  and  (not A266) );
 a87246a <=( a87245a  and  a87242a );
 a87249a <=( A298  and  (not A269) );
 a87253a <=( A302  and  A300 );
 a87254a <=( (not A299)  and  a87253a );
 a87255a <=( a87254a  and  a87249a );
 a87256a <=( a87255a  and  a87246a );
 a87259a <=( (not A168)  and  (not A169) );
 a87262a <=( A166  and  A167 );
 a87263a <=( a87262a  and  a87259a );
 a87266a <=( (not A200)  and  A199 );
 a87269a <=( A202  and  A201 );
 a87270a <=( a87269a  and  a87266a );
 a87271a <=( a87270a  and  a87263a );
 a87274a <=( A233  and  A232 );
 a87277a <=( (not A268)  and  A265 );
 a87278a <=( a87277a  and  a87274a );
 a87281a <=( A298  and  (not A269) );
 a87285a <=( A301  and  A300 );
 a87286a <=( (not A299)  and  a87285a );
 a87287a <=( a87286a  and  a87281a );
 a87288a <=( a87287a  and  a87278a );
 a87291a <=( (not A168)  and  (not A169) );
 a87294a <=( A166  and  A167 );
 a87295a <=( a87294a  and  a87291a );
 a87298a <=( (not A200)  and  A199 );
 a87301a <=( A202  and  A201 );
 a87302a <=( a87301a  and  a87298a );
 a87303a <=( a87302a  and  a87295a );
 a87306a <=( A233  and  A232 );
 a87309a <=( (not A268)  and  A265 );
 a87310a <=( a87309a  and  a87306a );
 a87313a <=( A298  and  (not A269) );
 a87317a <=( A302  and  A300 );
 a87318a <=( (not A299)  and  a87317a );
 a87319a <=( a87318a  and  a87313a );
 a87320a <=( a87319a  and  a87310a );
 a87323a <=( (not A168)  and  (not A169) );
 a87326a <=( A166  and  A167 );
 a87327a <=( a87326a  and  a87323a );
 a87330a <=( (not A200)  and  A199 );
 a87333a <=( A202  and  A201 );
 a87334a <=( a87333a  and  a87330a );
 a87335a <=( a87334a  and  a87327a );
 a87338a <=( (not A235)  and  (not A233) );
 a87341a <=( A265  and  (not A236) );
 a87342a <=( a87341a  and  a87338a );
 a87345a <=( A298  and  A266 );
 a87349a <=( A301  and  A300 );
 a87350a <=( (not A299)  and  a87349a );
 a87351a <=( a87350a  and  a87345a );
 a87352a <=( a87351a  and  a87342a );
 a87355a <=( (not A168)  and  (not A169) );
 a87358a <=( A166  and  A167 );
 a87359a <=( a87358a  and  a87355a );
 a87362a <=( (not A200)  and  A199 );
 a87365a <=( A202  and  A201 );
 a87366a <=( a87365a  and  a87362a );
 a87367a <=( a87366a  and  a87359a );
 a87370a <=( (not A235)  and  (not A233) );
 a87373a <=( A265  and  (not A236) );
 a87374a <=( a87373a  and  a87370a );
 a87377a <=( A298  and  A266 );
 a87381a <=( A302  and  A300 );
 a87382a <=( (not A299)  and  a87381a );
 a87383a <=( a87382a  and  a87377a );
 a87384a <=( a87383a  and  a87374a );
 a87387a <=( (not A168)  and  (not A169) );
 a87390a <=( A166  and  A167 );
 a87391a <=( a87390a  and  a87387a );
 a87394a <=( (not A200)  and  A199 );
 a87397a <=( A202  and  A201 );
 a87398a <=( a87397a  and  a87394a );
 a87399a <=( a87398a  and  a87391a );
 a87402a <=( (not A235)  and  (not A233) );
 a87405a <=( (not A266)  and  (not A236) );
 a87406a <=( a87405a  and  a87402a );
 a87409a <=( A298  and  (not A267) );
 a87413a <=( A301  and  A300 );
 a87414a <=( (not A299)  and  a87413a );
 a87415a <=( a87414a  and  a87409a );
 a87416a <=( a87415a  and  a87406a );
 a87419a <=( (not A168)  and  (not A169) );
 a87422a <=( A166  and  A167 );
 a87423a <=( a87422a  and  a87419a );
 a87426a <=( (not A200)  and  A199 );
 a87429a <=( A202  and  A201 );
 a87430a <=( a87429a  and  a87426a );
 a87431a <=( a87430a  and  a87423a );
 a87434a <=( (not A235)  and  (not A233) );
 a87437a <=( (not A266)  and  (not A236) );
 a87438a <=( a87437a  and  a87434a );
 a87441a <=( A298  and  (not A267) );
 a87445a <=( A302  and  A300 );
 a87446a <=( (not A299)  and  a87445a );
 a87447a <=( a87446a  and  a87441a );
 a87448a <=( a87447a  and  a87438a );
 a87451a <=( (not A168)  and  (not A169) );
 a87454a <=( A166  and  A167 );
 a87455a <=( a87454a  and  a87451a );
 a87458a <=( (not A200)  and  A199 );
 a87461a <=( A202  and  A201 );
 a87462a <=( a87461a  and  a87458a );
 a87463a <=( a87462a  and  a87455a );
 a87466a <=( (not A235)  and  (not A233) );
 a87469a <=( (not A265)  and  (not A236) );
 a87470a <=( a87469a  and  a87466a );
 a87473a <=( A298  and  (not A266) );
 a87477a <=( A301  and  A300 );
 a87478a <=( (not A299)  and  a87477a );
 a87479a <=( a87478a  and  a87473a );
 a87480a <=( a87479a  and  a87470a );
 a87483a <=( (not A168)  and  (not A169) );
 a87486a <=( A166  and  A167 );
 a87487a <=( a87486a  and  a87483a );
 a87490a <=( (not A200)  and  A199 );
 a87493a <=( A202  and  A201 );
 a87494a <=( a87493a  and  a87490a );
 a87495a <=( a87494a  and  a87487a );
 a87498a <=( (not A235)  and  (not A233) );
 a87501a <=( (not A265)  and  (not A236) );
 a87502a <=( a87501a  and  a87498a );
 a87505a <=( A298  and  (not A266) );
 a87509a <=( A302  and  A300 );
 a87510a <=( (not A299)  and  a87509a );
 a87511a <=( a87510a  and  a87505a );
 a87512a <=( a87511a  and  a87502a );
 a87515a <=( (not A168)  and  (not A169) );
 a87518a <=( A166  and  A167 );
 a87519a <=( a87518a  and  a87515a );
 a87522a <=( (not A200)  and  A199 );
 a87525a <=( A202  and  A201 );
 a87526a <=( a87525a  and  a87522a );
 a87527a <=( a87526a  and  a87519a );
 a87530a <=( (not A234)  and  (not A233) );
 a87533a <=( (not A268)  and  (not A266) );
 a87534a <=( a87533a  and  a87530a );
 a87537a <=( A298  and  (not A269) );
 a87541a <=( A301  and  A300 );
 a87542a <=( (not A299)  and  a87541a );
 a87543a <=( a87542a  and  a87537a );
 a87544a <=( a87543a  and  a87534a );
 a87547a <=( (not A168)  and  (not A169) );
 a87550a <=( A166  and  A167 );
 a87551a <=( a87550a  and  a87547a );
 a87554a <=( (not A200)  and  A199 );
 a87557a <=( A202  and  A201 );
 a87558a <=( a87557a  and  a87554a );
 a87559a <=( a87558a  and  a87551a );
 a87562a <=( (not A234)  and  (not A233) );
 a87565a <=( (not A268)  and  (not A266) );
 a87566a <=( a87565a  and  a87562a );
 a87569a <=( A298  and  (not A269) );
 a87573a <=( A302  and  A300 );
 a87574a <=( (not A299)  and  a87573a );
 a87575a <=( a87574a  and  a87569a );
 a87576a <=( a87575a  and  a87566a );
 a87579a <=( (not A168)  and  (not A169) );
 a87582a <=( A166  and  A167 );
 a87583a <=( a87582a  and  a87579a );
 a87586a <=( (not A200)  and  A199 );
 a87589a <=( A202  and  A201 );
 a87590a <=( a87589a  and  a87586a );
 a87591a <=( a87590a  and  a87583a );
 a87594a <=( (not A233)  and  (not A232) );
 a87597a <=( (not A268)  and  (not A266) );
 a87598a <=( a87597a  and  a87594a );
 a87601a <=( A298  and  (not A269) );
 a87605a <=( A301  and  A300 );
 a87606a <=( (not A299)  and  a87605a );
 a87607a <=( a87606a  and  a87601a );
 a87608a <=( a87607a  and  a87598a );
 a87611a <=( (not A168)  and  (not A169) );
 a87614a <=( A166  and  A167 );
 a87615a <=( a87614a  and  a87611a );
 a87618a <=( (not A200)  and  A199 );
 a87621a <=( A202  and  A201 );
 a87622a <=( a87621a  and  a87618a );
 a87623a <=( a87622a  and  a87615a );
 a87626a <=( (not A233)  and  (not A232) );
 a87629a <=( (not A268)  and  (not A266) );
 a87630a <=( a87629a  and  a87626a );
 a87633a <=( A298  and  (not A269) );
 a87637a <=( A302  and  A300 );
 a87638a <=( (not A299)  and  a87637a );
 a87639a <=( a87638a  and  a87633a );
 a87640a <=( a87639a  and  a87630a );
 a87643a <=( (not A168)  and  (not A169) );
 a87646a <=( A166  and  A167 );
 a87647a <=( a87646a  and  a87643a );
 a87650a <=( (not A200)  and  A199 );
 a87653a <=( A203  and  A201 );
 a87654a <=( a87653a  and  a87650a );
 a87655a <=( a87654a  and  a87647a );
 a87658a <=( A233  and  A232 );
 a87661a <=( (not A268)  and  A265 );
 a87662a <=( a87661a  and  a87658a );
 a87665a <=( A298  and  (not A269) );
 a87669a <=( A301  and  A300 );
 a87670a <=( (not A299)  and  a87669a );
 a87671a <=( a87670a  and  a87665a );
 a87672a <=( a87671a  and  a87662a );
 a87675a <=( (not A168)  and  (not A169) );
 a87678a <=( A166  and  A167 );
 a87679a <=( a87678a  and  a87675a );
 a87682a <=( (not A200)  and  A199 );
 a87685a <=( A203  and  A201 );
 a87686a <=( a87685a  and  a87682a );
 a87687a <=( a87686a  and  a87679a );
 a87690a <=( A233  and  A232 );
 a87693a <=( (not A268)  and  A265 );
 a87694a <=( a87693a  and  a87690a );
 a87697a <=( A298  and  (not A269) );
 a87701a <=( A302  and  A300 );
 a87702a <=( (not A299)  and  a87701a );
 a87703a <=( a87702a  and  a87697a );
 a87704a <=( a87703a  and  a87694a );
 a87707a <=( (not A168)  and  (not A169) );
 a87710a <=( A166  and  A167 );
 a87711a <=( a87710a  and  a87707a );
 a87714a <=( (not A200)  and  A199 );
 a87717a <=( A203  and  A201 );
 a87718a <=( a87717a  and  a87714a );
 a87719a <=( a87718a  and  a87711a );
 a87722a <=( (not A235)  and  (not A233) );
 a87725a <=( A265  and  (not A236) );
 a87726a <=( a87725a  and  a87722a );
 a87729a <=( A298  and  A266 );
 a87733a <=( A301  and  A300 );
 a87734a <=( (not A299)  and  a87733a );
 a87735a <=( a87734a  and  a87729a );
 a87736a <=( a87735a  and  a87726a );
 a87739a <=( (not A168)  and  (not A169) );
 a87742a <=( A166  and  A167 );
 a87743a <=( a87742a  and  a87739a );
 a87746a <=( (not A200)  and  A199 );
 a87749a <=( A203  and  A201 );
 a87750a <=( a87749a  and  a87746a );
 a87751a <=( a87750a  and  a87743a );
 a87754a <=( (not A235)  and  (not A233) );
 a87757a <=( A265  and  (not A236) );
 a87758a <=( a87757a  and  a87754a );
 a87761a <=( A298  and  A266 );
 a87765a <=( A302  and  A300 );
 a87766a <=( (not A299)  and  a87765a );
 a87767a <=( a87766a  and  a87761a );
 a87768a <=( a87767a  and  a87758a );
 a87771a <=( (not A168)  and  (not A169) );
 a87774a <=( A166  and  A167 );
 a87775a <=( a87774a  and  a87771a );
 a87778a <=( (not A200)  and  A199 );
 a87781a <=( A203  and  A201 );
 a87782a <=( a87781a  and  a87778a );
 a87783a <=( a87782a  and  a87775a );
 a87786a <=( (not A235)  and  (not A233) );
 a87789a <=( (not A266)  and  (not A236) );
 a87790a <=( a87789a  and  a87786a );
 a87793a <=( A298  and  (not A267) );
 a87797a <=( A301  and  A300 );
 a87798a <=( (not A299)  and  a87797a );
 a87799a <=( a87798a  and  a87793a );
 a87800a <=( a87799a  and  a87790a );
 a87803a <=( (not A168)  and  (not A169) );
 a87806a <=( A166  and  A167 );
 a87807a <=( a87806a  and  a87803a );
 a87810a <=( (not A200)  and  A199 );
 a87813a <=( A203  and  A201 );
 a87814a <=( a87813a  and  a87810a );
 a87815a <=( a87814a  and  a87807a );
 a87818a <=( (not A235)  and  (not A233) );
 a87821a <=( (not A266)  and  (not A236) );
 a87822a <=( a87821a  and  a87818a );
 a87825a <=( A298  and  (not A267) );
 a87829a <=( A302  and  A300 );
 a87830a <=( (not A299)  and  a87829a );
 a87831a <=( a87830a  and  a87825a );
 a87832a <=( a87831a  and  a87822a );
 a87835a <=( (not A168)  and  (not A169) );
 a87838a <=( A166  and  A167 );
 a87839a <=( a87838a  and  a87835a );
 a87842a <=( (not A200)  and  A199 );
 a87845a <=( A203  and  A201 );
 a87846a <=( a87845a  and  a87842a );
 a87847a <=( a87846a  and  a87839a );
 a87850a <=( (not A235)  and  (not A233) );
 a87853a <=( (not A265)  and  (not A236) );
 a87854a <=( a87853a  and  a87850a );
 a87857a <=( A298  and  (not A266) );
 a87861a <=( A301  and  A300 );
 a87862a <=( (not A299)  and  a87861a );
 a87863a <=( a87862a  and  a87857a );
 a87864a <=( a87863a  and  a87854a );
 a87867a <=( (not A168)  and  (not A169) );
 a87870a <=( A166  and  A167 );
 a87871a <=( a87870a  and  a87867a );
 a87874a <=( (not A200)  and  A199 );
 a87877a <=( A203  and  A201 );
 a87878a <=( a87877a  and  a87874a );
 a87879a <=( a87878a  and  a87871a );
 a87882a <=( (not A235)  and  (not A233) );
 a87885a <=( (not A265)  and  (not A236) );
 a87886a <=( a87885a  and  a87882a );
 a87889a <=( A298  and  (not A266) );
 a87893a <=( A302  and  A300 );
 a87894a <=( (not A299)  and  a87893a );
 a87895a <=( a87894a  and  a87889a );
 a87896a <=( a87895a  and  a87886a );
 a87899a <=( (not A168)  and  (not A169) );
 a87902a <=( A166  and  A167 );
 a87903a <=( a87902a  and  a87899a );
 a87906a <=( (not A200)  and  A199 );
 a87909a <=( A203  and  A201 );
 a87910a <=( a87909a  and  a87906a );
 a87911a <=( a87910a  and  a87903a );
 a87914a <=( (not A234)  and  (not A233) );
 a87917a <=( (not A268)  and  (not A266) );
 a87918a <=( a87917a  and  a87914a );
 a87921a <=( A298  and  (not A269) );
 a87925a <=( A301  and  A300 );
 a87926a <=( (not A299)  and  a87925a );
 a87927a <=( a87926a  and  a87921a );
 a87928a <=( a87927a  and  a87918a );
 a87931a <=( (not A168)  and  (not A169) );
 a87934a <=( A166  and  A167 );
 a87935a <=( a87934a  and  a87931a );
 a87938a <=( (not A200)  and  A199 );
 a87941a <=( A203  and  A201 );
 a87942a <=( a87941a  and  a87938a );
 a87943a <=( a87942a  and  a87935a );
 a87946a <=( (not A234)  and  (not A233) );
 a87949a <=( (not A268)  and  (not A266) );
 a87950a <=( a87949a  and  a87946a );
 a87953a <=( A298  and  (not A269) );
 a87957a <=( A302  and  A300 );
 a87958a <=( (not A299)  and  a87957a );
 a87959a <=( a87958a  and  a87953a );
 a87960a <=( a87959a  and  a87950a );
 a87963a <=( (not A168)  and  (not A169) );
 a87966a <=( A166  and  A167 );
 a87967a <=( a87966a  and  a87963a );
 a87970a <=( (not A200)  and  A199 );
 a87973a <=( A203  and  A201 );
 a87974a <=( a87973a  and  a87970a );
 a87975a <=( a87974a  and  a87967a );
 a87978a <=( (not A233)  and  (not A232) );
 a87981a <=( (not A268)  and  (not A266) );
 a87982a <=( a87981a  and  a87978a );
 a87985a <=( A298  and  (not A269) );
 a87989a <=( A301  and  A300 );
 a87990a <=( (not A299)  and  a87989a );
 a87991a <=( a87990a  and  a87985a );
 a87992a <=( a87991a  and  a87982a );
 a87995a <=( (not A168)  and  (not A169) );
 a87998a <=( A166  and  A167 );
 a87999a <=( a87998a  and  a87995a );
 a88002a <=( (not A200)  and  A199 );
 a88005a <=( A203  and  A201 );
 a88006a <=( a88005a  and  a88002a );
 a88007a <=( a88006a  and  a87999a );
 a88010a <=( (not A233)  and  (not A232) );
 a88013a <=( (not A268)  and  (not A266) );
 a88014a <=( a88013a  and  a88010a );
 a88017a <=( A298  and  (not A269) );
 a88021a <=( A302  and  A300 );
 a88022a <=( (not A299)  and  a88021a );
 a88023a <=( a88022a  and  a88017a );
 a88024a <=( a88023a  and  a88014a );
 a88027a <=( (not A169)  and  A170 );
 a88030a <=( (not A166)  and  A167 );
 a88031a <=( a88030a  and  a88027a );
 a88034a <=( (not A202)  and  (not A200) );
 a88037a <=( (not A233)  and  (not A203) );
 a88038a <=( a88037a  and  a88034a );
 a88039a <=( a88038a  and  a88031a );
 a88042a <=( (not A236)  and  (not A235) );
 a88045a <=( (not A268)  and  (not A266) );
 a88046a <=( a88045a  and  a88042a );
 a88049a <=( A298  and  (not A269) );
 a88053a <=( A301  and  A300 );
 a88054a <=( (not A299)  and  a88053a );
 a88055a <=( a88054a  and  a88049a );
 a88056a <=( a88055a  and  a88046a );
 a88059a <=( (not A169)  and  A170 );
 a88062a <=( (not A166)  and  A167 );
 a88063a <=( a88062a  and  a88059a );
 a88066a <=( (not A202)  and  (not A200) );
 a88069a <=( (not A233)  and  (not A203) );
 a88070a <=( a88069a  and  a88066a );
 a88071a <=( a88070a  and  a88063a );
 a88074a <=( (not A236)  and  (not A235) );
 a88077a <=( (not A268)  and  (not A266) );
 a88078a <=( a88077a  and  a88074a );
 a88081a <=( A298  and  (not A269) );
 a88085a <=( A302  and  A300 );
 a88086a <=( (not A299)  and  a88085a );
 a88087a <=( a88086a  and  a88081a );
 a88088a <=( a88087a  and  a88078a );
 a88091a <=( (not A169)  and  A170 );
 a88094a <=( A166  and  (not A167) );
 a88095a <=( a88094a  and  a88091a );
 a88098a <=( (not A202)  and  (not A200) );
 a88101a <=( (not A233)  and  (not A203) );
 a88102a <=( a88101a  and  a88098a );
 a88103a <=( a88102a  and  a88095a );
 a88106a <=( (not A236)  and  (not A235) );
 a88109a <=( (not A268)  and  (not A266) );
 a88110a <=( a88109a  and  a88106a );
 a88113a <=( A298  and  (not A269) );
 a88117a <=( A301  and  A300 );
 a88118a <=( (not A299)  and  a88117a );
 a88119a <=( a88118a  and  a88113a );
 a88120a <=( a88119a  and  a88110a );
 a88123a <=( (not A169)  and  A170 );
 a88126a <=( A166  and  (not A167) );
 a88127a <=( a88126a  and  a88123a );
 a88130a <=( (not A202)  and  (not A200) );
 a88133a <=( (not A233)  and  (not A203) );
 a88134a <=( a88133a  and  a88130a );
 a88135a <=( a88134a  and  a88127a );
 a88138a <=( (not A236)  and  (not A235) );
 a88141a <=( (not A268)  and  (not A266) );
 a88142a <=( a88141a  and  a88138a );
 a88145a <=( A298  and  (not A269) );
 a88149a <=( A302  and  A300 );
 a88150a <=( (not A299)  and  a88149a );
 a88151a <=( a88150a  and  a88145a );
 a88152a <=( a88151a  and  a88142a );
 a88155a <=( (not A169)  and  (not A170) );
 a88158a <=( A199  and  (not A168) );
 a88159a <=( a88158a  and  a88155a );
 a88162a <=( A201  and  (not A200) );
 a88165a <=( (not A233)  and  A202 );
 a88166a <=( a88165a  and  a88162a );
 a88167a <=( a88166a  and  a88159a );
 a88170a <=( (not A236)  and  (not A235) );
 a88173a <=( (not A268)  and  (not A266) );
 a88174a <=( a88173a  and  a88170a );
 a88177a <=( A298  and  (not A269) );
 a88181a <=( A301  and  A300 );
 a88182a <=( (not A299)  and  a88181a );
 a88183a <=( a88182a  and  a88177a );
 a88184a <=( a88183a  and  a88174a );
 a88187a <=( (not A169)  and  (not A170) );
 a88190a <=( A199  and  (not A168) );
 a88191a <=( a88190a  and  a88187a );
 a88194a <=( A201  and  (not A200) );
 a88197a <=( (not A233)  and  A202 );
 a88198a <=( a88197a  and  a88194a );
 a88199a <=( a88198a  and  a88191a );
 a88202a <=( (not A236)  and  (not A235) );
 a88205a <=( (not A268)  and  (not A266) );
 a88206a <=( a88205a  and  a88202a );
 a88209a <=( A298  and  (not A269) );
 a88213a <=( A302  and  A300 );
 a88214a <=( (not A299)  and  a88213a );
 a88215a <=( a88214a  and  a88209a );
 a88216a <=( a88215a  and  a88206a );
 a88219a <=( (not A169)  and  (not A170) );
 a88222a <=( A199  and  (not A168) );
 a88223a <=( a88222a  and  a88219a );
 a88226a <=( A201  and  (not A200) );
 a88229a <=( (not A233)  and  A203 );
 a88230a <=( a88229a  and  a88226a );
 a88231a <=( a88230a  and  a88223a );
 a88234a <=( (not A236)  and  (not A235) );
 a88237a <=( (not A268)  and  (not A266) );
 a88238a <=( a88237a  and  a88234a );
 a88241a <=( A298  and  (not A269) );
 a88245a <=( A301  and  A300 );
 a88246a <=( (not A299)  and  a88245a );
 a88247a <=( a88246a  and  a88241a );
 a88248a <=( a88247a  and  a88238a );
 a88251a <=( (not A169)  and  (not A170) );
 a88254a <=( A199  and  (not A168) );
 a88255a <=( a88254a  and  a88251a );
 a88258a <=( A201  and  (not A200) );
 a88261a <=( (not A233)  and  A203 );
 a88262a <=( a88261a  and  a88258a );
 a88263a <=( a88262a  and  a88255a );
 a88266a <=( (not A236)  and  (not A235) );
 a88269a <=( (not A268)  and  (not A266) );
 a88270a <=( a88269a  and  a88266a );
 a88273a <=( A298  and  (not A269) );
 a88277a <=( A302  and  A300 );
 a88278a <=( (not A299)  and  a88277a );
 a88279a <=( a88278a  and  a88273a );
 a88280a <=( a88279a  and  a88270a );
 a88283a <=( (not A168)  and  A169 );
 a88286a <=( (not A166)  and  A167 );
 a88287a <=( a88286a  and  a88283a );
 a88290a <=( (not A200)  and  A199 );
 a88294a <=( (not A233)  and  A202 );
 a88295a <=( A201  and  a88294a );
 a88296a <=( a88295a  and  a88290a );
 a88297a <=( a88296a  and  a88287a );
 a88300a <=( (not A236)  and  (not A235) );
 a88303a <=( (not A268)  and  (not A266) );
 a88304a <=( a88303a  and  a88300a );
 a88307a <=( A298  and  (not A269) );
 a88311a <=( A301  and  A300 );
 a88312a <=( (not A299)  and  a88311a );
 a88313a <=( a88312a  and  a88307a );
 a88314a <=( a88313a  and  a88304a );
 a88317a <=( (not A168)  and  A169 );
 a88320a <=( (not A166)  and  A167 );
 a88321a <=( a88320a  and  a88317a );
 a88324a <=( (not A200)  and  A199 );
 a88328a <=( (not A233)  and  A202 );
 a88329a <=( A201  and  a88328a );
 a88330a <=( a88329a  and  a88324a );
 a88331a <=( a88330a  and  a88321a );
 a88334a <=( (not A236)  and  (not A235) );
 a88337a <=( (not A268)  and  (not A266) );
 a88338a <=( a88337a  and  a88334a );
 a88341a <=( A298  and  (not A269) );
 a88345a <=( A302  and  A300 );
 a88346a <=( (not A299)  and  a88345a );
 a88347a <=( a88346a  and  a88341a );
 a88348a <=( a88347a  and  a88338a );
 a88351a <=( (not A168)  and  A169 );
 a88354a <=( (not A166)  and  A167 );
 a88355a <=( a88354a  and  a88351a );
 a88358a <=( (not A200)  and  A199 );
 a88362a <=( (not A233)  and  A203 );
 a88363a <=( A201  and  a88362a );
 a88364a <=( a88363a  and  a88358a );
 a88365a <=( a88364a  and  a88355a );
 a88368a <=( (not A236)  and  (not A235) );
 a88371a <=( (not A268)  and  (not A266) );
 a88372a <=( a88371a  and  a88368a );
 a88375a <=( A298  and  (not A269) );
 a88379a <=( A301  and  A300 );
 a88380a <=( (not A299)  and  a88379a );
 a88381a <=( a88380a  and  a88375a );
 a88382a <=( a88381a  and  a88372a );
 a88385a <=( (not A168)  and  A169 );
 a88388a <=( (not A166)  and  A167 );
 a88389a <=( a88388a  and  a88385a );
 a88392a <=( (not A200)  and  A199 );
 a88396a <=( (not A233)  and  A203 );
 a88397a <=( A201  and  a88396a );
 a88398a <=( a88397a  and  a88392a );
 a88399a <=( a88398a  and  a88389a );
 a88402a <=( (not A236)  and  (not A235) );
 a88405a <=( (not A268)  and  (not A266) );
 a88406a <=( a88405a  and  a88402a );
 a88409a <=( A298  and  (not A269) );
 a88413a <=( A302  and  A300 );
 a88414a <=( (not A299)  and  a88413a );
 a88415a <=( a88414a  and  a88409a );
 a88416a <=( a88415a  and  a88406a );
 a88419a <=( (not A168)  and  A169 );
 a88422a <=( A166  and  (not A167) );
 a88423a <=( a88422a  and  a88419a );
 a88426a <=( (not A200)  and  A199 );
 a88430a <=( (not A233)  and  A202 );
 a88431a <=( A201  and  a88430a );
 a88432a <=( a88431a  and  a88426a );
 a88433a <=( a88432a  and  a88423a );
 a88436a <=( (not A236)  and  (not A235) );
 a88439a <=( (not A268)  and  (not A266) );
 a88440a <=( a88439a  and  a88436a );
 a88443a <=( A298  and  (not A269) );
 a88447a <=( A301  and  A300 );
 a88448a <=( (not A299)  and  a88447a );
 a88449a <=( a88448a  and  a88443a );
 a88450a <=( a88449a  and  a88440a );
 a88453a <=( (not A168)  and  A169 );
 a88456a <=( A166  and  (not A167) );
 a88457a <=( a88456a  and  a88453a );
 a88460a <=( (not A200)  and  A199 );
 a88464a <=( (not A233)  and  A202 );
 a88465a <=( A201  and  a88464a );
 a88466a <=( a88465a  and  a88460a );
 a88467a <=( a88466a  and  a88457a );
 a88470a <=( (not A236)  and  (not A235) );
 a88473a <=( (not A268)  and  (not A266) );
 a88474a <=( a88473a  and  a88470a );
 a88477a <=( A298  and  (not A269) );
 a88481a <=( A302  and  A300 );
 a88482a <=( (not A299)  and  a88481a );
 a88483a <=( a88482a  and  a88477a );
 a88484a <=( a88483a  and  a88474a );
 a88487a <=( (not A168)  and  A169 );
 a88490a <=( A166  and  (not A167) );
 a88491a <=( a88490a  and  a88487a );
 a88494a <=( (not A200)  and  A199 );
 a88498a <=( (not A233)  and  A203 );
 a88499a <=( A201  and  a88498a );
 a88500a <=( a88499a  and  a88494a );
 a88501a <=( a88500a  and  a88491a );
 a88504a <=( (not A236)  and  (not A235) );
 a88507a <=( (not A268)  and  (not A266) );
 a88508a <=( a88507a  and  a88504a );
 a88511a <=( A298  and  (not A269) );
 a88515a <=( A301  and  A300 );
 a88516a <=( (not A299)  and  a88515a );
 a88517a <=( a88516a  and  a88511a );
 a88518a <=( a88517a  and  a88508a );
 a88521a <=( (not A168)  and  A169 );
 a88524a <=( A166  and  (not A167) );
 a88525a <=( a88524a  and  a88521a );
 a88528a <=( (not A200)  and  A199 );
 a88532a <=( (not A233)  and  A203 );
 a88533a <=( A201  and  a88532a );
 a88534a <=( a88533a  and  a88528a );
 a88535a <=( a88534a  and  a88525a );
 a88538a <=( (not A236)  and  (not A235) );
 a88541a <=( (not A268)  and  (not A266) );
 a88542a <=( a88541a  and  a88538a );
 a88545a <=( A298  and  (not A269) );
 a88549a <=( A302  and  A300 );
 a88550a <=( (not A299)  and  a88549a );
 a88551a <=( a88550a  and  a88545a );
 a88552a <=( a88551a  and  a88542a );
 a88555a <=( (not A168)  and  (not A169) );
 a88558a <=( A166  and  A167 );
 a88559a <=( a88558a  and  a88555a );
 a88562a <=( (not A200)  and  A199 );
 a88566a <=( (not A233)  and  A202 );
 a88567a <=( A201  and  a88566a );
 a88568a <=( a88567a  and  a88562a );
 a88569a <=( a88568a  and  a88559a );
 a88572a <=( (not A236)  and  (not A235) );
 a88575a <=( (not A268)  and  (not A266) );
 a88576a <=( a88575a  and  a88572a );
 a88579a <=( A298  and  (not A269) );
 a88583a <=( A301  and  A300 );
 a88584a <=( (not A299)  and  a88583a );
 a88585a <=( a88584a  and  a88579a );
 a88586a <=( a88585a  and  a88576a );
 a88589a <=( (not A168)  and  (not A169) );
 a88592a <=( A166  and  A167 );
 a88593a <=( a88592a  and  a88589a );
 a88596a <=( (not A200)  and  A199 );
 a88600a <=( (not A233)  and  A202 );
 a88601a <=( A201  and  a88600a );
 a88602a <=( a88601a  and  a88596a );
 a88603a <=( a88602a  and  a88593a );
 a88606a <=( (not A236)  and  (not A235) );
 a88609a <=( (not A268)  and  (not A266) );
 a88610a <=( a88609a  and  a88606a );
 a88613a <=( A298  and  (not A269) );
 a88617a <=( A302  and  A300 );
 a88618a <=( (not A299)  and  a88617a );
 a88619a <=( a88618a  and  a88613a );
 a88620a <=( a88619a  and  a88610a );
 a88623a <=( (not A168)  and  (not A169) );
 a88626a <=( A166  and  A167 );
 a88627a <=( a88626a  and  a88623a );
 a88630a <=( (not A200)  and  A199 );
 a88634a <=( (not A233)  and  A203 );
 a88635a <=( A201  and  a88634a );
 a88636a <=( a88635a  and  a88630a );
 a88637a <=( a88636a  and  a88627a );
 a88640a <=( (not A236)  and  (not A235) );
 a88643a <=( (not A268)  and  (not A266) );
 a88644a <=( a88643a  and  a88640a );
 a88647a <=( A298  and  (not A269) );
 a88651a <=( A301  and  A300 );
 a88652a <=( (not A299)  and  a88651a );
 a88653a <=( a88652a  and  a88647a );
 a88654a <=( a88653a  and  a88644a );
 a88657a <=( (not A168)  and  (not A169) );
 a88660a <=( A166  and  A167 );
 a88661a <=( a88660a  and  a88657a );
 a88664a <=( (not A200)  and  A199 );
 a88668a <=( (not A233)  and  A203 );
 a88669a <=( A201  and  a88668a );
 a88670a <=( a88669a  and  a88664a );
 a88671a <=( a88670a  and  a88661a );
 a88674a <=( (not A236)  and  (not A235) );
 a88677a <=( (not A268)  and  (not A266) );
 a88678a <=( a88677a  and  a88674a );
 a88681a <=( A298  and  (not A269) );
 a88685a <=( A302  and  A300 );
 a88686a <=( (not A299)  and  a88685a );
 a88687a <=( a88686a  and  a88681a );
 a88688a <=( a88687a  and  a88678a );


end x25_10x_behav;
