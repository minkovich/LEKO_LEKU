Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_18x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A41: buffer std_logic
);
end x25_18x;

architecture x25_18x_behav of x25_18x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a351a,a355a,a356a,a357a,a360a,a364a,a365a,a366a,a367a,a370a,a374a,a375a,a376a,a380a,a381a,a385a,a386a,a387a,a388a,a389a,a392a,a396a,a397a,a398a,a402a,a403a,a407a,a408a,a409a,a410a,a413a,a417a,a418a,a419a,a423a,a424a,a428a,a429a,a430a,a431a,a432a,a433a,a436a,a440a,a441a,a442a,a446a,a447a,a451a,a452a,a453a,a454a,a457a,a461a,a462a,a463a,a467a,a468a,a472a,a473a,a474a,a475a,a476a,a479a,a483a,a484a,a485a,a489a,a490a,a494a,a495a,a496a,a497a,a500a,a504a,a505a,a506a,a510a,a511a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a524a,a528a,a529a,a530a,a533a,a537a,a538a,a539a,a540a,a543a,a547a,a548a,a549a,a553a,a554a,a558a,a559a,a560a,a561a,a562a,a565a,a569a,a570a,a571a,a575a,a576a,a580a,a581a,a582a,a583a,a586a,a590a,a591a,a592a,a596a,a597a,a601a,a602a,a603a,a604a,a605a,a606a,a609a,a613a,a614a,a615a,a619a,a620a,a624a,a625a,a626a,a627a,a630a,a634a,a635a,a636a,a640a,a641a,a645a,a646a,a647a,a648a,a649a,a652a,a656a,a657a,a658a,a662a,a663a,a667a,a668a,a669a,a670a,a673a,a677a,a678a,a679a,a683a,a684a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a698a,a702a,a703a,a704a,a707a,a711a,a712a,a713a,a714a,a717a,a721a,a722a,a723a,a727a,a728a,a732a,a733a,a734a,a735a,a736a,a739a,a743a,a744a,a745a,a749a,a750a,a754a,a755a,a756a,a757a,a760a,a764a,a765a,a766a,a770a,a771a,a775a,a776a,a777a,a778a,a779a,a780a,a783a,a787a,a788a,a789a,a793a,a794a,a798a,a799a,a800a,a801a,a804a,a808a,a809a,a810a,a814a,a815a,a819a,a820a,a821a,a822a,a823a,a826a,a830a,a831a,a832a,a836a,a837a,a841a,a842a,a843a,a844a,a847a,a851a,a852a,a853a,a857a,a858a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a871a,a875a,a876a,a877a,a880a,a884a,a885a,a886a,a887a,a890a,a894a,a895a,a896a,a900a,a901a,a905a,a906a,a907a,a908a,a909a,a912a,a916a,a917a,a918a,a922a,a923a,a927a,a928a,a929a,a930a,a933a,a937a,a938a,a939a,a943a,a944a,a948a,a949a,a950a,a951a,a952a,a953a,a956a,a960a,a961a,a962a,a966a,a967a,a971a,a972a,a973a,a974a,a977a,a981a,a982a,a983a,a987a,a988a,a992a,a993a,a994a,a995a,a996a,a999a,a1003a,a1004a,a1005a,a1009a,a1010a,a1014a,a1015a,a1016a,a1017a,a1020a,a1024a,a1025a,a1026a,a1030a,a1031a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1049a,a1052a,a1055a,a1058a,a1061a,a1064a,a1067a,a1070a,a1073a,a1076a,a1079a,a1082a,a1085a,a1088a,a1091a,a1094a,a1097a,a1100a,a1103a,a1106a,a1110a,a1111a,a1115a,a1116a,a1120a,a1121a,a1125a,a1126a,a1130a,a1131a,a1135a,a1136a,a1140a,a1141a,a1145a,a1146a,a1150a,a1151a,a1155a,a1156a,a1160a,a1161a,a1165a,a1166a,a1170a,a1171a,a1175a,a1176a,a1180a,a1181a,a1185a,a1186a,a1190a,a1191a,a1195a,a1196a,a1200a,a1201a,a1205a,a1206a,a1210a,a1211a,a1215a,a1216a,a1220a,a1221a,a1225a,a1226a,a1230a,a1231a,a1235a,a1236a,a1240a,a1241a,a1245a,a1246a,a1250a,a1251a,a1255a,a1256a,a1260a,a1261a,a1265a,a1266a,a1270a,a1271a,a1275a,a1276a,a1280a,a1281a,a1285a,a1286a,a1290a,a1291a,a1295a,a1296a,a1300a,a1301a,a1305a,a1306a,a1310a,a1311a,a1315a,a1316a,a1320a,a1321a,a1325a,a1326a,a1330a,a1331a,a1335a,a1336a,a1340a,a1341a,a1345a,a1346a,a1350a,a1351a,a1355a,a1356a,a1360a,a1361a,a1365a,a1366a,a1370a,a1371a,a1375a,a1376a,a1380a,a1381a,a1385a,a1386a,a1390a,a1391a,a1395a,a1396a,a1400a,a1401a,a1405a,a1406a,a1410a,a1411a,a1415a,a1416a,a1420a,a1421a,a1425a,a1426a,a1430a,a1431a,a1435a,a1436a,a1440a,a1441a,a1445a,a1446a,a1450a,a1451a,a1455a,a1456a,a1460a,a1461a,a1465a,a1466a,a1470a,a1471a,a1474a,a1477a,a1478a,a1482a,a1483a,a1486a,a1489a,a1490a,a1494a,a1495a,a1498a,a1501a,a1502a,a1506a,a1507a,a1510a,a1513a,a1514a,a1518a,a1519a,a1522a,a1525a,a1526a,a1530a,a1531a,a1534a,a1537a,a1538a,a1542a,a1543a,a1546a,a1549a,a1550a,a1554a,a1555a,a1558a,a1561a,a1562a,a1565a,a1568a,a1569a,a1572a,a1575a,a1576a,a1579a,a1582a,a1583a,a1586a,a1589a,a1590a,a1593a,a1596a,a1597a,a1600a,a1603a,a1604a,a1607a,a1610a,a1611a,a1614a,a1617a,a1618a,a1621a,a1624a,a1625a,a1628a,a1631a,a1632a,a1635a,a1638a,a1639a,a1642a,a1645a,a1646a,a1649a,a1652a,a1653a,a1656a,a1659a,a1660a,a1663a,a1666a,a1667a,a1670a,a1673a,a1674a,a1677a,a1680a,a1681a,a1684a,a1687a,a1688a,a1691a,a1694a,a1695a,a1698a,a1701a,a1702a,a1705a,a1708a,a1709a,a1712a,a1715a,a1716a,a1719a,a1722a,a1723a,a1726a,a1729a,a1730a,a1733a,a1736a,a1737a,a1740a,a1743a,a1744a,a1747a,a1750a,a1751a,a1754a,a1757a,a1758a,a1761a,a1764a,a1765a,a1768a,a1771a,a1772a,a1775a,a1778a,a1779a,a1782a,a1785a,a1786a,a1789a,a1792a,a1793a,a1796a,a1799a,a1800a,a1803a,a1806a,a1807a,a1810a,a1813a,a1814a,a1817a,a1820a,a1821a,a1824a,a1827a,a1828a,a1831a,a1834a,a1835a,a1838a,a1841a,a1842a,a1845a,a1848a,a1849a,a1852a,a1855a,a1856a,a1859a,a1862a,a1863a,a1866a,a1869a,a1870a,a1873a,a1876a,a1877a,a1880a,a1883a,a1884a,a1887a,a1890a,a1891a,a1894a,a1897a,a1898a,a1901a,a1904a,a1905a,a1908a,a1911a,a1912a,a1915a,a1918a,a1919a,a1922a,a1925a,a1926a,a1929a,a1932a,a1933a,a1936a,a1939a,a1940a,a1943a,a1946a,a1947a,a1950a,a1953a,a1954a,a1957a,a1960a,a1961a,a1964a,a1967a,a1968a,a1971a,a1974a,a1975a,a1978a,a1981a,a1982a,a1985a,a1988a,a1989a,a1992a,a1995a,a1996a,a1999a,a2002a,a2003a,a2006a,a2009a,a2010a,a2013a,a2016a,a2017a,a2020a,a2023a,a2024a,a2027a,a2030a,a2031a,a2034a,a2037a,a2038a,a2041a,a2044a,a2045a,a2048a,a2051a,a2052a,a2055a,a2058a,a2059a,a2062a,a2065a,a2066a,a2069a,a2072a,a2073a,a2076a,a2079a,a2080a,a2083a,a2086a,a2087a,a2090a,a2093a,a2094a,a2097a,a2100a,a2101a,a2104a,a2107a,a2108a,a2111a,a2114a,a2115a,a2118a,a2121a,a2122a,a2125a,a2128a,a2129a,a2132a,a2135a,a2136a,a2139a,a2142a,a2143a,a2146a,a2149a,a2150a,a2153a,a2156a,a2157a,a2160a,a2163a,a2164a,a2167a,a2170a,a2171a,a2174a,a2177a,a2178a,a2181a,a2184a,a2185a,a2188a,a2191a,a2192a,a2195a,a2198a,a2199a,a2202a,a2205a,a2206a,a2209a,a2212a,a2213a,a2216a,a2219a,a2220a,a2223a,a2226a,a2227a,a2230a,a2233a,a2234a,a2237a,a2240a,a2241a,a2244a,a2247a,a2248a,a2251a,a2254a,a2255a,a2258a,a2261a,a2262a,a2265a,a2268a,a2269a,a2272a,a2275a,a2276a,a2279a,a2282a,a2283a,a2286a,a2289a,a2290a,a2293a,a2296a,a2297a,a2300a,a2303a,a2304a,a2307a,a2310a,a2311a,a2314a,a2317a,a2318a,a2321a,a2324a,a2325a,a2328a,a2331a,a2332a,a2335a,a2338a,a2339a,a2342a,a2345a,a2346a,a2349a,a2352a,a2353a,a2356a,a2359a,a2360a,a2363a,a2366a,a2367a,a2370a,a2373a,a2374a,a2377a,a2380a,a2381a,a2384a,a2387a,a2388a,a2391a,a2394a,a2395a,a2398a,a2401a,a2402a,a2405a,a2408a,a2409a,a2412a,a2415a,a2416a,a2419a,a2422a,a2423a,a2426a,a2429a,a2430a,a2433a,a2436a,a2437a,a2440a,a2443a,a2444a,a2447a,a2450a,a2451a,a2454a,a2457a,a2458a,a2461a,a2464a,a2465a,a2468a,a2471a,a2472a,a2475a,a2478a,a2479a,a2482a,a2485a,a2486a,a2489a,a2492a,a2493a,a2496a,a2499a,a2500a,a2503a,a2506a,a2507a,a2510a,a2513a,a2514a,a2517a,a2520a,a2521a,a2524a,a2527a,a2528a,a2531a,a2534a,a2535a,a2538a,a2541a,a2542a,a2545a,a2548a,a2549a,a2552a,a2555a,a2556a,a2559a,a2562a,a2563a,a2566a,a2569a,a2570a,a2573a,a2576a,a2577a,a2580a,a2583a,a2584a,a2587a,a2590a,a2591a,a2594a,a2597a,a2598a,a2601a,a2604a,a2605a,a2608a,a2611a,a2612a,a2615a,a2618a,a2619a,a2622a,a2625a,a2626a,a2629a,a2632a,a2633a,a2636a,a2639a,a2640a,a2643a,a2646a,a2647a,a2650a,a2653a,a2654a,a2657a,a2660a,a2661a,a2664a,a2667a,a2668a,a2671a,a2674a,a2675a,a2678a,a2681a,a2682a,a2685a,a2688a,a2689a,a2692a,a2695a,a2696a,a2699a,a2702a,a2703a,a2706a,a2709a,a2710a,a2713a,a2716a,a2717a,a2720a,a2723a,a2724a,a2727a,a2730a,a2731a,a2734a,a2737a,a2738a,a2741a,a2744a,a2745a,a2748a,a2752a,a2753a,a2754a,a2757a,a2760a,a2761a,a2764a,a2768a,a2769a,a2770a,a2773a,a2776a,a2777a,a2780a,a2784a,a2785a,a2786a,a2789a,a2792a,a2793a,a2796a,a2800a,a2801a,a2802a,a2805a,a2808a,a2809a,a2812a,a2816a,a2817a,a2818a,a2821a,a2824a,a2825a,a2828a,a2832a,a2833a,a2834a,a2837a,a2840a,a2841a,a2844a,a2848a,a2849a,a2850a,a2853a,a2856a,a2857a,a2860a,a2864a,a2865a,a2866a,a2869a,a2872a,a2873a,a2876a,a2880a,a2881a,a2882a,a2885a,a2888a,a2889a,a2892a,a2896a,a2897a,a2898a,a2901a,a2904a,a2905a,a2908a,a2912a,a2913a,a2914a,a2917a,a2920a,a2921a,a2924a,a2928a,a2929a,a2930a,a2933a,a2936a,a2937a,a2940a,a2944a,a2945a,a2946a,a2949a,a2952a,a2953a,a2956a,a2960a,a2961a,a2962a,a2965a,a2968a,a2969a,a2972a,a2976a,a2977a,a2978a,a2981a,a2984a,a2985a,a2988a,a2992a,a2993a,a2994a,a2997a,a3000a,a3001a,a3004a,a3008a,a3009a,a3010a,a3013a,a3016a,a3017a,a3020a,a3024a,a3025a,a3026a,a3029a,a3032a,a3033a,a3036a,a3040a,a3041a,a3042a,a3045a,a3048a,a3049a,a3052a,a3056a,a3057a,a3058a,a3061a,a3064a,a3065a,a3068a,a3072a,a3073a,a3074a,a3077a,a3080a,a3081a,a3084a,a3088a,a3089a,a3090a,a3093a,a3096a,a3097a,a3100a,a3104a,a3105a,a3106a,a3109a,a3112a,a3113a,a3116a,a3120a,a3121a,a3122a,a3125a,a3128a,a3129a,a3132a,a3136a,a3137a,a3138a,a3141a,a3144a,a3145a,a3148a,a3152a,a3153a,a3154a,a3157a,a3160a,a3161a,a3164a,a3168a,a3169a,a3170a,a3173a,a3176a,a3177a,a3180a,a3184a,a3185a,a3186a,a3189a,a3192a,a3193a,a3196a,a3200a,a3201a,a3202a,a3205a,a3208a,a3209a,a3212a,a3216a,a3217a,a3218a,a3221a,a3224a,a3225a,a3228a,a3232a,a3233a,a3234a,a3237a,a3240a,a3241a,a3244a,a3248a,a3249a,a3250a,a3253a,a3257a,a3258a,a3259a,a3262a,a3266a,a3267a,a3268a,a3271a,a3275a,a3276a,a3277a,a3280a,a3284a,a3285a,a3286a,a3289a,a3293a,a3294a,a3295a,a3298a,a3302a,a3303a,a3304a,a3307a,a3311a,a3312a,a3313a,a3316a,a3320a,a3321a,a3322a,a3325a,a3329a,a3330a,a3331a,a3334a,a3338a,a3339a,a3340a,a3343a,a3347a,a3348a,a3349a,a3352a,a3356a,a3357a,a3358a,a3361a,a3365a,a3366a,a3367a,a3370a,a3374a,a3375a,a3376a,a3379a,a3383a,a3384a,a3385a,a3388a,a3392a,a3393a,a3394a,a3397a,a3401a,a3402a,a3403a,a3406a,a3410a,a3411a,a3412a,a3415a,a3419a,a3420a,a3421a,a3424a,a3428a,a3429a,a3430a,a3433a,a3437a,a3438a,a3439a,a3442a,a3446a,a3447a,a3448a,a3451a,a3455a,a3456a,a3457a,a3460a,a3464a,a3465a,a3466a,a3469a,a3473a,a3474a,a3475a,a3478a,a3482a,a3483a,a3484a,a3487a,a3491a,a3492a,a3493a,a3496a,a3500a,a3501a,a3502a,a3505a,a3509a,a3510a,a3511a,a3514a,a3518a,a3519a,a3520a,a3523a,a3527a,a3528a,a3529a,a3532a,a3536a,a3537a,a3538a,a3541a,a3545a,a3546a,a3547a,a3550a,a3554a,a3555a,a3556a,a3559a,a3563a,a3564a,a3565a,a3568a,a3572a,a3573a,a3574a,a3577a,a3581a,a3582a,a3583a,a3586a,a3590a,a3591a,a3592a,a3595a,a3599a,a3600a,a3601a,a3604a,a3608a,a3609a,a3610a,a3613a,a3617a,a3618a,a3619a,a3622a,a3626a,a3627a,a3628a,a3631a,a3635a,a3636a,a3637a,a3640a,a3644a,a3645a,a3646a,a3649a,a3653a,a3654a,a3655a,a3658a,a3662a,a3663a,a3664a,a3667a,a3671a,a3672a,a3673a,a3676a,a3680a,a3681a,a3682a,a3685a,a3689a,a3690a,a3691a,a3694a,a3698a,a3699a,a3700a,a3703a,a3707a,a3708a,a3709a,a3712a,a3716a,a3717a,a3718a,a3721a,a3725a,a3726a,a3727a,a3730a,a3734a,a3735a,a3736a,a3739a,a3743a,a3744a,a3745a,a3748a,a3752a,a3753a,a3754a,a3757a,a3761a,a3762a,a3763a,a3766a,a3770a,a3771a,a3772a,a3775a,a3779a,a3780a,a3781a,a3784a,a3788a,a3789a,a3790a,a3793a,a3797a,a3798a,a3799a,a3802a,a3806a,a3807a,a3808a,a3811a,a3815a,a3816a,a3817a,a3820a,a3824a,a3825a,a3826a,a3829a,a3833a,a3834a,a3835a,a3838a,a3842a,a3843a,a3844a,a3847a,a3851a,a3852a,a3853a,a3856a,a3860a,a3861a,a3862a,a3865a,a3869a,a3870a,a3871a,a3874a,a3878a,a3879a,a3880a,a3883a,a3887a,a3888a,a3889a,a3892a,a3896a,a3897a,a3898a,a3901a,a3905a,a3906a,a3907a,a3910a,a3914a,a3915a,a3916a,a3919a,a3923a,a3924a,a3925a,a3928a,a3932a,a3933a,a3934a,a3937a,a3941a,a3942a,a3943a,a3946a,a3950a,a3951a,a3952a,a3955a,a3959a,a3960a,a3961a,a3964a,a3968a,a3969a,a3970a,a3973a,a3977a,a3978a,a3979a,a3982a,a3986a,a3987a,a3988a,a3991a,a3995a,a3996a,a3997a,a4000a,a4004a,a4005a,a4006a,a4009a,a4013a,a4014a,a4015a,a4018a,a4022a,a4023a,a4024a,a4027a,a4031a,a4032a,a4033a,a4036a,a4040a,a4041a,a4042a,a4045a,a4049a,a4050a,a4051a,a4054a,a4058a,a4059a,a4060a,a4063a,a4067a,a4068a,a4069a,a4072a,a4076a,a4077a,a4078a,a4081a,a4085a,a4086a,a4087a,a4090a,a4094a,a4095a,a4096a,a4099a,a4103a,a4104a,a4105a,a4108a,a4112a,a4113a,a4114a,a4117a,a4121a,a4122a,a4123a,a4126a,a4130a,a4131a,a4132a,a4135a,a4139a,a4140a,a4141a,a4144a,a4148a,a4149a,a4150a,a4153a,a4157a,a4158a,a4159a,a4162a,a4166a,a4167a,a4168a,a4171a,a4175a,a4176a,a4177a,a4180a,a4184a,a4185a,a4186a,a4189a,a4193a,a4194a,a4195a,a4198a,a4202a,a4203a,a4204a,a4207a,a4211a,a4212a,a4213a,a4216a,a4220a,a4221a,a4222a,a4225a,a4229a,a4230a,a4231a,a4234a,a4238a,a4239a,a4240a,a4243a,a4247a,a4248a,a4249a,a4252a,a4256a,a4257a,a4258a,a4261a,a4265a,a4266a,a4267a,a4270a,a4274a,a4275a,a4276a,a4279a,a4283a,a4284a,a4285a,a4288a,a4292a,a4293a,a4294a,a4297a,a4301a,a4302a,a4303a,a4306a,a4310a,a4311a,a4312a,a4315a,a4319a,a4320a,a4321a,a4324a,a4328a,a4329a,a4330a,a4333a,a4337a,a4338a,a4339a,a4342a,a4346a,a4347a,a4348a,a4351a,a4355a,a4356a,a4357a,a4360a,a4364a,a4365a,a4366a,a4369a,a4373a,a4374a,a4375a,a4378a,a4382a,a4383a,a4384a,a4387a,a4391a,a4392a,a4393a,a4396a,a4400a,a4401a,a4402a,a4405a,a4409a,a4410a,a4411a,a4414a,a4418a,a4419a,a4420a,a4423a,a4427a,a4428a,a4429a,a4432a,a4436a,a4437a,a4438a,a4441a,a4445a,a4446a,a4447a,a4450a,a4454a,a4455a,a4456a,a4459a,a4463a,a4464a,a4465a,a4468a,a4472a,a4473a,a4474a,a4477a,a4481a,a4482a,a4483a,a4486a,a4490a,a4491a,a4492a,a4495a,a4499a,a4500a,a4501a,a4504a,a4508a,a4509a,a4510a,a4513a,a4517a,a4518a,a4519a,a4522a,a4526a,a4527a,a4528a,a4531a,a4535a,a4536a,a4537a,a4540a,a4544a,a4545a,a4546a,a4549a,a4553a,a4554a,a4555a,a4558a,a4562a,a4563a,a4564a,a4567a,a4571a,a4572a,a4573a,a4576a,a4580a,a4581a,a4582a,a4585a,a4589a,a4590a,a4591a,a4594a,a4598a,a4599a,a4600a,a4603a,a4607a,a4608a,a4609a,a4612a,a4616a,a4617a,a4618a,a4621a,a4625a,a4626a,a4627a,a4630a,a4634a,a4635a,a4636a,a4639a,a4643a,a4644a,a4645a,a4648a,a4652a,a4653a,a4654a,a4657a,a4661a,a4662a,a4663a,a4666a,a4670a,a4671a,a4672a,a4675a,a4679a,a4680a,a4681a,a4684a,a4688a,a4689a,a4690a,a4693a,a4697a,a4698a,a4699a,a4702a,a4706a,a4707a,a4708a,a4711a,a4715a,a4716a,a4717a,a4720a,a4724a,a4725a,a4726a,a4729a,a4733a,a4734a,a4735a,a4738a,a4742a,a4743a,a4744a,a4747a,a4751a,a4752a,a4753a,a4756a,a4760a,a4761a,a4762a,a4765a,a4769a,a4770a,a4771a,a4774a,a4778a,a4779a,a4780a,a4783a,a4787a,a4788a,a4789a,a4792a,a4796a,a4797a,a4798a,a4801a,a4805a,a4806a,a4807a,a4810a,a4814a,a4815a,a4816a,a4819a,a4823a,a4824a,a4825a,a4828a,a4832a,a4833a,a4834a,a4837a,a4841a,a4842a,a4843a,a4846a,a4850a,a4851a,a4852a,a4855a,a4859a,a4860a,a4861a,a4864a,a4868a,a4869a,a4870a,a4873a,a4877a,a4878a,a4879a,a4882a,a4886a,a4887a,a4888a,a4891a,a4895a,a4896a,a4897a,a4900a,a4904a,a4905a,a4906a,a4909a,a4913a,a4914a,a4915a,a4918a,a4922a,a4923a,a4924a,a4927a,a4931a,a4932a,a4933a,a4936a,a4940a,a4941a,a4942a,a4945a,a4949a,a4950a,a4951a,a4954a,a4958a,a4959a,a4960a,a4963a,a4967a,a4968a,a4969a,a4972a,a4976a,a4977a,a4978a,a4981a,a4985a,a4986a,a4987a,a4991a,a4992a,a4996a,a4997a,a4998a,a5001a,a5005a,a5006a,a5007a,a5011a,a5012a,a5016a,a5017a,a5018a,a5021a,a5025a,a5026a,a5027a,a5031a,a5032a,a5036a,a5037a,a5038a,a5041a,a5045a,a5046a,a5047a,a5051a,a5052a,a5056a,a5057a,a5058a,a5061a,a5065a,a5066a,a5067a,a5071a,a5072a,a5076a,a5077a,a5078a,a5081a,a5085a,a5086a,a5087a,a5091a,a5092a,a5096a,a5097a,a5098a,a5101a,a5105a,a5106a,a5107a,a5111a,a5112a,a5116a,a5117a,a5118a,a5121a,a5125a,a5126a,a5127a,a5131a,a5132a,a5136a,a5137a,a5138a,a5141a,a5145a,a5146a,a5147a,a5151a,a5152a,a5156a,a5157a,a5158a,a5161a,a5165a,a5166a,a5167a,a5171a,a5172a,a5176a,a5177a,a5178a,a5181a,a5185a,a5186a,a5187a,a5191a,a5192a,a5196a,a5197a,a5198a,a5201a,a5205a,a5206a,a5207a,a5211a,a5212a,a5216a,a5217a,a5218a,a5221a,a5225a,a5226a,a5227a,a5231a,a5232a,a5236a,a5237a,a5238a,a5241a,a5245a,a5246a,a5247a,a5251a,a5252a,a5256a,a5257a,a5258a,a5261a,a5265a,a5266a,a5267a,a5271a,a5272a,a5276a,a5277a,a5278a,a5281a,a5285a,a5286a,a5287a,a5291a,a5292a,a5296a,a5297a,a5298a,a5301a,a5305a,a5306a,a5307a,a5311a,a5312a,a5316a,a5317a,a5318a,a5321a,a5325a,a5326a,a5327a,a5331a,a5332a,a5336a,a5337a,a5338a,a5341a,a5345a,a5346a,a5347a,a5351a,a5352a,a5356a,a5357a,a5358a,a5361a,a5365a,a5366a,a5367a,a5371a,a5372a,a5376a,a5377a,a5378a,a5381a,a5385a,a5386a,a5387a,a5391a,a5392a,a5396a,a5397a,a5398a,a5401a,a5405a,a5406a,a5407a,a5411a,a5412a,a5416a,a5417a,a5418a,a5421a,a5425a,a5426a,a5427a,a5431a,a5432a,a5436a,a5437a,a5438a,a5441a,a5445a,a5446a,a5447a,a5451a,a5452a,a5456a,a5457a,a5458a,a5461a,a5465a,a5466a,a5467a,a5471a,a5472a,a5476a,a5477a,a5478a,a5481a,a5485a,a5486a,a5487a,a5491a,a5492a,a5496a,a5497a,a5498a,a5501a,a5505a,a5506a,a5507a,a5511a,a5512a,a5516a,a5517a,a5518a,a5521a,a5525a,a5526a,a5527a,a5531a,a5532a,a5536a,a5537a,a5538a,a5541a,a5545a,a5546a,a5547a,a5551a,a5552a,a5556a,a5557a,a5558a,a5561a,a5565a,a5566a,a5567a,a5571a,a5572a,a5576a,a5577a,a5578a,a5581a,a5585a,a5586a,a5587a,a5591a,a5592a,a5596a,a5597a,a5598a,a5601a,a5605a,a5606a,a5607a,a5611a,a5612a,a5616a,a5617a,a5618a,a5622a,a5623a,a5627a,a5628a,a5629a,a5633a,a5634a,a5638a,a5639a,a5640a,a5644a,a5645a,a5649a,a5650a,a5651a,a5655a,a5656a,a5660a,a5661a,a5662a,a5666a,a5667a,a5671a,a5672a,a5673a,a5677a,a5678a,a5682a,a5683a,a5684a,a5688a,a5689a,a5693a,a5694a,a5695a,a5699a,a5700a,a5704a,a5705a,a5706a,a5710a,a5711a,a5715a,a5716a,a5717a,a5721a,a5722a,a5726a,a5727a,a5728a,a5732a,a5733a,a5737a,a5738a,a5739a,a5743a,a5744a,a5748a,a5749a,a5750a,a5754a,a5755a,a5759a,a5760a,a5761a,a5765a,a5766a,a5770a,a5771a,a5772a,a5776a,a5777a,a5781a,a5782a,a5783a,a5787a,a5788a,a5792a,a5793a,a5794a,a5798a,a5799a,a5803a,a5804a,a5805a,a5809a,a5810a,a5814a,a5815a,a5816a,a5820a,a5821a,a5825a,a5826a,a5827a,a5831a,a5832a,a5836a,a5837a,a5838a,a5842a,a5843a,a5847a,a5848a,a5849a,a5853a,a5854a,a5858a,a5859a,a5860a,a5864a,a5865a,a5869a,a5870a,a5871a,a5875a,a5876a,a5880a,a5881a,a5882a,a5886a,a5887a,a5891a,a5892a,a5893a,a5897a,a5898a,a5902a,a5903a,a5904a,a5908a,a5909a,a5913a,a5914a,a5915a,a5919a,a5920a,a5924a,a5925a,a5926a,a5930a,a5931a,a5935a,a5936a,a5937a,a5941a,a5942a,a5946a,a5947a,a5948a,a5952a,a5953a,a5957a,a5958a,a5959a,a5963a,a5964a,a5968a,a5969a,a5970a,a5974a,a5975a,a5979a,a5980a,a5981a,a5985a,a5986a,a5990a,a5991a,a5992a,a5996a,a5997a,a6001a,a6002a,a6003a,a6007a,a6008a,a6012a,a6013a,a6014a,a6018a,a6019a,a6023a,a6024a,a6025a,a6029a,a6030a,a6034a,a6035a,a6036a,a6040a,a6041a,a6045a,a6046a,a6047a,a6051a,a6052a,a6056a,a6057a,a6058a,a6062a,a6063a,a6067a,a6068a,a6069a,a6073a,a6074a,a6078a,a6079a,a6080a,a6084a,a6085a,a6089a,a6090a,a6091a,a6095a,a6096a,a6100a,a6101a,a6102a,a6106a,a6107a,a6111a,a6112a,a6113a,a6117a,a6118a,a6122a,a6123a,a6124a,a6128a,a6129a,a6133a,a6134a,a6135a,a6139a,a6140a,a6144a,a6145a,a6146a,a6150a,a6151a,a6155a,a6156a,a6157a,a6161a,a6162a,a6166a,a6167a,a6168a,a6172a,a6173a,a6177a,a6178a,a6179a,a6183a,a6184a,a6188a,a6189a,a6190a,a6194a,a6195a,a6199a,a6200a,a6201a,a6205a,a6206a,a6210a,a6211a,a6212a,a6216a,a6217a,a6221a,a6222a,a6223a,a6227a,a6228a,a6232a,a6233a,a6234a,a6238a,a6239a,a6243a,a6244a,a6245a,a6249a,a6250a,a6254a,a6255a,a6256a,a6260a,a6261a,a6265a,a6266a,a6267a,a6271a,a6272a,a6276a,a6277a,a6278a,a6282a,a6283a,a6287a,a6288a,a6289a,a6293a,a6294a,a6298a,a6299a,a6300a,a6304a,a6305a,a6309a,a6310a,a6311a,a6315a,a6316a,a6320a,a6321a,a6322a,a6326a,a6327a,a6331a,a6332a,a6333a,a6337a,a6338a,a6342a,a6343a,a6344a,a6348a,a6349a,a6353a,a6354a,a6355a,a6359a,a6360a,a6364a,a6365a,a6366a,a6370a,a6371a,a6375a,a6376a,a6377a,a6381a,a6382a,a6386a,a6387a,a6388a,a6392a,a6393a,a6397a,a6398a,a6399a,a6403a,a6404a,a6408a,a6409a,a6410a,a6414a,a6415a,a6419a,a6420a,a6421a,a6425a,a6426a,a6430a,a6431a,a6432a,a6436a,a6437a,a6441a,a6442a,a6443a,a6447a,a6448a,a6452a,a6453a,a6454a,a6458a,a6459a,a6463a,a6464a,a6465a,a6469a,a6470a,a6474a,a6475a,a6476a,a6480a,a6481a,a6485a,a6486a,a6487a,a6491a,a6492a,a6496a,a6497a,a6498a,a6502a,a6503a,a6507a,a6508a,a6509a,a6513a,a6514a,a6518a,a6519a,a6520a,a6524a,a6525a,a6529a,a6530a,a6531a,a6535a,a6536a,a6540a,a6541a,a6542a,a6546a,a6547a,a6551a,a6552a,a6553a,a6557a,a6558a,a6562a,a6563a,a6564a,a6568a,a6569a,a6573a,a6574a,a6575a,a6579a,a6580a,a6584a,a6585a,a6586a,a6590a,a6591a,a6595a,a6596a,a6597a,a6601a,a6602a,a6606a,a6607a,a6608a,a6612a,a6613a,a6617a,a6618a,a6619a,a6623a,a6624a,a6628a,a6629a,a6630a,a6634a,a6635a,a6639a,a6640a,a6641a,a6645a,a6646a,a6650a,a6651a,a6652a,a6656a,a6657a,a6661a,a6662a,a6663a,a6667a,a6668a,a6672a,a6673a,a6674a: std_logic;
begin

A41 <=( a1042a ) or ( a695a );
 a1a <=( a6674a  and  a6663a );
 a2a <=( a6652a  and  a6641a );
 a3a <=( a6630a  and  a6619a );
 a4a <=( a6608a  and  a6597a );
 a5a <=( a6586a  and  a6575a );
 a6a <=( a6564a  and  a6553a );
 a7a <=( a6542a  and  a6531a );
 a8a <=( a6520a  and  a6509a );
 a9a <=( a6498a  and  a6487a );
 a10a <=( a6476a  and  a6465a );
 a11a <=( a6454a  and  a6443a );
 a12a <=( a6432a  and  a6421a );
 a13a <=( a6410a  and  a6399a );
 a14a <=( a6388a  and  a6377a );
 a15a <=( a6366a  and  a6355a );
 a16a <=( a6344a  and  a6333a );
 a17a <=( a6322a  and  a6311a );
 a18a <=( a6300a  and  a6289a );
 a19a <=( a6278a  and  a6267a );
 a20a <=( a6256a  and  a6245a );
 a21a <=( a6234a  and  a6223a );
 a22a <=( a6212a  and  a6201a );
 a23a <=( a6190a  and  a6179a );
 a24a <=( a6168a  and  a6157a );
 a25a <=( a6146a  and  a6135a );
 a26a <=( a6124a  and  a6113a );
 a27a <=( a6102a  and  a6091a );
 a28a <=( a6080a  and  a6069a );
 a29a <=( a6058a  and  a6047a );
 a30a <=( a6036a  and  a6025a );
 a31a <=( a6014a  and  a6003a );
 a32a <=( a5992a  and  a5981a );
 a33a <=( a5970a  and  a5959a );
 a34a <=( a5948a  and  a5937a );
 a35a <=( a5926a  and  a5915a );
 a36a <=( a5904a  and  a5893a );
 a37a <=( a5882a  and  a5871a );
 a38a <=( a5860a  and  a5849a );
 a39a <=( a5838a  and  a5827a );
 a40a <=( a5816a  and  a5805a );
 a41a <=( a5794a  and  a5783a );
 a42a <=( a5772a  and  a5761a );
 a43a <=( a5750a  and  a5739a );
 a44a <=( a5728a  and  a5717a );
 a45a <=( a5706a  and  a5695a );
 a46a <=( a5684a  and  a5673a );
 a47a <=( a5662a  and  a5651a );
 a48a <=( a5640a  and  a5629a );
 a49a <=( a5618a  and  a5607a );
 a50a <=( a5598a  and  a5587a );
 a51a <=( a5578a  and  a5567a );
 a52a <=( a5558a  and  a5547a );
 a53a <=( a5538a  and  a5527a );
 a54a <=( a5518a  and  a5507a );
 a55a <=( a5498a  and  a5487a );
 a56a <=( a5478a  and  a5467a );
 a57a <=( a5458a  and  a5447a );
 a58a <=( a5438a  and  a5427a );
 a59a <=( a5418a  and  a5407a );
 a60a <=( a5398a  and  a5387a );
 a61a <=( a5378a  and  a5367a );
 a62a <=( a5358a  and  a5347a );
 a63a <=( a5338a  and  a5327a );
 a64a <=( a5318a  and  a5307a );
 a65a <=( a5298a  and  a5287a );
 a66a <=( a5278a  and  a5267a );
 a67a <=( a5258a  and  a5247a );
 a68a <=( a5238a  and  a5227a );
 a69a <=( a5218a  and  a5207a );
 a70a <=( a5198a  and  a5187a );
 a71a <=( a5178a  and  a5167a );
 a72a <=( a5158a  and  a5147a );
 a73a <=( a5138a  and  a5127a );
 a74a <=( a5118a  and  a5107a );
 a75a <=( a5098a  and  a5087a );
 a76a <=( a5078a  and  a5067a );
 a77a <=( a5058a  and  a5047a );
 a78a <=( a5038a  and  a5027a );
 a79a <=( a5018a  and  a5007a );
 a80a <=( a4998a  and  a4987a );
 a81a <=( a4978a  and  a4969a );
 a82a <=( a4960a  and  a4951a );
 a83a <=( a4942a  and  a4933a );
 a84a <=( a4924a  and  a4915a );
 a85a <=( a4906a  and  a4897a );
 a86a <=( a4888a  and  a4879a );
 a87a <=( a4870a  and  a4861a );
 a88a <=( a4852a  and  a4843a );
 a89a <=( a4834a  and  a4825a );
 a90a <=( a4816a  and  a4807a );
 a91a <=( a4798a  and  a4789a );
 a92a <=( a4780a  and  a4771a );
 a93a <=( a4762a  and  a4753a );
 a94a <=( a4744a  and  a4735a );
 a95a <=( a4726a  and  a4717a );
 a96a <=( a4708a  and  a4699a );
 a97a <=( a4690a  and  a4681a );
 a98a <=( a4672a  and  a4663a );
 a99a <=( a4654a  and  a4645a );
 a100a <=( a4636a  and  a4627a );
 a101a <=( a4618a  and  a4609a );
 a102a <=( a4600a  and  a4591a );
 a103a <=( a4582a  and  a4573a );
 a104a <=( a4564a  and  a4555a );
 a105a <=( a4546a  and  a4537a );
 a106a <=( a4528a  and  a4519a );
 a107a <=( a4510a  and  a4501a );
 a108a <=( a4492a  and  a4483a );
 a109a <=( a4474a  and  a4465a );
 a110a <=( a4456a  and  a4447a );
 a111a <=( a4438a  and  a4429a );
 a112a <=( a4420a  and  a4411a );
 a113a <=( a4402a  and  a4393a );
 a114a <=( a4384a  and  a4375a );
 a115a <=( a4366a  and  a4357a );
 a116a <=( a4348a  and  a4339a );
 a117a <=( a4330a  and  a4321a );
 a118a <=( a4312a  and  a4303a );
 a119a <=( a4294a  and  a4285a );
 a120a <=( a4276a  and  a4267a );
 a121a <=( a4258a  and  a4249a );
 a122a <=( a4240a  and  a4231a );
 a123a <=( a4222a  and  a4213a );
 a124a <=( a4204a  and  a4195a );
 a125a <=( a4186a  and  a4177a );
 a126a <=( a4168a  and  a4159a );
 a127a <=( a4150a  and  a4141a );
 a128a <=( a4132a  and  a4123a );
 a129a <=( a4114a  and  a4105a );
 a130a <=( a4096a  and  a4087a );
 a131a <=( a4078a  and  a4069a );
 a132a <=( a4060a  and  a4051a );
 a133a <=( a4042a  and  a4033a );
 a134a <=( a4024a  and  a4015a );
 a135a <=( a4006a  and  a3997a );
 a136a <=( a3988a  and  a3979a );
 a137a <=( a3970a  and  a3961a );
 a138a <=( a3952a  and  a3943a );
 a139a <=( a3934a  and  a3925a );
 a140a <=( a3916a  and  a3907a );
 a141a <=( a3898a  and  a3889a );
 a142a <=( a3880a  and  a3871a );
 a143a <=( a3862a  and  a3853a );
 a144a <=( a3844a  and  a3835a );
 a145a <=( a3826a  and  a3817a );
 a146a <=( a3808a  and  a3799a );
 a147a <=( a3790a  and  a3781a );
 a148a <=( a3772a  and  a3763a );
 a149a <=( a3754a  and  a3745a );
 a150a <=( a3736a  and  a3727a );
 a151a <=( a3718a  and  a3709a );
 a152a <=( a3700a  and  a3691a );
 a153a <=( a3682a  and  a3673a );
 a154a <=( a3664a  and  a3655a );
 a155a <=( a3646a  and  a3637a );
 a156a <=( a3628a  and  a3619a );
 a157a <=( a3610a  and  a3601a );
 a158a <=( a3592a  and  a3583a );
 a159a <=( a3574a  and  a3565a );
 a160a <=( a3556a  and  a3547a );
 a161a <=( a3538a  and  a3529a );
 a162a <=( a3520a  and  a3511a );
 a163a <=( a3502a  and  a3493a );
 a164a <=( a3484a  and  a3475a );
 a165a <=( a3466a  and  a3457a );
 a166a <=( a3448a  and  a3439a );
 a167a <=( a3430a  and  a3421a );
 a168a <=( a3412a  and  a3403a );
 a169a <=( a3394a  and  a3385a );
 a170a <=( a3376a  and  a3367a );
 a171a <=( a3358a  and  a3349a );
 a172a <=( a3340a  and  a3331a );
 a173a <=( a3322a  and  a3313a );
 a174a <=( a3304a  and  a3295a );
 a175a <=( a3286a  and  a3277a );
 a176a <=( a3268a  and  a3259a );
 a177a <=( a3250a  and  a3241a );
 a178a <=( a3234a  and  a3225a );
 a179a <=( a3218a  and  a3209a );
 a180a <=( a3202a  and  a3193a );
 a181a <=( a3186a  and  a3177a );
 a182a <=( a3170a  and  a3161a );
 a183a <=( a3154a  and  a3145a );
 a184a <=( a3138a  and  a3129a );
 a185a <=( a3122a  and  a3113a );
 a186a <=( a3106a  and  a3097a );
 a187a <=( a3090a  and  a3081a );
 a188a <=( a3074a  and  a3065a );
 a189a <=( a3058a  and  a3049a );
 a190a <=( a3042a  and  a3033a );
 a191a <=( a3026a  and  a3017a );
 a192a <=( a3010a  and  a3001a );
 a193a <=( a2994a  and  a2985a );
 a194a <=( a2978a  and  a2969a );
 a195a <=( a2962a  and  a2953a );
 a196a <=( a2946a  and  a2937a );
 a197a <=( a2930a  and  a2921a );
 a198a <=( a2914a  and  a2905a );
 a199a <=( a2898a  and  a2889a );
 a200a <=( a2882a  and  a2873a );
 a201a <=( a2866a  and  a2857a );
 a202a <=( a2850a  and  a2841a );
 a203a <=( a2834a  and  a2825a );
 a204a <=( a2818a  and  a2809a );
 a205a <=( a2802a  and  a2793a );
 a206a <=( a2786a  and  a2777a );
 a207a <=( a2770a  and  a2761a );
 a208a <=( a2754a  and  a2745a );
 a209a <=( a2738a  and  a2731a );
 a210a <=( a2724a  and  a2717a );
 a211a <=( a2710a  and  a2703a );
 a212a <=( a2696a  and  a2689a );
 a213a <=( a2682a  and  a2675a );
 a214a <=( a2668a  and  a2661a );
 a215a <=( a2654a  and  a2647a );
 a216a <=( a2640a  and  a2633a );
 a217a <=( a2626a  and  a2619a );
 a218a <=( a2612a  and  a2605a );
 a219a <=( a2598a  and  a2591a );
 a220a <=( a2584a  and  a2577a );
 a221a <=( a2570a  and  a2563a );
 a222a <=( a2556a  and  a2549a );
 a223a <=( a2542a  and  a2535a );
 a224a <=( a2528a  and  a2521a );
 a225a <=( a2514a  and  a2507a );
 a226a <=( a2500a  and  a2493a );
 a227a <=( a2486a  and  a2479a );
 a228a <=( a2472a  and  a2465a );
 a229a <=( a2458a  and  a2451a );
 a230a <=( a2444a  and  a2437a );
 a231a <=( a2430a  and  a2423a );
 a232a <=( a2416a  and  a2409a );
 a233a <=( a2402a  and  a2395a );
 a234a <=( a2388a  and  a2381a );
 a235a <=( a2374a  and  a2367a );
 a236a <=( a2360a  and  a2353a );
 a237a <=( a2346a  and  a2339a );
 a238a <=( a2332a  and  a2325a );
 a239a <=( a2318a  and  a2311a );
 a240a <=( a2304a  and  a2297a );
 a241a <=( a2290a  and  a2283a );
 a242a <=( a2276a  and  a2269a );
 a243a <=( a2262a  and  a2255a );
 a244a <=( a2248a  and  a2241a );
 a245a <=( a2234a  and  a2227a );
 a246a <=( a2220a  and  a2213a );
 a247a <=( a2206a  and  a2199a );
 a248a <=( a2192a  and  a2185a );
 a249a <=( a2178a  and  a2171a );
 a250a <=( a2164a  and  a2157a );
 a251a <=( a2150a  and  a2143a );
 a252a <=( a2136a  and  a2129a );
 a253a <=( a2122a  and  a2115a );
 a254a <=( a2108a  and  a2101a );
 a255a <=( a2094a  and  a2087a );
 a256a <=( a2080a  and  a2073a );
 a257a <=( a2066a  and  a2059a );
 a258a <=( a2052a  and  a2045a );
 a259a <=( a2038a  and  a2031a );
 a260a <=( a2024a  and  a2017a );
 a261a <=( a2010a  and  a2003a );
 a262a <=( a1996a  and  a1989a );
 a263a <=( a1982a  and  a1975a );
 a264a <=( a1968a  and  a1961a );
 a265a <=( a1954a  and  a1947a );
 a266a <=( a1940a  and  a1933a );
 a267a <=( a1926a  and  a1919a );
 a268a <=( a1912a  and  a1905a );
 a269a <=( a1898a  and  a1891a );
 a270a <=( a1884a  and  a1877a );
 a271a <=( a1870a  and  a1863a );
 a272a <=( a1856a  and  a1849a );
 a273a <=( a1842a  and  a1835a );
 a274a <=( a1828a  and  a1821a );
 a275a <=( a1814a  and  a1807a );
 a276a <=( a1800a  and  a1793a );
 a277a <=( a1786a  and  a1779a );
 a278a <=( a1772a  and  a1765a );
 a279a <=( a1758a  and  a1751a );
 a280a <=( a1744a  and  a1737a );
 a281a <=( a1730a  and  a1723a );
 a282a <=( a1716a  and  a1709a );
 a283a <=( a1702a  and  a1695a );
 a284a <=( a1688a  and  a1681a );
 a285a <=( a1674a  and  a1667a );
 a286a <=( a1660a  and  a1653a );
 a287a <=( a1646a  and  a1639a );
 a288a <=( a1632a  and  a1625a );
 a289a <=( a1618a  and  a1611a );
 a290a <=( a1604a  and  a1597a );
 a291a <=( a1590a  and  a1583a );
 a292a <=( a1576a  and  a1569a );
 a293a <=( a1562a  and  a1555a );
 a294a <=( a1550a  and  a1543a );
 a295a <=( a1538a  and  a1531a );
 a296a <=( a1526a  and  a1519a );
 a297a <=( a1514a  and  a1507a );
 a298a <=( a1502a  and  a1495a );
 a299a <=( a1490a  and  a1483a );
 a300a <=( a1478a  and  a1471a );
 a301a <=( a1466a  and  a1461a );
 a302a <=( a1456a  and  a1451a );
 a303a <=( a1446a  and  a1441a );
 a304a <=( a1436a  and  a1431a );
 a305a <=( a1426a  and  a1421a );
 a306a <=( a1416a  and  a1411a );
 a307a <=( a1406a  and  a1401a );
 a308a <=( a1396a  and  a1391a );
 a309a <=( a1386a  and  a1381a );
 a310a <=( a1376a  and  a1371a );
 a311a <=( a1366a  and  a1361a );
 a312a <=( a1356a  and  a1351a );
 a313a <=( a1346a  and  a1341a );
 a314a <=( a1336a  and  a1331a );
 a315a <=( a1326a  and  a1321a );
 a316a <=( a1316a  and  a1311a );
 a317a <=( a1306a  and  a1301a );
 a318a <=( a1296a  and  a1291a );
 a319a <=( a1286a  and  a1281a );
 a320a <=( a1276a  and  a1271a );
 a321a <=( a1266a  and  a1261a );
 a322a <=( a1256a  and  a1251a );
 a323a <=( a1246a  and  a1241a );
 a324a <=( a1236a  and  a1231a );
 a325a <=( a1226a  and  a1221a );
 a326a <=( a1216a  and  a1211a );
 a327a <=( a1206a  and  a1201a );
 a328a <=( a1196a  and  a1191a );
 a329a <=( a1186a  and  a1181a );
 a330a <=( a1176a  and  a1171a );
 a331a <=( a1166a  and  a1161a );
 a332a <=( a1156a  and  a1151a );
 a333a <=( a1146a  and  a1141a );
 a334a <=( a1136a  and  a1131a );
 a335a <=( a1126a  and  a1121a );
 a336a <=( a1116a  and  a1111a );
 a337a <=( a1106a  and  a1103a );
 a338a <=( a1100a  and  a1097a );
 a339a <=( a1094a  and  a1091a );
 a340a <=( a1088a  and  a1085a );
 a341a <=( a1082a  and  a1079a );
 a342a <=( a1076a  and  a1073a );
 a343a <=( a1070a  and  a1067a );
 a344a <=( a1064a  and  a1061a );
 a345a <=( a1058a  and  a1055a );
 a346a <=( a1052a  and  a1049a );
 a347a <=( A267  and  A266 );
 a348a <=( A267  and  A265 );
 a351a <=( a347a ) or ( a348a );
 a355a <=( a344a ) or ( a345a );
 a356a <=( a346a ) or ( a355a );
 a357a <=( a356a ) or ( a351a );
 a360a <=( a342a ) or ( a343a );
 a364a <=( a339a ) or ( a340a );
 a365a <=( a341a ) or ( a364a );
 a366a <=( a365a ) or ( a360a );
 a367a <=( a366a ) or ( a357a );
 a370a <=( a337a ) or ( a338a );
 a374a <=( a334a ) or ( a335a );
 a375a <=( a336a ) or ( a374a );
 a376a <=( a375a ) or ( a370a );
 a380a <=( a331a ) or ( a332a );
 a381a <=( a333a ) or ( a380a );
 a385a <=( a328a ) or ( a329a );
 a386a <=( a330a ) or ( a385a );
 a387a <=( a386a ) or ( a381a );
 a388a <=( a387a ) or ( a376a );
 a389a <=( a388a ) or ( a367a );
 a392a <=( a326a ) or ( a327a );
 a396a <=( a323a ) or ( a324a );
 a397a <=( a325a ) or ( a396a );
 a398a <=( a397a ) or ( a392a );
 a402a <=( a320a ) or ( a321a );
 a403a <=( a322a ) or ( a402a );
 a407a <=( a317a ) or ( a318a );
 a408a <=( a319a ) or ( a407a );
 a409a <=( a408a ) or ( a403a );
 a410a <=( a409a ) or ( a398a );
 a413a <=( a315a ) or ( a316a );
 a417a <=( a312a ) or ( a313a );
 a418a <=( a314a ) or ( a417a );
 a419a <=( a418a ) or ( a413a );
 a423a <=( a309a ) or ( a310a );
 a424a <=( a311a ) or ( a423a );
 a428a <=( a306a ) or ( a307a );
 a429a <=( a308a ) or ( a428a );
 a430a <=( a429a ) or ( a424a );
 a431a <=( a430a ) or ( a419a );
 a432a <=( a431a ) or ( a410a );
 a433a <=( a432a ) or ( a389a );
 a436a <=( a304a ) or ( a305a );
 a440a <=( a301a ) or ( a302a );
 a441a <=( a303a ) or ( a440a );
 a442a <=( a441a ) or ( a436a );
 a446a <=( a298a ) or ( a299a );
 a447a <=( a300a ) or ( a446a );
 a451a <=( a295a ) or ( a296a );
 a452a <=( a297a ) or ( a451a );
 a453a <=( a452a ) or ( a447a );
 a454a <=( a453a ) or ( a442a );
 a457a <=( a293a ) or ( a294a );
 a461a <=( a290a ) or ( a291a );
 a462a <=( a292a ) or ( a461a );
 a463a <=( a462a ) or ( a457a );
 a467a <=( a287a ) or ( a288a );
 a468a <=( a289a ) or ( a467a );
 a472a <=( a284a ) or ( a285a );
 a473a <=( a286a ) or ( a472a );
 a474a <=( a473a ) or ( a468a );
 a475a <=( a474a ) or ( a463a );
 a476a <=( a475a ) or ( a454a );
 a479a <=( a282a ) or ( a283a );
 a483a <=( a279a ) or ( a280a );
 a484a <=( a281a ) or ( a483a );
 a485a <=( a484a ) or ( a479a );
 a489a <=( a276a ) or ( a277a );
 a490a <=( a278a ) or ( a489a );
 a494a <=( a273a ) or ( a274a );
 a495a <=( a275a ) or ( a494a );
 a496a <=( a495a ) or ( a490a );
 a497a <=( a496a ) or ( a485a );
 a500a <=( a271a ) or ( a272a );
 a504a <=( a268a ) or ( a269a );
 a505a <=( a270a ) or ( a504a );
 a506a <=( a505a ) or ( a500a );
 a510a <=( a265a ) or ( a266a );
 a511a <=( a267a ) or ( a510a );
 a515a <=( a262a ) or ( a263a );
 a516a <=( a264a ) or ( a515a );
 a517a <=( a516a ) or ( a511a );
 a518a <=( a517a ) or ( a506a );
 a519a <=( a518a ) or ( a497a );
 a520a <=( a519a ) or ( a476a );
 a521a <=( a520a ) or ( a433a );
 a524a <=( a260a ) or ( a261a );
 a528a <=( a257a ) or ( a258a );
 a529a <=( a259a ) or ( a528a );
 a530a <=( a529a ) or ( a524a );
 a533a <=( a255a ) or ( a256a );
 a537a <=( a252a ) or ( a253a );
 a538a <=( a254a ) or ( a537a );
 a539a <=( a538a ) or ( a533a );
 a540a <=( a539a ) or ( a530a );
 a543a <=( a250a ) or ( a251a );
 a547a <=( a247a ) or ( a248a );
 a548a <=( a249a ) or ( a547a );
 a549a <=( a548a ) or ( a543a );
 a553a <=( a244a ) or ( a245a );
 a554a <=( a246a ) or ( a553a );
 a558a <=( a241a ) or ( a242a );
 a559a <=( a243a ) or ( a558a );
 a560a <=( a559a ) or ( a554a );
 a561a <=( a560a ) or ( a549a );
 a562a <=( a561a ) or ( a540a );
 a565a <=( a239a ) or ( a240a );
 a569a <=( a236a ) or ( a237a );
 a570a <=( a238a ) or ( a569a );
 a571a <=( a570a ) or ( a565a );
 a575a <=( a233a ) or ( a234a );
 a576a <=( a235a ) or ( a575a );
 a580a <=( a230a ) or ( a231a );
 a581a <=( a232a ) or ( a580a );
 a582a <=( a581a ) or ( a576a );
 a583a <=( a582a ) or ( a571a );
 a586a <=( a228a ) or ( a229a );
 a590a <=( a225a ) or ( a226a );
 a591a <=( a227a ) or ( a590a );
 a592a <=( a591a ) or ( a586a );
 a596a <=( a222a ) or ( a223a );
 a597a <=( a224a ) or ( a596a );
 a601a <=( a219a ) or ( a220a );
 a602a <=( a221a ) or ( a601a );
 a603a <=( a602a ) or ( a597a );
 a604a <=( a603a ) or ( a592a );
 a605a <=( a604a ) or ( a583a );
 a606a <=( a605a ) or ( a562a );
 a609a <=( a217a ) or ( a218a );
 a613a <=( a214a ) or ( a215a );
 a614a <=( a216a ) or ( a613a );
 a615a <=( a614a ) or ( a609a );
 a619a <=( a211a ) or ( a212a );
 a620a <=( a213a ) or ( a619a );
 a624a <=( a208a ) or ( a209a );
 a625a <=( a210a ) or ( a624a );
 a626a <=( a625a ) or ( a620a );
 a627a <=( a626a ) or ( a615a );
 a630a <=( a206a ) or ( a207a );
 a634a <=( a203a ) or ( a204a );
 a635a <=( a205a ) or ( a634a );
 a636a <=( a635a ) or ( a630a );
 a640a <=( a200a ) or ( a201a );
 a641a <=( a202a ) or ( a640a );
 a645a <=( a197a ) or ( a198a );
 a646a <=( a199a ) or ( a645a );
 a647a <=( a646a ) or ( a641a );
 a648a <=( a647a ) or ( a636a );
 a649a <=( a648a ) or ( a627a );
 a652a <=( a195a ) or ( a196a );
 a656a <=( a192a ) or ( a193a );
 a657a <=( a194a ) or ( a656a );
 a658a <=( a657a ) or ( a652a );
 a662a <=( a189a ) or ( a190a );
 a663a <=( a191a ) or ( a662a );
 a667a <=( a186a ) or ( a187a );
 a668a <=( a188a ) or ( a667a );
 a669a <=( a668a ) or ( a663a );
 a670a <=( a669a ) or ( a658a );
 a673a <=( a184a ) or ( a185a );
 a677a <=( a181a ) or ( a182a );
 a678a <=( a183a ) or ( a677a );
 a679a <=( a678a ) or ( a673a );
 a683a <=( a178a ) or ( a179a );
 a684a <=( a180a ) or ( a683a );
 a688a <=( a175a ) or ( a176a );
 a689a <=( a177a ) or ( a688a );
 a690a <=( a689a ) or ( a684a );
 a691a <=( a690a ) or ( a679a );
 a692a <=( a691a ) or ( a670a );
 a693a <=( a692a ) or ( a649a );
 a694a <=( a693a ) or ( a606a );
 a695a <=( a694a ) or ( a521a );
 a698a <=( a173a ) or ( a174a );
 a702a <=( a170a ) or ( a171a );
 a703a <=( a172a ) or ( a702a );
 a704a <=( a703a ) or ( a698a );
 a707a <=( a168a ) or ( a169a );
 a711a <=( a165a ) or ( a166a );
 a712a <=( a167a ) or ( a711a );
 a713a <=( a712a ) or ( a707a );
 a714a <=( a713a ) or ( a704a );
 a717a <=( a163a ) or ( a164a );
 a721a <=( a160a ) or ( a161a );
 a722a <=( a162a ) or ( a721a );
 a723a <=( a722a ) or ( a717a );
 a727a <=( a157a ) or ( a158a );
 a728a <=( a159a ) or ( a727a );
 a732a <=( a154a ) or ( a155a );
 a733a <=( a156a ) or ( a732a );
 a734a <=( a733a ) or ( a728a );
 a735a <=( a734a ) or ( a723a );
 a736a <=( a735a ) or ( a714a );
 a739a <=( a152a ) or ( a153a );
 a743a <=( a149a ) or ( a150a );
 a744a <=( a151a ) or ( a743a );
 a745a <=( a744a ) or ( a739a );
 a749a <=( a146a ) or ( a147a );
 a750a <=( a148a ) or ( a749a );
 a754a <=( a143a ) or ( a144a );
 a755a <=( a145a ) or ( a754a );
 a756a <=( a755a ) or ( a750a );
 a757a <=( a756a ) or ( a745a );
 a760a <=( a141a ) or ( a142a );
 a764a <=( a138a ) or ( a139a );
 a765a <=( a140a ) or ( a764a );
 a766a <=( a765a ) or ( a760a );
 a770a <=( a135a ) or ( a136a );
 a771a <=( a137a ) or ( a770a );
 a775a <=( a132a ) or ( a133a );
 a776a <=( a134a ) or ( a775a );
 a777a <=( a776a ) or ( a771a );
 a778a <=( a777a ) or ( a766a );
 a779a <=( a778a ) or ( a757a );
 a780a <=( a779a ) or ( a736a );
 a783a <=( a130a ) or ( a131a );
 a787a <=( a127a ) or ( a128a );
 a788a <=( a129a ) or ( a787a );
 a789a <=( a788a ) or ( a783a );
 a793a <=( a124a ) or ( a125a );
 a794a <=( a126a ) or ( a793a );
 a798a <=( a121a ) or ( a122a );
 a799a <=( a123a ) or ( a798a );
 a800a <=( a799a ) or ( a794a );
 a801a <=( a800a ) or ( a789a );
 a804a <=( a119a ) or ( a120a );
 a808a <=( a116a ) or ( a117a );
 a809a <=( a118a ) or ( a808a );
 a810a <=( a809a ) or ( a804a );
 a814a <=( a113a ) or ( a114a );
 a815a <=( a115a ) or ( a814a );
 a819a <=( a110a ) or ( a111a );
 a820a <=( a112a ) or ( a819a );
 a821a <=( a820a ) or ( a815a );
 a822a <=( a821a ) or ( a810a );
 a823a <=( a822a ) or ( a801a );
 a826a <=( a108a ) or ( a109a );
 a830a <=( a105a ) or ( a106a );
 a831a <=( a107a ) or ( a830a );
 a832a <=( a831a ) or ( a826a );
 a836a <=( a102a ) or ( a103a );
 a837a <=( a104a ) or ( a836a );
 a841a <=( a99a ) or ( a100a );
 a842a <=( a101a ) or ( a841a );
 a843a <=( a842a ) or ( a837a );
 a844a <=( a843a ) or ( a832a );
 a847a <=( a97a ) or ( a98a );
 a851a <=( a94a ) or ( a95a );
 a852a <=( a96a ) or ( a851a );
 a853a <=( a852a ) or ( a847a );
 a857a <=( a91a ) or ( a92a );
 a858a <=( a93a ) or ( a857a );
 a862a <=( a88a ) or ( a89a );
 a863a <=( a90a ) or ( a862a );
 a864a <=( a863a ) or ( a858a );
 a865a <=( a864a ) or ( a853a );
 a866a <=( a865a ) or ( a844a );
 a867a <=( a866a ) or ( a823a );
 a868a <=( a867a ) or ( a780a );
 a871a <=( a86a ) or ( a87a );
 a875a <=( a83a ) or ( a84a );
 a876a <=( a85a ) or ( a875a );
 a877a <=( a876a ) or ( a871a );
 a880a <=( a81a ) or ( a82a );
 a884a <=( a78a ) or ( a79a );
 a885a <=( a80a ) or ( a884a );
 a886a <=( a885a ) or ( a880a );
 a887a <=( a886a ) or ( a877a );
 a890a <=( a76a ) or ( a77a );
 a894a <=( a73a ) or ( a74a );
 a895a <=( a75a ) or ( a894a );
 a896a <=( a895a ) or ( a890a );
 a900a <=( a70a ) or ( a71a );
 a901a <=( a72a ) or ( a900a );
 a905a <=( a67a ) or ( a68a );
 a906a <=( a69a ) or ( a905a );
 a907a <=( a906a ) or ( a901a );
 a908a <=( a907a ) or ( a896a );
 a909a <=( a908a ) or ( a887a );
 a912a <=( a65a ) or ( a66a );
 a916a <=( a62a ) or ( a63a );
 a917a <=( a64a ) or ( a916a );
 a918a <=( a917a ) or ( a912a );
 a922a <=( a59a ) or ( a60a );
 a923a <=( a61a ) or ( a922a );
 a927a <=( a56a ) or ( a57a );
 a928a <=( a58a ) or ( a927a );
 a929a <=( a928a ) or ( a923a );
 a930a <=( a929a ) or ( a918a );
 a933a <=( a54a ) or ( a55a );
 a937a <=( a51a ) or ( a52a );
 a938a <=( a53a ) or ( a937a );
 a939a <=( a938a ) or ( a933a );
 a943a <=( a48a ) or ( a49a );
 a944a <=( a50a ) or ( a943a );
 a948a <=( a45a ) or ( a46a );
 a949a <=( a47a ) or ( a948a );
 a950a <=( a949a ) or ( a944a );
 a951a <=( a950a ) or ( a939a );
 a952a <=( a951a ) or ( a930a );
 a953a <=( a952a ) or ( a909a );
 a956a <=( a43a ) or ( a44a );
 a960a <=( a40a ) or ( a41a );
 a961a <=( a42a ) or ( a960a );
 a962a <=( a961a ) or ( a956a );
 a966a <=( a37a ) or ( a38a );
 a967a <=( a39a ) or ( a966a );
 a971a <=( a34a ) or ( a35a );
 a972a <=( a36a ) or ( a971a );
 a973a <=( a972a ) or ( a967a );
 a974a <=( a973a ) or ( a962a );
 a977a <=( a32a ) or ( a33a );
 a981a <=( a29a ) or ( a30a );
 a982a <=( a31a ) or ( a981a );
 a983a <=( a982a ) or ( a977a );
 a987a <=( a26a ) or ( a27a );
 a988a <=( a28a ) or ( a987a );
 a992a <=( a23a ) or ( a24a );
 a993a <=( a25a ) or ( a992a );
 a994a <=( a993a ) or ( a988a );
 a995a <=( a994a ) or ( a983a );
 a996a <=( a995a ) or ( a974a );
 a999a <=( a21a ) or ( a22a );
 a1003a <=( a18a ) or ( a19a );
 a1004a <=( a20a ) or ( a1003a );
 a1005a <=( a1004a ) or ( a999a );
 a1009a <=( a15a ) or ( a16a );
 a1010a <=( a17a ) or ( a1009a );
 a1014a <=( a12a ) or ( a13a );
 a1015a <=( a14a ) or ( a1014a );
 a1016a <=( a1015a ) or ( a1010a );
 a1017a <=( a1016a ) or ( a1005a );
 a1020a <=( a10a ) or ( a11a );
 a1024a <=( a7a ) or ( a8a );
 a1025a <=( a9a ) or ( a1024a );
 a1026a <=( a1025a ) or ( a1020a );
 a1030a <=( a4a ) or ( a5a );
 a1031a <=( a6a ) or ( a1030a );
 a1035a <=( a1a ) or ( a2a );
 a1036a <=( a3a ) or ( a1035a );
 a1037a <=( a1036a ) or ( a1031a );
 a1038a <=( a1037a ) or ( a1026a );
 a1039a <=( a1038a ) or ( a1017a );
 a1040a <=( a1039a ) or ( a996a );
 a1041a <=( a1040a ) or ( a953a );
 a1042a <=( a1041a ) or ( a868a );
 a1049a <=( A266  and  A265 );
 a1052a <=( (not A269)  and  A268 );
 a1055a <=( A266  and  (not A265) );
 a1058a <=( A269  and  (not A268) );
 a1061a <=( (not A266)  and  A265 );
 a1064a <=( A269  and  (not A268) );
 a1067a <=( (not A266)  and  (not A265) );
 a1070a <=( (not A269)  and  A268 );
 a1073a <=( A201  and  A199 );
 a1076a <=( A234  and  A232 );
 a1079a <=( A201  and  A199 );
 a1082a <=( A234  and  A233 );
 a1085a <=( A201  and  A200 );
 a1088a <=( A234  and  A232 );
 a1091a <=( A201  and  A200 );
 a1094a <=( A234  and  A233 );
 a1097a <=( (not A166)  and  A167 );
 a1100a <=( A234  and  A232 );
 a1103a <=( (not A166)  and  A167 );
 a1106a <=( A234  and  A233 );
 a1110a <=( A232  and  A201 );
 a1111a <=( A199  and  a1110a );
 a1115a <=( (not A236)  and  A235 );
 a1116a <=( A233  and  a1115a );
 a1120a <=( (not A232)  and  A201 );
 a1121a <=( A199  and  a1120a );
 a1125a <=( A236  and  (not A235) );
 a1126a <=( A233  and  a1125a );
 a1130a <=( A232  and  A201 );
 a1131a <=( A199  and  a1130a );
 a1135a <=( A236  and  (not A235) );
 a1136a <=( (not A233)  and  a1135a );
 a1140a <=( (not A232)  and  A201 );
 a1141a <=( A199  and  a1140a );
 a1145a <=( (not A236)  and  A235 );
 a1146a <=( (not A233)  and  a1145a );
 a1150a <=( A232  and  A201 );
 a1151a <=( A200  and  a1150a );
 a1155a <=( (not A236)  and  A235 );
 a1156a <=( A233  and  a1155a );
 a1160a <=( (not A232)  and  A201 );
 a1161a <=( A200  and  a1160a );
 a1165a <=( A236  and  (not A235) );
 a1166a <=( A233  and  a1165a );
 a1170a <=( A232  and  A201 );
 a1171a <=( A200  and  a1170a );
 a1175a <=( A236  and  (not A235) );
 a1176a <=( (not A233)  and  a1175a );
 a1180a <=( (not A232)  and  A201 );
 a1181a <=( A200  and  a1180a );
 a1185a <=( (not A236)  and  A235 );
 a1186a <=( (not A233)  and  a1185a );
 a1190a <=( A202  and  A200 );
 a1191a <=( A199  and  a1190a );
 a1195a <=( A234  and  A232 );
 a1196a <=( (not A203)  and  a1195a );
 a1200a <=( A202  and  A200 );
 a1201a <=( A199  and  a1200a );
 a1205a <=( A234  and  A233 );
 a1206a <=( (not A203)  and  a1205a );
 a1210a <=( (not A202)  and  A200 );
 a1211a <=( (not A199)  and  a1210a );
 a1215a <=( A234  and  A232 );
 a1216a <=( A203  and  a1215a );
 a1220a <=( (not A202)  and  A200 );
 a1221a <=( (not A199)  and  a1220a );
 a1225a <=( A234  and  A233 );
 a1226a <=( A203  and  a1225a );
 a1230a <=( (not A202)  and  (not A200) );
 a1231a <=( A199  and  a1230a );
 a1235a <=( A234  and  A232 );
 a1236a <=( A203  and  a1235a );
 a1240a <=( (not A202)  and  (not A200) );
 a1241a <=( A199  and  a1240a );
 a1245a <=( A234  and  A233 );
 a1246a <=( A203  and  a1245a );
 a1250a <=( A202  and  (not A200) );
 a1251a <=( (not A199)  and  a1250a );
 a1255a <=( A234  and  A232 );
 a1256a <=( (not A203)  and  a1255a );
 a1260a <=( A202  and  (not A200) );
 a1261a <=( (not A199)  and  a1260a );
 a1265a <=( A234  and  A233 );
 a1266a <=( (not A203)  and  a1265a );
 a1270a <=( A199  and  A166 );
 a1271a <=( A167  and  a1270a );
 a1275a <=( A300  and  A299 );
 a1276a <=( A201  and  a1275a );
 a1280a <=( A199  and  A166 );
 a1281a <=( A167  and  a1280a );
 a1285a <=( A300  and  A298 );
 a1286a <=( A201  and  a1285a );
 a1290a <=( A200  and  A166 );
 a1291a <=( A167  and  a1290a );
 a1295a <=( A300  and  A299 );
 a1296a <=( A201  and  a1295a );
 a1300a <=( A200  and  A166 );
 a1301a <=( A167  and  a1300a );
 a1305a <=( A300  and  A298 );
 a1306a <=( A201  and  a1305a );
 a1310a <=( A232  and  (not A166) );
 a1311a <=( A167  and  a1310a );
 a1315a <=( (not A236)  and  A235 );
 a1316a <=( A233  and  a1315a );
 a1320a <=( (not A232)  and  (not A166) );
 a1321a <=( A167  and  a1320a );
 a1325a <=( A236  and  (not A235) );
 a1326a <=( A233  and  a1325a );
 a1330a <=( A232  and  (not A166) );
 a1331a <=( A167  and  a1330a );
 a1335a <=( A236  and  (not A235) );
 a1336a <=( (not A233)  and  a1335a );
 a1340a <=( (not A232)  and  (not A166) );
 a1341a <=( A167  and  a1340a );
 a1345a <=( (not A236)  and  A235 );
 a1346a <=( (not A233)  and  a1345a );
 a1350a <=( A199  and  (not A166) );
 a1351a <=( (not A167)  and  a1350a );
 a1355a <=( A300  and  A299 );
 a1356a <=( A201  and  a1355a );
 a1360a <=( A199  and  (not A166) );
 a1361a <=( (not A167)  and  a1360a );
 a1365a <=( A300  and  A298 );
 a1366a <=( A201  and  a1365a );
 a1370a <=( A200  and  (not A166) );
 a1371a <=( (not A167)  and  a1370a );
 a1375a <=( A300  and  A299 );
 a1376a <=( A201  and  a1375a );
 a1380a <=( A200  and  (not A166) );
 a1381a <=( (not A167)  and  a1380a );
 a1385a <=( A300  and  A298 );
 a1386a <=( A201  and  a1385a );
 a1390a <=( A199  and  (not A167) );
 a1391a <=( (not A168)  and  a1390a );
 a1395a <=( A300  and  A299 );
 a1396a <=( A201  and  a1395a );
 a1400a <=( A199  and  (not A167) );
 a1401a <=( (not A168)  and  a1400a );
 a1405a <=( A300  and  A298 );
 a1406a <=( A201  and  a1405a );
 a1410a <=( A200  and  (not A167) );
 a1411a <=( (not A168)  and  a1410a );
 a1415a <=( A300  and  A299 );
 a1416a <=( A201  and  a1415a );
 a1420a <=( A200  and  (not A167) );
 a1421a <=( (not A168)  and  a1420a );
 a1425a <=( A300  and  A298 );
 a1426a <=( A201  and  a1425a );
 a1430a <=( (not A167)  and  A168 );
 a1431a <=( A170  and  a1430a );
 a1435a <=( A234  and  A232 );
 a1436a <=( A166  and  a1435a );
 a1440a <=( (not A167)  and  A168 );
 a1441a <=( A170  and  a1440a );
 a1445a <=( A234  and  A233 );
 a1446a <=( A166  and  a1445a );
 a1450a <=( (not A167)  and  A168 );
 a1451a <=( A169  and  a1450a );
 a1455a <=( A234  and  A232 );
 a1456a <=( A166  and  a1455a );
 a1460a <=( (not A167)  and  A168 );
 a1461a <=( A169  and  a1460a );
 a1465a <=( A234  and  A233 );
 a1466a <=( A166  and  a1465a );
 a1470a <=( (not A199)  and  (not A166) );
 a1471a <=( A167  and  a1470a );
 a1474a <=( (not A202)  and  (not A200) );
 a1477a <=( A300  and  A299 );
 a1478a <=( a1477a  and  a1474a );
 a1482a <=( (not A199)  and  (not A166) );
 a1483a <=( A167  and  a1482a );
 a1486a <=( (not A202)  and  (not A200) );
 a1489a <=( A300  and  A298 );
 a1490a <=( a1489a  and  a1486a );
 a1494a <=( (not A199)  and  (not A166) );
 a1495a <=( A167  and  a1494a );
 a1498a <=( A203  and  (not A200) );
 a1501a <=( A300  and  A299 );
 a1502a <=( a1501a  and  a1498a );
 a1506a <=( (not A199)  and  (not A166) );
 a1507a <=( A167  and  a1506a );
 a1510a <=( A203  and  (not A200) );
 a1513a <=( A300  and  A298 );
 a1514a <=( a1513a  and  a1510a );
 a1518a <=( (not A167)  and  (not A169) );
 a1519a <=( (not A170)  and  a1518a );
 a1522a <=( A201  and  A199 );
 a1525a <=( A300  and  A299 );
 a1526a <=( a1525a  and  a1522a );
 a1530a <=( (not A167)  and  (not A169) );
 a1531a <=( (not A170)  and  a1530a );
 a1534a <=( A201  and  A199 );
 a1537a <=( A300  and  A298 );
 a1538a <=( a1537a  and  a1534a );
 a1542a <=( (not A167)  and  (not A169) );
 a1543a <=( (not A170)  and  a1542a );
 a1546a <=( A201  and  A200 );
 a1549a <=( A300  and  A299 );
 a1550a <=( a1549a  and  a1546a );
 a1554a <=( (not A167)  and  (not A169) );
 a1555a <=( (not A170)  and  a1554a );
 a1558a <=( A201  and  A200 );
 a1561a <=( A300  and  A298 );
 a1562a <=( a1561a  and  a1558a );
 a1565a <=( A200  and  A199 );
 a1568a <=( (not A203)  and  A202 );
 a1569a <=( a1568a  and  a1565a );
 a1572a <=( A233  and  A232 );
 a1575a <=( (not A236)  and  A235 );
 a1576a <=( a1575a  and  a1572a );
 a1579a <=( A200  and  A199 );
 a1582a <=( (not A203)  and  A202 );
 a1583a <=( a1582a  and  a1579a );
 a1586a <=( A233  and  (not A232) );
 a1589a <=( A236  and  (not A235) );
 a1590a <=( a1589a  and  a1586a );
 a1593a <=( A200  and  A199 );
 a1596a <=( (not A203)  and  A202 );
 a1597a <=( a1596a  and  a1593a );
 a1600a <=( (not A233)  and  A232 );
 a1603a <=( A236  and  (not A235) );
 a1604a <=( a1603a  and  a1600a );
 a1607a <=( A200  and  A199 );
 a1610a <=( (not A203)  and  A202 );
 a1611a <=( a1610a  and  a1607a );
 a1614a <=( (not A233)  and  (not A232) );
 a1617a <=( (not A236)  and  A235 );
 a1618a <=( a1617a  and  a1614a );
 a1621a <=( A200  and  (not A199) );
 a1624a <=( A203  and  (not A202) );
 a1625a <=( a1624a  and  a1621a );
 a1628a <=( A233  and  A232 );
 a1631a <=( (not A236)  and  A235 );
 a1632a <=( a1631a  and  a1628a );
 a1635a <=( A200  and  (not A199) );
 a1638a <=( A203  and  (not A202) );
 a1639a <=( a1638a  and  a1635a );
 a1642a <=( A233  and  (not A232) );
 a1645a <=( A236  and  (not A235) );
 a1646a <=( a1645a  and  a1642a );
 a1649a <=( A200  and  (not A199) );
 a1652a <=( A203  and  (not A202) );
 a1653a <=( a1652a  and  a1649a );
 a1656a <=( (not A233)  and  A232 );
 a1659a <=( A236  and  (not A235) );
 a1660a <=( a1659a  and  a1656a );
 a1663a <=( A200  and  (not A199) );
 a1666a <=( A203  and  (not A202) );
 a1667a <=( a1666a  and  a1663a );
 a1670a <=( (not A233)  and  (not A232) );
 a1673a <=( (not A236)  and  A235 );
 a1674a <=( a1673a  and  a1670a );
 a1677a <=( (not A200)  and  A199 );
 a1680a <=( A203  and  (not A202) );
 a1681a <=( a1680a  and  a1677a );
 a1684a <=( A233  and  A232 );
 a1687a <=( (not A236)  and  A235 );
 a1688a <=( a1687a  and  a1684a );
 a1691a <=( (not A200)  and  A199 );
 a1694a <=( A203  and  (not A202) );
 a1695a <=( a1694a  and  a1691a );
 a1698a <=( A233  and  (not A232) );
 a1701a <=( A236  and  (not A235) );
 a1702a <=( a1701a  and  a1698a );
 a1705a <=( (not A200)  and  A199 );
 a1708a <=( A203  and  (not A202) );
 a1709a <=( a1708a  and  a1705a );
 a1712a <=( (not A233)  and  A232 );
 a1715a <=( A236  and  (not A235) );
 a1716a <=( a1715a  and  a1712a );
 a1719a <=( (not A200)  and  A199 );
 a1722a <=( A203  and  (not A202) );
 a1723a <=( a1722a  and  a1719a );
 a1726a <=( (not A233)  and  (not A232) );
 a1729a <=( (not A236)  and  A235 );
 a1730a <=( a1729a  and  a1726a );
 a1733a <=( (not A200)  and  (not A199) );
 a1736a <=( (not A203)  and  A202 );
 a1737a <=( a1736a  and  a1733a );
 a1740a <=( A233  and  A232 );
 a1743a <=( (not A236)  and  A235 );
 a1744a <=( a1743a  and  a1740a );
 a1747a <=( (not A200)  and  (not A199) );
 a1750a <=( (not A203)  and  A202 );
 a1751a <=( a1750a  and  a1747a );
 a1754a <=( A233  and  (not A232) );
 a1757a <=( A236  and  (not A235) );
 a1758a <=( a1757a  and  a1754a );
 a1761a <=( (not A200)  and  (not A199) );
 a1764a <=( (not A203)  and  A202 );
 a1765a <=( a1764a  and  a1761a );
 a1768a <=( (not A233)  and  A232 );
 a1771a <=( A236  and  (not A235) );
 a1772a <=( a1771a  and  a1768a );
 a1775a <=( (not A200)  and  (not A199) );
 a1778a <=( (not A203)  and  A202 );
 a1779a <=( a1778a  and  a1775a );
 a1782a <=( (not A233)  and  (not A232) );
 a1785a <=( (not A236)  and  A235 );
 a1786a <=( a1785a  and  a1782a );
 a1789a <=( A166  and  A167 );
 a1792a <=( A201  and  A199 );
 a1793a <=( a1792a  and  a1789a );
 a1796a <=( A299  and  A298 );
 a1799a <=( (not A302)  and  A301 );
 a1800a <=( a1799a  and  a1796a );
 a1803a <=( A166  and  A167 );
 a1806a <=( A201  and  A199 );
 a1807a <=( a1806a  and  a1803a );
 a1810a <=( (not A299)  and  A298 );
 a1813a <=( A302  and  (not A301) );
 a1814a <=( a1813a  and  a1810a );
 a1817a <=( A166  and  A167 );
 a1820a <=( A201  and  A199 );
 a1821a <=( a1820a  and  a1817a );
 a1824a <=( A299  and  (not A298) );
 a1827a <=( A302  and  (not A301) );
 a1828a <=( a1827a  and  a1824a );
 a1831a <=( A166  and  A167 );
 a1834a <=( A201  and  A199 );
 a1835a <=( a1834a  and  a1831a );
 a1838a <=( (not A299)  and  (not A298) );
 a1841a <=( (not A302)  and  A301 );
 a1842a <=( a1841a  and  a1838a );
 a1845a <=( A166  and  A167 );
 a1848a <=( A201  and  A200 );
 a1849a <=( a1848a  and  a1845a );
 a1852a <=( A299  and  A298 );
 a1855a <=( (not A302)  and  A301 );
 a1856a <=( a1855a  and  a1852a );
 a1859a <=( A166  and  A167 );
 a1862a <=( A201  and  A200 );
 a1863a <=( a1862a  and  a1859a );
 a1866a <=( (not A299)  and  A298 );
 a1869a <=( A302  and  (not A301) );
 a1870a <=( a1869a  and  a1866a );
 a1873a <=( A166  and  A167 );
 a1876a <=( A201  and  A200 );
 a1877a <=( a1876a  and  a1873a );
 a1880a <=( A299  and  (not A298) );
 a1883a <=( A302  and  (not A301) );
 a1884a <=( a1883a  and  a1880a );
 a1887a <=( A166  and  A167 );
 a1890a <=( A201  and  A200 );
 a1891a <=( a1890a  and  a1887a );
 a1894a <=( (not A299)  and  (not A298) );
 a1897a <=( (not A302)  and  A301 );
 a1898a <=( a1897a  and  a1894a );
 a1901a <=( A166  and  A167 );
 a1904a <=( A200  and  A199 );
 a1905a <=( a1904a  and  a1901a );
 a1908a <=( (not A203)  and  A202 );
 a1911a <=( A300  and  A299 );
 a1912a <=( a1911a  and  a1908a );
 a1915a <=( A166  and  A167 );
 a1918a <=( A200  and  A199 );
 a1919a <=( a1918a  and  a1915a );
 a1922a <=( (not A203)  and  A202 );
 a1925a <=( A300  and  A298 );
 a1926a <=( a1925a  and  a1922a );
 a1929a <=( A166  and  A167 );
 a1932a <=( A200  and  (not A199) );
 a1933a <=( a1932a  and  a1929a );
 a1936a <=( A203  and  (not A202) );
 a1939a <=( A300  and  A299 );
 a1940a <=( a1939a  and  a1936a );
 a1943a <=( A166  and  A167 );
 a1946a <=( A200  and  (not A199) );
 a1947a <=( a1946a  and  a1943a );
 a1950a <=( A203  and  (not A202) );
 a1953a <=( A300  and  A298 );
 a1954a <=( a1953a  and  a1950a );
 a1957a <=( A166  and  A167 );
 a1960a <=( (not A200)  and  A199 );
 a1961a <=( a1960a  and  a1957a );
 a1964a <=( A203  and  (not A202) );
 a1967a <=( A300  and  A299 );
 a1968a <=( a1967a  and  a1964a );
 a1971a <=( A166  and  A167 );
 a1974a <=( (not A200)  and  A199 );
 a1975a <=( a1974a  and  a1971a );
 a1978a <=( A203  and  (not A202) );
 a1981a <=( A300  and  A298 );
 a1982a <=( a1981a  and  a1978a );
 a1985a <=( A166  and  A167 );
 a1988a <=( (not A200)  and  (not A199) );
 a1989a <=( a1988a  and  a1985a );
 a1992a <=( (not A203)  and  A202 );
 a1995a <=( A300  and  A299 );
 a1996a <=( a1995a  and  a1992a );
 a1999a <=( A166  and  A167 );
 a2002a <=( (not A200)  and  (not A199) );
 a2003a <=( a2002a  and  a1999a );
 a2006a <=( (not A203)  and  A202 );
 a2009a <=( A300  and  A298 );
 a2010a <=( a2009a  and  a2006a );
 a2013a <=( (not A166)  and  A167 );
 a2016a <=( A200  and  A199 );
 a2017a <=( a2016a  and  a2013a );
 a2020a <=( (not A202)  and  (not A201) );
 a2023a <=( A300  and  A299 );
 a2024a <=( a2023a  and  a2020a );
 a2027a <=( (not A166)  and  A167 );
 a2030a <=( A200  and  A199 );
 a2031a <=( a2030a  and  a2027a );
 a2034a <=( (not A202)  and  (not A201) );
 a2037a <=( A300  and  A298 );
 a2038a <=( a2037a  and  a2034a );
 a2041a <=( (not A166)  and  A167 );
 a2044a <=( A200  and  A199 );
 a2045a <=( a2044a  and  a2041a );
 a2048a <=( A203  and  (not A201) );
 a2051a <=( A300  and  A299 );
 a2052a <=( a2051a  and  a2048a );
 a2055a <=( (not A166)  and  A167 );
 a2058a <=( A200  and  A199 );
 a2059a <=( a2058a  and  a2055a );
 a2062a <=( A203  and  (not A201) );
 a2065a <=( A300  and  A298 );
 a2066a <=( a2065a  and  a2062a );
 a2069a <=( (not A166)  and  A167 );
 a2072a <=( A200  and  (not A199) );
 a2073a <=( a2072a  and  a2069a );
 a2076a <=( A202  and  (not A201) );
 a2079a <=( A300  and  A299 );
 a2080a <=( a2079a  and  a2076a );
 a2083a <=( (not A166)  and  A167 );
 a2086a <=( A200  and  (not A199) );
 a2087a <=( a2086a  and  a2083a );
 a2090a <=( A202  and  (not A201) );
 a2093a <=( A300  and  A298 );
 a2094a <=( a2093a  and  a2090a );
 a2097a <=( (not A166)  and  A167 );
 a2100a <=( A200  and  (not A199) );
 a2101a <=( a2100a  and  a2097a );
 a2104a <=( (not A203)  and  (not A201) );
 a2107a <=( A300  and  A299 );
 a2108a <=( a2107a  and  a2104a );
 a2111a <=( (not A166)  and  A167 );
 a2114a <=( A200  and  (not A199) );
 a2115a <=( a2114a  and  a2111a );
 a2118a <=( (not A203)  and  (not A201) );
 a2121a <=( A300  and  A298 );
 a2122a <=( a2121a  and  a2118a );
 a2125a <=( (not A166)  and  A167 );
 a2128a <=( (not A200)  and  A199 );
 a2129a <=( a2128a  and  a2125a );
 a2132a <=( A202  and  (not A201) );
 a2135a <=( A300  and  A299 );
 a2136a <=( a2135a  and  a2132a );
 a2139a <=( (not A166)  and  A167 );
 a2142a <=( (not A200)  and  A199 );
 a2143a <=( a2142a  and  a2139a );
 a2146a <=( A202  and  (not A201) );
 a2149a <=( A300  and  A298 );
 a2150a <=( a2149a  and  a2146a );
 a2153a <=( (not A166)  and  A167 );
 a2156a <=( (not A200)  and  A199 );
 a2157a <=( a2156a  and  a2153a );
 a2160a <=( (not A203)  and  (not A201) );
 a2163a <=( A300  and  A299 );
 a2164a <=( a2163a  and  a2160a );
 a2167a <=( (not A166)  and  A167 );
 a2170a <=( (not A200)  and  A199 );
 a2171a <=( a2170a  and  a2167a );
 a2174a <=( (not A203)  and  (not A201) );
 a2177a <=( A300  and  A298 );
 a2178a <=( a2177a  and  a2174a );
 a2181a <=( (not A166)  and  (not A167) );
 a2184a <=( A201  and  A199 );
 a2185a <=( a2184a  and  a2181a );
 a2188a <=( A299  and  A298 );
 a2191a <=( (not A302)  and  A301 );
 a2192a <=( a2191a  and  a2188a );
 a2195a <=( (not A166)  and  (not A167) );
 a2198a <=( A201  and  A199 );
 a2199a <=( a2198a  and  a2195a );
 a2202a <=( (not A299)  and  A298 );
 a2205a <=( A302  and  (not A301) );
 a2206a <=( a2205a  and  a2202a );
 a2209a <=( (not A166)  and  (not A167) );
 a2212a <=( A201  and  A199 );
 a2213a <=( a2212a  and  a2209a );
 a2216a <=( A299  and  (not A298) );
 a2219a <=( A302  and  (not A301) );
 a2220a <=( a2219a  and  a2216a );
 a2223a <=( (not A166)  and  (not A167) );
 a2226a <=( A201  and  A199 );
 a2227a <=( a2226a  and  a2223a );
 a2230a <=( (not A299)  and  (not A298) );
 a2233a <=( (not A302)  and  A301 );
 a2234a <=( a2233a  and  a2230a );
 a2237a <=( (not A166)  and  (not A167) );
 a2240a <=( A201  and  A200 );
 a2241a <=( a2240a  and  a2237a );
 a2244a <=( A299  and  A298 );
 a2247a <=( (not A302)  and  A301 );
 a2248a <=( a2247a  and  a2244a );
 a2251a <=( (not A166)  and  (not A167) );
 a2254a <=( A201  and  A200 );
 a2255a <=( a2254a  and  a2251a );
 a2258a <=( (not A299)  and  A298 );
 a2261a <=( A302  and  (not A301) );
 a2262a <=( a2261a  and  a2258a );
 a2265a <=( (not A166)  and  (not A167) );
 a2268a <=( A201  and  A200 );
 a2269a <=( a2268a  and  a2265a );
 a2272a <=( A299  and  (not A298) );
 a2275a <=( A302  and  (not A301) );
 a2276a <=( a2275a  and  a2272a );
 a2279a <=( (not A166)  and  (not A167) );
 a2282a <=( A201  and  A200 );
 a2283a <=( a2282a  and  a2279a );
 a2286a <=( (not A299)  and  (not A298) );
 a2289a <=( (not A302)  and  A301 );
 a2290a <=( a2289a  and  a2286a );
 a2293a <=( (not A166)  and  (not A167) );
 a2296a <=( A200  and  A199 );
 a2297a <=( a2296a  and  a2293a );
 a2300a <=( (not A203)  and  A202 );
 a2303a <=( A300  and  A299 );
 a2304a <=( a2303a  and  a2300a );
 a2307a <=( (not A166)  and  (not A167) );
 a2310a <=( A200  and  A199 );
 a2311a <=( a2310a  and  a2307a );
 a2314a <=( (not A203)  and  A202 );
 a2317a <=( A300  and  A298 );
 a2318a <=( a2317a  and  a2314a );
 a2321a <=( (not A166)  and  (not A167) );
 a2324a <=( A200  and  (not A199) );
 a2325a <=( a2324a  and  a2321a );
 a2328a <=( A203  and  (not A202) );
 a2331a <=( A300  and  A299 );
 a2332a <=( a2331a  and  a2328a );
 a2335a <=( (not A166)  and  (not A167) );
 a2338a <=( A200  and  (not A199) );
 a2339a <=( a2338a  and  a2335a );
 a2342a <=( A203  and  (not A202) );
 a2345a <=( A300  and  A298 );
 a2346a <=( a2345a  and  a2342a );
 a2349a <=( (not A166)  and  (not A167) );
 a2352a <=( (not A200)  and  A199 );
 a2353a <=( a2352a  and  a2349a );
 a2356a <=( A203  and  (not A202) );
 a2359a <=( A300  and  A299 );
 a2360a <=( a2359a  and  a2356a );
 a2363a <=( (not A166)  and  (not A167) );
 a2366a <=( (not A200)  and  A199 );
 a2367a <=( a2366a  and  a2363a );
 a2370a <=( A203  and  (not A202) );
 a2373a <=( A300  and  A298 );
 a2374a <=( a2373a  and  a2370a );
 a2377a <=( (not A166)  and  (not A167) );
 a2380a <=( (not A200)  and  (not A199) );
 a2381a <=( a2380a  and  a2377a );
 a2384a <=( (not A203)  and  A202 );
 a2387a <=( A300  and  A299 );
 a2388a <=( a2387a  and  a2384a );
 a2391a <=( (not A166)  and  (not A167) );
 a2394a <=( (not A200)  and  (not A199) );
 a2395a <=( a2394a  and  a2391a );
 a2398a <=( (not A203)  and  A202 );
 a2401a <=( A300  and  A298 );
 a2402a <=( a2401a  and  a2398a );
 a2405a <=( (not A167)  and  (not A168) );
 a2408a <=( A201  and  A199 );
 a2409a <=( a2408a  and  a2405a );
 a2412a <=( A299  and  A298 );
 a2415a <=( (not A302)  and  A301 );
 a2416a <=( a2415a  and  a2412a );
 a2419a <=( (not A167)  and  (not A168) );
 a2422a <=( A201  and  A199 );
 a2423a <=( a2422a  and  a2419a );
 a2426a <=( (not A299)  and  A298 );
 a2429a <=( A302  and  (not A301) );
 a2430a <=( a2429a  and  a2426a );
 a2433a <=( (not A167)  and  (not A168) );
 a2436a <=( A201  and  A199 );
 a2437a <=( a2436a  and  a2433a );
 a2440a <=( A299  and  (not A298) );
 a2443a <=( A302  and  (not A301) );
 a2444a <=( a2443a  and  a2440a );
 a2447a <=( (not A167)  and  (not A168) );
 a2450a <=( A201  and  A199 );
 a2451a <=( a2450a  and  a2447a );
 a2454a <=( (not A299)  and  (not A298) );
 a2457a <=( (not A302)  and  A301 );
 a2458a <=( a2457a  and  a2454a );
 a2461a <=( (not A167)  and  (not A168) );
 a2464a <=( A201  and  A200 );
 a2465a <=( a2464a  and  a2461a );
 a2468a <=( A299  and  A298 );
 a2471a <=( (not A302)  and  A301 );
 a2472a <=( a2471a  and  a2468a );
 a2475a <=( (not A167)  and  (not A168) );
 a2478a <=( A201  and  A200 );
 a2479a <=( a2478a  and  a2475a );
 a2482a <=( (not A299)  and  A298 );
 a2485a <=( A302  and  (not A301) );
 a2486a <=( a2485a  and  a2482a );
 a2489a <=( (not A167)  and  (not A168) );
 a2492a <=( A201  and  A200 );
 a2493a <=( a2492a  and  a2489a );
 a2496a <=( A299  and  (not A298) );
 a2499a <=( A302  and  (not A301) );
 a2500a <=( a2499a  and  a2496a );
 a2503a <=( (not A167)  and  (not A168) );
 a2506a <=( A201  and  A200 );
 a2507a <=( a2506a  and  a2503a );
 a2510a <=( (not A299)  and  (not A298) );
 a2513a <=( (not A302)  and  A301 );
 a2514a <=( a2513a  and  a2510a );
 a2517a <=( (not A167)  and  (not A168) );
 a2520a <=( A200  and  A199 );
 a2521a <=( a2520a  and  a2517a );
 a2524a <=( (not A203)  and  A202 );
 a2527a <=( A300  and  A299 );
 a2528a <=( a2527a  and  a2524a );
 a2531a <=( (not A167)  and  (not A168) );
 a2534a <=( A200  and  A199 );
 a2535a <=( a2534a  and  a2531a );
 a2538a <=( (not A203)  and  A202 );
 a2541a <=( A300  and  A298 );
 a2542a <=( a2541a  and  a2538a );
 a2545a <=( (not A167)  and  (not A168) );
 a2548a <=( A200  and  (not A199) );
 a2549a <=( a2548a  and  a2545a );
 a2552a <=( A203  and  (not A202) );
 a2555a <=( A300  and  A299 );
 a2556a <=( a2555a  and  a2552a );
 a2559a <=( (not A167)  and  (not A168) );
 a2562a <=( A200  and  (not A199) );
 a2563a <=( a2562a  and  a2559a );
 a2566a <=( A203  and  (not A202) );
 a2569a <=( A300  and  A298 );
 a2570a <=( a2569a  and  a2566a );
 a2573a <=( (not A167)  and  (not A168) );
 a2576a <=( (not A200)  and  A199 );
 a2577a <=( a2576a  and  a2573a );
 a2580a <=( A203  and  (not A202) );
 a2583a <=( A300  and  A299 );
 a2584a <=( a2583a  and  a2580a );
 a2587a <=( (not A167)  and  (not A168) );
 a2590a <=( (not A200)  and  A199 );
 a2591a <=( a2590a  and  a2587a );
 a2594a <=( A203  and  (not A202) );
 a2597a <=( A300  and  A298 );
 a2598a <=( a2597a  and  a2594a );
 a2601a <=( (not A167)  and  (not A168) );
 a2604a <=( (not A200)  and  (not A199) );
 a2605a <=( a2604a  and  a2601a );
 a2608a <=( (not A203)  and  A202 );
 a2611a <=( A300  and  A299 );
 a2612a <=( a2611a  and  a2608a );
 a2615a <=( (not A167)  and  (not A168) );
 a2618a <=( (not A200)  and  (not A199) );
 a2619a <=( a2618a  and  a2615a );
 a2622a <=( (not A203)  and  A202 );
 a2625a <=( A300  and  A298 );
 a2626a <=( a2625a  and  a2622a );
 a2629a <=( A168  and  A170 );
 a2632a <=( A166  and  (not A167) );
 a2633a <=( a2632a  and  a2629a );
 a2636a <=( A233  and  A232 );
 a2639a <=( (not A236)  and  A235 );
 a2640a <=( a2639a  and  a2636a );
 a2643a <=( A168  and  A170 );
 a2646a <=( A166  and  (not A167) );
 a2647a <=( a2646a  and  a2643a );
 a2650a <=( A233  and  (not A232) );
 a2653a <=( A236  and  (not A235) );
 a2654a <=( a2653a  and  a2650a );
 a2657a <=( A168  and  A170 );
 a2660a <=( A166  and  (not A167) );
 a2661a <=( a2660a  and  a2657a );
 a2664a <=( (not A233)  and  A232 );
 a2667a <=( A236  and  (not A235) );
 a2668a <=( a2667a  and  a2664a );
 a2671a <=( A168  and  A170 );
 a2674a <=( A166  and  (not A167) );
 a2675a <=( a2674a  and  a2671a );
 a2678a <=( (not A233)  and  (not A232) );
 a2681a <=( (not A236)  and  A235 );
 a2682a <=( a2681a  and  a2678a );
 a2685a <=( A168  and  A169 );
 a2688a <=( A166  and  (not A167) );
 a2689a <=( a2688a  and  a2685a );
 a2692a <=( A233  and  A232 );
 a2695a <=( (not A236)  and  A235 );
 a2696a <=( a2695a  and  a2692a );
 a2699a <=( A168  and  A169 );
 a2702a <=( A166  and  (not A167) );
 a2703a <=( a2702a  and  a2699a );
 a2706a <=( A233  and  (not A232) );
 a2709a <=( A236  and  (not A235) );
 a2710a <=( a2709a  and  a2706a );
 a2713a <=( A168  and  A169 );
 a2716a <=( A166  and  (not A167) );
 a2717a <=( a2716a  and  a2713a );
 a2720a <=( (not A233)  and  A232 );
 a2723a <=( A236  and  (not A235) );
 a2724a <=( a2723a  and  a2720a );
 a2727a <=( A168  and  A169 );
 a2730a <=( A166  and  (not A167) );
 a2731a <=( a2730a  and  a2727a );
 a2734a <=( (not A233)  and  (not A232) );
 a2737a <=( (not A236)  and  A235 );
 a2738a <=( a2737a  and  a2734a );
 a2741a <=( (not A166)  and  A167 );
 a2744a <=( (not A200)  and  (not A199) );
 a2745a <=( a2744a  and  a2741a );
 a2748a <=( A298  and  (not A202) );
 a2752a <=( (not A302)  and  A301 );
 a2753a <=( A299  and  a2752a );
 a2754a <=( a2753a  and  a2748a );
 a2757a <=( (not A166)  and  A167 );
 a2760a <=( (not A200)  and  (not A199) );
 a2761a <=( a2760a  and  a2757a );
 a2764a <=( A298  and  (not A202) );
 a2768a <=( A302  and  (not A301) );
 a2769a <=( (not A299)  and  a2768a );
 a2770a <=( a2769a  and  a2764a );
 a2773a <=( (not A166)  and  A167 );
 a2776a <=( (not A200)  and  (not A199) );
 a2777a <=( a2776a  and  a2773a );
 a2780a <=( (not A298)  and  (not A202) );
 a2784a <=( A302  and  (not A301) );
 a2785a <=( A299  and  a2784a );
 a2786a <=( a2785a  and  a2780a );
 a2789a <=( (not A166)  and  A167 );
 a2792a <=( (not A200)  and  (not A199) );
 a2793a <=( a2792a  and  a2789a );
 a2796a <=( (not A298)  and  (not A202) );
 a2800a <=( (not A302)  and  A301 );
 a2801a <=( (not A299)  and  a2800a );
 a2802a <=( a2801a  and  a2796a );
 a2805a <=( (not A166)  and  A167 );
 a2808a <=( (not A200)  and  (not A199) );
 a2809a <=( a2808a  and  a2805a );
 a2812a <=( A298  and  A203 );
 a2816a <=( (not A302)  and  A301 );
 a2817a <=( A299  and  a2816a );
 a2818a <=( a2817a  and  a2812a );
 a2821a <=( (not A166)  and  A167 );
 a2824a <=( (not A200)  and  (not A199) );
 a2825a <=( a2824a  and  a2821a );
 a2828a <=( A298  and  A203 );
 a2832a <=( A302  and  (not A301) );
 a2833a <=( (not A299)  and  a2832a );
 a2834a <=( a2833a  and  a2828a );
 a2837a <=( (not A166)  and  A167 );
 a2840a <=( (not A200)  and  (not A199) );
 a2841a <=( a2840a  and  a2837a );
 a2844a <=( (not A298)  and  A203 );
 a2848a <=( A302  and  (not A301) );
 a2849a <=( A299  and  a2848a );
 a2850a <=( a2849a  and  a2844a );
 a2853a <=( (not A166)  and  A167 );
 a2856a <=( (not A200)  and  (not A199) );
 a2857a <=( a2856a  and  a2853a );
 a2860a <=( (not A298)  and  A203 );
 a2864a <=( (not A302)  and  A301 );
 a2865a <=( (not A299)  and  a2864a );
 a2866a <=( a2865a  and  a2860a );
 a2869a <=( A168  and  A170 );
 a2872a <=( A166  and  (not A167) );
 a2873a <=( a2872a  and  a2869a );
 a2876a <=( (not A200)  and  (not A199) );
 a2880a <=( A300  and  A299 );
 a2881a <=( (not A202)  and  a2880a );
 a2882a <=( a2881a  and  a2876a );
 a2885a <=( A168  and  A170 );
 a2888a <=( A166  and  (not A167) );
 a2889a <=( a2888a  and  a2885a );
 a2892a <=( (not A200)  and  (not A199) );
 a2896a <=( A300  and  A298 );
 a2897a <=( (not A202)  and  a2896a );
 a2898a <=( a2897a  and  a2892a );
 a2901a <=( A168  and  A170 );
 a2904a <=( A166  and  (not A167) );
 a2905a <=( a2904a  and  a2901a );
 a2908a <=( (not A200)  and  (not A199) );
 a2912a <=( A300  and  A299 );
 a2913a <=( A203  and  a2912a );
 a2914a <=( a2913a  and  a2908a );
 a2917a <=( A168  and  A170 );
 a2920a <=( A166  and  (not A167) );
 a2921a <=( a2920a  and  a2917a );
 a2924a <=( (not A200)  and  (not A199) );
 a2928a <=( A300  and  A298 );
 a2929a <=( A203  and  a2928a );
 a2930a <=( a2929a  and  a2924a );
 a2933a <=( A168  and  A169 );
 a2936a <=( A166  and  (not A167) );
 a2937a <=( a2936a  and  a2933a );
 a2940a <=( (not A200)  and  (not A199) );
 a2944a <=( A300  and  A299 );
 a2945a <=( (not A202)  and  a2944a );
 a2946a <=( a2945a  and  a2940a );
 a2949a <=( A168  and  A169 );
 a2952a <=( A166  and  (not A167) );
 a2953a <=( a2952a  and  a2949a );
 a2956a <=( (not A200)  and  (not A199) );
 a2960a <=( A300  and  A298 );
 a2961a <=( (not A202)  and  a2960a );
 a2962a <=( a2961a  and  a2956a );
 a2965a <=( A168  and  A169 );
 a2968a <=( A166  and  (not A167) );
 a2969a <=( a2968a  and  a2965a );
 a2972a <=( (not A200)  and  (not A199) );
 a2976a <=( A300  and  A299 );
 a2977a <=( A203  and  a2976a );
 a2978a <=( a2977a  and  a2972a );
 a2981a <=( A168  and  A169 );
 a2984a <=( A166  and  (not A167) );
 a2985a <=( a2984a  and  a2981a );
 a2988a <=( (not A200)  and  (not A199) );
 a2992a <=( A300  and  A298 );
 a2993a <=( A203  and  a2992a );
 a2994a <=( a2993a  and  a2988a );
 a2997a <=( (not A169)  and  (not A170) );
 a3000a <=( A199  and  (not A167) );
 a3001a <=( a3000a  and  a2997a );
 a3004a <=( A298  and  A201 );
 a3008a <=( (not A302)  and  A301 );
 a3009a <=( A299  and  a3008a );
 a3010a <=( a3009a  and  a3004a );
 a3013a <=( (not A169)  and  (not A170) );
 a3016a <=( A199  and  (not A167) );
 a3017a <=( a3016a  and  a3013a );
 a3020a <=( A298  and  A201 );
 a3024a <=( A302  and  (not A301) );
 a3025a <=( (not A299)  and  a3024a );
 a3026a <=( a3025a  and  a3020a );
 a3029a <=( (not A169)  and  (not A170) );
 a3032a <=( A199  and  (not A167) );
 a3033a <=( a3032a  and  a3029a );
 a3036a <=( (not A298)  and  A201 );
 a3040a <=( A302  and  (not A301) );
 a3041a <=( A299  and  a3040a );
 a3042a <=( a3041a  and  a3036a );
 a3045a <=( (not A169)  and  (not A170) );
 a3048a <=( A199  and  (not A167) );
 a3049a <=( a3048a  and  a3045a );
 a3052a <=( (not A298)  and  A201 );
 a3056a <=( (not A302)  and  A301 );
 a3057a <=( (not A299)  and  a3056a );
 a3058a <=( a3057a  and  a3052a );
 a3061a <=( (not A169)  and  (not A170) );
 a3064a <=( A200  and  (not A167) );
 a3065a <=( a3064a  and  a3061a );
 a3068a <=( A298  and  A201 );
 a3072a <=( (not A302)  and  A301 );
 a3073a <=( A299  and  a3072a );
 a3074a <=( a3073a  and  a3068a );
 a3077a <=( (not A169)  and  (not A170) );
 a3080a <=( A200  and  (not A167) );
 a3081a <=( a3080a  and  a3077a );
 a3084a <=( A298  and  A201 );
 a3088a <=( A302  and  (not A301) );
 a3089a <=( (not A299)  and  a3088a );
 a3090a <=( a3089a  and  a3084a );
 a3093a <=( (not A169)  and  (not A170) );
 a3096a <=( A200  and  (not A167) );
 a3097a <=( a3096a  and  a3093a );
 a3100a <=( (not A298)  and  A201 );
 a3104a <=( A302  and  (not A301) );
 a3105a <=( A299  and  a3104a );
 a3106a <=( a3105a  and  a3100a );
 a3109a <=( (not A169)  and  (not A170) );
 a3112a <=( A200  and  (not A167) );
 a3113a <=( a3112a  and  a3109a );
 a3116a <=( (not A298)  and  A201 );
 a3120a <=( (not A302)  and  A301 );
 a3121a <=( (not A299)  and  a3120a );
 a3122a <=( a3121a  and  a3116a );
 a3125a <=( (not A169)  and  (not A170) );
 a3128a <=( A199  and  (not A167) );
 a3129a <=( a3128a  and  a3125a );
 a3132a <=( A202  and  A200 );
 a3136a <=( A300  and  A299 );
 a3137a <=( (not A203)  and  a3136a );
 a3138a <=( a3137a  and  a3132a );
 a3141a <=( (not A169)  and  (not A170) );
 a3144a <=( A199  and  (not A167) );
 a3145a <=( a3144a  and  a3141a );
 a3148a <=( A202  and  A200 );
 a3152a <=( A300  and  A298 );
 a3153a <=( (not A203)  and  a3152a );
 a3154a <=( a3153a  and  a3148a );
 a3157a <=( (not A169)  and  (not A170) );
 a3160a <=( (not A199)  and  (not A167) );
 a3161a <=( a3160a  and  a3157a );
 a3164a <=( (not A202)  and  A200 );
 a3168a <=( A300  and  A299 );
 a3169a <=( A203  and  a3168a );
 a3170a <=( a3169a  and  a3164a );
 a3173a <=( (not A169)  and  (not A170) );
 a3176a <=( (not A199)  and  (not A167) );
 a3177a <=( a3176a  and  a3173a );
 a3180a <=( (not A202)  and  A200 );
 a3184a <=( A300  and  A298 );
 a3185a <=( A203  and  a3184a );
 a3186a <=( a3185a  and  a3180a );
 a3189a <=( (not A169)  and  (not A170) );
 a3192a <=( A199  and  (not A167) );
 a3193a <=( a3192a  and  a3189a );
 a3196a <=( (not A202)  and  (not A200) );
 a3200a <=( A300  and  A299 );
 a3201a <=( A203  and  a3200a );
 a3202a <=( a3201a  and  a3196a );
 a3205a <=( (not A169)  and  (not A170) );
 a3208a <=( A199  and  (not A167) );
 a3209a <=( a3208a  and  a3205a );
 a3212a <=( (not A202)  and  (not A200) );
 a3216a <=( A300  and  A298 );
 a3217a <=( A203  and  a3216a );
 a3218a <=( a3217a  and  a3212a );
 a3221a <=( (not A169)  and  (not A170) );
 a3224a <=( (not A199)  and  (not A167) );
 a3225a <=( a3224a  and  a3221a );
 a3228a <=( A202  and  (not A200) );
 a3232a <=( A300  and  A299 );
 a3233a <=( (not A203)  and  a3232a );
 a3234a <=( a3233a  and  a3228a );
 a3237a <=( (not A169)  and  (not A170) );
 a3240a <=( (not A199)  and  (not A167) );
 a3241a <=( a3240a  and  a3237a );
 a3244a <=( A202  and  (not A200) );
 a3248a <=( A300  and  A298 );
 a3249a <=( (not A203)  and  a3248a );
 a3250a <=( a3249a  and  a3244a );
 a3253a <=( A166  and  A167 );
 a3257a <=( A202  and  A200 );
 a3258a <=( A199  and  a3257a );
 a3259a <=( a3258a  and  a3253a );
 a3262a <=( A298  and  (not A203) );
 a3266a <=( (not A302)  and  A301 );
 a3267a <=( A299  and  a3266a );
 a3268a <=( a3267a  and  a3262a );
 a3271a <=( A166  and  A167 );
 a3275a <=( A202  and  A200 );
 a3276a <=( A199  and  a3275a );
 a3277a <=( a3276a  and  a3271a );
 a3280a <=( A298  and  (not A203) );
 a3284a <=( A302  and  (not A301) );
 a3285a <=( (not A299)  and  a3284a );
 a3286a <=( a3285a  and  a3280a );
 a3289a <=( A166  and  A167 );
 a3293a <=( A202  and  A200 );
 a3294a <=( A199  and  a3293a );
 a3295a <=( a3294a  and  a3289a );
 a3298a <=( (not A298)  and  (not A203) );
 a3302a <=( A302  and  (not A301) );
 a3303a <=( A299  and  a3302a );
 a3304a <=( a3303a  and  a3298a );
 a3307a <=( A166  and  A167 );
 a3311a <=( A202  and  A200 );
 a3312a <=( A199  and  a3311a );
 a3313a <=( a3312a  and  a3307a );
 a3316a <=( (not A298)  and  (not A203) );
 a3320a <=( (not A302)  and  A301 );
 a3321a <=( (not A299)  and  a3320a );
 a3322a <=( a3321a  and  a3316a );
 a3325a <=( A166  and  A167 );
 a3329a <=( (not A202)  and  A200 );
 a3330a <=( (not A199)  and  a3329a );
 a3331a <=( a3330a  and  a3325a );
 a3334a <=( A298  and  A203 );
 a3338a <=( (not A302)  and  A301 );
 a3339a <=( A299  and  a3338a );
 a3340a <=( a3339a  and  a3334a );
 a3343a <=( A166  and  A167 );
 a3347a <=( (not A202)  and  A200 );
 a3348a <=( (not A199)  and  a3347a );
 a3349a <=( a3348a  and  a3343a );
 a3352a <=( A298  and  A203 );
 a3356a <=( A302  and  (not A301) );
 a3357a <=( (not A299)  and  a3356a );
 a3358a <=( a3357a  and  a3352a );
 a3361a <=( A166  and  A167 );
 a3365a <=( (not A202)  and  A200 );
 a3366a <=( (not A199)  and  a3365a );
 a3367a <=( a3366a  and  a3361a );
 a3370a <=( (not A298)  and  A203 );
 a3374a <=( A302  and  (not A301) );
 a3375a <=( A299  and  a3374a );
 a3376a <=( a3375a  and  a3370a );
 a3379a <=( A166  and  A167 );
 a3383a <=( (not A202)  and  A200 );
 a3384a <=( (not A199)  and  a3383a );
 a3385a <=( a3384a  and  a3379a );
 a3388a <=( (not A298)  and  A203 );
 a3392a <=( (not A302)  and  A301 );
 a3393a <=( (not A299)  and  a3392a );
 a3394a <=( a3393a  and  a3388a );
 a3397a <=( A166  and  A167 );
 a3401a <=( (not A202)  and  (not A200) );
 a3402a <=( A199  and  a3401a );
 a3403a <=( a3402a  and  a3397a );
 a3406a <=( A298  and  A203 );
 a3410a <=( (not A302)  and  A301 );
 a3411a <=( A299  and  a3410a );
 a3412a <=( a3411a  and  a3406a );
 a3415a <=( A166  and  A167 );
 a3419a <=( (not A202)  and  (not A200) );
 a3420a <=( A199  and  a3419a );
 a3421a <=( a3420a  and  a3415a );
 a3424a <=( A298  and  A203 );
 a3428a <=( A302  and  (not A301) );
 a3429a <=( (not A299)  and  a3428a );
 a3430a <=( a3429a  and  a3424a );
 a3433a <=( A166  and  A167 );
 a3437a <=( (not A202)  and  (not A200) );
 a3438a <=( A199  and  a3437a );
 a3439a <=( a3438a  and  a3433a );
 a3442a <=( (not A298)  and  A203 );
 a3446a <=( A302  and  (not A301) );
 a3447a <=( A299  and  a3446a );
 a3448a <=( a3447a  and  a3442a );
 a3451a <=( A166  and  A167 );
 a3455a <=( (not A202)  and  (not A200) );
 a3456a <=( A199  and  a3455a );
 a3457a <=( a3456a  and  a3451a );
 a3460a <=( (not A298)  and  A203 );
 a3464a <=( (not A302)  and  A301 );
 a3465a <=( (not A299)  and  a3464a );
 a3466a <=( a3465a  and  a3460a );
 a3469a <=( A166  and  A167 );
 a3473a <=( A202  and  (not A200) );
 a3474a <=( (not A199)  and  a3473a );
 a3475a <=( a3474a  and  a3469a );
 a3478a <=( A298  and  (not A203) );
 a3482a <=( (not A302)  and  A301 );
 a3483a <=( A299  and  a3482a );
 a3484a <=( a3483a  and  a3478a );
 a3487a <=( A166  and  A167 );
 a3491a <=( A202  and  (not A200) );
 a3492a <=( (not A199)  and  a3491a );
 a3493a <=( a3492a  and  a3487a );
 a3496a <=( A298  and  (not A203) );
 a3500a <=( A302  and  (not A301) );
 a3501a <=( (not A299)  and  a3500a );
 a3502a <=( a3501a  and  a3496a );
 a3505a <=( A166  and  A167 );
 a3509a <=( A202  and  (not A200) );
 a3510a <=( (not A199)  and  a3509a );
 a3511a <=( a3510a  and  a3505a );
 a3514a <=( (not A298)  and  (not A203) );
 a3518a <=( A302  and  (not A301) );
 a3519a <=( A299  and  a3518a );
 a3520a <=( a3519a  and  a3514a );
 a3523a <=( A166  and  A167 );
 a3527a <=( A202  and  (not A200) );
 a3528a <=( (not A199)  and  a3527a );
 a3529a <=( a3528a  and  a3523a );
 a3532a <=( (not A298)  and  (not A203) );
 a3536a <=( (not A302)  and  A301 );
 a3537a <=( (not A299)  and  a3536a );
 a3538a <=( a3537a  and  a3532a );
 a3541a <=( (not A166)  and  A167 );
 a3545a <=( (not A201)  and  A200 );
 a3546a <=( A199  and  a3545a );
 a3547a <=( a3546a  and  a3541a );
 a3550a <=( A298  and  (not A202) );
 a3554a <=( (not A302)  and  A301 );
 a3555a <=( A299  and  a3554a );
 a3556a <=( a3555a  and  a3550a );
 a3559a <=( (not A166)  and  A167 );
 a3563a <=( (not A201)  and  A200 );
 a3564a <=( A199  and  a3563a );
 a3565a <=( a3564a  and  a3559a );
 a3568a <=( A298  and  (not A202) );
 a3572a <=( A302  and  (not A301) );
 a3573a <=( (not A299)  and  a3572a );
 a3574a <=( a3573a  and  a3568a );
 a3577a <=( (not A166)  and  A167 );
 a3581a <=( (not A201)  and  A200 );
 a3582a <=( A199  and  a3581a );
 a3583a <=( a3582a  and  a3577a );
 a3586a <=( (not A298)  and  (not A202) );
 a3590a <=( A302  and  (not A301) );
 a3591a <=( A299  and  a3590a );
 a3592a <=( a3591a  and  a3586a );
 a3595a <=( (not A166)  and  A167 );
 a3599a <=( (not A201)  and  A200 );
 a3600a <=( A199  and  a3599a );
 a3601a <=( a3600a  and  a3595a );
 a3604a <=( (not A298)  and  (not A202) );
 a3608a <=( (not A302)  and  A301 );
 a3609a <=( (not A299)  and  a3608a );
 a3610a <=( a3609a  and  a3604a );
 a3613a <=( (not A166)  and  A167 );
 a3617a <=( (not A201)  and  A200 );
 a3618a <=( A199  and  a3617a );
 a3619a <=( a3618a  and  a3613a );
 a3622a <=( A298  and  A203 );
 a3626a <=( (not A302)  and  A301 );
 a3627a <=( A299  and  a3626a );
 a3628a <=( a3627a  and  a3622a );
 a3631a <=( (not A166)  and  A167 );
 a3635a <=( (not A201)  and  A200 );
 a3636a <=( A199  and  a3635a );
 a3637a <=( a3636a  and  a3631a );
 a3640a <=( A298  and  A203 );
 a3644a <=( A302  and  (not A301) );
 a3645a <=( (not A299)  and  a3644a );
 a3646a <=( a3645a  and  a3640a );
 a3649a <=( (not A166)  and  A167 );
 a3653a <=( (not A201)  and  A200 );
 a3654a <=( A199  and  a3653a );
 a3655a <=( a3654a  and  a3649a );
 a3658a <=( (not A298)  and  A203 );
 a3662a <=( A302  and  (not A301) );
 a3663a <=( A299  and  a3662a );
 a3664a <=( a3663a  and  a3658a );
 a3667a <=( (not A166)  and  A167 );
 a3671a <=( (not A201)  and  A200 );
 a3672a <=( A199  and  a3671a );
 a3673a <=( a3672a  and  a3667a );
 a3676a <=( (not A298)  and  A203 );
 a3680a <=( (not A302)  and  A301 );
 a3681a <=( (not A299)  and  a3680a );
 a3682a <=( a3681a  and  a3676a );
 a3685a <=( (not A166)  and  A167 );
 a3689a <=( (not A201)  and  A200 );
 a3690a <=( (not A199)  and  a3689a );
 a3691a <=( a3690a  and  a3685a );
 a3694a <=( A298  and  A202 );
 a3698a <=( (not A302)  and  A301 );
 a3699a <=( A299  and  a3698a );
 a3700a <=( a3699a  and  a3694a );
 a3703a <=( (not A166)  and  A167 );
 a3707a <=( (not A201)  and  A200 );
 a3708a <=( (not A199)  and  a3707a );
 a3709a <=( a3708a  and  a3703a );
 a3712a <=( A298  and  A202 );
 a3716a <=( A302  and  (not A301) );
 a3717a <=( (not A299)  and  a3716a );
 a3718a <=( a3717a  and  a3712a );
 a3721a <=( (not A166)  and  A167 );
 a3725a <=( (not A201)  and  A200 );
 a3726a <=( (not A199)  and  a3725a );
 a3727a <=( a3726a  and  a3721a );
 a3730a <=( (not A298)  and  A202 );
 a3734a <=( A302  and  (not A301) );
 a3735a <=( A299  and  a3734a );
 a3736a <=( a3735a  and  a3730a );
 a3739a <=( (not A166)  and  A167 );
 a3743a <=( (not A201)  and  A200 );
 a3744a <=( (not A199)  and  a3743a );
 a3745a <=( a3744a  and  a3739a );
 a3748a <=( (not A298)  and  A202 );
 a3752a <=( (not A302)  and  A301 );
 a3753a <=( (not A299)  and  a3752a );
 a3754a <=( a3753a  and  a3748a );
 a3757a <=( (not A166)  and  A167 );
 a3761a <=( (not A201)  and  A200 );
 a3762a <=( (not A199)  and  a3761a );
 a3763a <=( a3762a  and  a3757a );
 a3766a <=( A298  and  (not A203) );
 a3770a <=( (not A302)  and  A301 );
 a3771a <=( A299  and  a3770a );
 a3772a <=( a3771a  and  a3766a );
 a3775a <=( (not A166)  and  A167 );
 a3779a <=( (not A201)  and  A200 );
 a3780a <=( (not A199)  and  a3779a );
 a3781a <=( a3780a  and  a3775a );
 a3784a <=( A298  and  (not A203) );
 a3788a <=( A302  and  (not A301) );
 a3789a <=( (not A299)  and  a3788a );
 a3790a <=( a3789a  and  a3784a );
 a3793a <=( (not A166)  and  A167 );
 a3797a <=( (not A201)  and  A200 );
 a3798a <=( (not A199)  and  a3797a );
 a3799a <=( a3798a  and  a3793a );
 a3802a <=( (not A298)  and  (not A203) );
 a3806a <=( A302  and  (not A301) );
 a3807a <=( A299  and  a3806a );
 a3808a <=( a3807a  and  a3802a );
 a3811a <=( (not A166)  and  A167 );
 a3815a <=( (not A201)  and  A200 );
 a3816a <=( (not A199)  and  a3815a );
 a3817a <=( a3816a  and  a3811a );
 a3820a <=( (not A298)  and  (not A203) );
 a3824a <=( (not A302)  and  A301 );
 a3825a <=( (not A299)  and  a3824a );
 a3826a <=( a3825a  and  a3820a );
 a3829a <=( (not A166)  and  A167 );
 a3833a <=( (not A201)  and  (not A200) );
 a3834a <=( A199  and  a3833a );
 a3835a <=( a3834a  and  a3829a );
 a3838a <=( A298  and  A202 );
 a3842a <=( (not A302)  and  A301 );
 a3843a <=( A299  and  a3842a );
 a3844a <=( a3843a  and  a3838a );
 a3847a <=( (not A166)  and  A167 );
 a3851a <=( (not A201)  and  (not A200) );
 a3852a <=( A199  and  a3851a );
 a3853a <=( a3852a  and  a3847a );
 a3856a <=( A298  and  A202 );
 a3860a <=( A302  and  (not A301) );
 a3861a <=( (not A299)  and  a3860a );
 a3862a <=( a3861a  and  a3856a );
 a3865a <=( (not A166)  and  A167 );
 a3869a <=( (not A201)  and  (not A200) );
 a3870a <=( A199  and  a3869a );
 a3871a <=( a3870a  and  a3865a );
 a3874a <=( (not A298)  and  A202 );
 a3878a <=( A302  and  (not A301) );
 a3879a <=( A299  and  a3878a );
 a3880a <=( a3879a  and  a3874a );
 a3883a <=( (not A166)  and  A167 );
 a3887a <=( (not A201)  and  (not A200) );
 a3888a <=( A199  and  a3887a );
 a3889a <=( a3888a  and  a3883a );
 a3892a <=( (not A298)  and  A202 );
 a3896a <=( (not A302)  and  A301 );
 a3897a <=( (not A299)  and  a3896a );
 a3898a <=( a3897a  and  a3892a );
 a3901a <=( (not A166)  and  A167 );
 a3905a <=( (not A201)  and  (not A200) );
 a3906a <=( A199  and  a3905a );
 a3907a <=( a3906a  and  a3901a );
 a3910a <=( A298  and  (not A203) );
 a3914a <=( (not A302)  and  A301 );
 a3915a <=( A299  and  a3914a );
 a3916a <=( a3915a  and  a3910a );
 a3919a <=( (not A166)  and  A167 );
 a3923a <=( (not A201)  and  (not A200) );
 a3924a <=( A199  and  a3923a );
 a3925a <=( a3924a  and  a3919a );
 a3928a <=( A298  and  (not A203) );
 a3932a <=( A302  and  (not A301) );
 a3933a <=( (not A299)  and  a3932a );
 a3934a <=( a3933a  and  a3928a );
 a3937a <=( (not A166)  and  A167 );
 a3941a <=( (not A201)  and  (not A200) );
 a3942a <=( A199  and  a3941a );
 a3943a <=( a3942a  and  a3937a );
 a3946a <=( (not A298)  and  (not A203) );
 a3950a <=( A302  and  (not A301) );
 a3951a <=( A299  and  a3950a );
 a3952a <=( a3951a  and  a3946a );
 a3955a <=( (not A166)  and  A167 );
 a3959a <=( (not A201)  and  (not A200) );
 a3960a <=( A199  and  a3959a );
 a3961a <=( a3960a  and  a3955a );
 a3964a <=( (not A298)  and  (not A203) );
 a3968a <=( (not A302)  and  A301 );
 a3969a <=( (not A299)  and  a3968a );
 a3970a <=( a3969a  and  a3964a );
 a3973a <=( (not A166)  and  (not A167) );
 a3977a <=( A202  and  A200 );
 a3978a <=( A199  and  a3977a );
 a3979a <=( a3978a  and  a3973a );
 a3982a <=( A298  and  (not A203) );
 a3986a <=( (not A302)  and  A301 );
 a3987a <=( A299  and  a3986a );
 a3988a <=( a3987a  and  a3982a );
 a3991a <=( (not A166)  and  (not A167) );
 a3995a <=( A202  and  A200 );
 a3996a <=( A199  and  a3995a );
 a3997a <=( a3996a  and  a3991a );
 a4000a <=( A298  and  (not A203) );
 a4004a <=( A302  and  (not A301) );
 a4005a <=( (not A299)  and  a4004a );
 a4006a <=( a4005a  and  a4000a );
 a4009a <=( (not A166)  and  (not A167) );
 a4013a <=( A202  and  A200 );
 a4014a <=( A199  and  a4013a );
 a4015a <=( a4014a  and  a4009a );
 a4018a <=( (not A298)  and  (not A203) );
 a4022a <=( A302  and  (not A301) );
 a4023a <=( A299  and  a4022a );
 a4024a <=( a4023a  and  a4018a );
 a4027a <=( (not A166)  and  (not A167) );
 a4031a <=( A202  and  A200 );
 a4032a <=( A199  and  a4031a );
 a4033a <=( a4032a  and  a4027a );
 a4036a <=( (not A298)  and  (not A203) );
 a4040a <=( (not A302)  and  A301 );
 a4041a <=( (not A299)  and  a4040a );
 a4042a <=( a4041a  and  a4036a );
 a4045a <=( (not A166)  and  (not A167) );
 a4049a <=( (not A202)  and  A200 );
 a4050a <=( (not A199)  and  a4049a );
 a4051a <=( a4050a  and  a4045a );
 a4054a <=( A298  and  A203 );
 a4058a <=( (not A302)  and  A301 );
 a4059a <=( A299  and  a4058a );
 a4060a <=( a4059a  and  a4054a );
 a4063a <=( (not A166)  and  (not A167) );
 a4067a <=( (not A202)  and  A200 );
 a4068a <=( (not A199)  and  a4067a );
 a4069a <=( a4068a  and  a4063a );
 a4072a <=( A298  and  A203 );
 a4076a <=( A302  and  (not A301) );
 a4077a <=( (not A299)  and  a4076a );
 a4078a <=( a4077a  and  a4072a );
 a4081a <=( (not A166)  and  (not A167) );
 a4085a <=( (not A202)  and  A200 );
 a4086a <=( (not A199)  and  a4085a );
 a4087a <=( a4086a  and  a4081a );
 a4090a <=( (not A298)  and  A203 );
 a4094a <=( A302  and  (not A301) );
 a4095a <=( A299  and  a4094a );
 a4096a <=( a4095a  and  a4090a );
 a4099a <=( (not A166)  and  (not A167) );
 a4103a <=( (not A202)  and  A200 );
 a4104a <=( (not A199)  and  a4103a );
 a4105a <=( a4104a  and  a4099a );
 a4108a <=( (not A298)  and  A203 );
 a4112a <=( (not A302)  and  A301 );
 a4113a <=( (not A299)  and  a4112a );
 a4114a <=( a4113a  and  a4108a );
 a4117a <=( (not A166)  and  (not A167) );
 a4121a <=( (not A202)  and  (not A200) );
 a4122a <=( A199  and  a4121a );
 a4123a <=( a4122a  and  a4117a );
 a4126a <=( A298  and  A203 );
 a4130a <=( (not A302)  and  A301 );
 a4131a <=( A299  and  a4130a );
 a4132a <=( a4131a  and  a4126a );
 a4135a <=( (not A166)  and  (not A167) );
 a4139a <=( (not A202)  and  (not A200) );
 a4140a <=( A199  and  a4139a );
 a4141a <=( a4140a  and  a4135a );
 a4144a <=( A298  and  A203 );
 a4148a <=( A302  and  (not A301) );
 a4149a <=( (not A299)  and  a4148a );
 a4150a <=( a4149a  and  a4144a );
 a4153a <=( (not A166)  and  (not A167) );
 a4157a <=( (not A202)  and  (not A200) );
 a4158a <=( A199  and  a4157a );
 a4159a <=( a4158a  and  a4153a );
 a4162a <=( (not A298)  and  A203 );
 a4166a <=( A302  and  (not A301) );
 a4167a <=( A299  and  a4166a );
 a4168a <=( a4167a  and  a4162a );
 a4171a <=( (not A166)  and  (not A167) );
 a4175a <=( (not A202)  and  (not A200) );
 a4176a <=( A199  and  a4175a );
 a4177a <=( a4176a  and  a4171a );
 a4180a <=( (not A298)  and  A203 );
 a4184a <=( (not A302)  and  A301 );
 a4185a <=( (not A299)  and  a4184a );
 a4186a <=( a4185a  and  a4180a );
 a4189a <=( (not A166)  and  (not A167) );
 a4193a <=( A202  and  (not A200) );
 a4194a <=( (not A199)  and  a4193a );
 a4195a <=( a4194a  and  a4189a );
 a4198a <=( A298  and  (not A203) );
 a4202a <=( (not A302)  and  A301 );
 a4203a <=( A299  and  a4202a );
 a4204a <=( a4203a  and  a4198a );
 a4207a <=( (not A166)  and  (not A167) );
 a4211a <=( A202  and  (not A200) );
 a4212a <=( (not A199)  and  a4211a );
 a4213a <=( a4212a  and  a4207a );
 a4216a <=( A298  and  (not A203) );
 a4220a <=( A302  and  (not A301) );
 a4221a <=( (not A299)  and  a4220a );
 a4222a <=( a4221a  and  a4216a );
 a4225a <=( (not A166)  and  (not A167) );
 a4229a <=( A202  and  (not A200) );
 a4230a <=( (not A199)  and  a4229a );
 a4231a <=( a4230a  and  a4225a );
 a4234a <=( (not A298)  and  (not A203) );
 a4238a <=( A302  and  (not A301) );
 a4239a <=( A299  and  a4238a );
 a4240a <=( a4239a  and  a4234a );
 a4243a <=( (not A166)  and  (not A167) );
 a4247a <=( A202  and  (not A200) );
 a4248a <=( (not A199)  and  a4247a );
 a4249a <=( a4248a  and  a4243a );
 a4252a <=( (not A298)  and  (not A203) );
 a4256a <=( (not A302)  and  A301 );
 a4257a <=( (not A299)  and  a4256a );
 a4258a <=( a4257a  and  a4252a );
 a4261a <=( (not A167)  and  (not A168) );
 a4265a <=( A202  and  A200 );
 a4266a <=( A199  and  a4265a );
 a4267a <=( a4266a  and  a4261a );
 a4270a <=( A298  and  (not A203) );
 a4274a <=( (not A302)  and  A301 );
 a4275a <=( A299  and  a4274a );
 a4276a <=( a4275a  and  a4270a );
 a4279a <=( (not A167)  and  (not A168) );
 a4283a <=( A202  and  A200 );
 a4284a <=( A199  and  a4283a );
 a4285a <=( a4284a  and  a4279a );
 a4288a <=( A298  and  (not A203) );
 a4292a <=( A302  and  (not A301) );
 a4293a <=( (not A299)  and  a4292a );
 a4294a <=( a4293a  and  a4288a );
 a4297a <=( (not A167)  and  (not A168) );
 a4301a <=( A202  and  A200 );
 a4302a <=( A199  and  a4301a );
 a4303a <=( a4302a  and  a4297a );
 a4306a <=( (not A298)  and  (not A203) );
 a4310a <=( A302  and  (not A301) );
 a4311a <=( A299  and  a4310a );
 a4312a <=( a4311a  and  a4306a );
 a4315a <=( (not A167)  and  (not A168) );
 a4319a <=( A202  and  A200 );
 a4320a <=( A199  and  a4319a );
 a4321a <=( a4320a  and  a4315a );
 a4324a <=( (not A298)  and  (not A203) );
 a4328a <=( (not A302)  and  A301 );
 a4329a <=( (not A299)  and  a4328a );
 a4330a <=( a4329a  and  a4324a );
 a4333a <=( (not A167)  and  (not A168) );
 a4337a <=( (not A202)  and  A200 );
 a4338a <=( (not A199)  and  a4337a );
 a4339a <=( a4338a  and  a4333a );
 a4342a <=( A298  and  A203 );
 a4346a <=( (not A302)  and  A301 );
 a4347a <=( A299  and  a4346a );
 a4348a <=( a4347a  and  a4342a );
 a4351a <=( (not A167)  and  (not A168) );
 a4355a <=( (not A202)  and  A200 );
 a4356a <=( (not A199)  and  a4355a );
 a4357a <=( a4356a  and  a4351a );
 a4360a <=( A298  and  A203 );
 a4364a <=( A302  and  (not A301) );
 a4365a <=( (not A299)  and  a4364a );
 a4366a <=( a4365a  and  a4360a );
 a4369a <=( (not A167)  and  (not A168) );
 a4373a <=( (not A202)  and  A200 );
 a4374a <=( (not A199)  and  a4373a );
 a4375a <=( a4374a  and  a4369a );
 a4378a <=( (not A298)  and  A203 );
 a4382a <=( A302  and  (not A301) );
 a4383a <=( A299  and  a4382a );
 a4384a <=( a4383a  and  a4378a );
 a4387a <=( (not A167)  and  (not A168) );
 a4391a <=( (not A202)  and  A200 );
 a4392a <=( (not A199)  and  a4391a );
 a4393a <=( a4392a  and  a4387a );
 a4396a <=( (not A298)  and  A203 );
 a4400a <=( (not A302)  and  A301 );
 a4401a <=( (not A299)  and  a4400a );
 a4402a <=( a4401a  and  a4396a );
 a4405a <=( (not A167)  and  (not A168) );
 a4409a <=( (not A202)  and  (not A200) );
 a4410a <=( A199  and  a4409a );
 a4411a <=( a4410a  and  a4405a );
 a4414a <=( A298  and  A203 );
 a4418a <=( (not A302)  and  A301 );
 a4419a <=( A299  and  a4418a );
 a4420a <=( a4419a  and  a4414a );
 a4423a <=( (not A167)  and  (not A168) );
 a4427a <=( (not A202)  and  (not A200) );
 a4428a <=( A199  and  a4427a );
 a4429a <=( a4428a  and  a4423a );
 a4432a <=( A298  and  A203 );
 a4436a <=( A302  and  (not A301) );
 a4437a <=( (not A299)  and  a4436a );
 a4438a <=( a4437a  and  a4432a );
 a4441a <=( (not A167)  and  (not A168) );
 a4445a <=( (not A202)  and  (not A200) );
 a4446a <=( A199  and  a4445a );
 a4447a <=( a4446a  and  a4441a );
 a4450a <=( (not A298)  and  A203 );
 a4454a <=( A302  and  (not A301) );
 a4455a <=( A299  and  a4454a );
 a4456a <=( a4455a  and  a4450a );
 a4459a <=( (not A167)  and  (not A168) );
 a4463a <=( (not A202)  and  (not A200) );
 a4464a <=( A199  and  a4463a );
 a4465a <=( a4464a  and  a4459a );
 a4468a <=( (not A298)  and  A203 );
 a4472a <=( (not A302)  and  A301 );
 a4473a <=( (not A299)  and  a4472a );
 a4474a <=( a4473a  and  a4468a );
 a4477a <=( (not A167)  and  (not A168) );
 a4481a <=( A202  and  (not A200) );
 a4482a <=( (not A199)  and  a4481a );
 a4483a <=( a4482a  and  a4477a );
 a4486a <=( A298  and  (not A203) );
 a4490a <=( (not A302)  and  A301 );
 a4491a <=( A299  and  a4490a );
 a4492a <=( a4491a  and  a4486a );
 a4495a <=( (not A167)  and  (not A168) );
 a4499a <=( A202  and  (not A200) );
 a4500a <=( (not A199)  and  a4499a );
 a4501a <=( a4500a  and  a4495a );
 a4504a <=( A298  and  (not A203) );
 a4508a <=( A302  and  (not A301) );
 a4509a <=( (not A299)  and  a4508a );
 a4510a <=( a4509a  and  a4504a );
 a4513a <=( (not A167)  and  (not A168) );
 a4517a <=( A202  and  (not A200) );
 a4518a <=( (not A199)  and  a4517a );
 a4519a <=( a4518a  and  a4513a );
 a4522a <=( (not A298)  and  (not A203) );
 a4526a <=( A302  and  (not A301) );
 a4527a <=( A299  and  a4526a );
 a4528a <=( a4527a  and  a4522a );
 a4531a <=( (not A167)  and  (not A168) );
 a4535a <=( A202  and  (not A200) );
 a4536a <=( (not A199)  and  a4535a );
 a4537a <=( a4536a  and  a4531a );
 a4540a <=( (not A298)  and  (not A203) );
 a4544a <=( (not A302)  and  A301 );
 a4545a <=( (not A299)  and  a4544a );
 a4546a <=( a4545a  and  a4540a );
 a4549a <=( A168  and  A170 );
 a4553a <=( A199  and  A166 );
 a4554a <=( (not A167)  and  a4553a );
 a4555a <=( a4554a  and  a4549a );
 a4558a <=( (not A201)  and  A200 );
 a4562a <=( A300  and  A299 );
 a4563a <=( (not A202)  and  a4562a );
 a4564a <=( a4563a  and  a4558a );
 a4567a <=( A168  and  A170 );
 a4571a <=( A199  and  A166 );
 a4572a <=( (not A167)  and  a4571a );
 a4573a <=( a4572a  and  a4567a );
 a4576a <=( (not A201)  and  A200 );
 a4580a <=( A300  and  A298 );
 a4581a <=( (not A202)  and  a4580a );
 a4582a <=( a4581a  and  a4576a );
 a4585a <=( A168  and  A170 );
 a4589a <=( A199  and  A166 );
 a4590a <=( (not A167)  and  a4589a );
 a4591a <=( a4590a  and  a4585a );
 a4594a <=( (not A201)  and  A200 );
 a4598a <=( A300  and  A299 );
 a4599a <=( A203  and  a4598a );
 a4600a <=( a4599a  and  a4594a );
 a4603a <=( A168  and  A170 );
 a4607a <=( A199  and  A166 );
 a4608a <=( (not A167)  and  a4607a );
 a4609a <=( a4608a  and  a4603a );
 a4612a <=( (not A201)  and  A200 );
 a4616a <=( A300  and  A298 );
 a4617a <=( A203  and  a4616a );
 a4618a <=( a4617a  and  a4612a );
 a4621a <=( A168  and  A170 );
 a4625a <=( (not A199)  and  A166 );
 a4626a <=( (not A167)  and  a4625a );
 a4627a <=( a4626a  and  a4621a );
 a4630a <=( (not A201)  and  A200 );
 a4634a <=( A300  and  A299 );
 a4635a <=( A202  and  a4634a );
 a4636a <=( a4635a  and  a4630a );
 a4639a <=( A168  and  A170 );
 a4643a <=( (not A199)  and  A166 );
 a4644a <=( (not A167)  and  a4643a );
 a4645a <=( a4644a  and  a4639a );
 a4648a <=( (not A201)  and  A200 );
 a4652a <=( A300  and  A298 );
 a4653a <=( A202  and  a4652a );
 a4654a <=( a4653a  and  a4648a );
 a4657a <=( A168  and  A170 );
 a4661a <=( (not A199)  and  A166 );
 a4662a <=( (not A167)  and  a4661a );
 a4663a <=( a4662a  and  a4657a );
 a4666a <=( (not A201)  and  A200 );
 a4670a <=( A300  and  A299 );
 a4671a <=( (not A203)  and  a4670a );
 a4672a <=( a4671a  and  a4666a );
 a4675a <=( A168  and  A170 );
 a4679a <=( (not A199)  and  A166 );
 a4680a <=( (not A167)  and  a4679a );
 a4681a <=( a4680a  and  a4675a );
 a4684a <=( (not A201)  and  A200 );
 a4688a <=( A300  and  A298 );
 a4689a <=( (not A203)  and  a4688a );
 a4690a <=( a4689a  and  a4684a );
 a4693a <=( A168  and  A170 );
 a4697a <=( A199  and  A166 );
 a4698a <=( (not A167)  and  a4697a );
 a4699a <=( a4698a  and  a4693a );
 a4702a <=( (not A201)  and  (not A200) );
 a4706a <=( A300  and  A299 );
 a4707a <=( A202  and  a4706a );
 a4708a <=( a4707a  and  a4702a );
 a4711a <=( A168  and  A170 );
 a4715a <=( A199  and  A166 );
 a4716a <=( (not A167)  and  a4715a );
 a4717a <=( a4716a  and  a4711a );
 a4720a <=( (not A201)  and  (not A200) );
 a4724a <=( A300  and  A298 );
 a4725a <=( A202  and  a4724a );
 a4726a <=( a4725a  and  a4720a );
 a4729a <=( A168  and  A170 );
 a4733a <=( A199  and  A166 );
 a4734a <=( (not A167)  and  a4733a );
 a4735a <=( a4734a  and  a4729a );
 a4738a <=( (not A201)  and  (not A200) );
 a4742a <=( A300  and  A299 );
 a4743a <=( (not A203)  and  a4742a );
 a4744a <=( a4743a  and  a4738a );
 a4747a <=( A168  and  A170 );
 a4751a <=( A199  and  A166 );
 a4752a <=( (not A167)  and  a4751a );
 a4753a <=( a4752a  and  a4747a );
 a4756a <=( (not A201)  and  (not A200) );
 a4760a <=( A300  and  A298 );
 a4761a <=( (not A203)  and  a4760a );
 a4762a <=( a4761a  and  a4756a );
 a4765a <=( A168  and  A169 );
 a4769a <=( A199  and  A166 );
 a4770a <=( (not A167)  and  a4769a );
 a4771a <=( a4770a  and  a4765a );
 a4774a <=( (not A201)  and  A200 );
 a4778a <=( A300  and  A299 );
 a4779a <=( (not A202)  and  a4778a );
 a4780a <=( a4779a  and  a4774a );
 a4783a <=( A168  and  A169 );
 a4787a <=( A199  and  A166 );
 a4788a <=( (not A167)  and  a4787a );
 a4789a <=( a4788a  and  a4783a );
 a4792a <=( (not A201)  and  A200 );
 a4796a <=( A300  and  A298 );
 a4797a <=( (not A202)  and  a4796a );
 a4798a <=( a4797a  and  a4792a );
 a4801a <=( A168  and  A169 );
 a4805a <=( A199  and  A166 );
 a4806a <=( (not A167)  and  a4805a );
 a4807a <=( a4806a  and  a4801a );
 a4810a <=( (not A201)  and  A200 );
 a4814a <=( A300  and  A299 );
 a4815a <=( A203  and  a4814a );
 a4816a <=( a4815a  and  a4810a );
 a4819a <=( A168  and  A169 );
 a4823a <=( A199  and  A166 );
 a4824a <=( (not A167)  and  a4823a );
 a4825a <=( a4824a  and  a4819a );
 a4828a <=( (not A201)  and  A200 );
 a4832a <=( A300  and  A298 );
 a4833a <=( A203  and  a4832a );
 a4834a <=( a4833a  and  a4828a );
 a4837a <=( A168  and  A169 );
 a4841a <=( (not A199)  and  A166 );
 a4842a <=( (not A167)  and  a4841a );
 a4843a <=( a4842a  and  a4837a );
 a4846a <=( (not A201)  and  A200 );
 a4850a <=( A300  and  A299 );
 a4851a <=( A202  and  a4850a );
 a4852a <=( a4851a  and  a4846a );
 a4855a <=( A168  and  A169 );
 a4859a <=( (not A199)  and  A166 );
 a4860a <=( (not A167)  and  a4859a );
 a4861a <=( a4860a  and  a4855a );
 a4864a <=( (not A201)  and  A200 );
 a4868a <=( A300  and  A298 );
 a4869a <=( A202  and  a4868a );
 a4870a <=( a4869a  and  a4864a );
 a4873a <=( A168  and  A169 );
 a4877a <=( (not A199)  and  A166 );
 a4878a <=( (not A167)  and  a4877a );
 a4879a <=( a4878a  and  a4873a );
 a4882a <=( (not A201)  and  A200 );
 a4886a <=( A300  and  A299 );
 a4887a <=( (not A203)  and  a4886a );
 a4888a <=( a4887a  and  a4882a );
 a4891a <=( A168  and  A169 );
 a4895a <=( (not A199)  and  A166 );
 a4896a <=( (not A167)  and  a4895a );
 a4897a <=( a4896a  and  a4891a );
 a4900a <=( (not A201)  and  A200 );
 a4904a <=( A300  and  A298 );
 a4905a <=( (not A203)  and  a4904a );
 a4906a <=( a4905a  and  a4900a );
 a4909a <=( A168  and  A169 );
 a4913a <=( A199  and  A166 );
 a4914a <=( (not A167)  and  a4913a );
 a4915a <=( a4914a  and  a4909a );
 a4918a <=( (not A201)  and  (not A200) );
 a4922a <=( A300  and  A299 );
 a4923a <=( A202  and  a4922a );
 a4924a <=( a4923a  and  a4918a );
 a4927a <=( A168  and  A169 );
 a4931a <=( A199  and  A166 );
 a4932a <=( (not A167)  and  a4931a );
 a4933a <=( a4932a  and  a4927a );
 a4936a <=( (not A201)  and  (not A200) );
 a4940a <=( A300  and  A298 );
 a4941a <=( A202  and  a4940a );
 a4942a <=( a4941a  and  a4936a );
 a4945a <=( A168  and  A169 );
 a4949a <=( A199  and  A166 );
 a4950a <=( (not A167)  and  a4949a );
 a4951a <=( a4950a  and  a4945a );
 a4954a <=( (not A201)  and  (not A200) );
 a4958a <=( A300  and  A299 );
 a4959a <=( (not A203)  and  a4958a );
 a4960a <=( a4959a  and  a4954a );
 a4963a <=( A168  and  A169 );
 a4967a <=( A199  and  A166 );
 a4968a <=( (not A167)  and  a4967a );
 a4969a <=( a4968a  and  a4963a );
 a4972a <=( (not A201)  and  (not A200) );
 a4976a <=( A300  and  A298 );
 a4977a <=( (not A203)  and  a4976a );
 a4978a <=( a4977a  and  a4972a );
 a4981a <=( A168  and  A170 );
 a4985a <=( (not A199)  and  A166 );
 a4986a <=( (not A167)  and  a4985a );
 a4987a <=( a4986a  and  a4981a );
 a4991a <=( A298  and  (not A202) );
 a4992a <=( (not A200)  and  a4991a );
 a4996a <=( (not A302)  and  A301 );
 a4997a <=( A299  and  a4996a );
 a4998a <=( a4997a  and  a4992a );
 a5001a <=( A168  and  A170 );
 a5005a <=( (not A199)  and  A166 );
 a5006a <=( (not A167)  and  a5005a );
 a5007a <=( a5006a  and  a5001a );
 a5011a <=( A298  and  (not A202) );
 a5012a <=( (not A200)  and  a5011a );
 a5016a <=( A302  and  (not A301) );
 a5017a <=( (not A299)  and  a5016a );
 a5018a <=( a5017a  and  a5012a );
 a5021a <=( A168  and  A170 );
 a5025a <=( (not A199)  and  A166 );
 a5026a <=( (not A167)  and  a5025a );
 a5027a <=( a5026a  and  a5021a );
 a5031a <=( (not A298)  and  (not A202) );
 a5032a <=( (not A200)  and  a5031a );
 a5036a <=( A302  and  (not A301) );
 a5037a <=( A299  and  a5036a );
 a5038a <=( a5037a  and  a5032a );
 a5041a <=( A168  and  A170 );
 a5045a <=( (not A199)  and  A166 );
 a5046a <=( (not A167)  and  a5045a );
 a5047a <=( a5046a  and  a5041a );
 a5051a <=( (not A298)  and  (not A202) );
 a5052a <=( (not A200)  and  a5051a );
 a5056a <=( (not A302)  and  A301 );
 a5057a <=( (not A299)  and  a5056a );
 a5058a <=( a5057a  and  a5052a );
 a5061a <=( A168  and  A170 );
 a5065a <=( (not A199)  and  A166 );
 a5066a <=( (not A167)  and  a5065a );
 a5067a <=( a5066a  and  a5061a );
 a5071a <=( A298  and  A203 );
 a5072a <=( (not A200)  and  a5071a );
 a5076a <=( (not A302)  and  A301 );
 a5077a <=( A299  and  a5076a );
 a5078a <=( a5077a  and  a5072a );
 a5081a <=( A168  and  A170 );
 a5085a <=( (not A199)  and  A166 );
 a5086a <=( (not A167)  and  a5085a );
 a5087a <=( a5086a  and  a5081a );
 a5091a <=( A298  and  A203 );
 a5092a <=( (not A200)  and  a5091a );
 a5096a <=( A302  and  (not A301) );
 a5097a <=( (not A299)  and  a5096a );
 a5098a <=( a5097a  and  a5092a );
 a5101a <=( A168  and  A170 );
 a5105a <=( (not A199)  and  A166 );
 a5106a <=( (not A167)  and  a5105a );
 a5107a <=( a5106a  and  a5101a );
 a5111a <=( (not A298)  and  A203 );
 a5112a <=( (not A200)  and  a5111a );
 a5116a <=( A302  and  (not A301) );
 a5117a <=( A299  and  a5116a );
 a5118a <=( a5117a  and  a5112a );
 a5121a <=( A168  and  A170 );
 a5125a <=( (not A199)  and  A166 );
 a5126a <=( (not A167)  and  a5125a );
 a5127a <=( a5126a  and  a5121a );
 a5131a <=( (not A298)  and  A203 );
 a5132a <=( (not A200)  and  a5131a );
 a5136a <=( (not A302)  and  A301 );
 a5137a <=( (not A299)  and  a5136a );
 a5138a <=( a5137a  and  a5132a );
 a5141a <=( A168  and  A169 );
 a5145a <=( (not A199)  and  A166 );
 a5146a <=( (not A167)  and  a5145a );
 a5147a <=( a5146a  and  a5141a );
 a5151a <=( A298  and  (not A202) );
 a5152a <=( (not A200)  and  a5151a );
 a5156a <=( (not A302)  and  A301 );
 a5157a <=( A299  and  a5156a );
 a5158a <=( a5157a  and  a5152a );
 a5161a <=( A168  and  A169 );
 a5165a <=( (not A199)  and  A166 );
 a5166a <=( (not A167)  and  a5165a );
 a5167a <=( a5166a  and  a5161a );
 a5171a <=( A298  and  (not A202) );
 a5172a <=( (not A200)  and  a5171a );
 a5176a <=( A302  and  (not A301) );
 a5177a <=( (not A299)  and  a5176a );
 a5178a <=( a5177a  and  a5172a );
 a5181a <=( A168  and  A169 );
 a5185a <=( (not A199)  and  A166 );
 a5186a <=( (not A167)  and  a5185a );
 a5187a <=( a5186a  and  a5181a );
 a5191a <=( (not A298)  and  (not A202) );
 a5192a <=( (not A200)  and  a5191a );
 a5196a <=( A302  and  (not A301) );
 a5197a <=( A299  and  a5196a );
 a5198a <=( a5197a  and  a5192a );
 a5201a <=( A168  and  A169 );
 a5205a <=( (not A199)  and  A166 );
 a5206a <=( (not A167)  and  a5205a );
 a5207a <=( a5206a  and  a5201a );
 a5211a <=( (not A298)  and  (not A202) );
 a5212a <=( (not A200)  and  a5211a );
 a5216a <=( (not A302)  and  A301 );
 a5217a <=( (not A299)  and  a5216a );
 a5218a <=( a5217a  and  a5212a );
 a5221a <=( A168  and  A169 );
 a5225a <=( (not A199)  and  A166 );
 a5226a <=( (not A167)  and  a5225a );
 a5227a <=( a5226a  and  a5221a );
 a5231a <=( A298  and  A203 );
 a5232a <=( (not A200)  and  a5231a );
 a5236a <=( (not A302)  and  A301 );
 a5237a <=( A299  and  a5236a );
 a5238a <=( a5237a  and  a5232a );
 a5241a <=( A168  and  A169 );
 a5245a <=( (not A199)  and  A166 );
 a5246a <=( (not A167)  and  a5245a );
 a5247a <=( a5246a  and  a5241a );
 a5251a <=( A298  and  A203 );
 a5252a <=( (not A200)  and  a5251a );
 a5256a <=( A302  and  (not A301) );
 a5257a <=( (not A299)  and  a5256a );
 a5258a <=( a5257a  and  a5252a );
 a5261a <=( A168  and  A169 );
 a5265a <=( (not A199)  and  A166 );
 a5266a <=( (not A167)  and  a5265a );
 a5267a <=( a5266a  and  a5261a );
 a5271a <=( (not A298)  and  A203 );
 a5272a <=( (not A200)  and  a5271a );
 a5276a <=( A302  and  (not A301) );
 a5277a <=( A299  and  a5276a );
 a5278a <=( a5277a  and  a5272a );
 a5281a <=( A168  and  A169 );
 a5285a <=( (not A199)  and  A166 );
 a5286a <=( (not A167)  and  a5285a );
 a5287a <=( a5286a  and  a5281a );
 a5291a <=( (not A298)  and  A203 );
 a5292a <=( (not A200)  and  a5291a );
 a5296a <=( (not A302)  and  A301 );
 a5297a <=( (not A299)  and  a5296a );
 a5298a <=( a5297a  and  a5292a );
 a5301a <=( (not A169)  and  (not A170) );
 a5305a <=( A200  and  A199 );
 a5306a <=( (not A167)  and  a5305a );
 a5307a <=( a5306a  and  a5301a );
 a5311a <=( A298  and  (not A203) );
 a5312a <=( A202  and  a5311a );
 a5316a <=( (not A302)  and  A301 );
 a5317a <=( A299  and  a5316a );
 a5318a <=( a5317a  and  a5312a );
 a5321a <=( (not A169)  and  (not A170) );
 a5325a <=( A200  and  A199 );
 a5326a <=( (not A167)  and  a5325a );
 a5327a <=( a5326a  and  a5321a );
 a5331a <=( A298  and  (not A203) );
 a5332a <=( A202  and  a5331a );
 a5336a <=( A302  and  (not A301) );
 a5337a <=( (not A299)  and  a5336a );
 a5338a <=( a5337a  and  a5332a );
 a5341a <=( (not A169)  and  (not A170) );
 a5345a <=( A200  and  A199 );
 a5346a <=( (not A167)  and  a5345a );
 a5347a <=( a5346a  and  a5341a );
 a5351a <=( (not A298)  and  (not A203) );
 a5352a <=( A202  and  a5351a );
 a5356a <=( A302  and  (not A301) );
 a5357a <=( A299  and  a5356a );
 a5358a <=( a5357a  and  a5352a );
 a5361a <=( (not A169)  and  (not A170) );
 a5365a <=( A200  and  A199 );
 a5366a <=( (not A167)  and  a5365a );
 a5367a <=( a5366a  and  a5361a );
 a5371a <=( (not A298)  and  (not A203) );
 a5372a <=( A202  and  a5371a );
 a5376a <=( (not A302)  and  A301 );
 a5377a <=( (not A299)  and  a5376a );
 a5378a <=( a5377a  and  a5372a );
 a5381a <=( (not A169)  and  (not A170) );
 a5385a <=( A200  and  (not A199) );
 a5386a <=( (not A167)  and  a5385a );
 a5387a <=( a5386a  and  a5381a );
 a5391a <=( A298  and  A203 );
 a5392a <=( (not A202)  and  a5391a );
 a5396a <=( (not A302)  and  A301 );
 a5397a <=( A299  and  a5396a );
 a5398a <=( a5397a  and  a5392a );
 a5401a <=( (not A169)  and  (not A170) );
 a5405a <=( A200  and  (not A199) );
 a5406a <=( (not A167)  and  a5405a );
 a5407a <=( a5406a  and  a5401a );
 a5411a <=( A298  and  A203 );
 a5412a <=( (not A202)  and  a5411a );
 a5416a <=( A302  and  (not A301) );
 a5417a <=( (not A299)  and  a5416a );
 a5418a <=( a5417a  and  a5412a );
 a5421a <=( (not A169)  and  (not A170) );
 a5425a <=( A200  and  (not A199) );
 a5426a <=( (not A167)  and  a5425a );
 a5427a <=( a5426a  and  a5421a );
 a5431a <=( (not A298)  and  A203 );
 a5432a <=( (not A202)  and  a5431a );
 a5436a <=( A302  and  (not A301) );
 a5437a <=( A299  and  a5436a );
 a5438a <=( a5437a  and  a5432a );
 a5441a <=( (not A169)  and  (not A170) );
 a5445a <=( A200  and  (not A199) );
 a5446a <=( (not A167)  and  a5445a );
 a5447a <=( a5446a  and  a5441a );
 a5451a <=( (not A298)  and  A203 );
 a5452a <=( (not A202)  and  a5451a );
 a5456a <=( (not A302)  and  A301 );
 a5457a <=( (not A299)  and  a5456a );
 a5458a <=( a5457a  and  a5452a );
 a5461a <=( (not A169)  and  (not A170) );
 a5465a <=( (not A200)  and  A199 );
 a5466a <=( (not A167)  and  a5465a );
 a5467a <=( a5466a  and  a5461a );
 a5471a <=( A298  and  A203 );
 a5472a <=( (not A202)  and  a5471a );
 a5476a <=( (not A302)  and  A301 );
 a5477a <=( A299  and  a5476a );
 a5478a <=( a5477a  and  a5472a );
 a5481a <=( (not A169)  and  (not A170) );
 a5485a <=( (not A200)  and  A199 );
 a5486a <=( (not A167)  and  a5485a );
 a5487a <=( a5486a  and  a5481a );
 a5491a <=( A298  and  A203 );
 a5492a <=( (not A202)  and  a5491a );
 a5496a <=( A302  and  (not A301) );
 a5497a <=( (not A299)  and  a5496a );
 a5498a <=( a5497a  and  a5492a );
 a5501a <=( (not A169)  and  (not A170) );
 a5505a <=( (not A200)  and  A199 );
 a5506a <=( (not A167)  and  a5505a );
 a5507a <=( a5506a  and  a5501a );
 a5511a <=( (not A298)  and  A203 );
 a5512a <=( (not A202)  and  a5511a );
 a5516a <=( A302  and  (not A301) );
 a5517a <=( A299  and  a5516a );
 a5518a <=( a5517a  and  a5512a );
 a5521a <=( (not A169)  and  (not A170) );
 a5525a <=( (not A200)  and  A199 );
 a5526a <=( (not A167)  and  a5525a );
 a5527a <=( a5526a  and  a5521a );
 a5531a <=( (not A298)  and  A203 );
 a5532a <=( (not A202)  and  a5531a );
 a5536a <=( (not A302)  and  A301 );
 a5537a <=( (not A299)  and  a5536a );
 a5538a <=( a5537a  and  a5532a );
 a5541a <=( (not A169)  and  (not A170) );
 a5545a <=( (not A200)  and  (not A199) );
 a5546a <=( (not A167)  and  a5545a );
 a5547a <=( a5546a  and  a5541a );
 a5551a <=( A298  and  (not A203) );
 a5552a <=( A202  and  a5551a );
 a5556a <=( (not A302)  and  A301 );
 a5557a <=( A299  and  a5556a );
 a5558a <=( a5557a  and  a5552a );
 a5561a <=( (not A169)  and  (not A170) );
 a5565a <=( (not A200)  and  (not A199) );
 a5566a <=( (not A167)  and  a5565a );
 a5567a <=( a5566a  and  a5561a );
 a5571a <=( A298  and  (not A203) );
 a5572a <=( A202  and  a5571a );
 a5576a <=( A302  and  (not A301) );
 a5577a <=( (not A299)  and  a5576a );
 a5578a <=( a5577a  and  a5572a );
 a5581a <=( (not A169)  and  (not A170) );
 a5585a <=( (not A200)  and  (not A199) );
 a5586a <=( (not A167)  and  a5585a );
 a5587a <=( a5586a  and  a5581a );
 a5591a <=( (not A298)  and  (not A203) );
 a5592a <=( A202  and  a5591a );
 a5596a <=( A302  and  (not A301) );
 a5597a <=( A299  and  a5596a );
 a5598a <=( a5597a  and  a5592a );
 a5601a <=( (not A169)  and  (not A170) );
 a5605a <=( (not A200)  and  (not A199) );
 a5606a <=( (not A167)  and  a5605a );
 a5607a <=( a5606a  and  a5601a );
 a5611a <=( (not A298)  and  (not A203) );
 a5612a <=( A202  and  a5611a );
 a5616a <=( (not A302)  and  A301 );
 a5617a <=( (not A299)  and  a5616a );
 a5618a <=( a5617a  and  a5612a );
 a5622a <=( (not A167)  and  A168 );
 a5623a <=( A170  and  a5622a );
 a5627a <=( A200  and  A199 );
 a5628a <=( A166  and  a5627a );
 a5629a <=( a5628a  and  a5623a );
 a5633a <=( A298  and  (not A202) );
 a5634a <=( (not A201)  and  a5633a );
 a5638a <=( (not A302)  and  A301 );
 a5639a <=( A299  and  a5638a );
 a5640a <=( a5639a  and  a5634a );
 a5644a <=( (not A167)  and  A168 );
 a5645a <=( A170  and  a5644a );
 a5649a <=( A200  and  A199 );
 a5650a <=( A166  and  a5649a );
 a5651a <=( a5650a  and  a5645a );
 a5655a <=( A298  and  (not A202) );
 a5656a <=( (not A201)  and  a5655a );
 a5660a <=( A302  and  (not A301) );
 a5661a <=( (not A299)  and  a5660a );
 a5662a <=( a5661a  and  a5656a );
 a5666a <=( (not A167)  and  A168 );
 a5667a <=( A170  and  a5666a );
 a5671a <=( A200  and  A199 );
 a5672a <=( A166  and  a5671a );
 a5673a <=( a5672a  and  a5667a );
 a5677a <=( (not A298)  and  (not A202) );
 a5678a <=( (not A201)  and  a5677a );
 a5682a <=( A302  and  (not A301) );
 a5683a <=( A299  and  a5682a );
 a5684a <=( a5683a  and  a5678a );
 a5688a <=( (not A167)  and  A168 );
 a5689a <=( A170  and  a5688a );
 a5693a <=( A200  and  A199 );
 a5694a <=( A166  and  a5693a );
 a5695a <=( a5694a  and  a5689a );
 a5699a <=( (not A298)  and  (not A202) );
 a5700a <=( (not A201)  and  a5699a );
 a5704a <=( (not A302)  and  A301 );
 a5705a <=( (not A299)  and  a5704a );
 a5706a <=( a5705a  and  a5700a );
 a5710a <=( (not A167)  and  A168 );
 a5711a <=( A170  and  a5710a );
 a5715a <=( A200  and  A199 );
 a5716a <=( A166  and  a5715a );
 a5717a <=( a5716a  and  a5711a );
 a5721a <=( A298  and  A203 );
 a5722a <=( (not A201)  and  a5721a );
 a5726a <=( (not A302)  and  A301 );
 a5727a <=( A299  and  a5726a );
 a5728a <=( a5727a  and  a5722a );
 a5732a <=( (not A167)  and  A168 );
 a5733a <=( A170  and  a5732a );
 a5737a <=( A200  and  A199 );
 a5738a <=( A166  and  a5737a );
 a5739a <=( a5738a  and  a5733a );
 a5743a <=( A298  and  A203 );
 a5744a <=( (not A201)  and  a5743a );
 a5748a <=( A302  and  (not A301) );
 a5749a <=( (not A299)  and  a5748a );
 a5750a <=( a5749a  and  a5744a );
 a5754a <=( (not A167)  and  A168 );
 a5755a <=( A170  and  a5754a );
 a5759a <=( A200  and  A199 );
 a5760a <=( A166  and  a5759a );
 a5761a <=( a5760a  and  a5755a );
 a5765a <=( (not A298)  and  A203 );
 a5766a <=( (not A201)  and  a5765a );
 a5770a <=( A302  and  (not A301) );
 a5771a <=( A299  and  a5770a );
 a5772a <=( a5771a  and  a5766a );
 a5776a <=( (not A167)  and  A168 );
 a5777a <=( A170  and  a5776a );
 a5781a <=( A200  and  A199 );
 a5782a <=( A166  and  a5781a );
 a5783a <=( a5782a  and  a5777a );
 a5787a <=( (not A298)  and  A203 );
 a5788a <=( (not A201)  and  a5787a );
 a5792a <=( (not A302)  and  A301 );
 a5793a <=( (not A299)  and  a5792a );
 a5794a <=( a5793a  and  a5788a );
 a5798a <=( (not A167)  and  A168 );
 a5799a <=( A170  and  a5798a );
 a5803a <=( A200  and  (not A199) );
 a5804a <=( A166  and  a5803a );
 a5805a <=( a5804a  and  a5799a );
 a5809a <=( A298  and  A202 );
 a5810a <=( (not A201)  and  a5809a );
 a5814a <=( (not A302)  and  A301 );
 a5815a <=( A299  and  a5814a );
 a5816a <=( a5815a  and  a5810a );
 a5820a <=( (not A167)  and  A168 );
 a5821a <=( A170  and  a5820a );
 a5825a <=( A200  and  (not A199) );
 a5826a <=( A166  and  a5825a );
 a5827a <=( a5826a  and  a5821a );
 a5831a <=( A298  and  A202 );
 a5832a <=( (not A201)  and  a5831a );
 a5836a <=( A302  and  (not A301) );
 a5837a <=( (not A299)  and  a5836a );
 a5838a <=( a5837a  and  a5832a );
 a5842a <=( (not A167)  and  A168 );
 a5843a <=( A170  and  a5842a );
 a5847a <=( A200  and  (not A199) );
 a5848a <=( A166  and  a5847a );
 a5849a <=( a5848a  and  a5843a );
 a5853a <=( (not A298)  and  A202 );
 a5854a <=( (not A201)  and  a5853a );
 a5858a <=( A302  and  (not A301) );
 a5859a <=( A299  and  a5858a );
 a5860a <=( a5859a  and  a5854a );
 a5864a <=( (not A167)  and  A168 );
 a5865a <=( A170  and  a5864a );
 a5869a <=( A200  and  (not A199) );
 a5870a <=( A166  and  a5869a );
 a5871a <=( a5870a  and  a5865a );
 a5875a <=( (not A298)  and  A202 );
 a5876a <=( (not A201)  and  a5875a );
 a5880a <=( (not A302)  and  A301 );
 a5881a <=( (not A299)  and  a5880a );
 a5882a <=( a5881a  and  a5876a );
 a5886a <=( (not A167)  and  A168 );
 a5887a <=( A170  and  a5886a );
 a5891a <=( A200  and  (not A199) );
 a5892a <=( A166  and  a5891a );
 a5893a <=( a5892a  and  a5887a );
 a5897a <=( A298  and  (not A203) );
 a5898a <=( (not A201)  and  a5897a );
 a5902a <=( (not A302)  and  A301 );
 a5903a <=( A299  and  a5902a );
 a5904a <=( a5903a  and  a5898a );
 a5908a <=( (not A167)  and  A168 );
 a5909a <=( A170  and  a5908a );
 a5913a <=( A200  and  (not A199) );
 a5914a <=( A166  and  a5913a );
 a5915a <=( a5914a  and  a5909a );
 a5919a <=( A298  and  (not A203) );
 a5920a <=( (not A201)  and  a5919a );
 a5924a <=( A302  and  (not A301) );
 a5925a <=( (not A299)  and  a5924a );
 a5926a <=( a5925a  and  a5920a );
 a5930a <=( (not A167)  and  A168 );
 a5931a <=( A170  and  a5930a );
 a5935a <=( A200  and  (not A199) );
 a5936a <=( A166  and  a5935a );
 a5937a <=( a5936a  and  a5931a );
 a5941a <=( (not A298)  and  (not A203) );
 a5942a <=( (not A201)  and  a5941a );
 a5946a <=( A302  and  (not A301) );
 a5947a <=( A299  and  a5946a );
 a5948a <=( a5947a  and  a5942a );
 a5952a <=( (not A167)  and  A168 );
 a5953a <=( A170  and  a5952a );
 a5957a <=( A200  and  (not A199) );
 a5958a <=( A166  and  a5957a );
 a5959a <=( a5958a  and  a5953a );
 a5963a <=( (not A298)  and  (not A203) );
 a5964a <=( (not A201)  and  a5963a );
 a5968a <=( (not A302)  and  A301 );
 a5969a <=( (not A299)  and  a5968a );
 a5970a <=( a5969a  and  a5964a );
 a5974a <=( (not A167)  and  A168 );
 a5975a <=( A170  and  a5974a );
 a5979a <=( (not A200)  and  A199 );
 a5980a <=( A166  and  a5979a );
 a5981a <=( a5980a  and  a5975a );
 a5985a <=( A298  and  A202 );
 a5986a <=( (not A201)  and  a5985a );
 a5990a <=( (not A302)  and  A301 );
 a5991a <=( A299  and  a5990a );
 a5992a <=( a5991a  and  a5986a );
 a5996a <=( (not A167)  and  A168 );
 a5997a <=( A170  and  a5996a );
 a6001a <=( (not A200)  and  A199 );
 a6002a <=( A166  and  a6001a );
 a6003a <=( a6002a  and  a5997a );
 a6007a <=( A298  and  A202 );
 a6008a <=( (not A201)  and  a6007a );
 a6012a <=( A302  and  (not A301) );
 a6013a <=( (not A299)  and  a6012a );
 a6014a <=( a6013a  and  a6008a );
 a6018a <=( (not A167)  and  A168 );
 a6019a <=( A170  and  a6018a );
 a6023a <=( (not A200)  and  A199 );
 a6024a <=( A166  and  a6023a );
 a6025a <=( a6024a  and  a6019a );
 a6029a <=( (not A298)  and  A202 );
 a6030a <=( (not A201)  and  a6029a );
 a6034a <=( A302  and  (not A301) );
 a6035a <=( A299  and  a6034a );
 a6036a <=( a6035a  and  a6030a );
 a6040a <=( (not A167)  and  A168 );
 a6041a <=( A170  and  a6040a );
 a6045a <=( (not A200)  and  A199 );
 a6046a <=( A166  and  a6045a );
 a6047a <=( a6046a  and  a6041a );
 a6051a <=( (not A298)  and  A202 );
 a6052a <=( (not A201)  and  a6051a );
 a6056a <=( (not A302)  and  A301 );
 a6057a <=( (not A299)  and  a6056a );
 a6058a <=( a6057a  and  a6052a );
 a6062a <=( (not A167)  and  A168 );
 a6063a <=( A170  and  a6062a );
 a6067a <=( (not A200)  and  A199 );
 a6068a <=( A166  and  a6067a );
 a6069a <=( a6068a  and  a6063a );
 a6073a <=( A298  and  (not A203) );
 a6074a <=( (not A201)  and  a6073a );
 a6078a <=( (not A302)  and  A301 );
 a6079a <=( A299  and  a6078a );
 a6080a <=( a6079a  and  a6074a );
 a6084a <=( (not A167)  and  A168 );
 a6085a <=( A170  and  a6084a );
 a6089a <=( (not A200)  and  A199 );
 a6090a <=( A166  and  a6089a );
 a6091a <=( a6090a  and  a6085a );
 a6095a <=( A298  and  (not A203) );
 a6096a <=( (not A201)  and  a6095a );
 a6100a <=( A302  and  (not A301) );
 a6101a <=( (not A299)  and  a6100a );
 a6102a <=( a6101a  and  a6096a );
 a6106a <=( (not A167)  and  A168 );
 a6107a <=( A170  and  a6106a );
 a6111a <=( (not A200)  and  A199 );
 a6112a <=( A166  and  a6111a );
 a6113a <=( a6112a  and  a6107a );
 a6117a <=( (not A298)  and  (not A203) );
 a6118a <=( (not A201)  and  a6117a );
 a6122a <=( A302  and  (not A301) );
 a6123a <=( A299  and  a6122a );
 a6124a <=( a6123a  and  a6118a );
 a6128a <=( (not A167)  and  A168 );
 a6129a <=( A170  and  a6128a );
 a6133a <=( (not A200)  and  A199 );
 a6134a <=( A166  and  a6133a );
 a6135a <=( a6134a  and  a6129a );
 a6139a <=( (not A298)  and  (not A203) );
 a6140a <=( (not A201)  and  a6139a );
 a6144a <=( (not A302)  and  A301 );
 a6145a <=( (not A299)  and  a6144a );
 a6146a <=( a6145a  and  a6140a );
 a6150a <=( (not A167)  and  A168 );
 a6151a <=( A169  and  a6150a );
 a6155a <=( A200  and  A199 );
 a6156a <=( A166  and  a6155a );
 a6157a <=( a6156a  and  a6151a );
 a6161a <=( A298  and  (not A202) );
 a6162a <=( (not A201)  and  a6161a );
 a6166a <=( (not A302)  and  A301 );
 a6167a <=( A299  and  a6166a );
 a6168a <=( a6167a  and  a6162a );
 a6172a <=( (not A167)  and  A168 );
 a6173a <=( A169  and  a6172a );
 a6177a <=( A200  and  A199 );
 a6178a <=( A166  and  a6177a );
 a6179a <=( a6178a  and  a6173a );
 a6183a <=( A298  and  (not A202) );
 a6184a <=( (not A201)  and  a6183a );
 a6188a <=( A302  and  (not A301) );
 a6189a <=( (not A299)  and  a6188a );
 a6190a <=( a6189a  and  a6184a );
 a6194a <=( (not A167)  and  A168 );
 a6195a <=( A169  and  a6194a );
 a6199a <=( A200  and  A199 );
 a6200a <=( A166  and  a6199a );
 a6201a <=( a6200a  and  a6195a );
 a6205a <=( (not A298)  and  (not A202) );
 a6206a <=( (not A201)  and  a6205a );
 a6210a <=( A302  and  (not A301) );
 a6211a <=( A299  and  a6210a );
 a6212a <=( a6211a  and  a6206a );
 a6216a <=( (not A167)  and  A168 );
 a6217a <=( A169  and  a6216a );
 a6221a <=( A200  and  A199 );
 a6222a <=( A166  and  a6221a );
 a6223a <=( a6222a  and  a6217a );
 a6227a <=( (not A298)  and  (not A202) );
 a6228a <=( (not A201)  and  a6227a );
 a6232a <=( (not A302)  and  A301 );
 a6233a <=( (not A299)  and  a6232a );
 a6234a <=( a6233a  and  a6228a );
 a6238a <=( (not A167)  and  A168 );
 a6239a <=( A169  and  a6238a );
 a6243a <=( A200  and  A199 );
 a6244a <=( A166  and  a6243a );
 a6245a <=( a6244a  and  a6239a );
 a6249a <=( A298  and  A203 );
 a6250a <=( (not A201)  and  a6249a );
 a6254a <=( (not A302)  and  A301 );
 a6255a <=( A299  and  a6254a );
 a6256a <=( a6255a  and  a6250a );
 a6260a <=( (not A167)  and  A168 );
 a6261a <=( A169  and  a6260a );
 a6265a <=( A200  and  A199 );
 a6266a <=( A166  and  a6265a );
 a6267a <=( a6266a  and  a6261a );
 a6271a <=( A298  and  A203 );
 a6272a <=( (not A201)  and  a6271a );
 a6276a <=( A302  and  (not A301) );
 a6277a <=( (not A299)  and  a6276a );
 a6278a <=( a6277a  and  a6272a );
 a6282a <=( (not A167)  and  A168 );
 a6283a <=( A169  and  a6282a );
 a6287a <=( A200  and  A199 );
 a6288a <=( A166  and  a6287a );
 a6289a <=( a6288a  and  a6283a );
 a6293a <=( (not A298)  and  A203 );
 a6294a <=( (not A201)  and  a6293a );
 a6298a <=( A302  and  (not A301) );
 a6299a <=( A299  and  a6298a );
 a6300a <=( a6299a  and  a6294a );
 a6304a <=( (not A167)  and  A168 );
 a6305a <=( A169  and  a6304a );
 a6309a <=( A200  and  A199 );
 a6310a <=( A166  and  a6309a );
 a6311a <=( a6310a  and  a6305a );
 a6315a <=( (not A298)  and  A203 );
 a6316a <=( (not A201)  and  a6315a );
 a6320a <=( (not A302)  and  A301 );
 a6321a <=( (not A299)  and  a6320a );
 a6322a <=( a6321a  and  a6316a );
 a6326a <=( (not A167)  and  A168 );
 a6327a <=( A169  and  a6326a );
 a6331a <=( A200  and  (not A199) );
 a6332a <=( A166  and  a6331a );
 a6333a <=( a6332a  and  a6327a );
 a6337a <=( A298  and  A202 );
 a6338a <=( (not A201)  and  a6337a );
 a6342a <=( (not A302)  and  A301 );
 a6343a <=( A299  and  a6342a );
 a6344a <=( a6343a  and  a6338a );
 a6348a <=( (not A167)  and  A168 );
 a6349a <=( A169  and  a6348a );
 a6353a <=( A200  and  (not A199) );
 a6354a <=( A166  and  a6353a );
 a6355a <=( a6354a  and  a6349a );
 a6359a <=( A298  and  A202 );
 a6360a <=( (not A201)  and  a6359a );
 a6364a <=( A302  and  (not A301) );
 a6365a <=( (not A299)  and  a6364a );
 a6366a <=( a6365a  and  a6360a );
 a6370a <=( (not A167)  and  A168 );
 a6371a <=( A169  and  a6370a );
 a6375a <=( A200  and  (not A199) );
 a6376a <=( A166  and  a6375a );
 a6377a <=( a6376a  and  a6371a );
 a6381a <=( (not A298)  and  A202 );
 a6382a <=( (not A201)  and  a6381a );
 a6386a <=( A302  and  (not A301) );
 a6387a <=( A299  and  a6386a );
 a6388a <=( a6387a  and  a6382a );
 a6392a <=( (not A167)  and  A168 );
 a6393a <=( A169  and  a6392a );
 a6397a <=( A200  and  (not A199) );
 a6398a <=( A166  and  a6397a );
 a6399a <=( a6398a  and  a6393a );
 a6403a <=( (not A298)  and  A202 );
 a6404a <=( (not A201)  and  a6403a );
 a6408a <=( (not A302)  and  A301 );
 a6409a <=( (not A299)  and  a6408a );
 a6410a <=( a6409a  and  a6404a );
 a6414a <=( (not A167)  and  A168 );
 a6415a <=( A169  and  a6414a );
 a6419a <=( A200  and  (not A199) );
 a6420a <=( A166  and  a6419a );
 a6421a <=( a6420a  and  a6415a );
 a6425a <=( A298  and  (not A203) );
 a6426a <=( (not A201)  and  a6425a );
 a6430a <=( (not A302)  and  A301 );
 a6431a <=( A299  and  a6430a );
 a6432a <=( a6431a  and  a6426a );
 a6436a <=( (not A167)  and  A168 );
 a6437a <=( A169  and  a6436a );
 a6441a <=( A200  and  (not A199) );
 a6442a <=( A166  and  a6441a );
 a6443a <=( a6442a  and  a6437a );
 a6447a <=( A298  and  (not A203) );
 a6448a <=( (not A201)  and  a6447a );
 a6452a <=( A302  and  (not A301) );
 a6453a <=( (not A299)  and  a6452a );
 a6454a <=( a6453a  and  a6448a );
 a6458a <=( (not A167)  and  A168 );
 a6459a <=( A169  and  a6458a );
 a6463a <=( A200  and  (not A199) );
 a6464a <=( A166  and  a6463a );
 a6465a <=( a6464a  and  a6459a );
 a6469a <=( (not A298)  and  (not A203) );
 a6470a <=( (not A201)  and  a6469a );
 a6474a <=( A302  and  (not A301) );
 a6475a <=( A299  and  a6474a );
 a6476a <=( a6475a  and  a6470a );
 a6480a <=( (not A167)  and  A168 );
 a6481a <=( A169  and  a6480a );
 a6485a <=( A200  and  (not A199) );
 a6486a <=( A166  and  a6485a );
 a6487a <=( a6486a  and  a6481a );
 a6491a <=( (not A298)  and  (not A203) );
 a6492a <=( (not A201)  and  a6491a );
 a6496a <=( (not A302)  and  A301 );
 a6497a <=( (not A299)  and  a6496a );
 a6498a <=( a6497a  and  a6492a );
 a6502a <=( (not A167)  and  A168 );
 a6503a <=( A169  and  a6502a );
 a6507a <=( (not A200)  and  A199 );
 a6508a <=( A166  and  a6507a );
 a6509a <=( a6508a  and  a6503a );
 a6513a <=( A298  and  A202 );
 a6514a <=( (not A201)  and  a6513a );
 a6518a <=( (not A302)  and  A301 );
 a6519a <=( A299  and  a6518a );
 a6520a <=( a6519a  and  a6514a );
 a6524a <=( (not A167)  and  A168 );
 a6525a <=( A169  and  a6524a );
 a6529a <=( (not A200)  and  A199 );
 a6530a <=( A166  and  a6529a );
 a6531a <=( a6530a  and  a6525a );
 a6535a <=( A298  and  A202 );
 a6536a <=( (not A201)  and  a6535a );
 a6540a <=( A302  and  (not A301) );
 a6541a <=( (not A299)  and  a6540a );
 a6542a <=( a6541a  and  a6536a );
 a6546a <=( (not A167)  and  A168 );
 a6547a <=( A169  and  a6546a );
 a6551a <=( (not A200)  and  A199 );
 a6552a <=( A166  and  a6551a );
 a6553a <=( a6552a  and  a6547a );
 a6557a <=( (not A298)  and  A202 );
 a6558a <=( (not A201)  and  a6557a );
 a6562a <=( A302  and  (not A301) );
 a6563a <=( A299  and  a6562a );
 a6564a <=( a6563a  and  a6558a );
 a6568a <=( (not A167)  and  A168 );
 a6569a <=( A169  and  a6568a );
 a6573a <=( (not A200)  and  A199 );
 a6574a <=( A166  and  a6573a );
 a6575a <=( a6574a  and  a6569a );
 a6579a <=( (not A298)  and  A202 );
 a6580a <=( (not A201)  and  a6579a );
 a6584a <=( (not A302)  and  A301 );
 a6585a <=( (not A299)  and  a6584a );
 a6586a <=( a6585a  and  a6580a );
 a6590a <=( (not A167)  and  A168 );
 a6591a <=( A169  and  a6590a );
 a6595a <=( (not A200)  and  A199 );
 a6596a <=( A166  and  a6595a );
 a6597a <=( a6596a  and  a6591a );
 a6601a <=( A298  and  (not A203) );
 a6602a <=( (not A201)  and  a6601a );
 a6606a <=( (not A302)  and  A301 );
 a6607a <=( A299  and  a6606a );
 a6608a <=( a6607a  and  a6602a );
 a6612a <=( (not A167)  and  A168 );
 a6613a <=( A169  and  a6612a );
 a6617a <=( (not A200)  and  A199 );
 a6618a <=( A166  and  a6617a );
 a6619a <=( a6618a  and  a6613a );
 a6623a <=( A298  and  (not A203) );
 a6624a <=( (not A201)  and  a6623a );
 a6628a <=( A302  and  (not A301) );
 a6629a <=( (not A299)  and  a6628a );
 a6630a <=( a6629a  and  a6624a );
 a6634a <=( (not A167)  and  A168 );
 a6635a <=( A169  and  a6634a );
 a6639a <=( (not A200)  and  A199 );
 a6640a <=( A166  and  a6639a );
 a6641a <=( a6640a  and  a6635a );
 a6645a <=( (not A298)  and  (not A203) );
 a6646a <=( (not A201)  and  a6645a );
 a6650a <=( A302  and  (not A301) );
 a6651a <=( A299  and  a6650a );
 a6652a <=( a6651a  and  a6646a );
 a6656a <=( (not A167)  and  A168 );
 a6657a <=( A169  and  a6656a );
 a6661a <=( (not A200)  and  A199 );
 a6662a <=( A166  and  a6661a );
 a6663a <=( a6662a  and  a6657a );
 a6667a <=( (not A298)  and  (not A203) );
 a6668a <=( (not A201)  and  a6667a );
 a6672a <=( (not A302)  and  A301 );
 a6673a <=( (not A299)  and  a6672a );
 a6674a <=( a6673a  and  a6668a );


end x25_18x_behav;
