Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_7x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A108: buffer std_logic
);
end x25_7x;

architecture x25_7x_behav of x25_7x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a460a,a461a,a464a,a467a,a468a,a469a,a473a,a474a,a477a,a480a,a481a,a482a,a483a,a487a,a488a,a491a,a494a,a495a,a496a,a500a,a501a,a504a,a507a,a508a,a509a,a510a,a511a,a515a,a516a,a519a,a522a,a523a,a524a,a528a,a529a,a532a,a535a,a536a,a537a,a538a,a542a,a543a,a546a,a549a,a550a,a551a,a554a,a557a,a558a,a561a,a564a,a565a,a566a,a567a,a568a,a569a,a573a,a574a,a577a,a580a,a581a,a582a,a586a,a587a,a590a,a593a,a594a,a595a,a596a,a600a,a601a,a604a,a607a,a608a,a609a,a613a,a614a,a617a,a620a,a621a,a622a,a623a,a624a,a628a,a629a,a632a,a635a,a636a,a637a,a641a,a642a,a645a,a648a,a649a,a650a,a651a,a655a,a656a,a659a,a662a,a663a,a664a,a667a,a670a,a671a,a674a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a687a,a688a,a691a,a694a,a695a,a696a,a700a,a701a,a704a,a707a,a708a,a709a,a710a,a714a,a715a,a718a,a721a,a722a,a723a,a727a,a728a,a731a,a734a,a735a,a736a,a737a,a738a,a742a,a743a,a746a,a749a,a750a,a751a,a755a,a756a,a759a,a762a,a763a,a764a,a765a,a769a,a770a,a773a,a776a,a777a,a778a,a781a,a784a,a785a,a788a,a791a,a792a,a793a,a794a,a795a,a796a,a800a,a801a,a804a,a807a,a808a,a809a,a813a,a814a,a817a,a820a,a821a,a822a,a823a,a827a,a828a,a831a,a834a,a835a,a836a,a840a,a841a,a844a,a847a,a848a,a849a,a850a,a851a,a855a,a856a,a859a,a862a,a863a,a864a,a868a,a869a,a872a,a875a,a876a,a877a,a878a,a882a,a883a,a886a,a889a,a890a,a891a,a894a,a897a,a898a,a901a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a915a,a916a,a919a,a922a,a923a,a924a,a928a,a929a,a932a,a935a,a936a,a937a,a938a,a942a,a943a,a946a,a949a,a950a,a951a,a955a,a956a,a959a,a962a,a963a,a964a,a965a,a966a,a970a,a971a,a974a,a977a,a978a,a979a,a983a,a984a,a987a,a990a,a991a,a992a,a993a,a997a,a998a,a1001a,a1004a,a1005a,a1006a,a1009a,a1012a,a1013a,a1016a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1028a,a1029a,a1032a,a1035a,a1036a,a1037a,a1041a,a1042a,a1045a,a1048a,a1049a,a1050a,a1051a,a1055a,a1056a,a1059a,a1062a,a1063a,a1064a,a1068a,a1069a,a1072a,a1075a,a1076a,a1077a,a1078a,a1079a,a1083a,a1084a,a1087a,a1090a,a1091a,a1092a,a1096a,a1097a,a1100a,a1103a,a1104a,a1105a,a1106a,a1110a,a1111a,a1114a,a1117a,a1118a,a1119a,a1122a,a1125a,a1126a,a1129a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1142a,a1143a,a1146a,a1149a,a1150a,a1151a,a1155a,a1156a,a1159a,a1162a,a1163a,a1164a,a1165a,a1169a,a1170a,a1173a,a1176a,a1177a,a1178a,a1182a,a1183a,a1186a,a1189a,a1190a,a1191a,a1192a,a1193a,a1197a,a1198a,a1201a,a1204a,a1205a,a1206a,a1210a,a1211a,a1214a,a1217a,a1218a,a1219a,a1220a,a1224a,a1225a,a1228a,a1231a,a1232a,a1233a,a1236a,a1239a,a1240a,a1243a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1255a,a1256a,a1259a,a1262a,a1263a,a1264a,a1268a,a1269a,a1272a,a1275a,a1276a,a1277a,a1278a,a1282a,a1283a,a1286a,a1289a,a1290a,a1291a,a1295a,a1296a,a1299a,a1302a,a1303a,a1304a,a1305a,a1306a,a1310a,a1311a,a1314a,a1317a,a1318a,a1319a,a1323a,a1324a,a1327a,a1330a,a1331a,a1332a,a1333a,a1337a,a1338a,a1341a,a1344a,a1345a,a1346a,a1349a,a1352a,a1353a,a1356a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1369a,a1373a,a1374a,a1377a,a1381a,a1382a,a1386a,a1387a,a1391a,a1392a,a1396a,a1397a,a1401a,a1402a,a1406a,a1407a,a1411a,a1412a,a1416a,a1417a,a1421a,a1422a,a1426a,a1427a,a1431a,a1432a,a1436a,a1437a,a1441a,a1442a,a1446a,a1447a,a1450a,a1453a,a1454a,a1458a,a1459a,a1462a,a1465a,a1466a,a1470a,a1471a,a1474a,a1477a,a1478a,a1482a,a1483a,a1486a,a1489a,a1490a,a1493a,a1496a,a1497a,a1500a,a1503a,a1504a,a1507a,a1510a,a1511a,a1514a,a1517a,a1518a,a1521a,a1524a,a1525a,a1528a,a1531a,a1532a,a1535a,a1538a,a1539a,a1542a,a1545a,a1546a,a1549a,a1552a,a1553a,a1556a,a1559a,a1560a,a1563a,a1566a,a1567a,a1570a,a1573a,a1574a,a1577a,a1580a,a1581a,a1584a,a1587a,a1588a,a1591a,a1594a,a1595a,a1598a,a1601a,a1602a,a1605a,a1608a,a1609a,a1612a,a1615a,a1616a,a1619a,a1622a,a1623a,a1626a,a1629a,a1630a,a1633a,a1636a,a1637a,a1640a,a1643a,a1644a,a1647a,a1650a,a1651a,a1654a,a1657a,a1658a,a1661a,a1664a,a1665a,a1668a,a1671a,a1672a,a1675a,a1678a,a1679a,a1682a,a1685a,a1686a,a1689a,a1692a,a1693a,a1696a,a1699a,a1700a,a1703a,a1706a,a1707a,a1710a,a1713a,a1714a,a1717a,a1720a,a1721a,a1724a,a1727a,a1728a,a1731a,a1734a,a1735a,a1738a,a1741a,a1742a,a1745a,a1748a,a1749a,a1752a,a1755a,a1756a,a1759a,a1762a,a1763a,a1766a,a1769a,a1770a,a1773a,a1776a,a1777a,a1780a,a1783a,a1784a,a1787a,a1790a,a1791a,a1794a,a1797a,a1798a,a1801a,a1804a,a1805a,a1808a,a1811a,a1812a,a1815a,a1818a,a1819a,a1822a,a1825a,a1826a,a1829a,a1832a,a1833a,a1836a,a1840a,a1841a,a1842a,a1845a,a1848a,a1849a,a1852a,a1856a,a1857a,a1858a,a1861a,a1864a,a1865a,a1868a,a1872a,a1873a,a1874a,a1877a,a1880a,a1881a,a1884a,a1888a,a1889a,a1890a,a1893a,a1897a,a1898a,a1899a,a1902a,a1906a,a1907a,a1908a,a1911a,a1915a,a1916a,a1917a,a1920a,a1924a,a1925a,a1926a,a1929a,a1933a,a1934a,a1935a,a1938a,a1942a,a1943a,a1944a,a1947a,a1951a,a1952a,a1953a,a1956a,a1960a,a1961a,a1962a,a1965a,a1969a,a1970a,a1971a,a1974a,a1978a,a1979a,a1980a,a1983a,a1987a,a1988a,a1989a,a1992a,a1996a,a1997a,a1998a,a2001a,a2005a,a2006a,a2007a,a2010a,a2014a,a2015a,a2016a,a2019a,a2023a,a2024a,a2025a,a2028a,a2032a,a2033a,a2034a,a2037a,a2041a,a2042a,a2043a,a2046a,a2050a,a2051a,a2052a,a2055a,a2059a,a2060a,a2061a,a2064a,a2068a,a2069a,a2070a,a2073a,a2077a,a2078a,a2079a,a2082a,a2086a,a2087a,a2088a,a2091a,a2095a,a2096a,a2097a,a2100a,a2104a,a2105a,a2106a,a2109a,a2113a,a2114a,a2115a,a2118a,a2122a,a2123a,a2124a,a2127a,a2131a,a2132a,a2133a,a2136a,a2140a,a2141a,a2142a,a2145a,a2149a,a2150a,a2151a,a2154a,a2158a,a2159a,a2160a,a2163a,a2167a,a2168a,a2169a,a2172a,a2176a,a2177a,a2178a,a2181a,a2185a,a2186a,a2187a,a2190a,a2194a,a2195a,a2196a,a2199a,a2203a,a2204a,a2205a,a2208a,a2212a,a2213a,a2214a,a2217a,a2221a,a2222a,a2223a,a2226a,a2230a,a2231a,a2232a,a2235a,a2239a,a2240a,a2241a,a2244a,a2248a,a2249a,a2250a,a2253a,a2257a,a2258a,a2259a,a2262a,a2266a,a2267a,a2268a,a2271a,a2275a,a2276a,a2277a,a2280a,a2284a,a2285a,a2286a,a2289a,a2293a,a2294a,a2295a,a2298a,a2302a,a2303a,a2304a,a2307a,a2311a,a2312a,a2313a,a2316a,a2320a,a2321a,a2322a,a2325a,a2329a,a2330a,a2331a,a2334a,a2338a,a2339a,a2340a,a2343a,a2347a,a2348a,a2349a,a2352a,a2356a,a2357a,a2358a,a2361a,a2365a,a2366a,a2367a,a2370a,a2374a,a2375a,a2376a,a2379a,a2383a,a2384a,a2385a,a2388a,a2392a,a2393a,a2394a,a2397a,a2401a,a2402a,a2403a,a2406a,a2410a,a2411a,a2412a,a2415a,a2419a,a2420a,a2421a,a2424a,a2428a,a2429a,a2430a,a2433a,a2437a,a2438a,a2439a,a2442a,a2446a,a2447a,a2448a,a2451a,a2455a,a2456a,a2457a,a2460a,a2464a,a2465a,a2466a,a2469a,a2473a,a2474a,a2475a,a2478a,a2482a,a2483a,a2484a,a2487a,a2491a,a2492a,a2493a,a2496a,a2500a,a2501a,a2502a,a2505a,a2509a,a2510a,a2511a,a2514a,a2518a,a2519a,a2520a,a2523a,a2527a,a2528a,a2529a,a2532a,a2536a,a2537a,a2538a,a2541a,a2545a,a2546a,a2547a,a2550a,a2554a,a2555a,a2556a,a2559a,a2563a,a2564a,a2565a,a2568a,a2572a,a2573a,a2574a,a2577a,a2581a,a2582a,a2583a,a2586a,a2590a,a2591a,a2592a,a2595a,a2599a,a2600a,a2601a,a2604a,a2608a,a2609a,a2610a,a2613a,a2617a,a2618a,a2619a,a2622a,a2626a,a2627a,a2628a,a2631a,a2635a,a2636a,a2637a,a2640a,a2644a,a2645a,a2646a,a2649a,a2653a,a2654a,a2655a,a2658a,a2662a,a2663a,a2664a,a2667a,a2671a,a2672a,a2673a,a2676a,a2680a,a2681a,a2682a,a2685a,a2689a,a2690a,a2691a,a2694a,a2698a,a2699a,a2700a,a2703a,a2707a,a2708a,a2709a,a2712a,a2716a,a2717a,a2718a,a2721a,a2725a,a2726a,a2727a,a2730a,a2734a,a2735a,a2736a,a2739a,a2743a,a2744a,a2745a,a2748a,a2752a,a2753a,a2754a,a2757a,a2761a,a2762a,a2763a,a2766a,a2770a,a2771a,a2772a,a2775a,a2779a,a2780a,a2781a,a2784a,a2788a,a2789a,a2790a,a2793a,a2797a,a2798a,a2799a,a2802a,a2806a,a2807a,a2808a,a2811a,a2815a,a2816a,a2817a,a2820a,a2824a,a2825a,a2826a,a2829a,a2833a,a2834a,a2835a,a2838a,a2842a,a2843a,a2844a,a2847a,a2851a,a2852a,a2853a,a2856a,a2860a,a2861a,a2862a,a2865a,a2869a,a2870a,a2871a,a2874a,a2878a,a2879a,a2880a,a2883a,a2887a,a2888a,a2889a,a2892a,a2896a,a2897a,a2898a,a2901a,a2905a,a2906a,a2907a,a2910a,a2914a,a2915a,a2916a,a2919a,a2923a,a2924a,a2925a,a2928a,a2932a,a2933a,a2934a,a2937a,a2941a,a2942a,a2943a,a2946a,a2950a,a2951a,a2952a,a2955a,a2959a,a2960a,a2961a,a2964a,a2968a,a2969a,a2970a,a2973a,a2977a,a2978a,a2979a,a2982a,a2986a,a2987a,a2988a,a2991a,a2995a,a2996a,a2997a,a3000a,a3004a,a3005a,a3006a,a3009a,a3013a,a3014a,a3015a,a3018a,a3022a,a3023a,a3024a,a3027a,a3031a,a3032a,a3033a,a3036a,a3040a,a3041a,a3042a,a3045a,a3049a,a3050a,a3051a,a3054a,a3058a,a3059a,a3060a,a3063a,a3067a,a3068a,a3069a,a3072a,a3076a,a3077a,a3078a,a3081a,a3085a,a3086a,a3087a,a3090a,a3094a,a3095a,a3096a,a3099a,a3103a,a3104a,a3105a,a3108a,a3112a,a3113a,a3114a,a3117a,a3121a,a3122a,a3123a,a3126a,a3130a,a3131a,a3132a,a3135a,a3139a,a3140a,a3141a,a3144a,a3148a,a3149a,a3150a,a3153a,a3157a,a3158a,a3159a,a3162a,a3166a,a3167a,a3168a,a3171a,a3175a,a3176a,a3177a,a3180a,a3184a,a3185a,a3186a,a3189a,a3193a,a3194a,a3195a,a3199a,a3200a,a3204a,a3205a,a3206a,a3209a,a3213a,a3214a,a3215a,a3219a,a3220a,a3224a,a3225a,a3226a,a3229a,a3233a,a3234a,a3235a,a3239a,a3240a,a3244a,a3245a,a3246a,a3249a,a3253a,a3254a,a3255a,a3259a,a3260a,a3264a,a3265a,a3266a,a3269a,a3273a,a3274a,a3275a,a3279a,a3280a,a3284a,a3285a,a3286a,a3289a,a3293a,a3294a,a3295a,a3299a,a3300a,a3304a,a3305a,a3306a,a3309a,a3313a,a3314a,a3315a,a3319a,a3320a,a3324a,a3325a,a3326a,a3329a,a3333a,a3334a,a3335a,a3339a,a3340a,a3344a,a3345a,a3346a,a3349a,a3353a,a3354a,a3355a,a3359a,a3360a,a3364a,a3365a,a3366a,a3369a,a3373a,a3374a,a3375a,a3379a,a3380a,a3384a,a3385a,a3386a,a3389a,a3393a,a3394a,a3395a,a3399a,a3400a,a3404a,a3405a,a3406a,a3409a,a3413a,a3414a,a3415a,a3419a,a3420a,a3424a,a3425a,a3426a,a3429a,a3433a,a3434a,a3435a,a3439a,a3440a,a3444a,a3445a,a3446a,a3449a,a3453a,a3454a,a3455a,a3459a,a3460a,a3464a,a3465a,a3466a,a3469a,a3473a,a3474a,a3475a,a3479a,a3480a,a3484a,a3485a,a3486a,a3489a,a3493a,a3494a,a3495a,a3499a,a3500a,a3504a,a3505a,a3506a,a3509a,a3513a,a3514a,a3515a,a3519a,a3520a,a3524a,a3525a,a3526a,a3529a,a3533a,a3534a,a3535a,a3539a,a3540a,a3544a,a3545a,a3546a,a3549a,a3553a,a3554a,a3555a,a3559a,a3560a,a3564a,a3565a,a3566a,a3569a,a3573a,a3574a,a3575a,a3579a,a3580a,a3584a,a3585a,a3586a,a3589a,a3593a,a3594a,a3595a,a3599a,a3600a,a3604a,a3605a,a3606a,a3609a,a3613a,a3614a,a3615a,a3619a,a3620a,a3624a,a3625a,a3626a,a3629a,a3633a,a3634a,a3635a,a3639a,a3640a,a3644a,a3645a,a3646a,a3649a,a3653a,a3654a,a3655a,a3659a,a3660a,a3664a,a3665a,a3666a,a3670a,a3671a,a3675a,a3676a,a3677a,a3681a,a3682a,a3686a,a3687a,a3688a,a3692a,a3693a,a3697a,a3698a,a3699a,a3703a,a3704a,a3708a,a3709a,a3710a,a3714a,a3715a,a3719a,a3720a,a3721a,a3725a,a3726a,a3730a,a3731a,a3732a,a3736a,a3737a,a3741a,a3742a,a3743a,a3747a,a3748a,a3752a,a3753a,a3754a,a3758a,a3759a,a3763a,a3764a,a3765a,a3769a,a3770a,a3774a,a3775a,a3776a,a3780a,a3781a,a3785a,a3786a,a3787a,a3791a,a3792a,a3796a,a3797a,a3798a,a3802a,a3803a,a3807a,a3808a,a3809a,a3813a,a3814a,a3818a,a3819a,a3820a,a3824a,a3825a,a3829a,a3830a,a3831a,a3835a,a3836a,a3840a,a3841a,a3842a,a3846a,a3847a,a3851a,a3852a,a3853a,a3857a,a3858a,a3862a,a3863a,a3864a,a3868a,a3869a,a3873a,a3874a,a3875a,a3879a,a3880a,a3884a,a3885a,a3886a,a3890a,a3891a,a3895a,a3896a,a3897a,a3901a,a3902a,a3906a,a3907a,a3908a,a3912a,a3913a,a3917a,a3918a,a3919a,a3923a,a3924a,a3928a,a3929a,a3930a,a3934a,a3935a,a3939a,a3940a,a3941a,a3945a,a3946a,a3950a,a3951a,a3952a,a3956a,a3957a,a3961a,a3962a,a3963a,a3967a,a3968a,a3972a,a3973a,a3974a,a3978a,a3979a,a3983a,a3984a,a3985a,a3989a,a3990a,a3994a,a3995a,a3996a,a4000a,a4001a,a4005a,a4006a,a4007a,a4011a,a4012a,a4016a,a4017a,a4018a,a4022a,a4023a,a4027a,a4028a,a4029a,a4033a,a4034a,a4038a,a4039a,a4040a,a4044a,a4045a,a4049a,a4050a,a4051a,a4055a,a4056a,a4060a,a4061a,a4062a,a4066a,a4067a,a4071a,a4072a,a4073a,a4077a,a4078a,a4082a,a4083a,a4084a,a4088a,a4089a,a4093a,a4094a,a4095a,a4099a,a4100a,a4104a,a4105a,a4106a,a4110a,a4111a,a4115a,a4116a,a4117a,a4121a,a4122a,a4126a,a4127a,a4128a,a4132a,a4133a,a4137a,a4138a,a4139a,a4143a,a4144a,a4148a,a4149a,a4150a,a4154a,a4155a,a4159a,a4160a,a4161a,a4165a,a4166a,a4170a,a4171a,a4172a,a4176a,a4177a,a4181a,a4182a,a4183a,a4187a,a4188a,a4192a,a4193a,a4194a,a4198a,a4199a,a4203a,a4204a,a4205a,a4209a,a4210a,a4214a,a4215a,a4216a,a4220a,a4221a,a4225a,a4226a,a4227a,a4231a,a4232a,a4236a,a4237a,a4238a,a4242a,a4243a,a4247a,a4248a,a4249a,a4253a,a4254a,a4258a,a4259a,a4260a,a4264a,a4265a,a4269a,a4270a,a4271a,a4275a,a4276a,a4280a,a4281a,a4282a,a4286a,a4287a,a4291a,a4292a,a4293a,a4297a,a4298a,a4302a,a4303a,a4304a,a4308a,a4309a,a4313a,a4314a,a4315a,a4319a,a4320a,a4324a,a4325a,a4326a,a4330a,a4331a,a4335a,a4336a,a4337a,a4341a,a4342a,a4346a,a4347a,a4348a,a4352a,a4353a,a4357a,a4358a,a4359a,a4363a,a4364a,a4368a,a4369a,a4370a,a4374a,a4375a,a4379a,a4380a,a4381a,a4385a,a4386a,a4390a,a4391a,a4392a,a4396a,a4397a,a4401a,a4402a,a4403a,a4407a,a4408a,a4412a,a4413a,a4414a,a4418a,a4419a,a4423a,a4424a,a4425a,a4429a,a4430a,a4434a,a4435a,a4436a,a4440a,a4441a,a4445a,a4446a,a4447a,a4451a,a4452a,a4456a,a4457a,a4458a,a4462a,a4463a,a4467a,a4468a,a4469a,a4473a,a4474a,a4478a,a4479a,a4480a,a4484a,a4485a,a4489a,a4490a,a4491a,a4495a,a4496a,a4500a,a4501a,a4502a,a4506a,a4507a,a4511a,a4512a,a4513a,a4517a,a4518a,a4522a,a4523a,a4524a,a4528a,a4529a,a4533a,a4534a,a4535a,a4539a,a4540a,a4544a,a4545a,a4546a,a4550a,a4551a,a4555a,a4556a,a4557a,a4561a,a4562a,a4566a,a4567a,a4568a,a4572a,a4573a,a4577a,a4578a,a4579a,a4583a,a4584a,a4588a,a4589a,a4590a,a4594a,a4595a,a4599a,a4600a,a4601a,a4605a,a4606a,a4610a,a4611a,a4612a,a4616a,a4617a,a4621a,a4622a,a4623a,a4627a,a4628a,a4632a,a4633a,a4634a,a4638a,a4639a,a4643a,a4644a,a4645a,a4649a,a4650a,a4654a,a4655a,a4656a,a4660a,a4661a,a4665a,a4666a,a4667a,a4671a,a4672a,a4676a,a4677a,a4678a,a4682a,a4683a,a4687a,a4688a,a4689a,a4693a,a4694a,a4698a,a4699a,a4700a,a4704a,a4705a,a4709a,a4710a,a4711a,a4715a,a4716a,a4720a,a4721a,a4722a,a4726a,a4727a,a4731a,a4732a,a4733a,a4737a,a4738a,a4742a,a4743a,a4744a,a4748a,a4749a,a4753a,a4754a,a4755a,a4759a,a4760a,a4764a,a4765a,a4766a,a4770a,a4771a,a4775a,a4776a,a4777a,a4781a,a4782a,a4786a,a4787a,a4788a,a4792a,a4793a,a4797a,a4798a,a4799a,a4803a,a4804a,a4808a,a4809a,a4810a,a4814a,a4815a,a4819a,a4820a,a4821a,a4825a,a4826a,a4830a,a4831a,a4832a,a4836a,a4837a,a4841a,a4842a,a4843a,a4847a,a4848a,a4852a,a4853a,a4854a,a4858a,a4859a,a4863a,a4864a,a4865a,a4869a,a4870a,a4874a,a4875a,a4876a,a4880a,a4881a,a4885a,a4886a,a4887a,a4891a,a4892a,a4896a,a4897a,a4898a,a4902a,a4903a,a4907a,a4908a,a4909a,a4913a,a4914a,a4918a,a4919a,a4920a,a4924a,a4925a,a4929a,a4930a,a4931a,a4935a,a4936a,a4940a,a4941a,a4942a,a4946a,a4947a,a4951a,a4952a,a4953a,a4957a,a4958a,a4962a,a4963a,a4964a,a4968a,a4969a,a4973a,a4974a,a4975a,a4979a,a4980a,a4984a,a4985a,a4986a,a4990a,a4991a,a4995a,a4996a,a4997a,a5001a,a5002a,a5006a,a5007a,a5008a,a5012a,a5013a,a5017a,a5018a,a5019a,a5023a,a5024a,a5028a,a5029a,a5030a,a5034a,a5035a,a5039a,a5040a,a5041a,a5045a,a5046a,a5050a,a5051a,a5052a,a5056a,a5057a,a5061a,a5062a,a5063a,a5067a,a5068a,a5072a,a5073a,a5074a,a5078a,a5079a,a5083a,a5084a,a5085a,a5089a,a5090a,a5094a,a5095a,a5096a,a5100a,a5101a,a5105a,a5106a,a5107a,a5111a,a5112a,a5116a,a5117a,a5118a,a5122a,a5123a,a5127a,a5128a,a5129a,a5133a,a5134a,a5138a,a5139a,a5140a,a5144a,a5145a,a5149a,a5150a,a5151a,a5155a,a5156a,a5160a,a5161a,a5162a,a5166a,a5167a,a5171a,a5172a,a5173a,a5177a,a5178a,a5182a,a5183a,a5184a,a5188a,a5189a,a5193a,a5194a,a5195a,a5199a,a5200a,a5204a,a5205a,a5206a,a5210a,a5211a,a5215a,a5216a,a5217a,a5221a,a5222a,a5226a,a5227a,a5228a,a5232a,a5233a,a5237a,a5238a,a5239a,a5243a,a5244a,a5248a,a5249a,a5250a,a5254a,a5255a,a5259a,a5260a,a5261a,a5265a,a5266a,a5270a,a5271a,a5272a,a5276a,a5277a,a5281a,a5282a,a5283a,a5287a,a5288a,a5292a,a5293a,a5294a,a5298a,a5299a,a5303a,a5304a,a5305a,a5309a,a5310a,a5314a,a5315a,a5316a,a5320a,a5321a,a5325a,a5326a,a5327a,a5331a,a5332a,a5336a,a5337a,a5338a,a5342a,a5343a,a5347a,a5348a,a5349a,a5353a,a5354a,a5358a,a5359a,a5360a,a5364a,a5365a,a5369a,a5370a,a5371a,a5375a,a5376a,a5380a,a5381a,a5382a,a5386a,a5387a,a5391a,a5392a,a5393a,a5397a,a5398a,a5402a,a5403a,a5404a,a5408a,a5409a,a5413a,a5414a,a5415a,a5419a,a5420a,a5424a,a5425a,a5426a,a5430a,a5431a,a5435a,a5436a,a5437a,a5441a,a5442a,a5446a,a5447a,a5448a,a5452a,a5453a,a5457a,a5458a,a5459a,a5463a,a5464a,a5468a,a5469a,a5470a,a5474a,a5475a,a5479a,a5480a,a5481a,a5485a,a5486a,a5490a,a5491a,a5492a,a5496a,a5497a,a5501a,a5502a,a5503a,a5507a,a5508a,a5512a,a5513a,a5514a,a5518a,a5519a,a5523a,a5524a,a5525a,a5529a,a5530a,a5534a,a5535a,a5536a,a5540a,a5541a,a5545a,a5546a,a5547a,a5551a,a5552a,a5556a,a5557a,a5558a,a5562a,a5563a,a5567a,a5568a,a5569a,a5573a,a5574a,a5578a,a5579a,a5580a,a5584a,a5585a,a5589a,a5590a,a5591a,a5595a,a5596a,a5600a,a5601a,a5602a,a5606a,a5607a,a5611a,a5612a,a5613a,a5617a,a5618a,a5622a,a5623a,a5624a,a5628a,a5629a,a5633a,a5634a,a5635a,a5639a,a5640a,a5644a,a5645a,a5646a,a5650a,a5651a,a5655a,a5656a,a5657a,a5661a,a5662a,a5666a,a5667a,a5668a,a5672a,a5673a,a5677a,a5678a,a5679a,a5683a,a5684a,a5688a,a5689a,a5690a,a5694a,a5695a,a5699a,a5700a,a5701a,a5705a,a5706a,a5710a,a5711a,a5712a,a5716a,a5717a,a5721a,a5722a,a5723a,a5727a,a5728a,a5732a,a5733a,a5734a,a5738a,a5739a,a5743a,a5744a,a5745a,a5749a,a5750a,a5754a,a5755a,a5756a,a5760a,a5761a,a5765a,a5766a,a5767a,a5771a,a5772a,a5776a,a5777a,a5778a,a5782a,a5783a,a5787a,a5788a,a5789a,a5793a,a5794a,a5798a,a5799a,a5800a,a5804a,a5805a,a5809a,a5810a,a5811a,a5815a,a5816a,a5820a,a5821a,a5822a,a5826a,a5827a,a5831a,a5832a,a5833a,a5837a,a5838a,a5842a,a5843a,a5844a,a5848a,a5849a,a5853a,a5854a,a5855a,a5859a,a5860a,a5864a,a5865a,a5866a,a5870a,a5871a,a5875a,a5876a,a5877a,a5881a,a5882a,a5886a,a5887a,a5888a,a5892a,a5893a,a5897a,a5898a,a5899a,a5903a,a5904a,a5908a,a5909a,a5910a,a5914a,a5915a,a5919a,a5920a,a5921a,a5925a,a5926a,a5930a,a5931a,a5932a,a5936a,a5937a,a5941a,a5942a,a5943a,a5947a,a5948a,a5952a,a5953a,a5954a,a5958a,a5959a,a5963a,a5964a,a5965a,a5969a,a5970a,a5974a,a5975a,a5976a,a5980a,a5981a,a5985a,a5986a,a5987a,a5991a,a5992a,a5996a,a5997a,a5998a,a6002a,a6003a,a6007a,a6008a,a6009a,a6013a,a6014a,a6018a,a6019a,a6020a,a6024a,a6025a,a6029a,a6030a,a6031a,a6035a,a6036a,a6040a,a6041a,a6042a,a6046a,a6047a,a6051a,a6052a,a6053a,a6057a,a6058a,a6062a,a6063a,a6064a,a6068a,a6069a,a6073a,a6074a,a6075a,a6079a,a6080a,a6084a,a6085a,a6086a,a6090a,a6091a,a6095a,a6096a,a6097a,a6101a,a6102a,a6106a,a6107a,a6108a,a6112a,a6113a,a6117a,a6118a,a6119a,a6123a,a6124a,a6128a,a6129a,a6130a,a6134a,a6135a,a6139a,a6140a,a6141a,a6145a,a6146a,a6150a,a6151a,a6152a,a6156a,a6157a,a6161a,a6162a,a6163a,a6167a,a6168a,a6172a,a6173a,a6174a,a6178a,a6179a,a6183a,a6184a,a6185a,a6189a,a6190a,a6194a,a6195a,a6196a,a6200a,a6201a,a6205a,a6206a,a6207a,a6211a,a6212a,a6216a,a6217a,a6218a,a6222a,a6223a,a6227a,a6228a,a6229a,a6233a,a6234a,a6238a,a6239a,a6240a,a6244a,a6245a,a6249a,a6250a,a6251a,a6255a,a6256a,a6260a,a6261a,a6262a,a6266a,a6267a,a6271a,a6272a,a6273a,a6277a,a6278a,a6282a,a6283a,a6284a,a6288a,a6289a,a6293a,a6294a,a6295a,a6299a,a6300a,a6304a,a6305a,a6306a,a6310a,a6311a,a6315a,a6316a,a6317a,a6321a,a6322a,a6326a,a6327a,a6328a,a6332a,a6333a,a6337a,a6338a,a6339a,a6343a,a6344a,a6348a,a6349a,a6350a,a6354a,a6355a,a6359a,a6360a,a6361a,a6365a,a6366a,a6370a,a6371a,a6372a,a6376a,a6377a,a6381a,a6382a,a6383a,a6387a,a6388a,a6392a,a6393a,a6394a,a6398a,a6399a,a6403a,a6404a,a6405a,a6409a,a6410a,a6414a,a6415a,a6416a,a6420a,a6421a,a6425a,a6426a,a6427a,a6431a,a6432a,a6436a,a6437a,a6438a,a6442a,a6443a,a6447a,a6448a,a6449a,a6453a,a6454a,a6458a,a6459a,a6460a,a6464a,a6465a,a6469a,a6470a,a6471a,a6475a,a6476a,a6480a,a6481a,a6482a,a6486a,a6487a,a6491a,a6492a,a6493a,a6497a,a6498a,a6502a,a6503a,a6504a,a6508a,a6509a,a6513a,a6514a,a6515a,a6519a,a6520a,a6524a,a6525a,a6526a,a6530a,a6531a,a6535a,a6536a,a6537a,a6541a,a6542a,a6546a,a6547a,a6548a,a6552a,a6553a,a6557a,a6558a,a6559a,a6563a,a6564a,a6568a,a6569a,a6570a,a6574a,a6575a,a6579a,a6580a,a6581a,a6585a,a6586a,a6590a,a6591a,a6592a,a6596a,a6597a,a6601a,a6602a,a6603a,a6607a,a6608a,a6612a,a6613a,a6614a,a6618a,a6619a,a6623a,a6624a,a6625a,a6629a,a6630a,a6634a,a6635a,a6636a,a6640a,a6641a,a6645a,a6646a,a6647a,a6651a,a6652a,a6656a,a6657a,a6658a,a6662a,a6663a,a6667a,a6668a,a6669a,a6673a,a6674a,a6678a,a6679a,a6680a,a6684a,a6685a,a6689a,a6690a,a6691a,a6695a,a6696a,a6700a,a6701a,a6702a,a6706a,a6707a,a6711a,a6712a,a6713a,a6717a,a6718a,a6722a,a6723a,a6724a,a6728a,a6729a,a6733a,a6734a,a6735a,a6739a,a6740a,a6744a,a6745a,a6746a,a6750a,a6751a,a6755a,a6756a,a6757a,a6761a,a6762a,a6766a,a6767a,a6768a,a6772a,a6773a,a6777a,a6778a,a6779a,a6783a,a6784a,a6788a,a6789a,a6790a,a6794a,a6795a,a6799a,a6800a,a6801a,a6805a,a6806a,a6810a,a6811a,a6812a,a6816a,a6817a,a6821a,a6822a,a6823a,a6827a,a6828a,a6832a,a6833a,a6834a,a6838a,a6839a,a6843a,a6844a,a6845a,a6849a,a6850a,a6853a,a6856a,a6857a,a6858a,a6862a,a6863a,a6867a,a6868a,a6869a,a6873a,a6874a,a6877a,a6880a,a6881a,a6882a,a6886a,a6887a,a6891a,a6892a,a6893a,a6897a,a6898a,a6901a,a6904a,a6905a,a6906a,a6910a,a6911a,a6915a,a6916a,a6917a,a6921a,a6922a,a6925a,a6928a,a6929a,a6930a,a6934a,a6935a,a6939a,a6940a,a6941a,a6945a,a6946a,a6949a,a6952a,a6953a,a6954a,a6958a,a6959a,a6963a,a6964a,a6965a,a6969a,a6970a,a6973a,a6976a,a6977a,a6978a,a6982a,a6983a,a6987a,a6988a,a6989a,a6993a,a6994a,a6997a,a7000a,a7001a,a7002a,a7006a,a7007a,a7011a,a7012a,a7013a,a7017a,a7018a,a7021a,a7024a,a7025a,a7026a,a7030a,a7031a,a7035a,a7036a,a7037a,a7041a,a7042a,a7045a,a7048a,a7049a,a7050a,a7054a,a7055a,a7059a,a7060a,a7061a,a7065a,a7066a,a7069a,a7072a,a7073a,a7074a,a7078a,a7079a,a7083a,a7084a,a7085a,a7089a,a7090a,a7093a,a7096a,a7097a,a7098a,a7102a,a7103a,a7107a,a7108a,a7109a,a7113a,a7114a,a7117a,a7120a,a7121a,a7122a,a7126a,a7127a,a7131a,a7132a,a7133a,a7137a,a7138a,a7141a,a7144a,a7145a,a7146a,a7150a,a7151a,a7155a,a7156a,a7157a,a7161a,a7162a,a7165a,a7168a,a7169a,a7170a,a7174a,a7175a,a7179a,a7180a,a7181a,a7185a,a7186a,a7189a,a7192a,a7193a,a7194a,a7198a,a7199a,a7203a,a7204a,a7205a,a7209a,a7210a,a7213a,a7216a,a7217a,a7218a,a7222a,a7223a,a7227a,a7228a,a7229a,a7233a,a7234a,a7237a,a7240a,a7241a,a7242a,a7246a,a7247a,a7251a,a7252a,a7253a,a7257a,a7258a,a7261a,a7264a,a7265a,a7266a,a7270a,a7271a,a7275a,a7276a,a7277a,a7281a,a7282a,a7285a,a7288a,a7289a,a7290a,a7294a,a7295a,a7299a,a7300a,a7301a,a7305a,a7306a,a7309a,a7312a,a7313a,a7314a,a7318a,a7319a,a7323a,a7324a,a7325a,a7329a,a7330a,a7333a,a7336a,a7337a,a7338a,a7342a,a7343a,a7347a,a7348a,a7349a,a7353a,a7354a,a7357a,a7360a,a7361a,a7362a,a7366a,a7367a,a7371a,a7372a,a7373a,a7377a,a7378a,a7381a,a7384a,a7385a,a7386a,a7390a,a7391a,a7395a,a7396a,a7397a,a7401a,a7402a,a7405a,a7408a,a7409a,a7410a,a7414a,a7415a,a7419a,a7420a,a7421a,a7425a,a7426a,a7429a,a7432a,a7433a,a7434a,a7438a,a7439a,a7443a,a7444a,a7445a,a7449a,a7450a,a7453a,a7456a,a7457a,a7458a,a7462a,a7463a,a7467a,a7468a,a7469a,a7473a,a7474a,a7477a,a7480a,a7481a,a7482a,a7486a,a7487a,a7491a,a7492a,a7493a,a7497a,a7498a,a7501a,a7504a,a7505a,a7506a,a7510a,a7511a,a7515a,a7516a,a7517a,a7521a,a7522a,a7525a,a7528a,a7529a,a7530a,a7534a,a7535a,a7539a,a7540a,a7541a,a7545a,a7546a,a7549a,a7552a,a7553a,a7554a,a7558a,a7559a,a7563a,a7564a,a7565a,a7569a,a7570a,a7573a,a7576a,a7577a,a7578a,a7582a,a7583a,a7587a,a7588a,a7589a,a7593a,a7594a,a7597a,a7600a,a7601a,a7602a,a7606a,a7607a,a7611a,a7612a,a7613a,a7617a,a7618a,a7621a,a7624a,a7625a,a7626a,a7630a,a7631a,a7635a,a7636a,a7637a,a7641a,a7642a,a7645a,a7648a,a7649a,a7650a,a7654a,a7655a,a7659a,a7660a,a7661a,a7665a,a7666a,a7669a,a7672a,a7673a,a7674a,a7678a,a7679a,a7683a,a7684a,a7685a,a7689a,a7690a,a7693a,a7696a,a7697a,a7698a,a7702a,a7703a,a7707a,a7708a,a7709a,a7713a,a7714a,a7717a,a7720a,a7721a,a7722a,a7726a,a7727a,a7731a,a7732a,a7733a,a7737a,a7738a,a7741a,a7744a,a7745a,a7746a,a7750a,a7751a,a7755a,a7756a,a7757a,a7761a,a7762a,a7765a,a7768a,a7769a,a7770a,a7774a,a7775a,a7779a,a7780a,a7781a,a7785a,a7786a,a7789a,a7792a,a7793a,a7794a,a7798a,a7799a,a7803a,a7804a,a7805a,a7809a,a7810a,a7813a,a7816a,a7817a,a7818a,a7822a,a7823a,a7827a,a7828a,a7829a,a7833a,a7834a,a7837a,a7840a,a7841a,a7842a,a7846a,a7847a,a7851a,a7852a,a7853a,a7857a,a7858a,a7861a,a7864a,a7865a,a7866a,a7870a,a7871a,a7875a,a7876a,a7877a,a7881a,a7882a,a7885a,a7888a,a7889a,a7890a,a7894a,a7895a,a7899a,a7900a,a7901a,a7905a,a7906a,a7909a,a7912a,a7913a,a7914a,a7918a,a7919a,a7923a,a7924a,a7925a,a7929a,a7930a,a7933a,a7936a,a7937a,a7938a,a7942a,a7943a,a7947a,a7948a,a7949a,a7953a,a7954a,a7957a,a7960a,a7961a,a7962a,a7966a,a7967a,a7971a,a7972a,a7973a,a7977a,a7978a,a7981a,a7984a,a7985a,a7986a,a7990a,a7991a,a7994a,a7997a,a7998a,a7999a,a8003a,a8004a,a8007a,a8010a,a8011a,a8012a,a8016a,a8017a,a8020a,a8023a,a8024a,a8025a,a8029a,a8030a,a8033a,a8036a,a8037a,a8038a,a8042a,a8043a,a8046a,a8049a,a8050a,a8051a,a8055a,a8056a,a8059a,a8062a,a8063a,a8064a,a8068a,a8069a,a8072a,a8075a,a8076a,a8077a,a8081a,a8082a,a8085a,a8088a,a8089a,a8090a,a8094a,a8095a,a8098a,a8101a,a8102a,a8103a,a8107a,a8108a,a8111a,a8114a,a8115a,a8116a,a8120a,a8121a,a8124a,a8127a,a8128a,a8129a,a8133a,a8134a,a8137a,a8140a,a8141a,a8142a,a8146a,a8147a,a8150a,a8153a,a8154a,a8155a,a8159a,a8160a,a8163a,a8166a,a8167a,a8168a,a8172a,a8173a,a8176a,a8179a,a8180a,a8181a,a8185a,a8186a,a8189a,a8192a,a8193a,a8194a,a8198a,a8199a,a8202a,a8205a,a8206a,a8207a,a8211a,a8212a,a8215a,a8218a,a8219a,a8220a,a8224a,a8225a,a8228a,a8231a,a8232a,a8233a,a8237a,a8238a,a8241a,a8244a,a8245a,a8246a,a8250a,a8251a,a8254a,a8257a,a8258a,a8259a,a8263a,a8264a,a8267a,a8270a,a8271a,a8272a,a8276a,a8277a,a8280a,a8283a,a8284a,a8285a,a8289a,a8290a,a8293a,a8296a,a8297a,a8298a,a8302a,a8303a,a8306a,a8309a,a8310a,a8311a,a8315a,a8316a,a8319a,a8322a,a8323a,a8324a,a8328a,a8329a,a8332a,a8335a,a8336a,a8337a,a8341a,a8342a,a8345a,a8348a,a8349a,a8350a,a8354a,a8355a,a8358a,a8361a,a8362a,a8363a,a8367a,a8368a,a8371a,a8374a,a8375a,a8376a,a8380a,a8381a,a8384a,a8387a,a8388a,a8389a,a8393a,a8394a,a8397a,a8400a,a8401a,a8402a,a8406a,a8407a,a8410a,a8413a,a8414a,a8415a,a8419a,a8420a,a8423a,a8426a,a8427a,a8428a,a8432a,a8433a,a8436a,a8439a,a8440a,a8441a,a8445a,a8446a,a8449a,a8452a,a8453a,a8454a,a8458a,a8459a,a8462a,a8465a,a8466a,a8467a,a8471a,a8472a,a8475a,a8478a,a8479a,a8480a,a8484a,a8485a,a8488a,a8491a,a8492a,a8493a,a8497a,a8498a,a8501a,a8504a,a8505a,a8506a,a8510a,a8511a,a8514a,a8517a,a8518a,a8519a,a8523a,a8524a,a8527a,a8530a,a8531a,a8532a,a8536a,a8537a,a8540a,a8543a,a8544a,a8545a,a8549a,a8550a,a8553a,a8556a,a8557a,a8558a,a8562a,a8563a,a8566a,a8569a,a8570a,a8571a,a8575a,a8576a,a8579a,a8582a,a8583a,a8584a,a8588a,a8589a,a8592a,a8595a,a8596a,a8597a,a8601a,a8602a,a8605a,a8608a,a8609a,a8610a,a8614a,a8615a,a8618a,a8621a,a8622a,a8623a,a8627a,a8628a,a8631a,a8634a,a8635a,a8636a,a8640a,a8641a,a8644a,a8647a,a8648a,a8649a,a8653a,a8654a,a8657a,a8660a,a8661a,a8662a,a8666a,a8667a,a8670a,a8673a,a8674a,a8675a,a8679a,a8680a,a8683a,a8686a,a8687a,a8688a,a8692a,a8693a,a8696a,a8699a,a8700a,a8701a,a8705a,a8706a,a8709a,a8712a,a8713a,a8714a,a8718a,a8719a,a8722a,a8725a,a8726a,a8727a,a8731a,a8732a,a8735a,a8738a,a8739a,a8740a,a8744a,a8745a,a8748a,a8751a,a8752a,a8753a,a8757a,a8758a,a8761a,a8764a,a8765a,a8766a,a8770a,a8771a,a8774a,a8777a,a8778a,a8779a,a8783a,a8784a,a8787a,a8790a,a8791a,a8792a,a8796a,a8797a,a8800a,a8803a,a8804a,a8805a,a8809a,a8810a,a8813a,a8816a,a8817a,a8818a,a8822a,a8823a,a8826a,a8829a,a8830a,a8831a,a8835a,a8836a,a8839a,a8842a,a8843a,a8844a,a8848a,a8849a,a8852a,a8855a,a8856a,a8857a,a8861a,a8862a,a8865a,a8868a,a8869a,a8870a,a8874a,a8875a,a8878a,a8881a,a8882a,a8883a,a8887a,a8888a,a8891a,a8894a,a8895a,a8896a,a8900a,a8901a,a8904a,a8907a,a8908a,a8909a,a8913a,a8914a,a8917a,a8920a,a8921a,a8922a,a8926a,a8927a,a8930a,a8933a,a8934a,a8935a,a8939a,a8940a,a8943a,a8946a,a8947a,a8948a,a8952a,a8953a,a8956a,a8959a,a8960a,a8961a,a8965a,a8966a,a8969a,a8972a,a8973a,a8974a,a8978a,a8979a,a8982a,a8985a,a8986a,a8987a,a8991a,a8992a,a8995a,a8998a,a8999a,a9000a,a9004a,a9005a,a9008a,a9011a,a9012a,a9013a,a9017a,a9018a,a9021a,a9024a,a9025a,a9026a,a9030a,a9031a,a9034a,a9037a,a9038a,a9039a,a9043a,a9044a,a9047a,a9050a,a9051a,a9052a,a9056a,a9057a,a9060a,a9063a,a9064a,a9065a,a9069a,a9070a,a9073a,a9076a,a9077a,a9078a,a9082a,a9083a,a9086a,a9089a,a9090a,a9091a,a9095a,a9096a,a9099a,a9102a,a9103a,a9104a,a9108a,a9109a,a9112a,a9115a,a9116a,a9117a,a9121a,a9122a,a9125a,a9128a,a9129a,a9130a,a9134a,a9135a,a9138a,a9141a,a9142a,a9143a,a9147a,a9148a,a9151a,a9154a,a9155a,a9156a,a9160a,a9161a,a9164a,a9167a,a9168a,a9169a,a9173a,a9174a,a9177a,a9180a,a9181a,a9182a,a9186a,a9187a,a9190a,a9193a,a9194a,a9195a,a9199a,a9200a,a9203a,a9206a,a9207a,a9208a,a9212a,a9213a,a9216a,a9219a,a9220a,a9221a,a9225a,a9226a,a9229a,a9232a,a9233a,a9234a,a9238a,a9239a,a9242a,a9245a,a9246a,a9247a,a9251a,a9252a,a9255a,a9258a,a9259a,a9260a,a9264a,a9265a,a9268a,a9271a,a9272a,a9273a,a9277a,a9278a,a9281a,a9284a,a9285a,a9286a,a9290a,a9291a,a9294a,a9297a,a9298a,a9299a,a9303a,a9304a,a9307a,a9310a,a9311a,a9312a,a9316a,a9317a,a9320a,a9323a,a9324a,a9325a,a9329a,a9330a,a9333a,a9336a,a9337a,a9338a,a9342a,a9343a,a9346a,a9349a,a9350a,a9351a,a9355a,a9356a,a9359a,a9362a,a9363a,a9364a,a9368a,a9369a,a9372a,a9375a,a9376a,a9377a,a9381a,a9382a,a9385a,a9388a,a9389a,a9390a,a9394a,a9395a,a9398a,a9401a,a9402a,a9403a,a9407a,a9408a,a9411a,a9414a,a9415a,a9416a,a9420a,a9421a,a9424a,a9427a,a9428a,a9429a,a9433a,a9434a,a9437a,a9440a,a9441a,a9442a,a9446a,a9447a,a9450a,a9453a,a9454a,a9455a,a9459a,a9460a,a9463a,a9466a,a9467a,a9468a,a9472a,a9473a,a9476a,a9479a,a9480a,a9481a,a9485a,a9486a,a9489a,a9492a,a9493a,a9494a,a9498a,a9499a,a9502a,a9505a,a9506a,a9507a,a9511a,a9512a,a9515a,a9518a,a9519a,a9520a,a9524a,a9525a,a9528a,a9531a,a9532a,a9533a,a9537a,a9538a,a9541a,a9544a,a9545a,a9546a,a9550a,a9551a,a9554a,a9557a,a9558a,a9559a,a9563a,a9564a,a9567a,a9570a,a9571a,a9572a,a9576a,a9577a,a9580a,a9583a,a9584a,a9585a,a9589a,a9590a,a9593a,a9596a,a9597a,a9598a,a9602a,a9603a,a9606a,a9609a,a9610a,a9611a,a9615a,a9616a,a9619a,a9622a,a9623a,a9624a,a9628a,a9629a,a9632a,a9635a,a9636a,a9637a,a9641a,a9642a,a9645a,a9648a,a9649a,a9650a,a9654a,a9655a,a9658a,a9661a,a9662a,a9663a,a9667a,a9668a,a9671a,a9674a,a9675a,a9676a,a9680a,a9681a,a9684a,a9687a,a9688a,a9689a,a9693a,a9694a,a9697a,a9700a,a9701a,a9702a,a9706a,a9707a,a9710a,a9713a,a9714a,a9715a,a9719a,a9720a,a9723a,a9726a,a9727a,a9728a,a9732a,a9733a,a9736a,a9739a,a9740a,a9741a,a9745a,a9746a,a9749a,a9752a,a9753a,a9754a,a9758a,a9759a,a9762a,a9765a,a9766a,a9767a,a9771a,a9772a,a9775a,a9778a,a9779a,a9780a,a9784a,a9785a,a9788a,a9791a,a9792a,a9793a,a9797a,a9798a,a9801a,a9804a,a9805a,a9806a,a9810a,a9811a,a9814a,a9817a,a9818a,a9819a,a9823a,a9824a,a9827a,a9830a,a9831a,a9832a,a9836a,a9837a,a9840a,a9843a,a9844a,a9845a,a9849a,a9850a,a9853a,a9856a,a9857a,a9858a,a9862a,a9863a,a9866a,a9869a,a9870a,a9871a,a9875a,a9876a,a9879a,a9882a,a9883a,a9884a,a9888a,a9889a,a9892a,a9895a,a9896a,a9897a,a9901a,a9902a,a9905a,a9908a,a9909a,a9910a,a9914a,a9915a,a9918a,a9921a,a9922a,a9923a,a9927a,a9928a,a9931a,a9934a,a9935a,a9936a,a9940a,a9941a,a9944a,a9947a,a9948a,a9949a,a9953a,a9954a,a9957a,a9960a,a9961a,a9962a,a9966a,a9967a,a9970a,a9973a,a9974a,a9975a,a9979a,a9980a,a9983a,a9986a,a9987a,a9988a,a9992a,a9993a,a9996a,a9999a,a10000a,a10001a,a10005a,a10006a,a10009a,a10012a,a10013a,a10014a,a10018a,a10019a,a10022a,a10025a,a10026a,a10027a,a10031a,a10032a,a10035a,a10038a,a10039a,a10040a,a10044a,a10045a,a10048a,a10051a,a10052a,a10053a,a10057a,a10058a,a10061a,a10064a,a10065a,a10066a,a10070a,a10071a,a10074a,a10077a,a10078a,a10079a,a10083a,a10084a,a10087a,a10090a,a10091a,a10092a,a10096a,a10097a,a10100a,a10103a,a10104a,a10105a,a10109a,a10110a,a10113a,a10116a,a10117a,a10118a,a10122a,a10123a,a10126a,a10129a,a10130a,a10131a,a10135a,a10136a,a10139a,a10142a,a10143a,a10144a,a10148a,a10149a,a10152a,a10155a,a10156a,a10157a,a10161a,a10162a,a10165a,a10168a,a10169a,a10170a,a10174a,a10175a,a10178a,a10181a,a10182a,a10183a,a10187a,a10188a,a10191a,a10194a,a10195a,a10196a,a10200a,a10201a,a10204a,a10207a,a10208a,a10209a,a10213a,a10214a,a10217a,a10220a,a10221a,a10222a,a10226a,a10227a,a10230a,a10233a,a10234a,a10235a,a10239a,a10240a,a10243a,a10246a,a10247a,a10248a,a10252a,a10253a,a10256a,a10259a,a10260a,a10261a,a10265a,a10266a,a10269a,a10272a,a10273a,a10274a,a10278a,a10279a,a10282a,a10285a,a10286a,a10287a,a10291a,a10292a,a10295a,a10298a,a10299a,a10300a,a10304a,a10305a,a10308a,a10311a,a10312a,a10313a,a10317a,a10318a,a10321a,a10324a,a10325a,a10326a,a10330a,a10331a,a10334a,a10337a,a10338a,a10339a,a10343a,a10344a,a10347a,a10350a,a10351a,a10352a,a10356a,a10357a,a10360a,a10363a,a10364a,a10365a,a10369a,a10370a,a10373a,a10376a,a10377a,a10378a,a10382a,a10383a,a10386a,a10389a,a10390a,a10391a,a10395a,a10396a,a10399a,a10402a,a10403a,a10404a,a10408a,a10409a,a10412a,a10415a,a10416a,a10417a,a10421a,a10422a,a10425a,a10428a,a10429a,a10430a,a10434a,a10435a,a10438a,a10441a,a10442a,a10443a,a10447a,a10448a,a10451a,a10454a,a10455a,a10456a,a10460a,a10461a,a10464a,a10467a,a10468a,a10469a,a10473a,a10474a,a10477a,a10480a,a10481a,a10482a,a10486a,a10487a,a10490a,a10493a,a10494a,a10495a,a10498a,a10501a,a10502a,a10505a,a10508a,a10509a,a10510a,a10514a,a10515a,a10518a,a10521a,a10522a,a10523a,a10526a,a10529a,a10530a,a10533a,a10536a,a10537a,a10538a,a10542a,a10543a,a10546a,a10549a,a10550a,a10551a,a10554a,a10557a,a10558a,a10561a,a10564a,a10565a,a10566a,a10570a,a10571a,a10574a,a10577a,a10578a,a10579a,a10582a,a10585a,a10586a,a10589a,a10592a,a10593a,a10594a,a10598a,a10599a,a10602a,a10605a,a10606a,a10607a,a10610a,a10613a,a10614a,a10617a,a10620a,a10621a,a10622a,a10626a,a10627a,a10630a,a10633a,a10634a,a10635a,a10638a,a10641a,a10642a,a10645a,a10648a,a10649a,a10650a,a10654a,a10655a,a10658a,a10661a,a10662a,a10663a,a10666a,a10669a,a10670a,a10673a,a10676a,a10677a,a10678a,a10682a,a10683a,a10686a,a10689a,a10690a,a10691a,a10694a,a10697a,a10698a,a10701a,a10704a,a10705a,a10706a,a10710a,a10711a,a10714a,a10717a,a10718a,a10719a,a10722a,a10725a,a10726a,a10729a,a10732a,a10733a,a10734a,a10738a,a10739a,a10742a,a10745a,a10746a,a10747a,a10750a,a10753a,a10754a,a10757a,a10760a,a10761a,a10762a,a10766a,a10767a,a10770a,a10773a,a10774a,a10775a,a10778a,a10781a,a10782a,a10785a,a10788a,a10789a,a10790a,a10794a,a10795a,a10798a,a10801a,a10802a,a10803a,a10806a,a10809a,a10810a,a10813a,a10816a,a10817a,a10818a,a10822a,a10823a,a10826a,a10829a,a10830a,a10831a,a10834a,a10837a,a10838a,a10841a,a10844a,a10845a,a10846a,a10850a,a10851a,a10854a,a10857a,a10858a,a10859a,a10862a,a10865a,a10866a,a10869a,a10872a,a10873a,a10874a,a10878a,a10879a,a10882a,a10885a,a10886a,a10887a,a10890a,a10893a,a10894a,a10897a,a10900a,a10901a,a10902a,a10906a,a10907a,a10910a,a10913a,a10914a,a10915a,a10918a,a10921a,a10922a,a10925a,a10928a,a10929a,a10930a,a10934a,a10935a,a10938a,a10941a,a10942a,a10943a,a10946a,a10949a,a10950a,a10953a,a10956a,a10957a,a10958a,a10962a,a10963a,a10966a,a10969a,a10970a,a10971a,a10974a,a10977a,a10978a,a10981a,a10984a,a10985a,a10986a,a10990a,a10991a,a10994a,a10997a,a10998a,a10999a,a11002a,a11005a,a11006a,a11009a,a11012a,a11013a,a11014a,a11018a,a11019a,a11022a,a11025a,a11026a,a11027a,a11030a,a11033a,a11034a,a11037a,a11040a,a11041a,a11042a,a11046a,a11047a,a11050a,a11053a,a11054a,a11055a,a11058a,a11061a,a11062a,a11065a,a11068a,a11069a,a11070a,a11074a,a11075a,a11078a,a11081a,a11082a,a11083a,a11086a,a11089a,a11090a,a11093a,a11096a,a11097a,a11098a,a11102a,a11103a,a11106a,a11109a,a11110a,a11111a,a11114a,a11117a,a11118a,a11121a,a11124a,a11125a,a11126a,a11130a,a11131a,a11134a,a11137a,a11138a,a11139a,a11142a,a11145a,a11146a,a11149a,a11152a,a11153a,a11154a,a11158a,a11159a,a11162a,a11165a,a11166a,a11167a,a11170a,a11173a,a11174a,a11177a,a11180a,a11181a,a11182a,a11186a,a11187a,a11190a,a11193a,a11194a,a11195a,a11198a,a11201a,a11202a,a11205a,a11208a,a11209a,a11210a,a11214a,a11215a,a11218a,a11221a,a11222a,a11223a,a11226a,a11229a,a11230a,a11233a,a11236a,a11237a,a11238a,a11242a,a11243a,a11246a,a11249a,a11250a,a11251a,a11254a,a11257a,a11258a,a11261a,a11264a,a11265a,a11266a,a11270a,a11271a,a11274a,a11277a,a11278a,a11279a,a11282a,a11285a,a11286a,a11289a,a11292a,a11293a,a11294a,a11298a,a11299a,a11302a,a11305a,a11306a,a11307a,a11310a,a11313a,a11314a,a11317a,a11320a,a11321a,a11322a,a11326a,a11327a,a11330a,a11333a,a11334a,a11335a,a11338a,a11341a,a11342a,a11345a,a11348a,a11349a,a11350a,a11354a,a11355a,a11358a,a11361a,a11362a,a11363a,a11366a,a11369a,a11370a,a11373a,a11376a,a11377a,a11378a: std_logic;
begin

A108 <=( a1366a ) or ( a911a );
 a1a <=( a11378a  and  a11363a );
 a2a <=( a11350a  and  a11335a );
 a3a <=( a11322a  and  a11307a );
 a4a <=( a11294a  and  a11279a );
 a5a <=( a11266a  and  a11251a );
 a6a <=( a11238a  and  a11223a );
 a7a <=( a11210a  and  a11195a );
 a8a <=( a11182a  and  a11167a );
 a9a <=( a11154a  and  a11139a );
 a10a <=( a11126a  and  a11111a );
 a11a <=( a11098a  and  a11083a );
 a12a <=( a11070a  and  a11055a );
 a13a <=( a11042a  and  a11027a );
 a14a <=( a11014a  and  a10999a );
 a15a <=( a10986a  and  a10971a );
 a16a <=( a10958a  and  a10943a );
 a17a <=( a10930a  and  a10915a );
 a18a <=( a10902a  and  a10887a );
 a19a <=( a10874a  and  a10859a );
 a20a <=( a10846a  and  a10831a );
 a21a <=( a10818a  and  a10803a );
 a22a <=( a10790a  and  a10775a );
 a23a <=( a10762a  and  a10747a );
 a24a <=( a10734a  and  a10719a );
 a25a <=( a10706a  and  a10691a );
 a26a <=( a10678a  and  a10663a );
 a27a <=( a10650a  and  a10635a );
 a28a <=( a10622a  and  a10607a );
 a29a <=( a10594a  and  a10579a );
 a30a <=( a10566a  and  a10551a );
 a31a <=( a10538a  and  a10523a );
 a32a <=( a10510a  and  a10495a );
 a33a <=( a10482a  and  a10469a );
 a34a <=( a10456a  and  a10443a );
 a35a <=( a10430a  and  a10417a );
 a36a <=( a10404a  and  a10391a );
 a37a <=( a10378a  and  a10365a );
 a38a <=( a10352a  and  a10339a );
 a39a <=( a10326a  and  a10313a );
 a40a <=( a10300a  and  a10287a );
 a41a <=( a10274a  and  a10261a );
 a42a <=( a10248a  and  a10235a );
 a43a <=( a10222a  and  a10209a );
 a44a <=( a10196a  and  a10183a );
 a45a <=( a10170a  and  a10157a );
 a46a <=( a10144a  and  a10131a );
 a47a <=( a10118a  and  a10105a );
 a48a <=( a10092a  and  a10079a );
 a49a <=( a10066a  and  a10053a );
 a50a <=( a10040a  and  a10027a );
 a51a <=( a10014a  and  a10001a );
 a52a <=( a9988a  and  a9975a );
 a53a <=( a9962a  and  a9949a );
 a54a <=( a9936a  and  a9923a );
 a55a <=( a9910a  and  a9897a );
 a56a <=( a9884a  and  a9871a );
 a57a <=( a9858a  and  a9845a );
 a58a <=( a9832a  and  a9819a );
 a59a <=( a9806a  and  a9793a );
 a60a <=( a9780a  and  a9767a );
 a61a <=( a9754a  and  a9741a );
 a62a <=( a9728a  and  a9715a );
 a63a <=( a9702a  and  a9689a );
 a64a <=( a9676a  and  a9663a );
 a65a <=( a9650a  and  a9637a );
 a66a <=( a9624a  and  a9611a );
 a67a <=( a9598a  and  a9585a );
 a68a <=( a9572a  and  a9559a );
 a69a <=( a9546a  and  a9533a );
 a70a <=( a9520a  and  a9507a );
 a71a <=( a9494a  and  a9481a );
 a72a <=( a9468a  and  a9455a );
 a73a <=( a9442a  and  a9429a );
 a74a <=( a9416a  and  a9403a );
 a75a <=( a9390a  and  a9377a );
 a76a <=( a9364a  and  a9351a );
 a77a <=( a9338a  and  a9325a );
 a78a <=( a9312a  and  a9299a );
 a79a <=( a9286a  and  a9273a );
 a80a <=( a9260a  and  a9247a );
 a81a <=( a9234a  and  a9221a );
 a82a <=( a9208a  and  a9195a );
 a83a <=( a9182a  and  a9169a );
 a84a <=( a9156a  and  a9143a );
 a85a <=( a9130a  and  a9117a );
 a86a <=( a9104a  and  a9091a );
 a87a <=( a9078a  and  a9065a );
 a88a <=( a9052a  and  a9039a );
 a89a <=( a9026a  and  a9013a );
 a90a <=( a9000a  and  a8987a );
 a91a <=( a8974a  and  a8961a );
 a92a <=( a8948a  and  a8935a );
 a93a <=( a8922a  and  a8909a );
 a94a <=( a8896a  and  a8883a );
 a95a <=( a8870a  and  a8857a );
 a96a <=( a8844a  and  a8831a );
 a97a <=( a8818a  and  a8805a );
 a98a <=( a8792a  and  a8779a );
 a99a <=( a8766a  and  a8753a );
 a100a <=( a8740a  and  a8727a );
 a101a <=( a8714a  and  a8701a );
 a102a <=( a8688a  and  a8675a );
 a103a <=( a8662a  and  a8649a );
 a104a <=( a8636a  and  a8623a );
 a105a <=( a8610a  and  a8597a );
 a106a <=( a8584a  and  a8571a );
 a107a <=( a8558a  and  a8545a );
 a108a <=( a8532a  and  a8519a );
 a109a <=( a8506a  and  a8493a );
 a110a <=( a8480a  and  a8467a );
 a111a <=( a8454a  and  a8441a );
 a112a <=( a8428a  and  a8415a );
 a113a <=( a8402a  and  a8389a );
 a114a <=( a8376a  and  a8363a );
 a115a <=( a8350a  and  a8337a );
 a116a <=( a8324a  and  a8311a );
 a117a <=( a8298a  and  a8285a );
 a118a <=( a8272a  and  a8259a );
 a119a <=( a8246a  and  a8233a );
 a120a <=( a8220a  and  a8207a );
 a121a <=( a8194a  and  a8181a );
 a122a <=( a8168a  and  a8155a );
 a123a <=( a8142a  and  a8129a );
 a124a <=( a8116a  and  a8103a );
 a125a <=( a8090a  and  a8077a );
 a126a <=( a8064a  and  a8051a );
 a127a <=( a8038a  and  a8025a );
 a128a <=( a8012a  and  a7999a );
 a129a <=( a7986a  and  a7973a );
 a130a <=( a7962a  and  a7949a );
 a131a <=( a7938a  and  a7925a );
 a132a <=( a7914a  and  a7901a );
 a133a <=( a7890a  and  a7877a );
 a134a <=( a7866a  and  a7853a );
 a135a <=( a7842a  and  a7829a );
 a136a <=( a7818a  and  a7805a );
 a137a <=( a7794a  and  a7781a );
 a138a <=( a7770a  and  a7757a );
 a139a <=( a7746a  and  a7733a );
 a140a <=( a7722a  and  a7709a );
 a141a <=( a7698a  and  a7685a );
 a142a <=( a7674a  and  a7661a );
 a143a <=( a7650a  and  a7637a );
 a144a <=( a7626a  and  a7613a );
 a145a <=( a7602a  and  a7589a );
 a146a <=( a7578a  and  a7565a );
 a147a <=( a7554a  and  a7541a );
 a148a <=( a7530a  and  a7517a );
 a149a <=( a7506a  and  a7493a );
 a150a <=( a7482a  and  a7469a );
 a151a <=( a7458a  and  a7445a );
 a152a <=( a7434a  and  a7421a );
 a153a <=( a7410a  and  a7397a );
 a154a <=( a7386a  and  a7373a );
 a155a <=( a7362a  and  a7349a );
 a156a <=( a7338a  and  a7325a );
 a157a <=( a7314a  and  a7301a );
 a158a <=( a7290a  and  a7277a );
 a159a <=( a7266a  and  a7253a );
 a160a <=( a7242a  and  a7229a );
 a161a <=( a7218a  and  a7205a );
 a162a <=( a7194a  and  a7181a );
 a163a <=( a7170a  and  a7157a );
 a164a <=( a7146a  and  a7133a );
 a165a <=( a7122a  and  a7109a );
 a166a <=( a7098a  and  a7085a );
 a167a <=( a7074a  and  a7061a );
 a168a <=( a7050a  and  a7037a );
 a169a <=( a7026a  and  a7013a );
 a170a <=( a7002a  and  a6989a );
 a171a <=( a6978a  and  a6965a );
 a172a <=( a6954a  and  a6941a );
 a173a <=( a6930a  and  a6917a );
 a174a <=( a6906a  and  a6893a );
 a175a <=( a6882a  and  a6869a );
 a176a <=( a6858a  and  a6845a );
 a177a <=( a6834a  and  a6823a );
 a178a <=( a6812a  and  a6801a );
 a179a <=( a6790a  and  a6779a );
 a180a <=( a6768a  and  a6757a );
 a181a <=( a6746a  and  a6735a );
 a182a <=( a6724a  and  a6713a );
 a183a <=( a6702a  and  a6691a );
 a184a <=( a6680a  and  a6669a );
 a185a <=( a6658a  and  a6647a );
 a186a <=( a6636a  and  a6625a );
 a187a <=( a6614a  and  a6603a );
 a188a <=( a6592a  and  a6581a );
 a189a <=( a6570a  and  a6559a );
 a190a <=( a6548a  and  a6537a );
 a191a <=( a6526a  and  a6515a );
 a192a <=( a6504a  and  a6493a );
 a193a <=( a6482a  and  a6471a );
 a194a <=( a6460a  and  a6449a );
 a195a <=( a6438a  and  a6427a );
 a196a <=( a6416a  and  a6405a );
 a197a <=( a6394a  and  a6383a );
 a198a <=( a6372a  and  a6361a );
 a199a <=( a6350a  and  a6339a );
 a200a <=( a6328a  and  a6317a );
 a201a <=( a6306a  and  a6295a );
 a202a <=( a6284a  and  a6273a );
 a203a <=( a6262a  and  a6251a );
 a204a <=( a6240a  and  a6229a );
 a205a <=( a6218a  and  a6207a );
 a206a <=( a6196a  and  a6185a );
 a207a <=( a6174a  and  a6163a );
 a208a <=( a6152a  and  a6141a );
 a209a <=( a6130a  and  a6119a );
 a210a <=( a6108a  and  a6097a );
 a211a <=( a6086a  and  a6075a );
 a212a <=( a6064a  and  a6053a );
 a213a <=( a6042a  and  a6031a );
 a214a <=( a6020a  and  a6009a );
 a215a <=( a5998a  and  a5987a );
 a216a <=( a5976a  and  a5965a );
 a217a <=( a5954a  and  a5943a );
 a218a <=( a5932a  and  a5921a );
 a219a <=( a5910a  and  a5899a );
 a220a <=( a5888a  and  a5877a );
 a221a <=( a5866a  and  a5855a );
 a222a <=( a5844a  and  a5833a );
 a223a <=( a5822a  and  a5811a );
 a224a <=( a5800a  and  a5789a );
 a225a <=( a5778a  and  a5767a );
 a226a <=( a5756a  and  a5745a );
 a227a <=( a5734a  and  a5723a );
 a228a <=( a5712a  and  a5701a );
 a229a <=( a5690a  and  a5679a );
 a230a <=( a5668a  and  a5657a );
 a231a <=( a5646a  and  a5635a );
 a232a <=( a5624a  and  a5613a );
 a233a <=( a5602a  and  a5591a );
 a234a <=( a5580a  and  a5569a );
 a235a <=( a5558a  and  a5547a );
 a236a <=( a5536a  and  a5525a );
 a237a <=( a5514a  and  a5503a );
 a238a <=( a5492a  and  a5481a );
 a239a <=( a5470a  and  a5459a );
 a240a <=( a5448a  and  a5437a );
 a241a <=( a5426a  and  a5415a );
 a242a <=( a5404a  and  a5393a );
 a243a <=( a5382a  and  a5371a );
 a244a <=( a5360a  and  a5349a );
 a245a <=( a5338a  and  a5327a );
 a246a <=( a5316a  and  a5305a );
 a247a <=( a5294a  and  a5283a );
 a248a <=( a5272a  and  a5261a );
 a249a <=( a5250a  and  a5239a );
 a250a <=( a5228a  and  a5217a );
 a251a <=( a5206a  and  a5195a );
 a252a <=( a5184a  and  a5173a );
 a253a <=( a5162a  and  a5151a );
 a254a <=( a5140a  and  a5129a );
 a255a <=( a5118a  and  a5107a );
 a256a <=( a5096a  and  a5085a );
 a257a <=( a5074a  and  a5063a );
 a258a <=( a5052a  and  a5041a );
 a259a <=( a5030a  and  a5019a );
 a260a <=( a5008a  and  a4997a );
 a261a <=( a4986a  and  a4975a );
 a262a <=( a4964a  and  a4953a );
 a263a <=( a4942a  and  a4931a );
 a264a <=( a4920a  and  a4909a );
 a265a <=( a4898a  and  a4887a );
 a266a <=( a4876a  and  a4865a );
 a267a <=( a4854a  and  a4843a );
 a268a <=( a4832a  and  a4821a );
 a269a <=( a4810a  and  a4799a );
 a270a <=( a4788a  and  a4777a );
 a271a <=( a4766a  and  a4755a );
 a272a <=( a4744a  and  a4733a );
 a273a <=( a4722a  and  a4711a );
 a274a <=( a4700a  and  a4689a );
 a275a <=( a4678a  and  a4667a );
 a276a <=( a4656a  and  a4645a );
 a277a <=( a4634a  and  a4623a );
 a278a <=( a4612a  and  a4601a );
 a279a <=( a4590a  and  a4579a );
 a280a <=( a4568a  and  a4557a );
 a281a <=( a4546a  and  a4535a );
 a282a <=( a4524a  and  a4513a );
 a283a <=( a4502a  and  a4491a );
 a284a <=( a4480a  and  a4469a );
 a285a <=( a4458a  and  a4447a );
 a286a <=( a4436a  and  a4425a );
 a287a <=( a4414a  and  a4403a );
 a288a <=( a4392a  and  a4381a );
 a289a <=( a4370a  and  a4359a );
 a290a <=( a4348a  and  a4337a );
 a291a <=( a4326a  and  a4315a );
 a292a <=( a4304a  and  a4293a );
 a293a <=( a4282a  and  a4271a );
 a294a <=( a4260a  and  a4249a );
 a295a <=( a4238a  and  a4227a );
 a296a <=( a4216a  and  a4205a );
 a297a <=( a4194a  and  a4183a );
 a298a <=( a4172a  and  a4161a );
 a299a <=( a4150a  and  a4139a );
 a300a <=( a4128a  and  a4117a );
 a301a <=( a4106a  and  a4095a );
 a302a <=( a4084a  and  a4073a );
 a303a <=( a4062a  and  a4051a );
 a304a <=( a4040a  and  a4029a );
 a305a <=( a4018a  and  a4007a );
 a306a <=( a3996a  and  a3985a );
 a307a <=( a3974a  and  a3963a );
 a308a <=( a3952a  and  a3941a );
 a309a <=( a3930a  and  a3919a );
 a310a <=( a3908a  and  a3897a );
 a311a <=( a3886a  and  a3875a );
 a312a <=( a3864a  and  a3853a );
 a313a <=( a3842a  and  a3831a );
 a314a <=( a3820a  and  a3809a );
 a315a <=( a3798a  and  a3787a );
 a316a <=( a3776a  and  a3765a );
 a317a <=( a3754a  and  a3743a );
 a318a <=( a3732a  and  a3721a );
 a319a <=( a3710a  and  a3699a );
 a320a <=( a3688a  and  a3677a );
 a321a <=( a3666a  and  a3655a );
 a322a <=( a3646a  and  a3635a );
 a323a <=( a3626a  and  a3615a );
 a324a <=( a3606a  and  a3595a );
 a325a <=( a3586a  and  a3575a );
 a326a <=( a3566a  and  a3555a );
 a327a <=( a3546a  and  a3535a );
 a328a <=( a3526a  and  a3515a );
 a329a <=( a3506a  and  a3495a );
 a330a <=( a3486a  and  a3475a );
 a331a <=( a3466a  and  a3455a );
 a332a <=( a3446a  and  a3435a );
 a333a <=( a3426a  and  a3415a );
 a334a <=( a3406a  and  a3395a );
 a335a <=( a3386a  and  a3375a );
 a336a <=( a3366a  and  a3355a );
 a337a <=( a3346a  and  a3335a );
 a338a <=( a3326a  and  a3315a );
 a339a <=( a3306a  and  a3295a );
 a340a <=( a3286a  and  a3275a );
 a341a <=( a3266a  and  a3255a );
 a342a <=( a3246a  and  a3235a );
 a343a <=( a3226a  and  a3215a );
 a344a <=( a3206a  and  a3195a );
 a345a <=( a3186a  and  a3177a );
 a346a <=( a3168a  and  a3159a );
 a347a <=( a3150a  and  a3141a );
 a348a <=( a3132a  and  a3123a );
 a349a <=( a3114a  and  a3105a );
 a350a <=( a3096a  and  a3087a );
 a351a <=( a3078a  and  a3069a );
 a352a <=( a3060a  and  a3051a );
 a353a <=( a3042a  and  a3033a );
 a354a <=( a3024a  and  a3015a );
 a355a <=( a3006a  and  a2997a );
 a356a <=( a2988a  and  a2979a );
 a357a <=( a2970a  and  a2961a );
 a358a <=( a2952a  and  a2943a );
 a359a <=( a2934a  and  a2925a );
 a360a <=( a2916a  and  a2907a );
 a361a <=( a2898a  and  a2889a );
 a362a <=( a2880a  and  a2871a );
 a363a <=( a2862a  and  a2853a );
 a364a <=( a2844a  and  a2835a );
 a365a <=( a2826a  and  a2817a );
 a366a <=( a2808a  and  a2799a );
 a367a <=( a2790a  and  a2781a );
 a368a <=( a2772a  and  a2763a );
 a369a <=( a2754a  and  a2745a );
 a370a <=( a2736a  and  a2727a );
 a371a <=( a2718a  and  a2709a );
 a372a <=( a2700a  and  a2691a );
 a373a <=( a2682a  and  a2673a );
 a374a <=( a2664a  and  a2655a );
 a375a <=( a2646a  and  a2637a );
 a376a <=( a2628a  and  a2619a );
 a377a <=( a2610a  and  a2601a );
 a378a <=( a2592a  and  a2583a );
 a379a <=( a2574a  and  a2565a );
 a380a <=( a2556a  and  a2547a );
 a381a <=( a2538a  and  a2529a );
 a382a <=( a2520a  and  a2511a );
 a383a <=( a2502a  and  a2493a );
 a384a <=( a2484a  and  a2475a );
 a385a <=( a2466a  and  a2457a );
 a386a <=( a2448a  and  a2439a );
 a387a <=( a2430a  and  a2421a );
 a388a <=( a2412a  and  a2403a );
 a389a <=( a2394a  and  a2385a );
 a390a <=( a2376a  and  a2367a );
 a391a <=( a2358a  and  a2349a );
 a392a <=( a2340a  and  a2331a );
 a393a <=( a2322a  and  a2313a );
 a394a <=( a2304a  and  a2295a );
 a395a <=( a2286a  and  a2277a );
 a396a <=( a2268a  and  a2259a );
 a397a <=( a2250a  and  a2241a );
 a398a <=( a2232a  and  a2223a );
 a399a <=( a2214a  and  a2205a );
 a400a <=( a2196a  and  a2187a );
 a401a <=( a2178a  and  a2169a );
 a402a <=( a2160a  and  a2151a );
 a403a <=( a2142a  and  a2133a );
 a404a <=( a2124a  and  a2115a );
 a405a <=( a2106a  and  a2097a );
 a406a <=( a2088a  and  a2079a );
 a407a <=( a2070a  and  a2061a );
 a408a <=( a2052a  and  a2043a );
 a409a <=( a2034a  and  a2025a );
 a410a <=( a2016a  and  a2007a );
 a411a <=( a1998a  and  a1989a );
 a412a <=( a1980a  and  a1971a );
 a413a <=( a1962a  and  a1953a );
 a414a <=( a1944a  and  a1935a );
 a415a <=( a1926a  and  a1917a );
 a416a <=( a1908a  and  a1899a );
 a417a <=( a1890a  and  a1881a );
 a418a <=( a1874a  and  a1865a );
 a419a <=( a1858a  and  a1849a );
 a420a <=( a1842a  and  a1833a );
 a421a <=( a1826a  and  a1819a );
 a422a <=( a1812a  and  a1805a );
 a423a <=( a1798a  and  a1791a );
 a424a <=( a1784a  and  a1777a );
 a425a <=( a1770a  and  a1763a );
 a426a <=( a1756a  and  a1749a );
 a427a <=( a1742a  and  a1735a );
 a428a <=( a1728a  and  a1721a );
 a429a <=( a1714a  and  a1707a );
 a430a <=( a1700a  and  a1693a );
 a431a <=( a1686a  and  a1679a );
 a432a <=( a1672a  and  a1665a );
 a433a <=( a1658a  and  a1651a );
 a434a <=( a1644a  and  a1637a );
 a435a <=( a1630a  and  a1623a );
 a436a <=( a1616a  and  a1609a );
 a437a <=( a1602a  and  a1595a );
 a438a <=( a1588a  and  a1581a );
 a439a <=( a1574a  and  a1567a );
 a440a <=( a1560a  and  a1553a );
 a441a <=( a1546a  and  a1539a );
 a442a <=( a1532a  and  a1525a );
 a443a <=( a1518a  and  a1511a );
 a444a <=( a1504a  and  a1497a );
 a445a <=( a1490a  and  a1483a );
 a446a <=( a1478a  and  a1471a );
 a447a <=( a1466a  and  a1459a );
 a448a <=( a1454a  and  a1447a );
 a449a <=( a1442a  and  a1437a );
 a450a <=( a1432a  and  a1427a );
 a451a <=( a1422a  and  a1417a );
 a452a <=( a1412a  and  a1407a );
 a453a <=( a1402a  and  a1397a );
 a454a <=( a1392a  and  a1387a );
 a455a <=( a1382a  and  a1377a );
 a456a <=( a1374a  and  a1369a );
 a460a <=( a454a ) or ( a455a );
 a461a <=( a456a ) or ( a460a );
 a464a <=( a452a ) or ( a453a );
 a467a <=( a450a ) or ( a451a );
 a468a <=( a467a ) or ( a464a );
 a469a <=( a468a ) or ( a461a );
 a473a <=( a447a ) or ( a448a );
 a474a <=( a449a ) or ( a473a );
 a477a <=( a445a ) or ( a446a );
 a480a <=( a443a ) or ( a444a );
 a481a <=( a480a ) or ( a477a );
 a482a <=( a481a ) or ( a474a );
 a483a <=( a482a ) or ( a469a );
 a487a <=( a440a ) or ( a441a );
 a488a <=( a442a ) or ( a487a );
 a491a <=( a438a ) or ( a439a );
 a494a <=( a436a ) or ( a437a );
 a495a <=( a494a ) or ( a491a );
 a496a <=( a495a ) or ( a488a );
 a500a <=( a433a ) or ( a434a );
 a501a <=( a435a ) or ( a500a );
 a504a <=( a431a ) or ( a432a );
 a507a <=( a429a ) or ( a430a );
 a508a <=( a507a ) or ( a504a );
 a509a <=( a508a ) or ( a501a );
 a510a <=( a509a ) or ( a496a );
 a511a <=( a510a ) or ( a483a );
 a515a <=( a426a ) or ( a427a );
 a516a <=( a428a ) or ( a515a );
 a519a <=( a424a ) or ( a425a );
 a522a <=( a422a ) or ( a423a );
 a523a <=( a522a ) or ( a519a );
 a524a <=( a523a ) or ( a516a );
 a528a <=( a419a ) or ( a420a );
 a529a <=( a421a ) or ( a528a );
 a532a <=( a417a ) or ( a418a );
 a535a <=( a415a ) or ( a416a );
 a536a <=( a535a ) or ( a532a );
 a537a <=( a536a ) or ( a529a );
 a538a <=( a537a ) or ( a524a );
 a542a <=( a412a ) or ( a413a );
 a543a <=( a414a ) or ( a542a );
 a546a <=( a410a ) or ( a411a );
 a549a <=( a408a ) or ( a409a );
 a550a <=( a549a ) or ( a546a );
 a551a <=( a550a ) or ( a543a );
 a554a <=( a406a ) or ( a407a );
 a557a <=( a404a ) or ( a405a );
 a558a <=( a557a ) or ( a554a );
 a561a <=( a402a ) or ( a403a );
 a564a <=( a400a ) or ( a401a );
 a565a <=( a564a ) or ( a561a );
 a566a <=( a565a ) or ( a558a );
 a567a <=( a566a ) or ( a551a );
 a568a <=( a567a ) or ( a538a );
 a569a <=( a568a ) or ( a511a );
 a573a <=( a397a ) or ( a398a );
 a574a <=( a399a ) or ( a573a );
 a577a <=( a395a ) or ( a396a );
 a580a <=( a393a ) or ( a394a );
 a581a <=( a580a ) or ( a577a );
 a582a <=( a581a ) or ( a574a );
 a586a <=( a390a ) or ( a391a );
 a587a <=( a392a ) or ( a586a );
 a590a <=( a388a ) or ( a389a );
 a593a <=( a386a ) or ( a387a );
 a594a <=( a593a ) or ( a590a );
 a595a <=( a594a ) or ( a587a );
 a596a <=( a595a ) or ( a582a );
 a600a <=( a383a ) or ( a384a );
 a601a <=( a385a ) or ( a600a );
 a604a <=( a381a ) or ( a382a );
 a607a <=( a379a ) or ( a380a );
 a608a <=( a607a ) or ( a604a );
 a609a <=( a608a ) or ( a601a );
 a613a <=( a376a ) or ( a377a );
 a614a <=( a378a ) or ( a613a );
 a617a <=( a374a ) or ( a375a );
 a620a <=( a372a ) or ( a373a );
 a621a <=( a620a ) or ( a617a );
 a622a <=( a621a ) or ( a614a );
 a623a <=( a622a ) or ( a609a );
 a624a <=( a623a ) or ( a596a );
 a628a <=( a369a ) or ( a370a );
 a629a <=( a371a ) or ( a628a );
 a632a <=( a367a ) or ( a368a );
 a635a <=( a365a ) or ( a366a );
 a636a <=( a635a ) or ( a632a );
 a637a <=( a636a ) or ( a629a );
 a641a <=( a362a ) or ( a363a );
 a642a <=( a364a ) or ( a641a );
 a645a <=( a360a ) or ( a361a );
 a648a <=( a358a ) or ( a359a );
 a649a <=( a648a ) or ( a645a );
 a650a <=( a649a ) or ( a642a );
 a651a <=( a650a ) or ( a637a );
 a655a <=( a355a ) or ( a356a );
 a656a <=( a357a ) or ( a655a );
 a659a <=( a353a ) or ( a354a );
 a662a <=( a351a ) or ( a352a );
 a663a <=( a662a ) or ( a659a );
 a664a <=( a663a ) or ( a656a );
 a667a <=( a349a ) or ( a350a );
 a670a <=( a347a ) or ( a348a );
 a671a <=( a670a ) or ( a667a );
 a674a <=( a345a ) or ( a346a );
 a677a <=( a343a ) or ( a344a );
 a678a <=( a677a ) or ( a674a );
 a679a <=( a678a ) or ( a671a );
 a680a <=( a679a ) or ( a664a );
 a681a <=( a680a ) or ( a651a );
 a682a <=( a681a ) or ( a624a );
 a683a <=( a682a ) or ( a569a );
 a687a <=( a340a ) or ( a341a );
 a688a <=( a342a ) or ( a687a );
 a691a <=( a338a ) or ( a339a );
 a694a <=( a336a ) or ( a337a );
 a695a <=( a694a ) or ( a691a );
 a696a <=( a695a ) or ( a688a );
 a700a <=( a333a ) or ( a334a );
 a701a <=( a335a ) or ( a700a );
 a704a <=( a331a ) or ( a332a );
 a707a <=( a329a ) or ( a330a );
 a708a <=( a707a ) or ( a704a );
 a709a <=( a708a ) or ( a701a );
 a710a <=( a709a ) or ( a696a );
 a714a <=( a326a ) or ( a327a );
 a715a <=( a328a ) or ( a714a );
 a718a <=( a324a ) or ( a325a );
 a721a <=( a322a ) or ( a323a );
 a722a <=( a721a ) or ( a718a );
 a723a <=( a722a ) or ( a715a );
 a727a <=( a319a ) or ( a320a );
 a728a <=( a321a ) or ( a727a );
 a731a <=( a317a ) or ( a318a );
 a734a <=( a315a ) or ( a316a );
 a735a <=( a734a ) or ( a731a );
 a736a <=( a735a ) or ( a728a );
 a737a <=( a736a ) or ( a723a );
 a738a <=( a737a ) or ( a710a );
 a742a <=( a312a ) or ( a313a );
 a743a <=( a314a ) or ( a742a );
 a746a <=( a310a ) or ( a311a );
 a749a <=( a308a ) or ( a309a );
 a750a <=( a749a ) or ( a746a );
 a751a <=( a750a ) or ( a743a );
 a755a <=( a305a ) or ( a306a );
 a756a <=( a307a ) or ( a755a );
 a759a <=( a303a ) or ( a304a );
 a762a <=( a301a ) or ( a302a );
 a763a <=( a762a ) or ( a759a );
 a764a <=( a763a ) or ( a756a );
 a765a <=( a764a ) or ( a751a );
 a769a <=( a298a ) or ( a299a );
 a770a <=( a300a ) or ( a769a );
 a773a <=( a296a ) or ( a297a );
 a776a <=( a294a ) or ( a295a );
 a777a <=( a776a ) or ( a773a );
 a778a <=( a777a ) or ( a770a );
 a781a <=( a292a ) or ( a293a );
 a784a <=( a290a ) or ( a291a );
 a785a <=( a784a ) or ( a781a );
 a788a <=( a288a ) or ( a289a );
 a791a <=( a286a ) or ( a287a );
 a792a <=( a791a ) or ( a788a );
 a793a <=( a792a ) or ( a785a );
 a794a <=( a793a ) or ( a778a );
 a795a <=( a794a ) or ( a765a );
 a796a <=( a795a ) or ( a738a );
 a800a <=( a283a ) or ( a284a );
 a801a <=( a285a ) or ( a800a );
 a804a <=( a281a ) or ( a282a );
 a807a <=( a279a ) or ( a280a );
 a808a <=( a807a ) or ( a804a );
 a809a <=( a808a ) or ( a801a );
 a813a <=( a276a ) or ( a277a );
 a814a <=( a278a ) or ( a813a );
 a817a <=( a274a ) or ( a275a );
 a820a <=( a272a ) or ( a273a );
 a821a <=( a820a ) or ( a817a );
 a822a <=( a821a ) or ( a814a );
 a823a <=( a822a ) or ( a809a );
 a827a <=( a269a ) or ( a270a );
 a828a <=( a271a ) or ( a827a );
 a831a <=( a267a ) or ( a268a );
 a834a <=( a265a ) or ( a266a );
 a835a <=( a834a ) or ( a831a );
 a836a <=( a835a ) or ( a828a );
 a840a <=( a262a ) or ( a263a );
 a841a <=( a264a ) or ( a840a );
 a844a <=( a260a ) or ( a261a );
 a847a <=( a258a ) or ( a259a );
 a848a <=( a847a ) or ( a844a );
 a849a <=( a848a ) or ( a841a );
 a850a <=( a849a ) or ( a836a );
 a851a <=( a850a ) or ( a823a );
 a855a <=( a255a ) or ( a256a );
 a856a <=( a257a ) or ( a855a );
 a859a <=( a253a ) or ( a254a );
 a862a <=( a251a ) or ( a252a );
 a863a <=( a862a ) or ( a859a );
 a864a <=( a863a ) or ( a856a );
 a868a <=( a248a ) or ( a249a );
 a869a <=( a250a ) or ( a868a );
 a872a <=( a246a ) or ( a247a );
 a875a <=( a244a ) or ( a245a );
 a876a <=( a875a ) or ( a872a );
 a877a <=( a876a ) or ( a869a );
 a878a <=( a877a ) or ( a864a );
 a882a <=( a241a ) or ( a242a );
 a883a <=( a243a ) or ( a882a );
 a886a <=( a239a ) or ( a240a );
 a889a <=( a237a ) or ( a238a );
 a890a <=( a889a ) or ( a886a );
 a891a <=( a890a ) or ( a883a );
 a894a <=( a235a ) or ( a236a );
 a897a <=( a233a ) or ( a234a );
 a898a <=( a897a ) or ( a894a );
 a901a <=( a231a ) or ( a232a );
 a904a <=( a229a ) or ( a230a );
 a905a <=( a904a ) or ( a901a );
 a906a <=( a905a ) or ( a898a );
 a907a <=( a906a ) or ( a891a );
 a908a <=( a907a ) or ( a878a );
 a909a <=( a908a ) or ( a851a );
 a910a <=( a909a ) or ( a796a );
 a911a <=( a910a ) or ( a683a );
 a915a <=( a226a ) or ( a227a );
 a916a <=( a228a ) or ( a915a );
 a919a <=( a224a ) or ( a225a );
 a922a <=( a222a ) or ( a223a );
 a923a <=( a922a ) or ( a919a );
 a924a <=( a923a ) or ( a916a );
 a928a <=( a219a ) or ( a220a );
 a929a <=( a221a ) or ( a928a );
 a932a <=( a217a ) or ( a218a );
 a935a <=( a215a ) or ( a216a );
 a936a <=( a935a ) or ( a932a );
 a937a <=( a936a ) or ( a929a );
 a938a <=( a937a ) or ( a924a );
 a942a <=( a212a ) or ( a213a );
 a943a <=( a214a ) or ( a942a );
 a946a <=( a210a ) or ( a211a );
 a949a <=( a208a ) or ( a209a );
 a950a <=( a949a ) or ( a946a );
 a951a <=( a950a ) or ( a943a );
 a955a <=( a205a ) or ( a206a );
 a956a <=( a207a ) or ( a955a );
 a959a <=( a203a ) or ( a204a );
 a962a <=( a201a ) or ( a202a );
 a963a <=( a962a ) or ( a959a );
 a964a <=( a963a ) or ( a956a );
 a965a <=( a964a ) or ( a951a );
 a966a <=( a965a ) or ( a938a );
 a970a <=( a198a ) or ( a199a );
 a971a <=( a200a ) or ( a970a );
 a974a <=( a196a ) or ( a197a );
 a977a <=( a194a ) or ( a195a );
 a978a <=( a977a ) or ( a974a );
 a979a <=( a978a ) or ( a971a );
 a983a <=( a191a ) or ( a192a );
 a984a <=( a193a ) or ( a983a );
 a987a <=( a189a ) or ( a190a );
 a990a <=( a187a ) or ( a188a );
 a991a <=( a990a ) or ( a987a );
 a992a <=( a991a ) or ( a984a );
 a993a <=( a992a ) or ( a979a );
 a997a <=( a184a ) or ( a185a );
 a998a <=( a186a ) or ( a997a );
 a1001a <=( a182a ) or ( a183a );
 a1004a <=( a180a ) or ( a181a );
 a1005a <=( a1004a ) or ( a1001a );
 a1006a <=( a1005a ) or ( a998a );
 a1009a <=( a178a ) or ( a179a );
 a1012a <=( a176a ) or ( a177a );
 a1013a <=( a1012a ) or ( a1009a );
 a1016a <=( a174a ) or ( a175a );
 a1019a <=( a172a ) or ( a173a );
 a1020a <=( a1019a ) or ( a1016a );
 a1021a <=( a1020a ) or ( a1013a );
 a1022a <=( a1021a ) or ( a1006a );
 a1023a <=( a1022a ) or ( a993a );
 a1024a <=( a1023a ) or ( a966a );
 a1028a <=( a169a ) or ( a170a );
 a1029a <=( a171a ) or ( a1028a );
 a1032a <=( a167a ) or ( a168a );
 a1035a <=( a165a ) or ( a166a );
 a1036a <=( a1035a ) or ( a1032a );
 a1037a <=( a1036a ) or ( a1029a );
 a1041a <=( a162a ) or ( a163a );
 a1042a <=( a164a ) or ( a1041a );
 a1045a <=( a160a ) or ( a161a );
 a1048a <=( a158a ) or ( a159a );
 a1049a <=( a1048a ) or ( a1045a );
 a1050a <=( a1049a ) or ( a1042a );
 a1051a <=( a1050a ) or ( a1037a );
 a1055a <=( a155a ) or ( a156a );
 a1056a <=( a157a ) or ( a1055a );
 a1059a <=( a153a ) or ( a154a );
 a1062a <=( a151a ) or ( a152a );
 a1063a <=( a1062a ) or ( a1059a );
 a1064a <=( a1063a ) or ( a1056a );
 a1068a <=( a148a ) or ( a149a );
 a1069a <=( a150a ) or ( a1068a );
 a1072a <=( a146a ) or ( a147a );
 a1075a <=( a144a ) or ( a145a );
 a1076a <=( a1075a ) or ( a1072a );
 a1077a <=( a1076a ) or ( a1069a );
 a1078a <=( a1077a ) or ( a1064a );
 a1079a <=( a1078a ) or ( a1051a );
 a1083a <=( a141a ) or ( a142a );
 a1084a <=( a143a ) or ( a1083a );
 a1087a <=( a139a ) or ( a140a );
 a1090a <=( a137a ) or ( a138a );
 a1091a <=( a1090a ) or ( a1087a );
 a1092a <=( a1091a ) or ( a1084a );
 a1096a <=( a134a ) or ( a135a );
 a1097a <=( a136a ) or ( a1096a );
 a1100a <=( a132a ) or ( a133a );
 a1103a <=( a130a ) or ( a131a );
 a1104a <=( a1103a ) or ( a1100a );
 a1105a <=( a1104a ) or ( a1097a );
 a1106a <=( a1105a ) or ( a1092a );
 a1110a <=( a127a ) or ( a128a );
 a1111a <=( a129a ) or ( a1110a );
 a1114a <=( a125a ) or ( a126a );
 a1117a <=( a123a ) or ( a124a );
 a1118a <=( a1117a ) or ( a1114a );
 a1119a <=( a1118a ) or ( a1111a );
 a1122a <=( a121a ) or ( a122a );
 a1125a <=( a119a ) or ( a120a );
 a1126a <=( a1125a ) or ( a1122a );
 a1129a <=( a117a ) or ( a118a );
 a1132a <=( a115a ) or ( a116a );
 a1133a <=( a1132a ) or ( a1129a );
 a1134a <=( a1133a ) or ( a1126a );
 a1135a <=( a1134a ) or ( a1119a );
 a1136a <=( a1135a ) or ( a1106a );
 a1137a <=( a1136a ) or ( a1079a );
 a1138a <=( a1137a ) or ( a1024a );
 a1142a <=( a112a ) or ( a113a );
 a1143a <=( a114a ) or ( a1142a );
 a1146a <=( a110a ) or ( a111a );
 a1149a <=( a108a ) or ( a109a );
 a1150a <=( a1149a ) or ( a1146a );
 a1151a <=( a1150a ) or ( a1143a );
 a1155a <=( a105a ) or ( a106a );
 a1156a <=( a107a ) or ( a1155a );
 a1159a <=( a103a ) or ( a104a );
 a1162a <=( a101a ) or ( a102a );
 a1163a <=( a1162a ) or ( a1159a );
 a1164a <=( a1163a ) or ( a1156a );
 a1165a <=( a1164a ) or ( a1151a );
 a1169a <=( a98a ) or ( a99a );
 a1170a <=( a100a ) or ( a1169a );
 a1173a <=( a96a ) or ( a97a );
 a1176a <=( a94a ) or ( a95a );
 a1177a <=( a1176a ) or ( a1173a );
 a1178a <=( a1177a ) or ( a1170a );
 a1182a <=( a91a ) or ( a92a );
 a1183a <=( a93a ) or ( a1182a );
 a1186a <=( a89a ) or ( a90a );
 a1189a <=( a87a ) or ( a88a );
 a1190a <=( a1189a ) or ( a1186a );
 a1191a <=( a1190a ) or ( a1183a );
 a1192a <=( a1191a ) or ( a1178a );
 a1193a <=( a1192a ) or ( a1165a );
 a1197a <=( a84a ) or ( a85a );
 a1198a <=( a86a ) or ( a1197a );
 a1201a <=( a82a ) or ( a83a );
 a1204a <=( a80a ) or ( a81a );
 a1205a <=( a1204a ) or ( a1201a );
 a1206a <=( a1205a ) or ( a1198a );
 a1210a <=( a77a ) or ( a78a );
 a1211a <=( a79a ) or ( a1210a );
 a1214a <=( a75a ) or ( a76a );
 a1217a <=( a73a ) or ( a74a );
 a1218a <=( a1217a ) or ( a1214a );
 a1219a <=( a1218a ) or ( a1211a );
 a1220a <=( a1219a ) or ( a1206a );
 a1224a <=( a70a ) or ( a71a );
 a1225a <=( a72a ) or ( a1224a );
 a1228a <=( a68a ) or ( a69a );
 a1231a <=( a66a ) or ( a67a );
 a1232a <=( a1231a ) or ( a1228a );
 a1233a <=( a1232a ) or ( a1225a );
 a1236a <=( a64a ) or ( a65a );
 a1239a <=( a62a ) or ( a63a );
 a1240a <=( a1239a ) or ( a1236a );
 a1243a <=( a60a ) or ( a61a );
 a1246a <=( a58a ) or ( a59a );
 a1247a <=( a1246a ) or ( a1243a );
 a1248a <=( a1247a ) or ( a1240a );
 a1249a <=( a1248a ) or ( a1233a );
 a1250a <=( a1249a ) or ( a1220a );
 a1251a <=( a1250a ) or ( a1193a );
 a1255a <=( a55a ) or ( a56a );
 a1256a <=( a57a ) or ( a1255a );
 a1259a <=( a53a ) or ( a54a );
 a1262a <=( a51a ) or ( a52a );
 a1263a <=( a1262a ) or ( a1259a );
 a1264a <=( a1263a ) or ( a1256a );
 a1268a <=( a48a ) or ( a49a );
 a1269a <=( a50a ) or ( a1268a );
 a1272a <=( a46a ) or ( a47a );
 a1275a <=( a44a ) or ( a45a );
 a1276a <=( a1275a ) or ( a1272a );
 a1277a <=( a1276a ) or ( a1269a );
 a1278a <=( a1277a ) or ( a1264a );
 a1282a <=( a41a ) or ( a42a );
 a1283a <=( a43a ) or ( a1282a );
 a1286a <=( a39a ) or ( a40a );
 a1289a <=( a37a ) or ( a38a );
 a1290a <=( a1289a ) or ( a1286a );
 a1291a <=( a1290a ) or ( a1283a );
 a1295a <=( a34a ) or ( a35a );
 a1296a <=( a36a ) or ( a1295a );
 a1299a <=( a32a ) or ( a33a );
 a1302a <=( a30a ) or ( a31a );
 a1303a <=( a1302a ) or ( a1299a );
 a1304a <=( a1303a ) or ( a1296a );
 a1305a <=( a1304a ) or ( a1291a );
 a1306a <=( a1305a ) or ( a1278a );
 a1310a <=( a27a ) or ( a28a );
 a1311a <=( a29a ) or ( a1310a );
 a1314a <=( a25a ) or ( a26a );
 a1317a <=( a23a ) or ( a24a );
 a1318a <=( a1317a ) or ( a1314a );
 a1319a <=( a1318a ) or ( a1311a );
 a1323a <=( a20a ) or ( a21a );
 a1324a <=( a22a ) or ( a1323a );
 a1327a <=( a18a ) or ( a19a );
 a1330a <=( a16a ) or ( a17a );
 a1331a <=( a1330a ) or ( a1327a );
 a1332a <=( a1331a ) or ( a1324a );
 a1333a <=( a1332a ) or ( a1319a );
 a1337a <=( a13a ) or ( a14a );
 a1338a <=( a15a ) or ( a1337a );
 a1341a <=( a11a ) or ( a12a );
 a1344a <=( a9a ) or ( a10a );
 a1345a <=( a1344a ) or ( a1341a );
 a1346a <=( a1345a ) or ( a1338a );
 a1349a <=( a7a ) or ( a8a );
 a1352a <=( a5a ) or ( a6a );
 a1353a <=( a1352a ) or ( a1349a );
 a1356a <=( a3a ) or ( a4a );
 a1359a <=( a1a ) or ( a2a );
 a1360a <=( a1359a ) or ( a1356a );
 a1361a <=( a1360a ) or ( a1353a );
 a1362a <=( a1361a ) or ( a1346a );
 a1363a <=( a1362a ) or ( a1333a );
 a1364a <=( a1363a ) or ( a1306a );
 a1365a <=( a1364a ) or ( a1251a );
 a1366a <=( a1365a ) or ( a1138a );
 a1369a <=( (not A167)  and  A170 );
 a1373a <=( A200  and  (not A199) );
 a1374a <=( (not A166)  and  a1373a );
 a1377a <=( (not A167)  and  (not A169) );
 a1381a <=( A200  and  (not A199) );
 a1382a <=( (not A166)  and  a1381a );
 a1386a <=( A167  and  (not A168) );
 a1387a <=( A170  and  a1386a );
 a1391a <=( A200  and  (not A199) );
 a1392a <=( A166  and  a1391a );
 a1396a <=( A167  and  (not A168) );
 a1397a <=( (not A170)  and  a1396a );
 a1401a <=( A200  and  (not A199) );
 a1402a <=( (not A166)  and  a1401a );
 a1406a <=( (not A167)  and  (not A168) );
 a1407a <=( (not A170)  and  a1406a );
 a1411a <=( A200  and  (not A199) );
 a1412a <=( A166  and  a1411a );
 a1416a <=( A167  and  (not A168) );
 a1417a <=( A169  and  a1416a );
 a1421a <=( A200  and  (not A199) );
 a1422a <=( (not A166)  and  a1421a );
 a1426a <=( (not A167)  and  (not A168) );
 a1427a <=( A169  and  a1426a );
 a1431a <=( A200  and  (not A199) );
 a1432a <=( A166  and  a1431a );
 a1436a <=( A167  and  (not A168) );
 a1437a <=( (not A169)  and  a1436a );
 a1441a <=( A200  and  (not A199) );
 a1442a <=( A166  and  a1441a );
 a1446a <=( (not A166)  and  (not A167) );
 a1447a <=( A170  and  a1446a );
 a1450a <=( (not A200)  and  A199 );
 a1453a <=( A202  and  A201 );
 a1454a <=( a1453a  and  a1450a );
 a1458a <=( (not A166)  and  (not A167) );
 a1459a <=( A170  and  a1458a );
 a1462a <=( (not A200)  and  A199 );
 a1465a <=( A203  and  A201 );
 a1466a <=( a1465a  and  a1462a );
 a1470a <=( (not A166)  and  (not A167) );
 a1471a <=( (not A169)  and  a1470a );
 a1474a <=( (not A200)  and  A199 );
 a1477a <=( A202  and  A201 );
 a1478a <=( a1477a  and  a1474a );
 a1482a <=( (not A166)  and  (not A167) );
 a1483a <=( (not A169)  and  a1482a );
 a1486a <=( (not A200)  and  A199 );
 a1489a <=( A203  and  A201 );
 a1490a <=( a1489a  and  a1486a );
 a1493a <=( A166  and  A168 );
 a1496a <=( (not A201)  and  A199 );
 a1497a <=( a1496a  and  a1493a );
 a1500a <=( A233  and  (not A232) );
 a1503a <=( A299  and  (not A298) );
 a1504a <=( a1503a  and  a1500a );
 a1507a <=( A166  and  A168 );
 a1510a <=( (not A201)  and  A199 );
 a1511a <=( a1510a  and  a1507a );
 a1514a <=( A233  and  (not A232) );
 a1517a <=( A266  and  (not A265) );
 a1518a <=( a1517a  and  a1514a );
 a1521a <=( A166  and  A168 );
 a1524a <=( A200  and  A199 );
 a1525a <=( a1524a  and  a1521a );
 a1528a <=( A233  and  (not A232) );
 a1531a <=( A299  and  (not A298) );
 a1532a <=( a1531a  and  a1528a );
 a1535a <=( A166  and  A168 );
 a1538a <=( A200  and  A199 );
 a1539a <=( a1538a  and  a1535a );
 a1542a <=( A233  and  (not A232) );
 a1545a <=( A266  and  (not A265) );
 a1546a <=( a1545a  and  a1542a );
 a1549a <=( A166  and  A168 );
 a1552a <=( (not A200)  and  (not A199) );
 a1553a <=( a1552a  and  a1549a );
 a1556a <=( A233  and  (not A232) );
 a1559a <=( A299  and  (not A298) );
 a1560a <=( a1559a  and  a1556a );
 a1563a <=( A166  and  A168 );
 a1566a <=( (not A200)  and  (not A199) );
 a1567a <=( a1566a  and  a1563a );
 a1570a <=( A233  and  (not A232) );
 a1573a <=( A266  and  (not A265) );
 a1574a <=( a1573a  and  a1570a );
 a1577a <=( A167  and  A168 );
 a1580a <=( (not A201)  and  A199 );
 a1581a <=( a1580a  and  a1577a );
 a1584a <=( A233  and  (not A232) );
 a1587a <=( A299  and  (not A298) );
 a1588a <=( a1587a  and  a1584a );
 a1591a <=( A167  and  A168 );
 a1594a <=( (not A201)  and  A199 );
 a1595a <=( a1594a  and  a1591a );
 a1598a <=( A233  and  (not A232) );
 a1601a <=( A266  and  (not A265) );
 a1602a <=( a1601a  and  a1598a );
 a1605a <=( A167  and  A168 );
 a1608a <=( A200  and  A199 );
 a1609a <=( a1608a  and  a1605a );
 a1612a <=( A233  and  (not A232) );
 a1615a <=( A299  and  (not A298) );
 a1616a <=( a1615a  and  a1612a );
 a1619a <=( A167  and  A168 );
 a1622a <=( A200  and  A199 );
 a1623a <=( a1622a  and  a1619a );
 a1626a <=( A233  and  (not A232) );
 a1629a <=( A266  and  (not A265) );
 a1630a <=( a1629a  and  a1626a );
 a1633a <=( A167  and  A168 );
 a1636a <=( (not A200)  and  (not A199) );
 a1637a <=( a1636a  and  a1633a );
 a1640a <=( A233  and  (not A232) );
 a1643a <=( A299  and  (not A298) );
 a1644a <=( a1643a  and  a1640a );
 a1647a <=( A167  and  A168 );
 a1650a <=( (not A200)  and  (not A199) );
 a1651a <=( a1650a  and  a1647a );
 a1654a <=( A233  and  (not A232) );
 a1657a <=( A266  and  (not A265) );
 a1658a <=( a1657a  and  a1654a );
 a1661a <=( (not A168)  and  A170 );
 a1664a <=( A166  and  A167 );
 a1665a <=( a1664a  and  a1661a );
 a1668a <=( (not A200)  and  A199 );
 a1671a <=( A202  and  A201 );
 a1672a <=( a1671a  and  a1668a );
 a1675a <=( (not A168)  and  A170 );
 a1678a <=( A166  and  A167 );
 a1679a <=( a1678a  and  a1675a );
 a1682a <=( (not A200)  and  A199 );
 a1685a <=( A203  and  A201 );
 a1686a <=( a1685a  and  a1682a );
 a1689a <=( (not A168)  and  (not A170) );
 a1692a <=( (not A166)  and  A167 );
 a1693a <=( a1692a  and  a1689a );
 a1696a <=( (not A200)  and  A199 );
 a1699a <=( A202  and  A201 );
 a1700a <=( a1699a  and  a1696a );
 a1703a <=( (not A168)  and  (not A170) );
 a1706a <=( (not A166)  and  A167 );
 a1707a <=( a1706a  and  a1703a );
 a1710a <=( (not A200)  and  A199 );
 a1713a <=( A203  and  A201 );
 a1714a <=( a1713a  and  a1710a );
 a1717a <=( (not A168)  and  (not A170) );
 a1720a <=( A166  and  (not A167) );
 a1721a <=( a1720a  and  a1717a );
 a1724a <=( (not A200)  and  A199 );
 a1727a <=( A202  and  A201 );
 a1728a <=( a1727a  and  a1724a );
 a1731a <=( (not A168)  and  (not A170) );
 a1734a <=( A166  and  (not A167) );
 a1735a <=( a1734a  and  a1731a );
 a1738a <=( (not A200)  and  A199 );
 a1741a <=( A203  and  A201 );
 a1742a <=( a1741a  and  a1738a );
 a1745a <=( (not A168)  and  A169 );
 a1748a <=( (not A166)  and  A167 );
 a1749a <=( a1748a  and  a1745a );
 a1752a <=( (not A200)  and  A199 );
 a1755a <=( A202  and  A201 );
 a1756a <=( a1755a  and  a1752a );
 a1759a <=( (not A168)  and  A169 );
 a1762a <=( (not A166)  and  A167 );
 a1763a <=( a1762a  and  a1759a );
 a1766a <=( (not A200)  and  A199 );
 a1769a <=( A203  and  A201 );
 a1770a <=( a1769a  and  a1766a );
 a1773a <=( (not A168)  and  A169 );
 a1776a <=( A166  and  (not A167) );
 a1777a <=( a1776a  and  a1773a );
 a1780a <=( (not A200)  and  A199 );
 a1783a <=( A202  and  A201 );
 a1784a <=( a1783a  and  a1780a );
 a1787a <=( (not A168)  and  A169 );
 a1790a <=( A166  and  (not A167) );
 a1791a <=( a1790a  and  a1787a );
 a1794a <=( (not A200)  and  A199 );
 a1797a <=( A203  and  A201 );
 a1798a <=( a1797a  and  a1794a );
 a1801a <=( (not A168)  and  (not A169) );
 a1804a <=( A166  and  A167 );
 a1805a <=( a1804a  and  a1801a );
 a1808a <=( (not A200)  and  A199 );
 a1811a <=( A202  and  A201 );
 a1812a <=( a1811a  and  a1808a );
 a1815a <=( (not A168)  and  (not A169) );
 a1818a <=( A166  and  A167 );
 a1819a <=( a1818a  and  a1815a );
 a1822a <=( (not A200)  and  A199 );
 a1825a <=( A203  and  A201 );
 a1826a <=( a1825a  and  a1822a );
 a1829a <=( A166  and  A168 );
 a1832a <=( (not A202)  and  A199 );
 a1833a <=( a1832a  and  a1829a );
 a1836a <=( (not A232)  and  (not A203) );
 a1840a <=( A299  and  (not A298) );
 a1841a <=( A233  and  a1840a );
 a1842a <=( a1841a  and  a1836a );
 a1845a <=( A166  and  A168 );
 a1848a <=( (not A202)  and  A199 );
 a1849a <=( a1848a  and  a1845a );
 a1852a <=( (not A232)  and  (not A203) );
 a1856a <=( A266  and  (not A265) );
 a1857a <=( A233  and  a1856a );
 a1858a <=( a1857a  and  a1852a );
 a1861a <=( A167  and  A168 );
 a1864a <=( (not A202)  and  A199 );
 a1865a <=( a1864a  and  a1861a );
 a1868a <=( (not A232)  and  (not A203) );
 a1872a <=( A299  and  (not A298) );
 a1873a <=( A233  and  a1872a );
 a1874a <=( a1873a  and  a1868a );
 a1877a <=( A167  and  A168 );
 a1880a <=( (not A202)  and  A199 );
 a1881a <=( a1880a  and  a1877a );
 a1884a <=( (not A232)  and  (not A203) );
 a1888a <=( A266  and  (not A265) );
 a1889a <=( A233  and  a1888a );
 a1890a <=( a1889a  and  a1884a );
 a1893a <=( A166  and  A168 );
 a1897a <=( (not A232)  and  (not A201) );
 a1898a <=( A199  and  a1897a );
 a1899a <=( a1898a  and  a1893a );
 a1902a <=( A298  and  A233 );
 a1906a <=( A301  and  A300 );
 a1907a <=( (not A299)  and  a1906a );
 a1908a <=( a1907a  and  a1902a );
 a1911a <=( A166  and  A168 );
 a1915a <=( (not A232)  and  (not A201) );
 a1916a <=( A199  and  a1915a );
 a1917a <=( a1916a  and  a1911a );
 a1920a <=( A298  and  A233 );
 a1924a <=( A302  and  A300 );
 a1925a <=( (not A299)  and  a1924a );
 a1926a <=( a1925a  and  a1920a );
 a1929a <=( A166  and  A168 );
 a1933a <=( (not A232)  and  (not A201) );
 a1934a <=( A199  and  a1933a );
 a1935a <=( a1934a  and  a1929a );
 a1938a <=( A265  and  A233 );
 a1942a <=( A268  and  A267 );
 a1943a <=( (not A266)  and  a1942a );
 a1944a <=( a1943a  and  a1938a );
 a1947a <=( A166  and  A168 );
 a1951a <=( (not A232)  and  (not A201) );
 a1952a <=( A199  and  a1951a );
 a1953a <=( a1952a  and  a1947a );
 a1956a <=( A265  and  A233 );
 a1960a <=( A269  and  A267 );
 a1961a <=( (not A266)  and  a1960a );
 a1962a <=( a1961a  and  a1956a );
 a1965a <=( A166  and  A168 );
 a1969a <=( A232  and  (not A201) );
 a1970a <=( A199  and  a1969a );
 a1971a <=( a1970a  and  a1965a );
 a1974a <=( A234  and  (not A233) );
 a1978a <=( A299  and  (not A298) );
 a1979a <=( A235  and  a1978a );
 a1980a <=( a1979a  and  a1974a );
 a1983a <=( A166  and  A168 );
 a1987a <=( A232  and  (not A201) );
 a1988a <=( A199  and  a1987a );
 a1989a <=( a1988a  and  a1983a );
 a1992a <=( A234  and  (not A233) );
 a1996a <=( A266  and  (not A265) );
 a1997a <=( A235  and  a1996a );
 a1998a <=( a1997a  and  a1992a );
 a2001a <=( A166  and  A168 );
 a2005a <=( A232  and  (not A201) );
 a2006a <=( A199  and  a2005a );
 a2007a <=( a2006a  and  a2001a );
 a2010a <=( A234  and  (not A233) );
 a2014a <=( A299  and  (not A298) );
 a2015a <=( A236  and  a2014a );
 a2016a <=( a2015a  and  a2010a );
 a2019a <=( A166  and  A168 );
 a2023a <=( A232  and  (not A201) );
 a2024a <=( A199  and  a2023a );
 a2025a <=( a2024a  and  a2019a );
 a2028a <=( A234  and  (not A233) );
 a2032a <=( A266  and  (not A265) );
 a2033a <=( A236  and  a2032a );
 a2034a <=( a2033a  and  a2028a );
 a2037a <=( A166  and  A168 );
 a2041a <=( (not A232)  and  A200 );
 a2042a <=( A199  and  a2041a );
 a2043a <=( a2042a  and  a2037a );
 a2046a <=( A298  and  A233 );
 a2050a <=( A301  and  A300 );
 a2051a <=( (not A299)  and  a2050a );
 a2052a <=( a2051a  and  a2046a );
 a2055a <=( A166  and  A168 );
 a2059a <=( (not A232)  and  A200 );
 a2060a <=( A199  and  a2059a );
 a2061a <=( a2060a  and  a2055a );
 a2064a <=( A298  and  A233 );
 a2068a <=( A302  and  A300 );
 a2069a <=( (not A299)  and  a2068a );
 a2070a <=( a2069a  and  a2064a );
 a2073a <=( A166  and  A168 );
 a2077a <=( (not A232)  and  A200 );
 a2078a <=( A199  and  a2077a );
 a2079a <=( a2078a  and  a2073a );
 a2082a <=( A265  and  A233 );
 a2086a <=( A268  and  A267 );
 a2087a <=( (not A266)  and  a2086a );
 a2088a <=( a2087a  and  a2082a );
 a2091a <=( A166  and  A168 );
 a2095a <=( (not A232)  and  A200 );
 a2096a <=( A199  and  a2095a );
 a2097a <=( a2096a  and  a2091a );
 a2100a <=( A265  and  A233 );
 a2104a <=( A269  and  A267 );
 a2105a <=( (not A266)  and  a2104a );
 a2106a <=( a2105a  and  a2100a );
 a2109a <=( A166  and  A168 );
 a2113a <=( A232  and  A200 );
 a2114a <=( A199  and  a2113a );
 a2115a <=( a2114a  and  a2109a );
 a2118a <=( A234  and  (not A233) );
 a2122a <=( A299  and  (not A298) );
 a2123a <=( A235  and  a2122a );
 a2124a <=( a2123a  and  a2118a );
 a2127a <=( A166  and  A168 );
 a2131a <=( A232  and  A200 );
 a2132a <=( A199  and  a2131a );
 a2133a <=( a2132a  and  a2127a );
 a2136a <=( A234  and  (not A233) );
 a2140a <=( A266  and  (not A265) );
 a2141a <=( A235  and  a2140a );
 a2142a <=( a2141a  and  a2136a );
 a2145a <=( A166  and  A168 );
 a2149a <=( A232  and  A200 );
 a2150a <=( A199  and  a2149a );
 a2151a <=( a2150a  and  a2145a );
 a2154a <=( A234  and  (not A233) );
 a2158a <=( A299  and  (not A298) );
 a2159a <=( A236  and  a2158a );
 a2160a <=( a2159a  and  a2154a );
 a2163a <=( A166  and  A168 );
 a2167a <=( A232  and  A200 );
 a2168a <=( A199  and  a2167a );
 a2169a <=( a2168a  and  a2163a );
 a2172a <=( A234  and  (not A233) );
 a2176a <=( A266  and  (not A265) );
 a2177a <=( A236  and  a2176a );
 a2178a <=( a2177a  and  a2172a );
 a2181a <=( A166  and  A168 );
 a2185a <=( (not A232)  and  (not A200) );
 a2186a <=( (not A199)  and  a2185a );
 a2187a <=( a2186a  and  a2181a );
 a2190a <=( A298  and  A233 );
 a2194a <=( A301  and  A300 );
 a2195a <=( (not A299)  and  a2194a );
 a2196a <=( a2195a  and  a2190a );
 a2199a <=( A166  and  A168 );
 a2203a <=( (not A232)  and  (not A200) );
 a2204a <=( (not A199)  and  a2203a );
 a2205a <=( a2204a  and  a2199a );
 a2208a <=( A298  and  A233 );
 a2212a <=( A302  and  A300 );
 a2213a <=( (not A299)  and  a2212a );
 a2214a <=( a2213a  and  a2208a );
 a2217a <=( A166  and  A168 );
 a2221a <=( (not A232)  and  (not A200) );
 a2222a <=( (not A199)  and  a2221a );
 a2223a <=( a2222a  and  a2217a );
 a2226a <=( A265  and  A233 );
 a2230a <=( A268  and  A267 );
 a2231a <=( (not A266)  and  a2230a );
 a2232a <=( a2231a  and  a2226a );
 a2235a <=( A166  and  A168 );
 a2239a <=( (not A232)  and  (not A200) );
 a2240a <=( (not A199)  and  a2239a );
 a2241a <=( a2240a  and  a2235a );
 a2244a <=( A265  and  A233 );
 a2248a <=( A269  and  A267 );
 a2249a <=( (not A266)  and  a2248a );
 a2250a <=( a2249a  and  a2244a );
 a2253a <=( A166  and  A168 );
 a2257a <=( A232  and  (not A200) );
 a2258a <=( (not A199)  and  a2257a );
 a2259a <=( a2258a  and  a2253a );
 a2262a <=( A234  and  (not A233) );
 a2266a <=( A299  and  (not A298) );
 a2267a <=( A235  and  a2266a );
 a2268a <=( a2267a  and  a2262a );
 a2271a <=( A166  and  A168 );
 a2275a <=( A232  and  (not A200) );
 a2276a <=( (not A199)  and  a2275a );
 a2277a <=( a2276a  and  a2271a );
 a2280a <=( A234  and  (not A233) );
 a2284a <=( A266  and  (not A265) );
 a2285a <=( A235  and  a2284a );
 a2286a <=( a2285a  and  a2280a );
 a2289a <=( A166  and  A168 );
 a2293a <=( A232  and  (not A200) );
 a2294a <=( (not A199)  and  a2293a );
 a2295a <=( a2294a  and  a2289a );
 a2298a <=( A234  and  (not A233) );
 a2302a <=( A299  and  (not A298) );
 a2303a <=( A236  and  a2302a );
 a2304a <=( a2303a  and  a2298a );
 a2307a <=( A166  and  A168 );
 a2311a <=( A232  and  (not A200) );
 a2312a <=( (not A199)  and  a2311a );
 a2313a <=( a2312a  and  a2307a );
 a2316a <=( A234  and  (not A233) );
 a2320a <=( A266  and  (not A265) );
 a2321a <=( A236  and  a2320a );
 a2322a <=( a2321a  and  a2316a );
 a2325a <=( A167  and  A168 );
 a2329a <=( (not A232)  and  (not A201) );
 a2330a <=( A199  and  a2329a );
 a2331a <=( a2330a  and  a2325a );
 a2334a <=( A298  and  A233 );
 a2338a <=( A301  and  A300 );
 a2339a <=( (not A299)  and  a2338a );
 a2340a <=( a2339a  and  a2334a );
 a2343a <=( A167  and  A168 );
 a2347a <=( (not A232)  and  (not A201) );
 a2348a <=( A199  and  a2347a );
 a2349a <=( a2348a  and  a2343a );
 a2352a <=( A298  and  A233 );
 a2356a <=( A302  and  A300 );
 a2357a <=( (not A299)  and  a2356a );
 a2358a <=( a2357a  and  a2352a );
 a2361a <=( A167  and  A168 );
 a2365a <=( (not A232)  and  (not A201) );
 a2366a <=( A199  and  a2365a );
 a2367a <=( a2366a  and  a2361a );
 a2370a <=( A265  and  A233 );
 a2374a <=( A268  and  A267 );
 a2375a <=( (not A266)  and  a2374a );
 a2376a <=( a2375a  and  a2370a );
 a2379a <=( A167  and  A168 );
 a2383a <=( (not A232)  and  (not A201) );
 a2384a <=( A199  and  a2383a );
 a2385a <=( a2384a  and  a2379a );
 a2388a <=( A265  and  A233 );
 a2392a <=( A269  and  A267 );
 a2393a <=( (not A266)  and  a2392a );
 a2394a <=( a2393a  and  a2388a );
 a2397a <=( A167  and  A168 );
 a2401a <=( A232  and  (not A201) );
 a2402a <=( A199  and  a2401a );
 a2403a <=( a2402a  and  a2397a );
 a2406a <=( A234  and  (not A233) );
 a2410a <=( A299  and  (not A298) );
 a2411a <=( A235  and  a2410a );
 a2412a <=( a2411a  and  a2406a );
 a2415a <=( A167  and  A168 );
 a2419a <=( A232  and  (not A201) );
 a2420a <=( A199  and  a2419a );
 a2421a <=( a2420a  and  a2415a );
 a2424a <=( A234  and  (not A233) );
 a2428a <=( A266  and  (not A265) );
 a2429a <=( A235  and  a2428a );
 a2430a <=( a2429a  and  a2424a );
 a2433a <=( A167  and  A168 );
 a2437a <=( A232  and  (not A201) );
 a2438a <=( A199  and  a2437a );
 a2439a <=( a2438a  and  a2433a );
 a2442a <=( A234  and  (not A233) );
 a2446a <=( A299  and  (not A298) );
 a2447a <=( A236  and  a2446a );
 a2448a <=( a2447a  and  a2442a );
 a2451a <=( A167  and  A168 );
 a2455a <=( A232  and  (not A201) );
 a2456a <=( A199  and  a2455a );
 a2457a <=( a2456a  and  a2451a );
 a2460a <=( A234  and  (not A233) );
 a2464a <=( A266  and  (not A265) );
 a2465a <=( A236  and  a2464a );
 a2466a <=( a2465a  and  a2460a );
 a2469a <=( A167  and  A168 );
 a2473a <=( (not A232)  and  A200 );
 a2474a <=( A199  and  a2473a );
 a2475a <=( a2474a  and  a2469a );
 a2478a <=( A298  and  A233 );
 a2482a <=( A301  and  A300 );
 a2483a <=( (not A299)  and  a2482a );
 a2484a <=( a2483a  and  a2478a );
 a2487a <=( A167  and  A168 );
 a2491a <=( (not A232)  and  A200 );
 a2492a <=( A199  and  a2491a );
 a2493a <=( a2492a  and  a2487a );
 a2496a <=( A298  and  A233 );
 a2500a <=( A302  and  A300 );
 a2501a <=( (not A299)  and  a2500a );
 a2502a <=( a2501a  and  a2496a );
 a2505a <=( A167  and  A168 );
 a2509a <=( (not A232)  and  A200 );
 a2510a <=( A199  and  a2509a );
 a2511a <=( a2510a  and  a2505a );
 a2514a <=( A265  and  A233 );
 a2518a <=( A268  and  A267 );
 a2519a <=( (not A266)  and  a2518a );
 a2520a <=( a2519a  and  a2514a );
 a2523a <=( A167  and  A168 );
 a2527a <=( (not A232)  and  A200 );
 a2528a <=( A199  and  a2527a );
 a2529a <=( a2528a  and  a2523a );
 a2532a <=( A265  and  A233 );
 a2536a <=( A269  and  A267 );
 a2537a <=( (not A266)  and  a2536a );
 a2538a <=( a2537a  and  a2532a );
 a2541a <=( A167  and  A168 );
 a2545a <=( A232  and  A200 );
 a2546a <=( A199  and  a2545a );
 a2547a <=( a2546a  and  a2541a );
 a2550a <=( A234  and  (not A233) );
 a2554a <=( A299  and  (not A298) );
 a2555a <=( A235  and  a2554a );
 a2556a <=( a2555a  and  a2550a );
 a2559a <=( A167  and  A168 );
 a2563a <=( A232  and  A200 );
 a2564a <=( A199  and  a2563a );
 a2565a <=( a2564a  and  a2559a );
 a2568a <=( A234  and  (not A233) );
 a2572a <=( A266  and  (not A265) );
 a2573a <=( A235  and  a2572a );
 a2574a <=( a2573a  and  a2568a );
 a2577a <=( A167  and  A168 );
 a2581a <=( A232  and  A200 );
 a2582a <=( A199  and  a2581a );
 a2583a <=( a2582a  and  a2577a );
 a2586a <=( A234  and  (not A233) );
 a2590a <=( A299  and  (not A298) );
 a2591a <=( A236  and  a2590a );
 a2592a <=( a2591a  and  a2586a );
 a2595a <=( A167  and  A168 );
 a2599a <=( A232  and  A200 );
 a2600a <=( A199  and  a2599a );
 a2601a <=( a2600a  and  a2595a );
 a2604a <=( A234  and  (not A233) );
 a2608a <=( A266  and  (not A265) );
 a2609a <=( A236  and  a2608a );
 a2610a <=( a2609a  and  a2604a );
 a2613a <=( A167  and  A168 );
 a2617a <=( (not A232)  and  (not A200) );
 a2618a <=( (not A199)  and  a2617a );
 a2619a <=( a2618a  and  a2613a );
 a2622a <=( A298  and  A233 );
 a2626a <=( A301  and  A300 );
 a2627a <=( (not A299)  and  a2626a );
 a2628a <=( a2627a  and  a2622a );
 a2631a <=( A167  and  A168 );
 a2635a <=( (not A232)  and  (not A200) );
 a2636a <=( (not A199)  and  a2635a );
 a2637a <=( a2636a  and  a2631a );
 a2640a <=( A298  and  A233 );
 a2644a <=( A302  and  A300 );
 a2645a <=( (not A299)  and  a2644a );
 a2646a <=( a2645a  and  a2640a );
 a2649a <=( A167  and  A168 );
 a2653a <=( (not A232)  and  (not A200) );
 a2654a <=( (not A199)  and  a2653a );
 a2655a <=( a2654a  and  a2649a );
 a2658a <=( A265  and  A233 );
 a2662a <=( A268  and  A267 );
 a2663a <=( (not A266)  and  a2662a );
 a2664a <=( a2663a  and  a2658a );
 a2667a <=( A167  and  A168 );
 a2671a <=( (not A232)  and  (not A200) );
 a2672a <=( (not A199)  and  a2671a );
 a2673a <=( a2672a  and  a2667a );
 a2676a <=( A265  and  A233 );
 a2680a <=( A269  and  A267 );
 a2681a <=( (not A266)  and  a2680a );
 a2682a <=( a2681a  and  a2676a );
 a2685a <=( A167  and  A168 );
 a2689a <=( A232  and  (not A200) );
 a2690a <=( (not A199)  and  a2689a );
 a2691a <=( a2690a  and  a2685a );
 a2694a <=( A234  and  (not A233) );
 a2698a <=( A299  and  (not A298) );
 a2699a <=( A235  and  a2698a );
 a2700a <=( a2699a  and  a2694a );
 a2703a <=( A167  and  A168 );
 a2707a <=( A232  and  (not A200) );
 a2708a <=( (not A199)  and  a2707a );
 a2709a <=( a2708a  and  a2703a );
 a2712a <=( A234  and  (not A233) );
 a2716a <=( A266  and  (not A265) );
 a2717a <=( A235  and  a2716a );
 a2718a <=( a2717a  and  a2712a );
 a2721a <=( A167  and  A168 );
 a2725a <=( A232  and  (not A200) );
 a2726a <=( (not A199)  and  a2725a );
 a2727a <=( a2726a  and  a2721a );
 a2730a <=( A234  and  (not A233) );
 a2734a <=( A299  and  (not A298) );
 a2735a <=( A236  and  a2734a );
 a2736a <=( a2735a  and  a2730a );
 a2739a <=( A167  and  A168 );
 a2743a <=( A232  and  (not A200) );
 a2744a <=( (not A199)  and  a2743a );
 a2745a <=( a2744a  and  a2739a );
 a2748a <=( A234  and  (not A233) );
 a2752a <=( A266  and  (not A265) );
 a2753a <=( A236  and  a2752a );
 a2754a <=( a2753a  and  a2748a );
 a2757a <=( A169  and  (not A170) );
 a2761a <=( A199  and  A166 );
 a2762a <=( A167  and  a2761a );
 a2763a <=( a2762a  and  a2757a );
 a2766a <=( (not A232)  and  (not A201) );
 a2770a <=( A299  and  (not A298) );
 a2771a <=( A233  and  a2770a );
 a2772a <=( a2771a  and  a2766a );
 a2775a <=( A169  and  (not A170) );
 a2779a <=( A199  and  A166 );
 a2780a <=( A167  and  a2779a );
 a2781a <=( a2780a  and  a2775a );
 a2784a <=( (not A232)  and  (not A201) );
 a2788a <=( A266  and  (not A265) );
 a2789a <=( A233  and  a2788a );
 a2790a <=( a2789a  and  a2784a );
 a2793a <=( A169  and  (not A170) );
 a2797a <=( A199  and  A166 );
 a2798a <=( A167  and  a2797a );
 a2799a <=( a2798a  and  a2793a );
 a2802a <=( (not A232)  and  A200 );
 a2806a <=( A299  and  (not A298) );
 a2807a <=( A233  and  a2806a );
 a2808a <=( a2807a  and  a2802a );
 a2811a <=( A169  and  (not A170) );
 a2815a <=( A199  and  A166 );
 a2816a <=( A167  and  a2815a );
 a2817a <=( a2816a  and  a2811a );
 a2820a <=( (not A232)  and  A200 );
 a2824a <=( A266  and  (not A265) );
 a2825a <=( A233  and  a2824a );
 a2826a <=( a2825a  and  a2820a );
 a2829a <=( A169  and  (not A170) );
 a2833a <=( (not A199)  and  A166 );
 a2834a <=( A167  and  a2833a );
 a2835a <=( a2834a  and  a2829a );
 a2838a <=( (not A232)  and  (not A200) );
 a2842a <=( A299  and  (not A298) );
 a2843a <=( A233  and  a2842a );
 a2844a <=( a2843a  and  a2838a );
 a2847a <=( A169  and  (not A170) );
 a2851a <=( (not A199)  and  A166 );
 a2852a <=( A167  and  a2851a );
 a2853a <=( a2852a  and  a2847a );
 a2856a <=( (not A232)  and  (not A200) );
 a2860a <=( A266  and  (not A265) );
 a2861a <=( A233  and  a2860a );
 a2862a <=( a2861a  and  a2856a );
 a2865a <=( A169  and  (not A170) );
 a2869a <=( A199  and  (not A166) );
 a2870a <=( (not A167)  and  a2869a );
 a2871a <=( a2870a  and  a2865a );
 a2874a <=( (not A232)  and  (not A201) );
 a2878a <=( A299  and  (not A298) );
 a2879a <=( A233  and  a2878a );
 a2880a <=( a2879a  and  a2874a );
 a2883a <=( A169  and  (not A170) );
 a2887a <=( A199  and  (not A166) );
 a2888a <=( (not A167)  and  a2887a );
 a2889a <=( a2888a  and  a2883a );
 a2892a <=( (not A232)  and  (not A201) );
 a2896a <=( A266  and  (not A265) );
 a2897a <=( A233  and  a2896a );
 a2898a <=( a2897a  and  a2892a );
 a2901a <=( A169  and  (not A170) );
 a2905a <=( A199  and  (not A166) );
 a2906a <=( (not A167)  and  a2905a );
 a2907a <=( a2906a  and  a2901a );
 a2910a <=( (not A232)  and  A200 );
 a2914a <=( A299  and  (not A298) );
 a2915a <=( A233  and  a2914a );
 a2916a <=( a2915a  and  a2910a );
 a2919a <=( A169  and  (not A170) );
 a2923a <=( A199  and  (not A166) );
 a2924a <=( (not A167)  and  a2923a );
 a2925a <=( a2924a  and  a2919a );
 a2928a <=( (not A232)  and  A200 );
 a2932a <=( A266  and  (not A265) );
 a2933a <=( A233  and  a2932a );
 a2934a <=( a2933a  and  a2928a );
 a2937a <=( A169  and  (not A170) );
 a2941a <=( (not A199)  and  (not A166) );
 a2942a <=( (not A167)  and  a2941a );
 a2943a <=( a2942a  and  a2937a );
 a2946a <=( (not A232)  and  (not A200) );
 a2950a <=( A299  and  (not A298) );
 a2951a <=( A233  and  a2950a );
 a2952a <=( a2951a  and  a2946a );
 a2955a <=( A169  and  (not A170) );
 a2959a <=( (not A199)  and  (not A166) );
 a2960a <=( (not A167)  and  a2959a );
 a2961a <=( a2960a  and  a2955a );
 a2964a <=( (not A232)  and  (not A200) );
 a2968a <=( A266  and  (not A265) );
 a2969a <=( A233  and  a2968a );
 a2970a <=( a2969a  and  a2964a );
 a2973a <=( (not A169)  and  A170 );
 a2977a <=( A199  and  (not A166) );
 a2978a <=( A167  and  a2977a );
 a2979a <=( a2978a  and  a2973a );
 a2982a <=( (not A232)  and  (not A201) );
 a2986a <=( A299  and  (not A298) );
 a2987a <=( A233  and  a2986a );
 a2988a <=( a2987a  and  a2982a );
 a2991a <=( (not A169)  and  A170 );
 a2995a <=( A199  and  (not A166) );
 a2996a <=( A167  and  a2995a );
 a2997a <=( a2996a  and  a2991a );
 a3000a <=( (not A232)  and  (not A201) );
 a3004a <=( A266  and  (not A265) );
 a3005a <=( A233  and  a3004a );
 a3006a <=( a3005a  and  a3000a );
 a3009a <=( (not A169)  and  A170 );
 a3013a <=( A199  and  (not A166) );
 a3014a <=( A167  and  a3013a );
 a3015a <=( a3014a  and  a3009a );
 a3018a <=( (not A232)  and  A200 );
 a3022a <=( A299  and  (not A298) );
 a3023a <=( A233  and  a3022a );
 a3024a <=( a3023a  and  a3018a );
 a3027a <=( (not A169)  and  A170 );
 a3031a <=( A199  and  (not A166) );
 a3032a <=( A167  and  a3031a );
 a3033a <=( a3032a  and  a3027a );
 a3036a <=( (not A232)  and  A200 );
 a3040a <=( A266  and  (not A265) );
 a3041a <=( A233  and  a3040a );
 a3042a <=( a3041a  and  a3036a );
 a3045a <=( (not A169)  and  A170 );
 a3049a <=( (not A199)  and  (not A166) );
 a3050a <=( A167  and  a3049a );
 a3051a <=( a3050a  and  a3045a );
 a3054a <=( (not A232)  and  (not A200) );
 a3058a <=( A299  and  (not A298) );
 a3059a <=( A233  and  a3058a );
 a3060a <=( a3059a  and  a3054a );
 a3063a <=( (not A169)  and  A170 );
 a3067a <=( (not A199)  and  (not A166) );
 a3068a <=( A167  and  a3067a );
 a3069a <=( a3068a  and  a3063a );
 a3072a <=( (not A232)  and  (not A200) );
 a3076a <=( A266  and  (not A265) );
 a3077a <=( A233  and  a3076a );
 a3078a <=( a3077a  and  a3072a );
 a3081a <=( (not A169)  and  A170 );
 a3085a <=( A199  and  A166 );
 a3086a <=( (not A167)  and  a3085a );
 a3087a <=( a3086a  and  a3081a );
 a3090a <=( (not A232)  and  (not A201) );
 a3094a <=( A299  and  (not A298) );
 a3095a <=( A233  and  a3094a );
 a3096a <=( a3095a  and  a3090a );
 a3099a <=( (not A169)  and  A170 );
 a3103a <=( A199  and  A166 );
 a3104a <=( (not A167)  and  a3103a );
 a3105a <=( a3104a  and  a3099a );
 a3108a <=( (not A232)  and  (not A201) );
 a3112a <=( A266  and  (not A265) );
 a3113a <=( A233  and  a3112a );
 a3114a <=( a3113a  and  a3108a );
 a3117a <=( (not A169)  and  A170 );
 a3121a <=( A199  and  A166 );
 a3122a <=( (not A167)  and  a3121a );
 a3123a <=( a3122a  and  a3117a );
 a3126a <=( (not A232)  and  A200 );
 a3130a <=( A299  and  (not A298) );
 a3131a <=( A233  and  a3130a );
 a3132a <=( a3131a  and  a3126a );
 a3135a <=( (not A169)  and  A170 );
 a3139a <=( A199  and  A166 );
 a3140a <=( (not A167)  and  a3139a );
 a3141a <=( a3140a  and  a3135a );
 a3144a <=( (not A232)  and  A200 );
 a3148a <=( A266  and  (not A265) );
 a3149a <=( A233  and  a3148a );
 a3150a <=( a3149a  and  a3144a );
 a3153a <=( (not A169)  and  A170 );
 a3157a <=( (not A199)  and  A166 );
 a3158a <=( (not A167)  and  a3157a );
 a3159a <=( a3158a  and  a3153a );
 a3162a <=( (not A232)  and  (not A200) );
 a3166a <=( A299  and  (not A298) );
 a3167a <=( A233  and  a3166a );
 a3168a <=( a3167a  and  a3162a );
 a3171a <=( (not A169)  and  A170 );
 a3175a <=( (not A199)  and  A166 );
 a3176a <=( (not A167)  and  a3175a );
 a3177a <=( a3176a  and  a3171a );
 a3180a <=( (not A232)  and  (not A200) );
 a3184a <=( A266  and  (not A265) );
 a3185a <=( A233  and  a3184a );
 a3186a <=( a3185a  and  a3180a );
 a3189a <=( A166  and  A168 );
 a3193a <=( (not A203)  and  (not A202) );
 a3194a <=( A199  and  a3193a );
 a3195a <=( a3194a  and  a3189a );
 a3199a <=( A298  and  A233 );
 a3200a <=( (not A232)  and  a3199a );
 a3204a <=( A301  and  A300 );
 a3205a <=( (not A299)  and  a3204a );
 a3206a <=( a3205a  and  a3200a );
 a3209a <=( A166  and  A168 );
 a3213a <=( (not A203)  and  (not A202) );
 a3214a <=( A199  and  a3213a );
 a3215a <=( a3214a  and  a3209a );
 a3219a <=( A298  and  A233 );
 a3220a <=( (not A232)  and  a3219a );
 a3224a <=( A302  and  A300 );
 a3225a <=( (not A299)  and  a3224a );
 a3226a <=( a3225a  and  a3220a );
 a3229a <=( A166  and  A168 );
 a3233a <=( (not A203)  and  (not A202) );
 a3234a <=( A199  and  a3233a );
 a3235a <=( a3234a  and  a3229a );
 a3239a <=( A265  and  A233 );
 a3240a <=( (not A232)  and  a3239a );
 a3244a <=( A268  and  A267 );
 a3245a <=( (not A266)  and  a3244a );
 a3246a <=( a3245a  and  a3240a );
 a3249a <=( A166  and  A168 );
 a3253a <=( (not A203)  and  (not A202) );
 a3254a <=( A199  and  a3253a );
 a3255a <=( a3254a  and  a3249a );
 a3259a <=( A265  and  A233 );
 a3260a <=( (not A232)  and  a3259a );
 a3264a <=( A269  and  A267 );
 a3265a <=( (not A266)  and  a3264a );
 a3266a <=( a3265a  and  a3260a );
 a3269a <=( A166  and  A168 );
 a3273a <=( (not A203)  and  (not A202) );
 a3274a <=( A199  and  a3273a );
 a3275a <=( a3274a  and  a3269a );
 a3279a <=( A234  and  (not A233) );
 a3280a <=( A232  and  a3279a );
 a3284a <=( A299  and  (not A298) );
 a3285a <=( A235  and  a3284a );
 a3286a <=( a3285a  and  a3280a );
 a3289a <=( A166  and  A168 );
 a3293a <=( (not A203)  and  (not A202) );
 a3294a <=( A199  and  a3293a );
 a3295a <=( a3294a  and  a3289a );
 a3299a <=( A234  and  (not A233) );
 a3300a <=( A232  and  a3299a );
 a3304a <=( A266  and  (not A265) );
 a3305a <=( A235  and  a3304a );
 a3306a <=( a3305a  and  a3300a );
 a3309a <=( A166  and  A168 );
 a3313a <=( (not A203)  and  (not A202) );
 a3314a <=( A199  and  a3313a );
 a3315a <=( a3314a  and  a3309a );
 a3319a <=( A234  and  (not A233) );
 a3320a <=( A232  and  a3319a );
 a3324a <=( A299  and  (not A298) );
 a3325a <=( A236  and  a3324a );
 a3326a <=( a3325a  and  a3320a );
 a3329a <=( A166  and  A168 );
 a3333a <=( (not A203)  and  (not A202) );
 a3334a <=( A199  and  a3333a );
 a3335a <=( a3334a  and  a3329a );
 a3339a <=( A234  and  (not A233) );
 a3340a <=( A232  and  a3339a );
 a3344a <=( A266  and  (not A265) );
 a3345a <=( A236  and  a3344a );
 a3346a <=( a3345a  and  a3340a );
 a3349a <=( A167  and  A168 );
 a3353a <=( (not A203)  and  (not A202) );
 a3354a <=( A199  and  a3353a );
 a3355a <=( a3354a  and  a3349a );
 a3359a <=( A298  and  A233 );
 a3360a <=( (not A232)  and  a3359a );
 a3364a <=( A301  and  A300 );
 a3365a <=( (not A299)  and  a3364a );
 a3366a <=( a3365a  and  a3360a );
 a3369a <=( A167  and  A168 );
 a3373a <=( (not A203)  and  (not A202) );
 a3374a <=( A199  and  a3373a );
 a3375a <=( a3374a  and  a3369a );
 a3379a <=( A298  and  A233 );
 a3380a <=( (not A232)  and  a3379a );
 a3384a <=( A302  and  A300 );
 a3385a <=( (not A299)  and  a3384a );
 a3386a <=( a3385a  and  a3380a );
 a3389a <=( A167  and  A168 );
 a3393a <=( (not A203)  and  (not A202) );
 a3394a <=( A199  and  a3393a );
 a3395a <=( a3394a  and  a3389a );
 a3399a <=( A265  and  A233 );
 a3400a <=( (not A232)  and  a3399a );
 a3404a <=( A268  and  A267 );
 a3405a <=( (not A266)  and  a3404a );
 a3406a <=( a3405a  and  a3400a );
 a3409a <=( A167  and  A168 );
 a3413a <=( (not A203)  and  (not A202) );
 a3414a <=( A199  and  a3413a );
 a3415a <=( a3414a  and  a3409a );
 a3419a <=( A265  and  A233 );
 a3420a <=( (not A232)  and  a3419a );
 a3424a <=( A269  and  A267 );
 a3425a <=( (not A266)  and  a3424a );
 a3426a <=( a3425a  and  a3420a );
 a3429a <=( A167  and  A168 );
 a3433a <=( (not A203)  and  (not A202) );
 a3434a <=( A199  and  a3433a );
 a3435a <=( a3434a  and  a3429a );
 a3439a <=( A234  and  (not A233) );
 a3440a <=( A232  and  a3439a );
 a3444a <=( A299  and  (not A298) );
 a3445a <=( A235  and  a3444a );
 a3446a <=( a3445a  and  a3440a );
 a3449a <=( A167  and  A168 );
 a3453a <=( (not A203)  and  (not A202) );
 a3454a <=( A199  and  a3453a );
 a3455a <=( a3454a  and  a3449a );
 a3459a <=( A234  and  (not A233) );
 a3460a <=( A232  and  a3459a );
 a3464a <=( A266  and  (not A265) );
 a3465a <=( A235  and  a3464a );
 a3466a <=( a3465a  and  a3460a );
 a3469a <=( A167  and  A168 );
 a3473a <=( (not A203)  and  (not A202) );
 a3474a <=( A199  and  a3473a );
 a3475a <=( a3474a  and  a3469a );
 a3479a <=( A234  and  (not A233) );
 a3480a <=( A232  and  a3479a );
 a3484a <=( A299  and  (not A298) );
 a3485a <=( A236  and  a3484a );
 a3486a <=( a3485a  and  a3480a );
 a3489a <=( A167  and  A168 );
 a3493a <=( (not A203)  and  (not A202) );
 a3494a <=( A199  and  a3493a );
 a3495a <=( a3494a  and  a3489a );
 a3499a <=( A234  and  (not A233) );
 a3500a <=( A232  and  a3499a );
 a3504a <=( A266  and  (not A265) );
 a3505a <=( A236  and  a3504a );
 a3506a <=( a3505a  and  a3500a );
 a3509a <=( A169  and  (not A170) );
 a3513a <=( A199  and  A166 );
 a3514a <=( A167  and  a3513a );
 a3515a <=( a3514a  and  a3509a );
 a3519a <=( (not A232)  and  (not A203) );
 a3520a <=( (not A202)  and  a3519a );
 a3524a <=( A299  and  (not A298) );
 a3525a <=( A233  and  a3524a );
 a3526a <=( a3525a  and  a3520a );
 a3529a <=( A169  and  (not A170) );
 a3533a <=( A199  and  A166 );
 a3534a <=( A167  and  a3533a );
 a3535a <=( a3534a  and  a3529a );
 a3539a <=( (not A232)  and  (not A203) );
 a3540a <=( (not A202)  and  a3539a );
 a3544a <=( A266  and  (not A265) );
 a3545a <=( A233  and  a3544a );
 a3546a <=( a3545a  and  a3540a );
 a3549a <=( A169  and  (not A170) );
 a3553a <=( A199  and  (not A166) );
 a3554a <=( (not A167)  and  a3553a );
 a3555a <=( a3554a  and  a3549a );
 a3559a <=( (not A232)  and  (not A203) );
 a3560a <=( (not A202)  and  a3559a );
 a3564a <=( A299  and  (not A298) );
 a3565a <=( A233  and  a3564a );
 a3566a <=( a3565a  and  a3560a );
 a3569a <=( A169  and  (not A170) );
 a3573a <=( A199  and  (not A166) );
 a3574a <=( (not A167)  and  a3573a );
 a3575a <=( a3574a  and  a3569a );
 a3579a <=( (not A232)  and  (not A203) );
 a3580a <=( (not A202)  and  a3579a );
 a3584a <=( A266  and  (not A265) );
 a3585a <=( A233  and  a3584a );
 a3586a <=( a3585a  and  a3580a );
 a3589a <=( (not A169)  and  A170 );
 a3593a <=( A199  and  (not A166) );
 a3594a <=( A167  and  a3593a );
 a3595a <=( a3594a  and  a3589a );
 a3599a <=( (not A232)  and  (not A203) );
 a3600a <=( (not A202)  and  a3599a );
 a3604a <=( A299  and  (not A298) );
 a3605a <=( A233  and  a3604a );
 a3606a <=( a3605a  and  a3600a );
 a3609a <=( (not A169)  and  A170 );
 a3613a <=( A199  and  (not A166) );
 a3614a <=( A167  and  a3613a );
 a3615a <=( a3614a  and  a3609a );
 a3619a <=( (not A232)  and  (not A203) );
 a3620a <=( (not A202)  and  a3619a );
 a3624a <=( A266  and  (not A265) );
 a3625a <=( A233  and  a3624a );
 a3626a <=( a3625a  and  a3620a );
 a3629a <=( (not A169)  and  A170 );
 a3633a <=( A199  and  A166 );
 a3634a <=( (not A167)  and  a3633a );
 a3635a <=( a3634a  and  a3629a );
 a3639a <=( (not A232)  and  (not A203) );
 a3640a <=( (not A202)  and  a3639a );
 a3644a <=( A299  and  (not A298) );
 a3645a <=( A233  and  a3644a );
 a3646a <=( a3645a  and  a3640a );
 a3649a <=( (not A169)  and  A170 );
 a3653a <=( A199  and  A166 );
 a3654a <=( (not A167)  and  a3653a );
 a3655a <=( a3654a  and  a3649a );
 a3659a <=( (not A232)  and  (not A203) );
 a3660a <=( (not A202)  and  a3659a );
 a3664a <=( A266  and  (not A265) );
 a3665a <=( A233  and  a3664a );
 a3666a <=( a3665a  and  a3660a );
 a3670a <=( A199  and  A166 );
 a3671a <=( A168  and  a3670a );
 a3675a <=( (not A233)  and  A232 );
 a3676a <=( (not A201)  and  a3675a );
 a3677a <=( a3676a  and  a3671a );
 a3681a <=( A298  and  A235 );
 a3682a <=( A234  and  a3681a );
 a3686a <=( A301  and  A300 );
 a3687a <=( (not A299)  and  a3686a );
 a3688a <=( a3687a  and  a3682a );
 a3692a <=( A199  and  A166 );
 a3693a <=( A168  and  a3692a );
 a3697a <=( (not A233)  and  A232 );
 a3698a <=( (not A201)  and  a3697a );
 a3699a <=( a3698a  and  a3693a );
 a3703a <=( A298  and  A235 );
 a3704a <=( A234  and  a3703a );
 a3708a <=( A302  and  A300 );
 a3709a <=( (not A299)  and  a3708a );
 a3710a <=( a3709a  and  a3704a );
 a3714a <=( A199  and  A166 );
 a3715a <=( A168  and  a3714a );
 a3719a <=( (not A233)  and  A232 );
 a3720a <=( (not A201)  and  a3719a );
 a3721a <=( a3720a  and  a3715a );
 a3725a <=( A265  and  A235 );
 a3726a <=( A234  and  a3725a );
 a3730a <=( A268  and  A267 );
 a3731a <=( (not A266)  and  a3730a );
 a3732a <=( a3731a  and  a3726a );
 a3736a <=( A199  and  A166 );
 a3737a <=( A168  and  a3736a );
 a3741a <=( (not A233)  and  A232 );
 a3742a <=( (not A201)  and  a3741a );
 a3743a <=( a3742a  and  a3737a );
 a3747a <=( A265  and  A235 );
 a3748a <=( A234  and  a3747a );
 a3752a <=( A269  and  A267 );
 a3753a <=( (not A266)  and  a3752a );
 a3754a <=( a3753a  and  a3748a );
 a3758a <=( A199  and  A166 );
 a3759a <=( A168  and  a3758a );
 a3763a <=( (not A233)  and  A232 );
 a3764a <=( (not A201)  and  a3763a );
 a3765a <=( a3764a  and  a3759a );
 a3769a <=( A298  and  A236 );
 a3770a <=( A234  and  a3769a );
 a3774a <=( A301  and  A300 );
 a3775a <=( (not A299)  and  a3774a );
 a3776a <=( a3775a  and  a3770a );
 a3780a <=( A199  and  A166 );
 a3781a <=( A168  and  a3780a );
 a3785a <=( (not A233)  and  A232 );
 a3786a <=( (not A201)  and  a3785a );
 a3787a <=( a3786a  and  a3781a );
 a3791a <=( A298  and  A236 );
 a3792a <=( A234  and  a3791a );
 a3796a <=( A302  and  A300 );
 a3797a <=( (not A299)  and  a3796a );
 a3798a <=( a3797a  and  a3792a );
 a3802a <=( A199  and  A166 );
 a3803a <=( A168  and  a3802a );
 a3807a <=( (not A233)  and  A232 );
 a3808a <=( (not A201)  and  a3807a );
 a3809a <=( a3808a  and  a3803a );
 a3813a <=( A265  and  A236 );
 a3814a <=( A234  and  a3813a );
 a3818a <=( A268  and  A267 );
 a3819a <=( (not A266)  and  a3818a );
 a3820a <=( a3819a  and  a3814a );
 a3824a <=( A199  and  A166 );
 a3825a <=( A168  and  a3824a );
 a3829a <=( (not A233)  and  A232 );
 a3830a <=( (not A201)  and  a3829a );
 a3831a <=( a3830a  and  a3825a );
 a3835a <=( A265  and  A236 );
 a3836a <=( A234  and  a3835a );
 a3840a <=( A269  and  A267 );
 a3841a <=( (not A266)  and  a3840a );
 a3842a <=( a3841a  and  a3836a );
 a3846a <=( A199  and  A166 );
 a3847a <=( A168  and  a3846a );
 a3851a <=( (not A233)  and  A232 );
 a3852a <=( A200  and  a3851a );
 a3853a <=( a3852a  and  a3847a );
 a3857a <=( A298  and  A235 );
 a3858a <=( A234  and  a3857a );
 a3862a <=( A301  and  A300 );
 a3863a <=( (not A299)  and  a3862a );
 a3864a <=( a3863a  and  a3858a );
 a3868a <=( A199  and  A166 );
 a3869a <=( A168  and  a3868a );
 a3873a <=( (not A233)  and  A232 );
 a3874a <=( A200  and  a3873a );
 a3875a <=( a3874a  and  a3869a );
 a3879a <=( A298  and  A235 );
 a3880a <=( A234  and  a3879a );
 a3884a <=( A302  and  A300 );
 a3885a <=( (not A299)  and  a3884a );
 a3886a <=( a3885a  and  a3880a );
 a3890a <=( A199  and  A166 );
 a3891a <=( A168  and  a3890a );
 a3895a <=( (not A233)  and  A232 );
 a3896a <=( A200  and  a3895a );
 a3897a <=( a3896a  and  a3891a );
 a3901a <=( A265  and  A235 );
 a3902a <=( A234  and  a3901a );
 a3906a <=( A268  and  A267 );
 a3907a <=( (not A266)  and  a3906a );
 a3908a <=( a3907a  and  a3902a );
 a3912a <=( A199  and  A166 );
 a3913a <=( A168  and  a3912a );
 a3917a <=( (not A233)  and  A232 );
 a3918a <=( A200  and  a3917a );
 a3919a <=( a3918a  and  a3913a );
 a3923a <=( A265  and  A235 );
 a3924a <=( A234  and  a3923a );
 a3928a <=( A269  and  A267 );
 a3929a <=( (not A266)  and  a3928a );
 a3930a <=( a3929a  and  a3924a );
 a3934a <=( A199  and  A166 );
 a3935a <=( A168  and  a3934a );
 a3939a <=( (not A233)  and  A232 );
 a3940a <=( A200  and  a3939a );
 a3941a <=( a3940a  and  a3935a );
 a3945a <=( A298  and  A236 );
 a3946a <=( A234  and  a3945a );
 a3950a <=( A301  and  A300 );
 a3951a <=( (not A299)  and  a3950a );
 a3952a <=( a3951a  and  a3946a );
 a3956a <=( A199  and  A166 );
 a3957a <=( A168  and  a3956a );
 a3961a <=( (not A233)  and  A232 );
 a3962a <=( A200  and  a3961a );
 a3963a <=( a3962a  and  a3957a );
 a3967a <=( A298  and  A236 );
 a3968a <=( A234  and  a3967a );
 a3972a <=( A302  and  A300 );
 a3973a <=( (not A299)  and  a3972a );
 a3974a <=( a3973a  and  a3968a );
 a3978a <=( A199  and  A166 );
 a3979a <=( A168  and  a3978a );
 a3983a <=( (not A233)  and  A232 );
 a3984a <=( A200  and  a3983a );
 a3985a <=( a3984a  and  a3979a );
 a3989a <=( A265  and  A236 );
 a3990a <=( A234  and  a3989a );
 a3994a <=( A268  and  A267 );
 a3995a <=( (not A266)  and  a3994a );
 a3996a <=( a3995a  and  a3990a );
 a4000a <=( A199  and  A166 );
 a4001a <=( A168  and  a4000a );
 a4005a <=( (not A233)  and  A232 );
 a4006a <=( A200  and  a4005a );
 a4007a <=( a4006a  and  a4001a );
 a4011a <=( A265  and  A236 );
 a4012a <=( A234  and  a4011a );
 a4016a <=( A269  and  A267 );
 a4017a <=( (not A266)  and  a4016a );
 a4018a <=( a4017a  and  a4012a );
 a4022a <=( (not A199)  and  A166 );
 a4023a <=( A168  and  a4022a );
 a4027a <=( (not A233)  and  A232 );
 a4028a <=( (not A200)  and  a4027a );
 a4029a <=( a4028a  and  a4023a );
 a4033a <=( A298  and  A235 );
 a4034a <=( A234  and  a4033a );
 a4038a <=( A301  and  A300 );
 a4039a <=( (not A299)  and  a4038a );
 a4040a <=( a4039a  and  a4034a );
 a4044a <=( (not A199)  and  A166 );
 a4045a <=( A168  and  a4044a );
 a4049a <=( (not A233)  and  A232 );
 a4050a <=( (not A200)  and  a4049a );
 a4051a <=( a4050a  and  a4045a );
 a4055a <=( A298  and  A235 );
 a4056a <=( A234  and  a4055a );
 a4060a <=( A302  and  A300 );
 a4061a <=( (not A299)  and  a4060a );
 a4062a <=( a4061a  and  a4056a );
 a4066a <=( (not A199)  and  A166 );
 a4067a <=( A168  and  a4066a );
 a4071a <=( (not A233)  and  A232 );
 a4072a <=( (not A200)  and  a4071a );
 a4073a <=( a4072a  and  a4067a );
 a4077a <=( A265  and  A235 );
 a4078a <=( A234  and  a4077a );
 a4082a <=( A268  and  A267 );
 a4083a <=( (not A266)  and  a4082a );
 a4084a <=( a4083a  and  a4078a );
 a4088a <=( (not A199)  and  A166 );
 a4089a <=( A168  and  a4088a );
 a4093a <=( (not A233)  and  A232 );
 a4094a <=( (not A200)  and  a4093a );
 a4095a <=( a4094a  and  a4089a );
 a4099a <=( A265  and  A235 );
 a4100a <=( A234  and  a4099a );
 a4104a <=( A269  and  A267 );
 a4105a <=( (not A266)  and  a4104a );
 a4106a <=( a4105a  and  a4100a );
 a4110a <=( (not A199)  and  A166 );
 a4111a <=( A168  and  a4110a );
 a4115a <=( (not A233)  and  A232 );
 a4116a <=( (not A200)  and  a4115a );
 a4117a <=( a4116a  and  a4111a );
 a4121a <=( A298  and  A236 );
 a4122a <=( A234  and  a4121a );
 a4126a <=( A301  and  A300 );
 a4127a <=( (not A299)  and  a4126a );
 a4128a <=( a4127a  and  a4122a );
 a4132a <=( (not A199)  and  A166 );
 a4133a <=( A168  and  a4132a );
 a4137a <=( (not A233)  and  A232 );
 a4138a <=( (not A200)  and  a4137a );
 a4139a <=( a4138a  and  a4133a );
 a4143a <=( A298  and  A236 );
 a4144a <=( A234  and  a4143a );
 a4148a <=( A302  and  A300 );
 a4149a <=( (not A299)  and  a4148a );
 a4150a <=( a4149a  and  a4144a );
 a4154a <=( (not A199)  and  A166 );
 a4155a <=( A168  and  a4154a );
 a4159a <=( (not A233)  and  A232 );
 a4160a <=( (not A200)  and  a4159a );
 a4161a <=( a4160a  and  a4155a );
 a4165a <=( A265  and  A236 );
 a4166a <=( A234  and  a4165a );
 a4170a <=( A268  and  A267 );
 a4171a <=( (not A266)  and  a4170a );
 a4172a <=( a4171a  and  a4166a );
 a4176a <=( (not A199)  and  A166 );
 a4177a <=( A168  and  a4176a );
 a4181a <=( (not A233)  and  A232 );
 a4182a <=( (not A200)  and  a4181a );
 a4183a <=( a4182a  and  a4177a );
 a4187a <=( A265  and  A236 );
 a4188a <=( A234  and  a4187a );
 a4192a <=( A269  and  A267 );
 a4193a <=( (not A266)  and  a4192a );
 a4194a <=( a4193a  and  a4188a );
 a4198a <=( A199  and  A167 );
 a4199a <=( A168  and  a4198a );
 a4203a <=( (not A233)  and  A232 );
 a4204a <=( (not A201)  and  a4203a );
 a4205a <=( a4204a  and  a4199a );
 a4209a <=( A298  and  A235 );
 a4210a <=( A234  and  a4209a );
 a4214a <=( A301  and  A300 );
 a4215a <=( (not A299)  and  a4214a );
 a4216a <=( a4215a  and  a4210a );
 a4220a <=( A199  and  A167 );
 a4221a <=( A168  and  a4220a );
 a4225a <=( (not A233)  and  A232 );
 a4226a <=( (not A201)  and  a4225a );
 a4227a <=( a4226a  and  a4221a );
 a4231a <=( A298  and  A235 );
 a4232a <=( A234  and  a4231a );
 a4236a <=( A302  and  A300 );
 a4237a <=( (not A299)  and  a4236a );
 a4238a <=( a4237a  and  a4232a );
 a4242a <=( A199  and  A167 );
 a4243a <=( A168  and  a4242a );
 a4247a <=( (not A233)  and  A232 );
 a4248a <=( (not A201)  and  a4247a );
 a4249a <=( a4248a  and  a4243a );
 a4253a <=( A265  and  A235 );
 a4254a <=( A234  and  a4253a );
 a4258a <=( A268  and  A267 );
 a4259a <=( (not A266)  and  a4258a );
 a4260a <=( a4259a  and  a4254a );
 a4264a <=( A199  and  A167 );
 a4265a <=( A168  and  a4264a );
 a4269a <=( (not A233)  and  A232 );
 a4270a <=( (not A201)  and  a4269a );
 a4271a <=( a4270a  and  a4265a );
 a4275a <=( A265  and  A235 );
 a4276a <=( A234  and  a4275a );
 a4280a <=( A269  and  A267 );
 a4281a <=( (not A266)  and  a4280a );
 a4282a <=( a4281a  and  a4276a );
 a4286a <=( A199  and  A167 );
 a4287a <=( A168  and  a4286a );
 a4291a <=( (not A233)  and  A232 );
 a4292a <=( (not A201)  and  a4291a );
 a4293a <=( a4292a  and  a4287a );
 a4297a <=( A298  and  A236 );
 a4298a <=( A234  and  a4297a );
 a4302a <=( A301  and  A300 );
 a4303a <=( (not A299)  and  a4302a );
 a4304a <=( a4303a  and  a4298a );
 a4308a <=( A199  and  A167 );
 a4309a <=( A168  and  a4308a );
 a4313a <=( (not A233)  and  A232 );
 a4314a <=( (not A201)  and  a4313a );
 a4315a <=( a4314a  and  a4309a );
 a4319a <=( A298  and  A236 );
 a4320a <=( A234  and  a4319a );
 a4324a <=( A302  and  A300 );
 a4325a <=( (not A299)  and  a4324a );
 a4326a <=( a4325a  and  a4320a );
 a4330a <=( A199  and  A167 );
 a4331a <=( A168  and  a4330a );
 a4335a <=( (not A233)  and  A232 );
 a4336a <=( (not A201)  and  a4335a );
 a4337a <=( a4336a  and  a4331a );
 a4341a <=( A265  and  A236 );
 a4342a <=( A234  and  a4341a );
 a4346a <=( A268  and  A267 );
 a4347a <=( (not A266)  and  a4346a );
 a4348a <=( a4347a  and  a4342a );
 a4352a <=( A199  and  A167 );
 a4353a <=( A168  and  a4352a );
 a4357a <=( (not A233)  and  A232 );
 a4358a <=( (not A201)  and  a4357a );
 a4359a <=( a4358a  and  a4353a );
 a4363a <=( A265  and  A236 );
 a4364a <=( A234  and  a4363a );
 a4368a <=( A269  and  A267 );
 a4369a <=( (not A266)  and  a4368a );
 a4370a <=( a4369a  and  a4364a );
 a4374a <=( A199  and  A167 );
 a4375a <=( A168  and  a4374a );
 a4379a <=( (not A233)  and  A232 );
 a4380a <=( A200  and  a4379a );
 a4381a <=( a4380a  and  a4375a );
 a4385a <=( A298  and  A235 );
 a4386a <=( A234  and  a4385a );
 a4390a <=( A301  and  A300 );
 a4391a <=( (not A299)  and  a4390a );
 a4392a <=( a4391a  and  a4386a );
 a4396a <=( A199  and  A167 );
 a4397a <=( A168  and  a4396a );
 a4401a <=( (not A233)  and  A232 );
 a4402a <=( A200  and  a4401a );
 a4403a <=( a4402a  and  a4397a );
 a4407a <=( A298  and  A235 );
 a4408a <=( A234  and  a4407a );
 a4412a <=( A302  and  A300 );
 a4413a <=( (not A299)  and  a4412a );
 a4414a <=( a4413a  and  a4408a );
 a4418a <=( A199  and  A167 );
 a4419a <=( A168  and  a4418a );
 a4423a <=( (not A233)  and  A232 );
 a4424a <=( A200  and  a4423a );
 a4425a <=( a4424a  and  a4419a );
 a4429a <=( A265  and  A235 );
 a4430a <=( A234  and  a4429a );
 a4434a <=( A268  and  A267 );
 a4435a <=( (not A266)  and  a4434a );
 a4436a <=( a4435a  and  a4430a );
 a4440a <=( A199  and  A167 );
 a4441a <=( A168  and  a4440a );
 a4445a <=( (not A233)  and  A232 );
 a4446a <=( A200  and  a4445a );
 a4447a <=( a4446a  and  a4441a );
 a4451a <=( A265  and  A235 );
 a4452a <=( A234  and  a4451a );
 a4456a <=( A269  and  A267 );
 a4457a <=( (not A266)  and  a4456a );
 a4458a <=( a4457a  and  a4452a );
 a4462a <=( A199  and  A167 );
 a4463a <=( A168  and  a4462a );
 a4467a <=( (not A233)  and  A232 );
 a4468a <=( A200  and  a4467a );
 a4469a <=( a4468a  and  a4463a );
 a4473a <=( A298  and  A236 );
 a4474a <=( A234  and  a4473a );
 a4478a <=( A301  and  A300 );
 a4479a <=( (not A299)  and  a4478a );
 a4480a <=( a4479a  and  a4474a );
 a4484a <=( A199  and  A167 );
 a4485a <=( A168  and  a4484a );
 a4489a <=( (not A233)  and  A232 );
 a4490a <=( A200  and  a4489a );
 a4491a <=( a4490a  and  a4485a );
 a4495a <=( A298  and  A236 );
 a4496a <=( A234  and  a4495a );
 a4500a <=( A302  and  A300 );
 a4501a <=( (not A299)  and  a4500a );
 a4502a <=( a4501a  and  a4496a );
 a4506a <=( A199  and  A167 );
 a4507a <=( A168  and  a4506a );
 a4511a <=( (not A233)  and  A232 );
 a4512a <=( A200  and  a4511a );
 a4513a <=( a4512a  and  a4507a );
 a4517a <=( A265  and  A236 );
 a4518a <=( A234  and  a4517a );
 a4522a <=( A268  and  A267 );
 a4523a <=( (not A266)  and  a4522a );
 a4524a <=( a4523a  and  a4518a );
 a4528a <=( A199  and  A167 );
 a4529a <=( A168  and  a4528a );
 a4533a <=( (not A233)  and  A232 );
 a4534a <=( A200  and  a4533a );
 a4535a <=( a4534a  and  a4529a );
 a4539a <=( A265  and  A236 );
 a4540a <=( A234  and  a4539a );
 a4544a <=( A269  and  A267 );
 a4545a <=( (not A266)  and  a4544a );
 a4546a <=( a4545a  and  a4540a );
 a4550a <=( (not A199)  and  A167 );
 a4551a <=( A168  and  a4550a );
 a4555a <=( (not A233)  and  A232 );
 a4556a <=( (not A200)  and  a4555a );
 a4557a <=( a4556a  and  a4551a );
 a4561a <=( A298  and  A235 );
 a4562a <=( A234  and  a4561a );
 a4566a <=( A301  and  A300 );
 a4567a <=( (not A299)  and  a4566a );
 a4568a <=( a4567a  and  a4562a );
 a4572a <=( (not A199)  and  A167 );
 a4573a <=( A168  and  a4572a );
 a4577a <=( (not A233)  and  A232 );
 a4578a <=( (not A200)  and  a4577a );
 a4579a <=( a4578a  and  a4573a );
 a4583a <=( A298  and  A235 );
 a4584a <=( A234  and  a4583a );
 a4588a <=( A302  and  A300 );
 a4589a <=( (not A299)  and  a4588a );
 a4590a <=( a4589a  and  a4584a );
 a4594a <=( (not A199)  and  A167 );
 a4595a <=( A168  and  a4594a );
 a4599a <=( (not A233)  and  A232 );
 a4600a <=( (not A200)  and  a4599a );
 a4601a <=( a4600a  and  a4595a );
 a4605a <=( A265  and  A235 );
 a4606a <=( A234  and  a4605a );
 a4610a <=( A268  and  A267 );
 a4611a <=( (not A266)  and  a4610a );
 a4612a <=( a4611a  and  a4606a );
 a4616a <=( (not A199)  and  A167 );
 a4617a <=( A168  and  a4616a );
 a4621a <=( (not A233)  and  A232 );
 a4622a <=( (not A200)  and  a4621a );
 a4623a <=( a4622a  and  a4617a );
 a4627a <=( A265  and  A235 );
 a4628a <=( A234  and  a4627a );
 a4632a <=( A269  and  A267 );
 a4633a <=( (not A266)  and  a4632a );
 a4634a <=( a4633a  and  a4628a );
 a4638a <=( (not A199)  and  A167 );
 a4639a <=( A168  and  a4638a );
 a4643a <=( (not A233)  and  A232 );
 a4644a <=( (not A200)  and  a4643a );
 a4645a <=( a4644a  and  a4639a );
 a4649a <=( A298  and  A236 );
 a4650a <=( A234  and  a4649a );
 a4654a <=( A301  and  A300 );
 a4655a <=( (not A299)  and  a4654a );
 a4656a <=( a4655a  and  a4650a );
 a4660a <=( (not A199)  and  A167 );
 a4661a <=( A168  and  a4660a );
 a4665a <=( (not A233)  and  A232 );
 a4666a <=( (not A200)  and  a4665a );
 a4667a <=( a4666a  and  a4661a );
 a4671a <=( A298  and  A236 );
 a4672a <=( A234  and  a4671a );
 a4676a <=( A302  and  A300 );
 a4677a <=( (not A299)  and  a4676a );
 a4678a <=( a4677a  and  a4672a );
 a4682a <=( (not A199)  and  A167 );
 a4683a <=( A168  and  a4682a );
 a4687a <=( (not A233)  and  A232 );
 a4688a <=( (not A200)  and  a4687a );
 a4689a <=( a4688a  and  a4683a );
 a4693a <=( A265  and  A236 );
 a4694a <=( A234  and  a4693a );
 a4698a <=( A268  and  A267 );
 a4699a <=( (not A266)  and  a4698a );
 a4700a <=( a4699a  and  a4694a );
 a4704a <=( (not A199)  and  A167 );
 a4705a <=( A168  and  a4704a );
 a4709a <=( (not A233)  and  A232 );
 a4710a <=( (not A200)  and  a4709a );
 a4711a <=( a4710a  and  a4705a );
 a4715a <=( A265  and  A236 );
 a4716a <=( A234  and  a4715a );
 a4720a <=( A269  and  A267 );
 a4721a <=( (not A266)  and  a4720a );
 a4722a <=( a4721a  and  a4716a );
 a4726a <=( A167  and  A169 );
 a4727a <=( (not A170)  and  a4726a );
 a4731a <=( (not A201)  and  A199 );
 a4732a <=( A166  and  a4731a );
 a4733a <=( a4732a  and  a4727a );
 a4737a <=( A298  and  A233 );
 a4738a <=( (not A232)  and  a4737a );
 a4742a <=( A301  and  A300 );
 a4743a <=( (not A299)  and  a4742a );
 a4744a <=( a4743a  and  a4738a );
 a4748a <=( A167  and  A169 );
 a4749a <=( (not A170)  and  a4748a );
 a4753a <=( (not A201)  and  A199 );
 a4754a <=( A166  and  a4753a );
 a4755a <=( a4754a  and  a4749a );
 a4759a <=( A298  and  A233 );
 a4760a <=( (not A232)  and  a4759a );
 a4764a <=( A302  and  A300 );
 a4765a <=( (not A299)  and  a4764a );
 a4766a <=( a4765a  and  a4760a );
 a4770a <=( A167  and  A169 );
 a4771a <=( (not A170)  and  a4770a );
 a4775a <=( (not A201)  and  A199 );
 a4776a <=( A166  and  a4775a );
 a4777a <=( a4776a  and  a4771a );
 a4781a <=( A265  and  A233 );
 a4782a <=( (not A232)  and  a4781a );
 a4786a <=( A268  and  A267 );
 a4787a <=( (not A266)  and  a4786a );
 a4788a <=( a4787a  and  a4782a );
 a4792a <=( A167  and  A169 );
 a4793a <=( (not A170)  and  a4792a );
 a4797a <=( (not A201)  and  A199 );
 a4798a <=( A166  and  a4797a );
 a4799a <=( a4798a  and  a4793a );
 a4803a <=( A265  and  A233 );
 a4804a <=( (not A232)  and  a4803a );
 a4808a <=( A269  and  A267 );
 a4809a <=( (not A266)  and  a4808a );
 a4810a <=( a4809a  and  a4804a );
 a4814a <=( A167  and  A169 );
 a4815a <=( (not A170)  and  a4814a );
 a4819a <=( (not A201)  and  A199 );
 a4820a <=( A166  and  a4819a );
 a4821a <=( a4820a  and  a4815a );
 a4825a <=( A234  and  (not A233) );
 a4826a <=( A232  and  a4825a );
 a4830a <=( A299  and  (not A298) );
 a4831a <=( A235  and  a4830a );
 a4832a <=( a4831a  and  a4826a );
 a4836a <=( A167  and  A169 );
 a4837a <=( (not A170)  and  a4836a );
 a4841a <=( (not A201)  and  A199 );
 a4842a <=( A166  and  a4841a );
 a4843a <=( a4842a  and  a4837a );
 a4847a <=( A234  and  (not A233) );
 a4848a <=( A232  and  a4847a );
 a4852a <=( A266  and  (not A265) );
 a4853a <=( A235  and  a4852a );
 a4854a <=( a4853a  and  a4848a );
 a4858a <=( A167  and  A169 );
 a4859a <=( (not A170)  and  a4858a );
 a4863a <=( (not A201)  and  A199 );
 a4864a <=( A166  and  a4863a );
 a4865a <=( a4864a  and  a4859a );
 a4869a <=( A234  and  (not A233) );
 a4870a <=( A232  and  a4869a );
 a4874a <=( A299  and  (not A298) );
 a4875a <=( A236  and  a4874a );
 a4876a <=( a4875a  and  a4870a );
 a4880a <=( A167  and  A169 );
 a4881a <=( (not A170)  and  a4880a );
 a4885a <=( (not A201)  and  A199 );
 a4886a <=( A166  and  a4885a );
 a4887a <=( a4886a  and  a4881a );
 a4891a <=( A234  and  (not A233) );
 a4892a <=( A232  and  a4891a );
 a4896a <=( A266  and  (not A265) );
 a4897a <=( A236  and  a4896a );
 a4898a <=( a4897a  and  a4892a );
 a4902a <=( A167  and  A169 );
 a4903a <=( (not A170)  and  a4902a );
 a4907a <=( A200  and  A199 );
 a4908a <=( A166  and  a4907a );
 a4909a <=( a4908a  and  a4903a );
 a4913a <=( A298  and  A233 );
 a4914a <=( (not A232)  and  a4913a );
 a4918a <=( A301  and  A300 );
 a4919a <=( (not A299)  and  a4918a );
 a4920a <=( a4919a  and  a4914a );
 a4924a <=( A167  and  A169 );
 a4925a <=( (not A170)  and  a4924a );
 a4929a <=( A200  and  A199 );
 a4930a <=( A166  and  a4929a );
 a4931a <=( a4930a  and  a4925a );
 a4935a <=( A298  and  A233 );
 a4936a <=( (not A232)  and  a4935a );
 a4940a <=( A302  and  A300 );
 a4941a <=( (not A299)  and  a4940a );
 a4942a <=( a4941a  and  a4936a );
 a4946a <=( A167  and  A169 );
 a4947a <=( (not A170)  and  a4946a );
 a4951a <=( A200  and  A199 );
 a4952a <=( A166  and  a4951a );
 a4953a <=( a4952a  and  a4947a );
 a4957a <=( A265  and  A233 );
 a4958a <=( (not A232)  and  a4957a );
 a4962a <=( A268  and  A267 );
 a4963a <=( (not A266)  and  a4962a );
 a4964a <=( a4963a  and  a4958a );
 a4968a <=( A167  and  A169 );
 a4969a <=( (not A170)  and  a4968a );
 a4973a <=( A200  and  A199 );
 a4974a <=( A166  and  a4973a );
 a4975a <=( a4974a  and  a4969a );
 a4979a <=( A265  and  A233 );
 a4980a <=( (not A232)  and  a4979a );
 a4984a <=( A269  and  A267 );
 a4985a <=( (not A266)  and  a4984a );
 a4986a <=( a4985a  and  a4980a );
 a4990a <=( A167  and  A169 );
 a4991a <=( (not A170)  and  a4990a );
 a4995a <=( A200  and  A199 );
 a4996a <=( A166  and  a4995a );
 a4997a <=( a4996a  and  a4991a );
 a5001a <=( A234  and  (not A233) );
 a5002a <=( A232  and  a5001a );
 a5006a <=( A299  and  (not A298) );
 a5007a <=( A235  and  a5006a );
 a5008a <=( a5007a  and  a5002a );
 a5012a <=( A167  and  A169 );
 a5013a <=( (not A170)  and  a5012a );
 a5017a <=( A200  and  A199 );
 a5018a <=( A166  and  a5017a );
 a5019a <=( a5018a  and  a5013a );
 a5023a <=( A234  and  (not A233) );
 a5024a <=( A232  and  a5023a );
 a5028a <=( A266  and  (not A265) );
 a5029a <=( A235  and  a5028a );
 a5030a <=( a5029a  and  a5024a );
 a5034a <=( A167  and  A169 );
 a5035a <=( (not A170)  and  a5034a );
 a5039a <=( A200  and  A199 );
 a5040a <=( A166  and  a5039a );
 a5041a <=( a5040a  and  a5035a );
 a5045a <=( A234  and  (not A233) );
 a5046a <=( A232  and  a5045a );
 a5050a <=( A299  and  (not A298) );
 a5051a <=( A236  and  a5050a );
 a5052a <=( a5051a  and  a5046a );
 a5056a <=( A167  and  A169 );
 a5057a <=( (not A170)  and  a5056a );
 a5061a <=( A200  and  A199 );
 a5062a <=( A166  and  a5061a );
 a5063a <=( a5062a  and  a5057a );
 a5067a <=( A234  and  (not A233) );
 a5068a <=( A232  and  a5067a );
 a5072a <=( A266  and  (not A265) );
 a5073a <=( A236  and  a5072a );
 a5074a <=( a5073a  and  a5068a );
 a5078a <=( A167  and  A169 );
 a5079a <=( (not A170)  and  a5078a );
 a5083a <=( (not A200)  and  (not A199) );
 a5084a <=( A166  and  a5083a );
 a5085a <=( a5084a  and  a5079a );
 a5089a <=( A298  and  A233 );
 a5090a <=( (not A232)  and  a5089a );
 a5094a <=( A301  and  A300 );
 a5095a <=( (not A299)  and  a5094a );
 a5096a <=( a5095a  and  a5090a );
 a5100a <=( A167  and  A169 );
 a5101a <=( (not A170)  and  a5100a );
 a5105a <=( (not A200)  and  (not A199) );
 a5106a <=( A166  and  a5105a );
 a5107a <=( a5106a  and  a5101a );
 a5111a <=( A298  and  A233 );
 a5112a <=( (not A232)  and  a5111a );
 a5116a <=( A302  and  A300 );
 a5117a <=( (not A299)  and  a5116a );
 a5118a <=( a5117a  and  a5112a );
 a5122a <=( A167  and  A169 );
 a5123a <=( (not A170)  and  a5122a );
 a5127a <=( (not A200)  and  (not A199) );
 a5128a <=( A166  and  a5127a );
 a5129a <=( a5128a  and  a5123a );
 a5133a <=( A265  and  A233 );
 a5134a <=( (not A232)  and  a5133a );
 a5138a <=( A268  and  A267 );
 a5139a <=( (not A266)  and  a5138a );
 a5140a <=( a5139a  and  a5134a );
 a5144a <=( A167  and  A169 );
 a5145a <=( (not A170)  and  a5144a );
 a5149a <=( (not A200)  and  (not A199) );
 a5150a <=( A166  and  a5149a );
 a5151a <=( a5150a  and  a5145a );
 a5155a <=( A265  and  A233 );
 a5156a <=( (not A232)  and  a5155a );
 a5160a <=( A269  and  A267 );
 a5161a <=( (not A266)  and  a5160a );
 a5162a <=( a5161a  and  a5156a );
 a5166a <=( A167  and  A169 );
 a5167a <=( (not A170)  and  a5166a );
 a5171a <=( (not A200)  and  (not A199) );
 a5172a <=( A166  and  a5171a );
 a5173a <=( a5172a  and  a5167a );
 a5177a <=( A234  and  (not A233) );
 a5178a <=( A232  and  a5177a );
 a5182a <=( A299  and  (not A298) );
 a5183a <=( A235  and  a5182a );
 a5184a <=( a5183a  and  a5178a );
 a5188a <=( A167  and  A169 );
 a5189a <=( (not A170)  and  a5188a );
 a5193a <=( (not A200)  and  (not A199) );
 a5194a <=( A166  and  a5193a );
 a5195a <=( a5194a  and  a5189a );
 a5199a <=( A234  and  (not A233) );
 a5200a <=( A232  and  a5199a );
 a5204a <=( A266  and  (not A265) );
 a5205a <=( A235  and  a5204a );
 a5206a <=( a5205a  and  a5200a );
 a5210a <=( A167  and  A169 );
 a5211a <=( (not A170)  and  a5210a );
 a5215a <=( (not A200)  and  (not A199) );
 a5216a <=( A166  and  a5215a );
 a5217a <=( a5216a  and  a5211a );
 a5221a <=( A234  and  (not A233) );
 a5222a <=( A232  and  a5221a );
 a5226a <=( A299  and  (not A298) );
 a5227a <=( A236  and  a5226a );
 a5228a <=( a5227a  and  a5222a );
 a5232a <=( A167  and  A169 );
 a5233a <=( (not A170)  and  a5232a );
 a5237a <=( (not A200)  and  (not A199) );
 a5238a <=( A166  and  a5237a );
 a5239a <=( a5238a  and  a5233a );
 a5243a <=( A234  and  (not A233) );
 a5244a <=( A232  and  a5243a );
 a5248a <=( A266  and  (not A265) );
 a5249a <=( A236  and  a5248a );
 a5250a <=( a5249a  and  a5244a );
 a5254a <=( (not A167)  and  A169 );
 a5255a <=( (not A170)  and  a5254a );
 a5259a <=( (not A201)  and  A199 );
 a5260a <=( (not A166)  and  a5259a );
 a5261a <=( a5260a  and  a5255a );
 a5265a <=( A298  and  A233 );
 a5266a <=( (not A232)  and  a5265a );
 a5270a <=( A301  and  A300 );
 a5271a <=( (not A299)  and  a5270a );
 a5272a <=( a5271a  and  a5266a );
 a5276a <=( (not A167)  and  A169 );
 a5277a <=( (not A170)  and  a5276a );
 a5281a <=( (not A201)  and  A199 );
 a5282a <=( (not A166)  and  a5281a );
 a5283a <=( a5282a  and  a5277a );
 a5287a <=( A298  and  A233 );
 a5288a <=( (not A232)  and  a5287a );
 a5292a <=( A302  and  A300 );
 a5293a <=( (not A299)  and  a5292a );
 a5294a <=( a5293a  and  a5288a );
 a5298a <=( (not A167)  and  A169 );
 a5299a <=( (not A170)  and  a5298a );
 a5303a <=( (not A201)  and  A199 );
 a5304a <=( (not A166)  and  a5303a );
 a5305a <=( a5304a  and  a5299a );
 a5309a <=( A265  and  A233 );
 a5310a <=( (not A232)  and  a5309a );
 a5314a <=( A268  and  A267 );
 a5315a <=( (not A266)  and  a5314a );
 a5316a <=( a5315a  and  a5310a );
 a5320a <=( (not A167)  and  A169 );
 a5321a <=( (not A170)  and  a5320a );
 a5325a <=( (not A201)  and  A199 );
 a5326a <=( (not A166)  and  a5325a );
 a5327a <=( a5326a  and  a5321a );
 a5331a <=( A265  and  A233 );
 a5332a <=( (not A232)  and  a5331a );
 a5336a <=( A269  and  A267 );
 a5337a <=( (not A266)  and  a5336a );
 a5338a <=( a5337a  and  a5332a );
 a5342a <=( (not A167)  and  A169 );
 a5343a <=( (not A170)  and  a5342a );
 a5347a <=( (not A201)  and  A199 );
 a5348a <=( (not A166)  and  a5347a );
 a5349a <=( a5348a  and  a5343a );
 a5353a <=( A234  and  (not A233) );
 a5354a <=( A232  and  a5353a );
 a5358a <=( A299  and  (not A298) );
 a5359a <=( A235  and  a5358a );
 a5360a <=( a5359a  and  a5354a );
 a5364a <=( (not A167)  and  A169 );
 a5365a <=( (not A170)  and  a5364a );
 a5369a <=( (not A201)  and  A199 );
 a5370a <=( (not A166)  and  a5369a );
 a5371a <=( a5370a  and  a5365a );
 a5375a <=( A234  and  (not A233) );
 a5376a <=( A232  and  a5375a );
 a5380a <=( A266  and  (not A265) );
 a5381a <=( A235  and  a5380a );
 a5382a <=( a5381a  and  a5376a );
 a5386a <=( (not A167)  and  A169 );
 a5387a <=( (not A170)  and  a5386a );
 a5391a <=( (not A201)  and  A199 );
 a5392a <=( (not A166)  and  a5391a );
 a5393a <=( a5392a  and  a5387a );
 a5397a <=( A234  and  (not A233) );
 a5398a <=( A232  and  a5397a );
 a5402a <=( A299  and  (not A298) );
 a5403a <=( A236  and  a5402a );
 a5404a <=( a5403a  and  a5398a );
 a5408a <=( (not A167)  and  A169 );
 a5409a <=( (not A170)  and  a5408a );
 a5413a <=( (not A201)  and  A199 );
 a5414a <=( (not A166)  and  a5413a );
 a5415a <=( a5414a  and  a5409a );
 a5419a <=( A234  and  (not A233) );
 a5420a <=( A232  and  a5419a );
 a5424a <=( A266  and  (not A265) );
 a5425a <=( A236  and  a5424a );
 a5426a <=( a5425a  and  a5420a );
 a5430a <=( (not A167)  and  A169 );
 a5431a <=( (not A170)  and  a5430a );
 a5435a <=( A200  and  A199 );
 a5436a <=( (not A166)  and  a5435a );
 a5437a <=( a5436a  and  a5431a );
 a5441a <=( A298  and  A233 );
 a5442a <=( (not A232)  and  a5441a );
 a5446a <=( A301  and  A300 );
 a5447a <=( (not A299)  and  a5446a );
 a5448a <=( a5447a  and  a5442a );
 a5452a <=( (not A167)  and  A169 );
 a5453a <=( (not A170)  and  a5452a );
 a5457a <=( A200  and  A199 );
 a5458a <=( (not A166)  and  a5457a );
 a5459a <=( a5458a  and  a5453a );
 a5463a <=( A298  and  A233 );
 a5464a <=( (not A232)  and  a5463a );
 a5468a <=( A302  and  A300 );
 a5469a <=( (not A299)  and  a5468a );
 a5470a <=( a5469a  and  a5464a );
 a5474a <=( (not A167)  and  A169 );
 a5475a <=( (not A170)  and  a5474a );
 a5479a <=( A200  and  A199 );
 a5480a <=( (not A166)  and  a5479a );
 a5481a <=( a5480a  and  a5475a );
 a5485a <=( A265  and  A233 );
 a5486a <=( (not A232)  and  a5485a );
 a5490a <=( A268  and  A267 );
 a5491a <=( (not A266)  and  a5490a );
 a5492a <=( a5491a  and  a5486a );
 a5496a <=( (not A167)  and  A169 );
 a5497a <=( (not A170)  and  a5496a );
 a5501a <=( A200  and  A199 );
 a5502a <=( (not A166)  and  a5501a );
 a5503a <=( a5502a  and  a5497a );
 a5507a <=( A265  and  A233 );
 a5508a <=( (not A232)  and  a5507a );
 a5512a <=( A269  and  A267 );
 a5513a <=( (not A266)  and  a5512a );
 a5514a <=( a5513a  and  a5508a );
 a5518a <=( (not A167)  and  A169 );
 a5519a <=( (not A170)  and  a5518a );
 a5523a <=( A200  and  A199 );
 a5524a <=( (not A166)  and  a5523a );
 a5525a <=( a5524a  and  a5519a );
 a5529a <=( A234  and  (not A233) );
 a5530a <=( A232  and  a5529a );
 a5534a <=( A299  and  (not A298) );
 a5535a <=( A235  and  a5534a );
 a5536a <=( a5535a  and  a5530a );
 a5540a <=( (not A167)  and  A169 );
 a5541a <=( (not A170)  and  a5540a );
 a5545a <=( A200  and  A199 );
 a5546a <=( (not A166)  and  a5545a );
 a5547a <=( a5546a  and  a5541a );
 a5551a <=( A234  and  (not A233) );
 a5552a <=( A232  and  a5551a );
 a5556a <=( A266  and  (not A265) );
 a5557a <=( A235  and  a5556a );
 a5558a <=( a5557a  and  a5552a );
 a5562a <=( (not A167)  and  A169 );
 a5563a <=( (not A170)  and  a5562a );
 a5567a <=( A200  and  A199 );
 a5568a <=( (not A166)  and  a5567a );
 a5569a <=( a5568a  and  a5563a );
 a5573a <=( A234  and  (not A233) );
 a5574a <=( A232  and  a5573a );
 a5578a <=( A299  and  (not A298) );
 a5579a <=( A236  and  a5578a );
 a5580a <=( a5579a  and  a5574a );
 a5584a <=( (not A167)  and  A169 );
 a5585a <=( (not A170)  and  a5584a );
 a5589a <=( A200  and  A199 );
 a5590a <=( (not A166)  and  a5589a );
 a5591a <=( a5590a  and  a5585a );
 a5595a <=( A234  and  (not A233) );
 a5596a <=( A232  and  a5595a );
 a5600a <=( A266  and  (not A265) );
 a5601a <=( A236  and  a5600a );
 a5602a <=( a5601a  and  a5596a );
 a5606a <=( (not A167)  and  A169 );
 a5607a <=( (not A170)  and  a5606a );
 a5611a <=( (not A200)  and  (not A199) );
 a5612a <=( (not A166)  and  a5611a );
 a5613a <=( a5612a  and  a5607a );
 a5617a <=( A298  and  A233 );
 a5618a <=( (not A232)  and  a5617a );
 a5622a <=( A301  and  A300 );
 a5623a <=( (not A299)  and  a5622a );
 a5624a <=( a5623a  and  a5618a );
 a5628a <=( (not A167)  and  A169 );
 a5629a <=( (not A170)  and  a5628a );
 a5633a <=( (not A200)  and  (not A199) );
 a5634a <=( (not A166)  and  a5633a );
 a5635a <=( a5634a  and  a5629a );
 a5639a <=( A298  and  A233 );
 a5640a <=( (not A232)  and  a5639a );
 a5644a <=( A302  and  A300 );
 a5645a <=( (not A299)  and  a5644a );
 a5646a <=( a5645a  and  a5640a );
 a5650a <=( (not A167)  and  A169 );
 a5651a <=( (not A170)  and  a5650a );
 a5655a <=( (not A200)  and  (not A199) );
 a5656a <=( (not A166)  and  a5655a );
 a5657a <=( a5656a  and  a5651a );
 a5661a <=( A265  and  A233 );
 a5662a <=( (not A232)  and  a5661a );
 a5666a <=( A268  and  A267 );
 a5667a <=( (not A266)  and  a5666a );
 a5668a <=( a5667a  and  a5662a );
 a5672a <=( (not A167)  and  A169 );
 a5673a <=( (not A170)  and  a5672a );
 a5677a <=( (not A200)  and  (not A199) );
 a5678a <=( (not A166)  and  a5677a );
 a5679a <=( a5678a  and  a5673a );
 a5683a <=( A265  and  A233 );
 a5684a <=( (not A232)  and  a5683a );
 a5688a <=( A269  and  A267 );
 a5689a <=( (not A266)  and  a5688a );
 a5690a <=( a5689a  and  a5684a );
 a5694a <=( (not A167)  and  A169 );
 a5695a <=( (not A170)  and  a5694a );
 a5699a <=( (not A200)  and  (not A199) );
 a5700a <=( (not A166)  and  a5699a );
 a5701a <=( a5700a  and  a5695a );
 a5705a <=( A234  and  (not A233) );
 a5706a <=( A232  and  a5705a );
 a5710a <=( A299  and  (not A298) );
 a5711a <=( A235  and  a5710a );
 a5712a <=( a5711a  and  a5706a );
 a5716a <=( (not A167)  and  A169 );
 a5717a <=( (not A170)  and  a5716a );
 a5721a <=( (not A200)  and  (not A199) );
 a5722a <=( (not A166)  and  a5721a );
 a5723a <=( a5722a  and  a5717a );
 a5727a <=( A234  and  (not A233) );
 a5728a <=( A232  and  a5727a );
 a5732a <=( A266  and  (not A265) );
 a5733a <=( A235  and  a5732a );
 a5734a <=( a5733a  and  a5728a );
 a5738a <=( (not A167)  and  A169 );
 a5739a <=( (not A170)  and  a5738a );
 a5743a <=( (not A200)  and  (not A199) );
 a5744a <=( (not A166)  and  a5743a );
 a5745a <=( a5744a  and  a5739a );
 a5749a <=( A234  and  (not A233) );
 a5750a <=( A232  and  a5749a );
 a5754a <=( A299  and  (not A298) );
 a5755a <=( A236  and  a5754a );
 a5756a <=( a5755a  and  a5750a );
 a5760a <=( (not A167)  and  A169 );
 a5761a <=( (not A170)  and  a5760a );
 a5765a <=( (not A200)  and  (not A199) );
 a5766a <=( (not A166)  and  a5765a );
 a5767a <=( a5766a  and  a5761a );
 a5771a <=( A234  and  (not A233) );
 a5772a <=( A232  and  a5771a );
 a5776a <=( A266  and  (not A265) );
 a5777a <=( A236  and  a5776a );
 a5778a <=( a5777a  and  a5772a );
 a5782a <=( A167  and  (not A169) );
 a5783a <=( A170  and  a5782a );
 a5787a <=( (not A201)  and  A199 );
 a5788a <=( (not A166)  and  a5787a );
 a5789a <=( a5788a  and  a5783a );
 a5793a <=( A298  and  A233 );
 a5794a <=( (not A232)  and  a5793a );
 a5798a <=( A301  and  A300 );
 a5799a <=( (not A299)  and  a5798a );
 a5800a <=( a5799a  and  a5794a );
 a5804a <=( A167  and  (not A169) );
 a5805a <=( A170  and  a5804a );
 a5809a <=( (not A201)  and  A199 );
 a5810a <=( (not A166)  and  a5809a );
 a5811a <=( a5810a  and  a5805a );
 a5815a <=( A298  and  A233 );
 a5816a <=( (not A232)  and  a5815a );
 a5820a <=( A302  and  A300 );
 a5821a <=( (not A299)  and  a5820a );
 a5822a <=( a5821a  and  a5816a );
 a5826a <=( A167  and  (not A169) );
 a5827a <=( A170  and  a5826a );
 a5831a <=( (not A201)  and  A199 );
 a5832a <=( (not A166)  and  a5831a );
 a5833a <=( a5832a  and  a5827a );
 a5837a <=( A265  and  A233 );
 a5838a <=( (not A232)  and  a5837a );
 a5842a <=( A268  and  A267 );
 a5843a <=( (not A266)  and  a5842a );
 a5844a <=( a5843a  and  a5838a );
 a5848a <=( A167  and  (not A169) );
 a5849a <=( A170  and  a5848a );
 a5853a <=( (not A201)  and  A199 );
 a5854a <=( (not A166)  and  a5853a );
 a5855a <=( a5854a  and  a5849a );
 a5859a <=( A265  and  A233 );
 a5860a <=( (not A232)  and  a5859a );
 a5864a <=( A269  and  A267 );
 a5865a <=( (not A266)  and  a5864a );
 a5866a <=( a5865a  and  a5860a );
 a5870a <=( A167  and  (not A169) );
 a5871a <=( A170  and  a5870a );
 a5875a <=( (not A201)  and  A199 );
 a5876a <=( (not A166)  and  a5875a );
 a5877a <=( a5876a  and  a5871a );
 a5881a <=( A234  and  (not A233) );
 a5882a <=( A232  and  a5881a );
 a5886a <=( A299  and  (not A298) );
 a5887a <=( A235  and  a5886a );
 a5888a <=( a5887a  and  a5882a );
 a5892a <=( A167  and  (not A169) );
 a5893a <=( A170  and  a5892a );
 a5897a <=( (not A201)  and  A199 );
 a5898a <=( (not A166)  and  a5897a );
 a5899a <=( a5898a  and  a5893a );
 a5903a <=( A234  and  (not A233) );
 a5904a <=( A232  and  a5903a );
 a5908a <=( A266  and  (not A265) );
 a5909a <=( A235  and  a5908a );
 a5910a <=( a5909a  and  a5904a );
 a5914a <=( A167  and  (not A169) );
 a5915a <=( A170  and  a5914a );
 a5919a <=( (not A201)  and  A199 );
 a5920a <=( (not A166)  and  a5919a );
 a5921a <=( a5920a  and  a5915a );
 a5925a <=( A234  and  (not A233) );
 a5926a <=( A232  and  a5925a );
 a5930a <=( A299  and  (not A298) );
 a5931a <=( A236  and  a5930a );
 a5932a <=( a5931a  and  a5926a );
 a5936a <=( A167  and  (not A169) );
 a5937a <=( A170  and  a5936a );
 a5941a <=( (not A201)  and  A199 );
 a5942a <=( (not A166)  and  a5941a );
 a5943a <=( a5942a  and  a5937a );
 a5947a <=( A234  and  (not A233) );
 a5948a <=( A232  and  a5947a );
 a5952a <=( A266  and  (not A265) );
 a5953a <=( A236  and  a5952a );
 a5954a <=( a5953a  and  a5948a );
 a5958a <=( A167  and  (not A169) );
 a5959a <=( A170  and  a5958a );
 a5963a <=( A200  and  A199 );
 a5964a <=( (not A166)  and  a5963a );
 a5965a <=( a5964a  and  a5959a );
 a5969a <=( A298  and  A233 );
 a5970a <=( (not A232)  and  a5969a );
 a5974a <=( A301  and  A300 );
 a5975a <=( (not A299)  and  a5974a );
 a5976a <=( a5975a  and  a5970a );
 a5980a <=( A167  and  (not A169) );
 a5981a <=( A170  and  a5980a );
 a5985a <=( A200  and  A199 );
 a5986a <=( (not A166)  and  a5985a );
 a5987a <=( a5986a  and  a5981a );
 a5991a <=( A298  and  A233 );
 a5992a <=( (not A232)  and  a5991a );
 a5996a <=( A302  and  A300 );
 a5997a <=( (not A299)  and  a5996a );
 a5998a <=( a5997a  and  a5992a );
 a6002a <=( A167  and  (not A169) );
 a6003a <=( A170  and  a6002a );
 a6007a <=( A200  and  A199 );
 a6008a <=( (not A166)  and  a6007a );
 a6009a <=( a6008a  and  a6003a );
 a6013a <=( A265  and  A233 );
 a6014a <=( (not A232)  and  a6013a );
 a6018a <=( A268  and  A267 );
 a6019a <=( (not A266)  and  a6018a );
 a6020a <=( a6019a  and  a6014a );
 a6024a <=( A167  and  (not A169) );
 a6025a <=( A170  and  a6024a );
 a6029a <=( A200  and  A199 );
 a6030a <=( (not A166)  and  a6029a );
 a6031a <=( a6030a  and  a6025a );
 a6035a <=( A265  and  A233 );
 a6036a <=( (not A232)  and  a6035a );
 a6040a <=( A269  and  A267 );
 a6041a <=( (not A266)  and  a6040a );
 a6042a <=( a6041a  and  a6036a );
 a6046a <=( A167  and  (not A169) );
 a6047a <=( A170  and  a6046a );
 a6051a <=( A200  and  A199 );
 a6052a <=( (not A166)  and  a6051a );
 a6053a <=( a6052a  and  a6047a );
 a6057a <=( A234  and  (not A233) );
 a6058a <=( A232  and  a6057a );
 a6062a <=( A299  and  (not A298) );
 a6063a <=( A235  and  a6062a );
 a6064a <=( a6063a  and  a6058a );
 a6068a <=( A167  and  (not A169) );
 a6069a <=( A170  and  a6068a );
 a6073a <=( A200  and  A199 );
 a6074a <=( (not A166)  and  a6073a );
 a6075a <=( a6074a  and  a6069a );
 a6079a <=( A234  and  (not A233) );
 a6080a <=( A232  and  a6079a );
 a6084a <=( A266  and  (not A265) );
 a6085a <=( A235  and  a6084a );
 a6086a <=( a6085a  and  a6080a );
 a6090a <=( A167  and  (not A169) );
 a6091a <=( A170  and  a6090a );
 a6095a <=( A200  and  A199 );
 a6096a <=( (not A166)  and  a6095a );
 a6097a <=( a6096a  and  a6091a );
 a6101a <=( A234  and  (not A233) );
 a6102a <=( A232  and  a6101a );
 a6106a <=( A299  and  (not A298) );
 a6107a <=( A236  and  a6106a );
 a6108a <=( a6107a  and  a6102a );
 a6112a <=( A167  and  (not A169) );
 a6113a <=( A170  and  a6112a );
 a6117a <=( A200  and  A199 );
 a6118a <=( (not A166)  and  a6117a );
 a6119a <=( a6118a  and  a6113a );
 a6123a <=( A234  and  (not A233) );
 a6124a <=( A232  and  a6123a );
 a6128a <=( A266  and  (not A265) );
 a6129a <=( A236  and  a6128a );
 a6130a <=( a6129a  and  a6124a );
 a6134a <=( A167  and  (not A169) );
 a6135a <=( A170  and  a6134a );
 a6139a <=( (not A200)  and  (not A199) );
 a6140a <=( (not A166)  and  a6139a );
 a6141a <=( a6140a  and  a6135a );
 a6145a <=( A298  and  A233 );
 a6146a <=( (not A232)  and  a6145a );
 a6150a <=( A301  and  A300 );
 a6151a <=( (not A299)  and  a6150a );
 a6152a <=( a6151a  and  a6146a );
 a6156a <=( A167  and  (not A169) );
 a6157a <=( A170  and  a6156a );
 a6161a <=( (not A200)  and  (not A199) );
 a6162a <=( (not A166)  and  a6161a );
 a6163a <=( a6162a  and  a6157a );
 a6167a <=( A298  and  A233 );
 a6168a <=( (not A232)  and  a6167a );
 a6172a <=( A302  and  A300 );
 a6173a <=( (not A299)  and  a6172a );
 a6174a <=( a6173a  and  a6168a );
 a6178a <=( A167  and  (not A169) );
 a6179a <=( A170  and  a6178a );
 a6183a <=( (not A200)  and  (not A199) );
 a6184a <=( (not A166)  and  a6183a );
 a6185a <=( a6184a  and  a6179a );
 a6189a <=( A265  and  A233 );
 a6190a <=( (not A232)  and  a6189a );
 a6194a <=( A268  and  A267 );
 a6195a <=( (not A266)  and  a6194a );
 a6196a <=( a6195a  and  a6190a );
 a6200a <=( A167  and  (not A169) );
 a6201a <=( A170  and  a6200a );
 a6205a <=( (not A200)  and  (not A199) );
 a6206a <=( (not A166)  and  a6205a );
 a6207a <=( a6206a  and  a6201a );
 a6211a <=( A265  and  A233 );
 a6212a <=( (not A232)  and  a6211a );
 a6216a <=( A269  and  A267 );
 a6217a <=( (not A266)  and  a6216a );
 a6218a <=( a6217a  and  a6212a );
 a6222a <=( A167  and  (not A169) );
 a6223a <=( A170  and  a6222a );
 a6227a <=( (not A200)  and  (not A199) );
 a6228a <=( (not A166)  and  a6227a );
 a6229a <=( a6228a  and  a6223a );
 a6233a <=( A234  and  (not A233) );
 a6234a <=( A232  and  a6233a );
 a6238a <=( A299  and  (not A298) );
 a6239a <=( A235  and  a6238a );
 a6240a <=( a6239a  and  a6234a );
 a6244a <=( A167  and  (not A169) );
 a6245a <=( A170  and  a6244a );
 a6249a <=( (not A200)  and  (not A199) );
 a6250a <=( (not A166)  and  a6249a );
 a6251a <=( a6250a  and  a6245a );
 a6255a <=( A234  and  (not A233) );
 a6256a <=( A232  and  a6255a );
 a6260a <=( A266  and  (not A265) );
 a6261a <=( A235  and  a6260a );
 a6262a <=( a6261a  and  a6256a );
 a6266a <=( A167  and  (not A169) );
 a6267a <=( A170  and  a6266a );
 a6271a <=( (not A200)  and  (not A199) );
 a6272a <=( (not A166)  and  a6271a );
 a6273a <=( a6272a  and  a6267a );
 a6277a <=( A234  and  (not A233) );
 a6278a <=( A232  and  a6277a );
 a6282a <=( A299  and  (not A298) );
 a6283a <=( A236  and  a6282a );
 a6284a <=( a6283a  and  a6278a );
 a6288a <=( A167  and  (not A169) );
 a6289a <=( A170  and  a6288a );
 a6293a <=( (not A200)  and  (not A199) );
 a6294a <=( (not A166)  and  a6293a );
 a6295a <=( a6294a  and  a6289a );
 a6299a <=( A234  and  (not A233) );
 a6300a <=( A232  and  a6299a );
 a6304a <=( A266  and  (not A265) );
 a6305a <=( A236  and  a6304a );
 a6306a <=( a6305a  and  a6300a );
 a6310a <=( (not A167)  and  (not A169) );
 a6311a <=( A170  and  a6310a );
 a6315a <=( (not A201)  and  A199 );
 a6316a <=( A166  and  a6315a );
 a6317a <=( a6316a  and  a6311a );
 a6321a <=( A298  and  A233 );
 a6322a <=( (not A232)  and  a6321a );
 a6326a <=( A301  and  A300 );
 a6327a <=( (not A299)  and  a6326a );
 a6328a <=( a6327a  and  a6322a );
 a6332a <=( (not A167)  and  (not A169) );
 a6333a <=( A170  and  a6332a );
 a6337a <=( (not A201)  and  A199 );
 a6338a <=( A166  and  a6337a );
 a6339a <=( a6338a  and  a6333a );
 a6343a <=( A298  and  A233 );
 a6344a <=( (not A232)  and  a6343a );
 a6348a <=( A302  and  A300 );
 a6349a <=( (not A299)  and  a6348a );
 a6350a <=( a6349a  and  a6344a );
 a6354a <=( (not A167)  and  (not A169) );
 a6355a <=( A170  and  a6354a );
 a6359a <=( (not A201)  and  A199 );
 a6360a <=( A166  and  a6359a );
 a6361a <=( a6360a  and  a6355a );
 a6365a <=( A265  and  A233 );
 a6366a <=( (not A232)  and  a6365a );
 a6370a <=( A268  and  A267 );
 a6371a <=( (not A266)  and  a6370a );
 a6372a <=( a6371a  and  a6366a );
 a6376a <=( (not A167)  and  (not A169) );
 a6377a <=( A170  and  a6376a );
 a6381a <=( (not A201)  and  A199 );
 a6382a <=( A166  and  a6381a );
 a6383a <=( a6382a  and  a6377a );
 a6387a <=( A265  and  A233 );
 a6388a <=( (not A232)  and  a6387a );
 a6392a <=( A269  and  A267 );
 a6393a <=( (not A266)  and  a6392a );
 a6394a <=( a6393a  and  a6388a );
 a6398a <=( (not A167)  and  (not A169) );
 a6399a <=( A170  and  a6398a );
 a6403a <=( (not A201)  and  A199 );
 a6404a <=( A166  and  a6403a );
 a6405a <=( a6404a  and  a6399a );
 a6409a <=( A234  and  (not A233) );
 a6410a <=( A232  and  a6409a );
 a6414a <=( A299  and  (not A298) );
 a6415a <=( A235  and  a6414a );
 a6416a <=( a6415a  and  a6410a );
 a6420a <=( (not A167)  and  (not A169) );
 a6421a <=( A170  and  a6420a );
 a6425a <=( (not A201)  and  A199 );
 a6426a <=( A166  and  a6425a );
 a6427a <=( a6426a  and  a6421a );
 a6431a <=( A234  and  (not A233) );
 a6432a <=( A232  and  a6431a );
 a6436a <=( A266  and  (not A265) );
 a6437a <=( A235  and  a6436a );
 a6438a <=( a6437a  and  a6432a );
 a6442a <=( (not A167)  and  (not A169) );
 a6443a <=( A170  and  a6442a );
 a6447a <=( (not A201)  and  A199 );
 a6448a <=( A166  and  a6447a );
 a6449a <=( a6448a  and  a6443a );
 a6453a <=( A234  and  (not A233) );
 a6454a <=( A232  and  a6453a );
 a6458a <=( A299  and  (not A298) );
 a6459a <=( A236  and  a6458a );
 a6460a <=( a6459a  and  a6454a );
 a6464a <=( (not A167)  and  (not A169) );
 a6465a <=( A170  and  a6464a );
 a6469a <=( (not A201)  and  A199 );
 a6470a <=( A166  and  a6469a );
 a6471a <=( a6470a  and  a6465a );
 a6475a <=( A234  and  (not A233) );
 a6476a <=( A232  and  a6475a );
 a6480a <=( A266  and  (not A265) );
 a6481a <=( A236  and  a6480a );
 a6482a <=( a6481a  and  a6476a );
 a6486a <=( (not A167)  and  (not A169) );
 a6487a <=( A170  and  a6486a );
 a6491a <=( A200  and  A199 );
 a6492a <=( A166  and  a6491a );
 a6493a <=( a6492a  and  a6487a );
 a6497a <=( A298  and  A233 );
 a6498a <=( (not A232)  and  a6497a );
 a6502a <=( A301  and  A300 );
 a6503a <=( (not A299)  and  a6502a );
 a6504a <=( a6503a  and  a6498a );
 a6508a <=( (not A167)  and  (not A169) );
 a6509a <=( A170  and  a6508a );
 a6513a <=( A200  and  A199 );
 a6514a <=( A166  and  a6513a );
 a6515a <=( a6514a  and  a6509a );
 a6519a <=( A298  and  A233 );
 a6520a <=( (not A232)  and  a6519a );
 a6524a <=( A302  and  A300 );
 a6525a <=( (not A299)  and  a6524a );
 a6526a <=( a6525a  and  a6520a );
 a6530a <=( (not A167)  and  (not A169) );
 a6531a <=( A170  and  a6530a );
 a6535a <=( A200  and  A199 );
 a6536a <=( A166  and  a6535a );
 a6537a <=( a6536a  and  a6531a );
 a6541a <=( A265  and  A233 );
 a6542a <=( (not A232)  and  a6541a );
 a6546a <=( A268  and  A267 );
 a6547a <=( (not A266)  and  a6546a );
 a6548a <=( a6547a  and  a6542a );
 a6552a <=( (not A167)  and  (not A169) );
 a6553a <=( A170  and  a6552a );
 a6557a <=( A200  and  A199 );
 a6558a <=( A166  and  a6557a );
 a6559a <=( a6558a  and  a6553a );
 a6563a <=( A265  and  A233 );
 a6564a <=( (not A232)  and  a6563a );
 a6568a <=( A269  and  A267 );
 a6569a <=( (not A266)  and  a6568a );
 a6570a <=( a6569a  and  a6564a );
 a6574a <=( (not A167)  and  (not A169) );
 a6575a <=( A170  and  a6574a );
 a6579a <=( A200  and  A199 );
 a6580a <=( A166  and  a6579a );
 a6581a <=( a6580a  and  a6575a );
 a6585a <=( A234  and  (not A233) );
 a6586a <=( A232  and  a6585a );
 a6590a <=( A299  and  (not A298) );
 a6591a <=( A235  and  a6590a );
 a6592a <=( a6591a  and  a6586a );
 a6596a <=( (not A167)  and  (not A169) );
 a6597a <=( A170  and  a6596a );
 a6601a <=( A200  and  A199 );
 a6602a <=( A166  and  a6601a );
 a6603a <=( a6602a  and  a6597a );
 a6607a <=( A234  and  (not A233) );
 a6608a <=( A232  and  a6607a );
 a6612a <=( A266  and  (not A265) );
 a6613a <=( A235  and  a6612a );
 a6614a <=( a6613a  and  a6608a );
 a6618a <=( (not A167)  and  (not A169) );
 a6619a <=( A170  and  a6618a );
 a6623a <=( A200  and  A199 );
 a6624a <=( A166  and  a6623a );
 a6625a <=( a6624a  and  a6619a );
 a6629a <=( A234  and  (not A233) );
 a6630a <=( A232  and  a6629a );
 a6634a <=( A299  and  (not A298) );
 a6635a <=( A236  and  a6634a );
 a6636a <=( a6635a  and  a6630a );
 a6640a <=( (not A167)  and  (not A169) );
 a6641a <=( A170  and  a6640a );
 a6645a <=( A200  and  A199 );
 a6646a <=( A166  and  a6645a );
 a6647a <=( a6646a  and  a6641a );
 a6651a <=( A234  and  (not A233) );
 a6652a <=( A232  and  a6651a );
 a6656a <=( A266  and  (not A265) );
 a6657a <=( A236  and  a6656a );
 a6658a <=( a6657a  and  a6652a );
 a6662a <=( (not A167)  and  (not A169) );
 a6663a <=( A170  and  a6662a );
 a6667a <=( (not A200)  and  (not A199) );
 a6668a <=( A166  and  a6667a );
 a6669a <=( a6668a  and  a6663a );
 a6673a <=( A298  and  A233 );
 a6674a <=( (not A232)  and  a6673a );
 a6678a <=( A301  and  A300 );
 a6679a <=( (not A299)  and  a6678a );
 a6680a <=( a6679a  and  a6674a );
 a6684a <=( (not A167)  and  (not A169) );
 a6685a <=( A170  and  a6684a );
 a6689a <=( (not A200)  and  (not A199) );
 a6690a <=( A166  and  a6689a );
 a6691a <=( a6690a  and  a6685a );
 a6695a <=( A298  and  A233 );
 a6696a <=( (not A232)  and  a6695a );
 a6700a <=( A302  and  A300 );
 a6701a <=( (not A299)  and  a6700a );
 a6702a <=( a6701a  and  a6696a );
 a6706a <=( (not A167)  and  (not A169) );
 a6707a <=( A170  and  a6706a );
 a6711a <=( (not A200)  and  (not A199) );
 a6712a <=( A166  and  a6711a );
 a6713a <=( a6712a  and  a6707a );
 a6717a <=( A265  and  A233 );
 a6718a <=( (not A232)  and  a6717a );
 a6722a <=( A268  and  A267 );
 a6723a <=( (not A266)  and  a6722a );
 a6724a <=( a6723a  and  a6718a );
 a6728a <=( (not A167)  and  (not A169) );
 a6729a <=( A170  and  a6728a );
 a6733a <=( (not A200)  and  (not A199) );
 a6734a <=( A166  and  a6733a );
 a6735a <=( a6734a  and  a6729a );
 a6739a <=( A265  and  A233 );
 a6740a <=( (not A232)  and  a6739a );
 a6744a <=( A269  and  A267 );
 a6745a <=( (not A266)  and  a6744a );
 a6746a <=( a6745a  and  a6740a );
 a6750a <=( (not A167)  and  (not A169) );
 a6751a <=( A170  and  a6750a );
 a6755a <=( (not A200)  and  (not A199) );
 a6756a <=( A166  and  a6755a );
 a6757a <=( a6756a  and  a6751a );
 a6761a <=( A234  and  (not A233) );
 a6762a <=( A232  and  a6761a );
 a6766a <=( A299  and  (not A298) );
 a6767a <=( A235  and  a6766a );
 a6768a <=( a6767a  and  a6762a );
 a6772a <=( (not A167)  and  (not A169) );
 a6773a <=( A170  and  a6772a );
 a6777a <=( (not A200)  and  (not A199) );
 a6778a <=( A166  and  a6777a );
 a6779a <=( a6778a  and  a6773a );
 a6783a <=( A234  and  (not A233) );
 a6784a <=( A232  and  a6783a );
 a6788a <=( A266  and  (not A265) );
 a6789a <=( A235  and  a6788a );
 a6790a <=( a6789a  and  a6784a );
 a6794a <=( (not A167)  and  (not A169) );
 a6795a <=( A170  and  a6794a );
 a6799a <=( (not A200)  and  (not A199) );
 a6800a <=( A166  and  a6799a );
 a6801a <=( a6800a  and  a6795a );
 a6805a <=( A234  and  (not A233) );
 a6806a <=( A232  and  a6805a );
 a6810a <=( A299  and  (not A298) );
 a6811a <=( A236  and  a6810a );
 a6812a <=( a6811a  and  a6806a );
 a6816a <=( (not A167)  and  (not A169) );
 a6817a <=( A170  and  a6816a );
 a6821a <=( (not A200)  and  (not A199) );
 a6822a <=( A166  and  a6821a );
 a6823a <=( a6822a  and  a6817a );
 a6827a <=( A234  and  (not A233) );
 a6828a <=( A232  and  a6827a );
 a6832a <=( A266  and  (not A265) );
 a6833a <=( A236  and  a6832a );
 a6834a <=( a6833a  and  a6828a );
 a6838a <=( A199  and  A166 );
 a6839a <=( A168  and  a6838a );
 a6843a <=( A232  and  (not A203) );
 a6844a <=( (not A202)  and  a6843a );
 a6845a <=( a6844a  and  a6839a );
 a6849a <=( A235  and  A234 );
 a6850a <=( (not A233)  and  a6849a );
 a6853a <=( (not A299)  and  A298 );
 a6856a <=( A301  and  A300 );
 a6857a <=( a6856a  and  a6853a );
 a6858a <=( a6857a  and  a6850a );
 a6862a <=( A199  and  A166 );
 a6863a <=( A168  and  a6862a );
 a6867a <=( A232  and  (not A203) );
 a6868a <=( (not A202)  and  a6867a );
 a6869a <=( a6868a  and  a6863a );
 a6873a <=( A235  and  A234 );
 a6874a <=( (not A233)  and  a6873a );
 a6877a <=( (not A299)  and  A298 );
 a6880a <=( A302  and  A300 );
 a6881a <=( a6880a  and  a6877a );
 a6882a <=( a6881a  and  a6874a );
 a6886a <=( A199  and  A166 );
 a6887a <=( A168  and  a6886a );
 a6891a <=( A232  and  (not A203) );
 a6892a <=( (not A202)  and  a6891a );
 a6893a <=( a6892a  and  a6887a );
 a6897a <=( A235  and  A234 );
 a6898a <=( (not A233)  and  a6897a );
 a6901a <=( (not A266)  and  A265 );
 a6904a <=( A268  and  A267 );
 a6905a <=( a6904a  and  a6901a );
 a6906a <=( a6905a  and  a6898a );
 a6910a <=( A199  and  A166 );
 a6911a <=( A168  and  a6910a );
 a6915a <=( A232  and  (not A203) );
 a6916a <=( (not A202)  and  a6915a );
 a6917a <=( a6916a  and  a6911a );
 a6921a <=( A235  and  A234 );
 a6922a <=( (not A233)  and  a6921a );
 a6925a <=( (not A266)  and  A265 );
 a6928a <=( A269  and  A267 );
 a6929a <=( a6928a  and  a6925a );
 a6930a <=( a6929a  and  a6922a );
 a6934a <=( A199  and  A166 );
 a6935a <=( A168  and  a6934a );
 a6939a <=( A232  and  (not A203) );
 a6940a <=( (not A202)  and  a6939a );
 a6941a <=( a6940a  and  a6935a );
 a6945a <=( A236  and  A234 );
 a6946a <=( (not A233)  and  a6945a );
 a6949a <=( (not A299)  and  A298 );
 a6952a <=( A301  and  A300 );
 a6953a <=( a6952a  and  a6949a );
 a6954a <=( a6953a  and  a6946a );
 a6958a <=( A199  and  A166 );
 a6959a <=( A168  and  a6958a );
 a6963a <=( A232  and  (not A203) );
 a6964a <=( (not A202)  and  a6963a );
 a6965a <=( a6964a  and  a6959a );
 a6969a <=( A236  and  A234 );
 a6970a <=( (not A233)  and  a6969a );
 a6973a <=( (not A299)  and  A298 );
 a6976a <=( A302  and  A300 );
 a6977a <=( a6976a  and  a6973a );
 a6978a <=( a6977a  and  a6970a );
 a6982a <=( A199  and  A166 );
 a6983a <=( A168  and  a6982a );
 a6987a <=( A232  and  (not A203) );
 a6988a <=( (not A202)  and  a6987a );
 a6989a <=( a6988a  and  a6983a );
 a6993a <=( A236  and  A234 );
 a6994a <=( (not A233)  and  a6993a );
 a6997a <=( (not A266)  and  A265 );
 a7000a <=( A268  and  A267 );
 a7001a <=( a7000a  and  a6997a );
 a7002a <=( a7001a  and  a6994a );
 a7006a <=( A199  and  A166 );
 a7007a <=( A168  and  a7006a );
 a7011a <=( A232  and  (not A203) );
 a7012a <=( (not A202)  and  a7011a );
 a7013a <=( a7012a  and  a7007a );
 a7017a <=( A236  and  A234 );
 a7018a <=( (not A233)  and  a7017a );
 a7021a <=( (not A266)  and  A265 );
 a7024a <=( A269  and  A267 );
 a7025a <=( a7024a  and  a7021a );
 a7026a <=( a7025a  and  a7018a );
 a7030a <=( A199  and  A167 );
 a7031a <=( A168  and  a7030a );
 a7035a <=( A232  and  (not A203) );
 a7036a <=( (not A202)  and  a7035a );
 a7037a <=( a7036a  and  a7031a );
 a7041a <=( A235  and  A234 );
 a7042a <=( (not A233)  and  a7041a );
 a7045a <=( (not A299)  and  A298 );
 a7048a <=( A301  and  A300 );
 a7049a <=( a7048a  and  a7045a );
 a7050a <=( a7049a  and  a7042a );
 a7054a <=( A199  and  A167 );
 a7055a <=( A168  and  a7054a );
 a7059a <=( A232  and  (not A203) );
 a7060a <=( (not A202)  and  a7059a );
 a7061a <=( a7060a  and  a7055a );
 a7065a <=( A235  and  A234 );
 a7066a <=( (not A233)  and  a7065a );
 a7069a <=( (not A299)  and  A298 );
 a7072a <=( A302  and  A300 );
 a7073a <=( a7072a  and  a7069a );
 a7074a <=( a7073a  and  a7066a );
 a7078a <=( A199  and  A167 );
 a7079a <=( A168  and  a7078a );
 a7083a <=( A232  and  (not A203) );
 a7084a <=( (not A202)  and  a7083a );
 a7085a <=( a7084a  and  a7079a );
 a7089a <=( A235  and  A234 );
 a7090a <=( (not A233)  and  a7089a );
 a7093a <=( (not A266)  and  A265 );
 a7096a <=( A268  and  A267 );
 a7097a <=( a7096a  and  a7093a );
 a7098a <=( a7097a  and  a7090a );
 a7102a <=( A199  and  A167 );
 a7103a <=( A168  and  a7102a );
 a7107a <=( A232  and  (not A203) );
 a7108a <=( (not A202)  and  a7107a );
 a7109a <=( a7108a  and  a7103a );
 a7113a <=( A235  and  A234 );
 a7114a <=( (not A233)  and  a7113a );
 a7117a <=( (not A266)  and  A265 );
 a7120a <=( A269  and  A267 );
 a7121a <=( a7120a  and  a7117a );
 a7122a <=( a7121a  and  a7114a );
 a7126a <=( A199  and  A167 );
 a7127a <=( A168  and  a7126a );
 a7131a <=( A232  and  (not A203) );
 a7132a <=( (not A202)  and  a7131a );
 a7133a <=( a7132a  and  a7127a );
 a7137a <=( A236  and  A234 );
 a7138a <=( (not A233)  and  a7137a );
 a7141a <=( (not A299)  and  A298 );
 a7144a <=( A301  and  A300 );
 a7145a <=( a7144a  and  a7141a );
 a7146a <=( a7145a  and  a7138a );
 a7150a <=( A199  and  A167 );
 a7151a <=( A168  and  a7150a );
 a7155a <=( A232  and  (not A203) );
 a7156a <=( (not A202)  and  a7155a );
 a7157a <=( a7156a  and  a7151a );
 a7161a <=( A236  and  A234 );
 a7162a <=( (not A233)  and  a7161a );
 a7165a <=( (not A299)  and  A298 );
 a7168a <=( A302  and  A300 );
 a7169a <=( a7168a  and  a7165a );
 a7170a <=( a7169a  and  a7162a );
 a7174a <=( A199  and  A167 );
 a7175a <=( A168  and  a7174a );
 a7179a <=( A232  and  (not A203) );
 a7180a <=( (not A202)  and  a7179a );
 a7181a <=( a7180a  and  a7175a );
 a7185a <=( A236  and  A234 );
 a7186a <=( (not A233)  and  a7185a );
 a7189a <=( (not A266)  and  A265 );
 a7192a <=( A268  and  A267 );
 a7193a <=( a7192a  and  a7189a );
 a7194a <=( a7193a  and  a7186a );
 a7198a <=( A199  and  A167 );
 a7199a <=( A168  and  a7198a );
 a7203a <=( A232  and  (not A203) );
 a7204a <=( (not A202)  and  a7203a );
 a7205a <=( a7204a  and  a7199a );
 a7209a <=( A236  and  A234 );
 a7210a <=( (not A233)  and  a7209a );
 a7213a <=( (not A266)  and  A265 );
 a7216a <=( A269  and  A267 );
 a7217a <=( a7216a  and  a7213a );
 a7218a <=( a7217a  and  a7210a );
 a7222a <=( A167  and  A169 );
 a7223a <=( (not A170)  and  a7222a );
 a7227a <=( (not A202)  and  A199 );
 a7228a <=( A166  and  a7227a );
 a7229a <=( a7228a  and  a7223a );
 a7233a <=( A233  and  (not A232) );
 a7234a <=( (not A203)  and  a7233a );
 a7237a <=( (not A299)  and  A298 );
 a7240a <=( A301  and  A300 );
 a7241a <=( a7240a  and  a7237a );
 a7242a <=( a7241a  and  a7234a );
 a7246a <=( A167  and  A169 );
 a7247a <=( (not A170)  and  a7246a );
 a7251a <=( (not A202)  and  A199 );
 a7252a <=( A166  and  a7251a );
 a7253a <=( a7252a  and  a7247a );
 a7257a <=( A233  and  (not A232) );
 a7258a <=( (not A203)  and  a7257a );
 a7261a <=( (not A299)  and  A298 );
 a7264a <=( A302  and  A300 );
 a7265a <=( a7264a  and  a7261a );
 a7266a <=( a7265a  and  a7258a );
 a7270a <=( A167  and  A169 );
 a7271a <=( (not A170)  and  a7270a );
 a7275a <=( (not A202)  and  A199 );
 a7276a <=( A166  and  a7275a );
 a7277a <=( a7276a  and  a7271a );
 a7281a <=( A233  and  (not A232) );
 a7282a <=( (not A203)  and  a7281a );
 a7285a <=( (not A266)  and  A265 );
 a7288a <=( A268  and  A267 );
 a7289a <=( a7288a  and  a7285a );
 a7290a <=( a7289a  and  a7282a );
 a7294a <=( A167  and  A169 );
 a7295a <=( (not A170)  and  a7294a );
 a7299a <=( (not A202)  and  A199 );
 a7300a <=( A166  and  a7299a );
 a7301a <=( a7300a  and  a7295a );
 a7305a <=( A233  and  (not A232) );
 a7306a <=( (not A203)  and  a7305a );
 a7309a <=( (not A266)  and  A265 );
 a7312a <=( A269  and  A267 );
 a7313a <=( a7312a  and  a7309a );
 a7314a <=( a7313a  and  a7306a );
 a7318a <=( A167  and  A169 );
 a7319a <=( (not A170)  and  a7318a );
 a7323a <=( (not A202)  and  A199 );
 a7324a <=( A166  and  a7323a );
 a7325a <=( a7324a  and  a7319a );
 a7329a <=( (not A233)  and  A232 );
 a7330a <=( (not A203)  and  a7329a );
 a7333a <=( A235  and  A234 );
 a7336a <=( A299  and  (not A298) );
 a7337a <=( a7336a  and  a7333a );
 a7338a <=( a7337a  and  a7330a );
 a7342a <=( A167  and  A169 );
 a7343a <=( (not A170)  and  a7342a );
 a7347a <=( (not A202)  and  A199 );
 a7348a <=( A166  and  a7347a );
 a7349a <=( a7348a  and  a7343a );
 a7353a <=( (not A233)  and  A232 );
 a7354a <=( (not A203)  and  a7353a );
 a7357a <=( A235  and  A234 );
 a7360a <=( A266  and  (not A265) );
 a7361a <=( a7360a  and  a7357a );
 a7362a <=( a7361a  and  a7354a );
 a7366a <=( A167  and  A169 );
 a7367a <=( (not A170)  and  a7366a );
 a7371a <=( (not A202)  and  A199 );
 a7372a <=( A166  and  a7371a );
 a7373a <=( a7372a  and  a7367a );
 a7377a <=( (not A233)  and  A232 );
 a7378a <=( (not A203)  and  a7377a );
 a7381a <=( A236  and  A234 );
 a7384a <=( A299  and  (not A298) );
 a7385a <=( a7384a  and  a7381a );
 a7386a <=( a7385a  and  a7378a );
 a7390a <=( A167  and  A169 );
 a7391a <=( (not A170)  and  a7390a );
 a7395a <=( (not A202)  and  A199 );
 a7396a <=( A166  and  a7395a );
 a7397a <=( a7396a  and  a7391a );
 a7401a <=( (not A233)  and  A232 );
 a7402a <=( (not A203)  and  a7401a );
 a7405a <=( A236  and  A234 );
 a7408a <=( A266  and  (not A265) );
 a7409a <=( a7408a  and  a7405a );
 a7410a <=( a7409a  and  a7402a );
 a7414a <=( (not A167)  and  A169 );
 a7415a <=( (not A170)  and  a7414a );
 a7419a <=( (not A202)  and  A199 );
 a7420a <=( (not A166)  and  a7419a );
 a7421a <=( a7420a  and  a7415a );
 a7425a <=( A233  and  (not A232) );
 a7426a <=( (not A203)  and  a7425a );
 a7429a <=( (not A299)  and  A298 );
 a7432a <=( A301  and  A300 );
 a7433a <=( a7432a  and  a7429a );
 a7434a <=( a7433a  and  a7426a );
 a7438a <=( (not A167)  and  A169 );
 a7439a <=( (not A170)  and  a7438a );
 a7443a <=( (not A202)  and  A199 );
 a7444a <=( (not A166)  and  a7443a );
 a7445a <=( a7444a  and  a7439a );
 a7449a <=( A233  and  (not A232) );
 a7450a <=( (not A203)  and  a7449a );
 a7453a <=( (not A299)  and  A298 );
 a7456a <=( A302  and  A300 );
 a7457a <=( a7456a  and  a7453a );
 a7458a <=( a7457a  and  a7450a );
 a7462a <=( (not A167)  and  A169 );
 a7463a <=( (not A170)  and  a7462a );
 a7467a <=( (not A202)  and  A199 );
 a7468a <=( (not A166)  and  a7467a );
 a7469a <=( a7468a  and  a7463a );
 a7473a <=( A233  and  (not A232) );
 a7474a <=( (not A203)  and  a7473a );
 a7477a <=( (not A266)  and  A265 );
 a7480a <=( A268  and  A267 );
 a7481a <=( a7480a  and  a7477a );
 a7482a <=( a7481a  and  a7474a );
 a7486a <=( (not A167)  and  A169 );
 a7487a <=( (not A170)  and  a7486a );
 a7491a <=( (not A202)  and  A199 );
 a7492a <=( (not A166)  and  a7491a );
 a7493a <=( a7492a  and  a7487a );
 a7497a <=( A233  and  (not A232) );
 a7498a <=( (not A203)  and  a7497a );
 a7501a <=( (not A266)  and  A265 );
 a7504a <=( A269  and  A267 );
 a7505a <=( a7504a  and  a7501a );
 a7506a <=( a7505a  and  a7498a );
 a7510a <=( (not A167)  and  A169 );
 a7511a <=( (not A170)  and  a7510a );
 a7515a <=( (not A202)  and  A199 );
 a7516a <=( (not A166)  and  a7515a );
 a7517a <=( a7516a  and  a7511a );
 a7521a <=( (not A233)  and  A232 );
 a7522a <=( (not A203)  and  a7521a );
 a7525a <=( A235  and  A234 );
 a7528a <=( A299  and  (not A298) );
 a7529a <=( a7528a  and  a7525a );
 a7530a <=( a7529a  and  a7522a );
 a7534a <=( (not A167)  and  A169 );
 a7535a <=( (not A170)  and  a7534a );
 a7539a <=( (not A202)  and  A199 );
 a7540a <=( (not A166)  and  a7539a );
 a7541a <=( a7540a  and  a7535a );
 a7545a <=( (not A233)  and  A232 );
 a7546a <=( (not A203)  and  a7545a );
 a7549a <=( A235  and  A234 );
 a7552a <=( A266  and  (not A265) );
 a7553a <=( a7552a  and  a7549a );
 a7554a <=( a7553a  and  a7546a );
 a7558a <=( (not A167)  and  A169 );
 a7559a <=( (not A170)  and  a7558a );
 a7563a <=( (not A202)  and  A199 );
 a7564a <=( (not A166)  and  a7563a );
 a7565a <=( a7564a  and  a7559a );
 a7569a <=( (not A233)  and  A232 );
 a7570a <=( (not A203)  and  a7569a );
 a7573a <=( A236  and  A234 );
 a7576a <=( A299  and  (not A298) );
 a7577a <=( a7576a  and  a7573a );
 a7578a <=( a7577a  and  a7570a );
 a7582a <=( (not A167)  and  A169 );
 a7583a <=( (not A170)  and  a7582a );
 a7587a <=( (not A202)  and  A199 );
 a7588a <=( (not A166)  and  a7587a );
 a7589a <=( a7588a  and  a7583a );
 a7593a <=( (not A233)  and  A232 );
 a7594a <=( (not A203)  and  a7593a );
 a7597a <=( A236  and  A234 );
 a7600a <=( A266  and  (not A265) );
 a7601a <=( a7600a  and  a7597a );
 a7602a <=( a7601a  and  a7594a );
 a7606a <=( A167  and  (not A169) );
 a7607a <=( A170  and  a7606a );
 a7611a <=( (not A202)  and  A199 );
 a7612a <=( (not A166)  and  a7611a );
 a7613a <=( a7612a  and  a7607a );
 a7617a <=( A233  and  (not A232) );
 a7618a <=( (not A203)  and  a7617a );
 a7621a <=( (not A299)  and  A298 );
 a7624a <=( A301  and  A300 );
 a7625a <=( a7624a  and  a7621a );
 a7626a <=( a7625a  and  a7618a );
 a7630a <=( A167  and  (not A169) );
 a7631a <=( A170  and  a7630a );
 a7635a <=( (not A202)  and  A199 );
 a7636a <=( (not A166)  and  a7635a );
 a7637a <=( a7636a  and  a7631a );
 a7641a <=( A233  and  (not A232) );
 a7642a <=( (not A203)  and  a7641a );
 a7645a <=( (not A299)  and  A298 );
 a7648a <=( A302  and  A300 );
 a7649a <=( a7648a  and  a7645a );
 a7650a <=( a7649a  and  a7642a );
 a7654a <=( A167  and  (not A169) );
 a7655a <=( A170  and  a7654a );
 a7659a <=( (not A202)  and  A199 );
 a7660a <=( (not A166)  and  a7659a );
 a7661a <=( a7660a  and  a7655a );
 a7665a <=( A233  and  (not A232) );
 a7666a <=( (not A203)  and  a7665a );
 a7669a <=( (not A266)  and  A265 );
 a7672a <=( A268  and  A267 );
 a7673a <=( a7672a  and  a7669a );
 a7674a <=( a7673a  and  a7666a );
 a7678a <=( A167  and  (not A169) );
 a7679a <=( A170  and  a7678a );
 a7683a <=( (not A202)  and  A199 );
 a7684a <=( (not A166)  and  a7683a );
 a7685a <=( a7684a  and  a7679a );
 a7689a <=( A233  and  (not A232) );
 a7690a <=( (not A203)  and  a7689a );
 a7693a <=( (not A266)  and  A265 );
 a7696a <=( A269  and  A267 );
 a7697a <=( a7696a  and  a7693a );
 a7698a <=( a7697a  and  a7690a );
 a7702a <=( A167  and  (not A169) );
 a7703a <=( A170  and  a7702a );
 a7707a <=( (not A202)  and  A199 );
 a7708a <=( (not A166)  and  a7707a );
 a7709a <=( a7708a  and  a7703a );
 a7713a <=( (not A233)  and  A232 );
 a7714a <=( (not A203)  and  a7713a );
 a7717a <=( A235  and  A234 );
 a7720a <=( A299  and  (not A298) );
 a7721a <=( a7720a  and  a7717a );
 a7722a <=( a7721a  and  a7714a );
 a7726a <=( A167  and  (not A169) );
 a7727a <=( A170  and  a7726a );
 a7731a <=( (not A202)  and  A199 );
 a7732a <=( (not A166)  and  a7731a );
 a7733a <=( a7732a  and  a7727a );
 a7737a <=( (not A233)  and  A232 );
 a7738a <=( (not A203)  and  a7737a );
 a7741a <=( A235  and  A234 );
 a7744a <=( A266  and  (not A265) );
 a7745a <=( a7744a  and  a7741a );
 a7746a <=( a7745a  and  a7738a );
 a7750a <=( A167  and  (not A169) );
 a7751a <=( A170  and  a7750a );
 a7755a <=( (not A202)  and  A199 );
 a7756a <=( (not A166)  and  a7755a );
 a7757a <=( a7756a  and  a7751a );
 a7761a <=( (not A233)  and  A232 );
 a7762a <=( (not A203)  and  a7761a );
 a7765a <=( A236  and  A234 );
 a7768a <=( A299  and  (not A298) );
 a7769a <=( a7768a  and  a7765a );
 a7770a <=( a7769a  and  a7762a );
 a7774a <=( A167  and  (not A169) );
 a7775a <=( A170  and  a7774a );
 a7779a <=( (not A202)  and  A199 );
 a7780a <=( (not A166)  and  a7779a );
 a7781a <=( a7780a  and  a7775a );
 a7785a <=( (not A233)  and  A232 );
 a7786a <=( (not A203)  and  a7785a );
 a7789a <=( A236  and  A234 );
 a7792a <=( A266  and  (not A265) );
 a7793a <=( a7792a  and  a7789a );
 a7794a <=( a7793a  and  a7786a );
 a7798a <=( (not A167)  and  (not A169) );
 a7799a <=( A170  and  a7798a );
 a7803a <=( (not A202)  and  A199 );
 a7804a <=( A166  and  a7803a );
 a7805a <=( a7804a  and  a7799a );
 a7809a <=( A233  and  (not A232) );
 a7810a <=( (not A203)  and  a7809a );
 a7813a <=( (not A299)  and  A298 );
 a7816a <=( A301  and  A300 );
 a7817a <=( a7816a  and  a7813a );
 a7818a <=( a7817a  and  a7810a );
 a7822a <=( (not A167)  and  (not A169) );
 a7823a <=( A170  and  a7822a );
 a7827a <=( (not A202)  and  A199 );
 a7828a <=( A166  and  a7827a );
 a7829a <=( a7828a  and  a7823a );
 a7833a <=( A233  and  (not A232) );
 a7834a <=( (not A203)  and  a7833a );
 a7837a <=( (not A299)  and  A298 );
 a7840a <=( A302  and  A300 );
 a7841a <=( a7840a  and  a7837a );
 a7842a <=( a7841a  and  a7834a );
 a7846a <=( (not A167)  and  (not A169) );
 a7847a <=( A170  and  a7846a );
 a7851a <=( (not A202)  and  A199 );
 a7852a <=( A166  and  a7851a );
 a7853a <=( a7852a  and  a7847a );
 a7857a <=( A233  and  (not A232) );
 a7858a <=( (not A203)  and  a7857a );
 a7861a <=( (not A266)  and  A265 );
 a7864a <=( A268  and  A267 );
 a7865a <=( a7864a  and  a7861a );
 a7866a <=( a7865a  and  a7858a );
 a7870a <=( (not A167)  and  (not A169) );
 a7871a <=( A170  and  a7870a );
 a7875a <=( (not A202)  and  A199 );
 a7876a <=( A166  and  a7875a );
 a7877a <=( a7876a  and  a7871a );
 a7881a <=( A233  and  (not A232) );
 a7882a <=( (not A203)  and  a7881a );
 a7885a <=( (not A266)  and  A265 );
 a7888a <=( A269  and  A267 );
 a7889a <=( a7888a  and  a7885a );
 a7890a <=( a7889a  and  a7882a );
 a7894a <=( (not A167)  and  (not A169) );
 a7895a <=( A170  and  a7894a );
 a7899a <=( (not A202)  and  A199 );
 a7900a <=( A166  and  a7899a );
 a7901a <=( a7900a  and  a7895a );
 a7905a <=( (not A233)  and  A232 );
 a7906a <=( (not A203)  and  a7905a );
 a7909a <=( A235  and  A234 );
 a7912a <=( A299  and  (not A298) );
 a7913a <=( a7912a  and  a7909a );
 a7914a <=( a7913a  and  a7906a );
 a7918a <=( (not A167)  and  (not A169) );
 a7919a <=( A170  and  a7918a );
 a7923a <=( (not A202)  and  A199 );
 a7924a <=( A166  and  a7923a );
 a7925a <=( a7924a  and  a7919a );
 a7929a <=( (not A233)  and  A232 );
 a7930a <=( (not A203)  and  a7929a );
 a7933a <=( A235  and  A234 );
 a7936a <=( A266  and  (not A265) );
 a7937a <=( a7936a  and  a7933a );
 a7938a <=( a7937a  and  a7930a );
 a7942a <=( (not A167)  and  (not A169) );
 a7943a <=( A170  and  a7942a );
 a7947a <=( (not A202)  and  A199 );
 a7948a <=( A166  and  a7947a );
 a7949a <=( a7948a  and  a7943a );
 a7953a <=( (not A233)  and  A232 );
 a7954a <=( (not A203)  and  a7953a );
 a7957a <=( A236  and  A234 );
 a7960a <=( A299  and  (not A298) );
 a7961a <=( a7960a  and  a7957a );
 a7962a <=( a7961a  and  a7954a );
 a7966a <=( (not A167)  and  (not A169) );
 a7967a <=( A170  and  a7966a );
 a7971a <=( (not A202)  and  A199 );
 a7972a <=( A166  and  a7971a );
 a7973a <=( a7972a  and  a7967a );
 a7977a <=( (not A233)  and  A232 );
 a7978a <=( (not A203)  and  a7977a );
 a7981a <=( A236  and  A234 );
 a7984a <=( A266  and  (not A265) );
 a7985a <=( a7984a  and  a7981a );
 a7986a <=( a7985a  and  a7978a );
 a7990a <=( A167  and  A169 );
 a7991a <=( (not A170)  and  a7990a );
 a7994a <=( A199  and  A166 );
 a7997a <=( A232  and  (not A201) );
 a7998a <=( a7997a  and  a7994a );
 a7999a <=( a7998a  and  a7991a );
 a8003a <=( A235  and  A234 );
 a8004a <=( (not A233)  and  a8003a );
 a8007a <=( (not A299)  and  A298 );
 a8010a <=( A301  and  A300 );
 a8011a <=( a8010a  and  a8007a );
 a8012a <=( a8011a  and  a8004a );
 a8016a <=( A167  and  A169 );
 a8017a <=( (not A170)  and  a8016a );
 a8020a <=( A199  and  A166 );
 a8023a <=( A232  and  (not A201) );
 a8024a <=( a8023a  and  a8020a );
 a8025a <=( a8024a  and  a8017a );
 a8029a <=( A235  and  A234 );
 a8030a <=( (not A233)  and  a8029a );
 a8033a <=( (not A299)  and  A298 );
 a8036a <=( A302  and  A300 );
 a8037a <=( a8036a  and  a8033a );
 a8038a <=( a8037a  and  a8030a );
 a8042a <=( A167  and  A169 );
 a8043a <=( (not A170)  and  a8042a );
 a8046a <=( A199  and  A166 );
 a8049a <=( A232  and  (not A201) );
 a8050a <=( a8049a  and  a8046a );
 a8051a <=( a8050a  and  a8043a );
 a8055a <=( A235  and  A234 );
 a8056a <=( (not A233)  and  a8055a );
 a8059a <=( (not A266)  and  A265 );
 a8062a <=( A268  and  A267 );
 a8063a <=( a8062a  and  a8059a );
 a8064a <=( a8063a  and  a8056a );
 a8068a <=( A167  and  A169 );
 a8069a <=( (not A170)  and  a8068a );
 a8072a <=( A199  and  A166 );
 a8075a <=( A232  and  (not A201) );
 a8076a <=( a8075a  and  a8072a );
 a8077a <=( a8076a  and  a8069a );
 a8081a <=( A235  and  A234 );
 a8082a <=( (not A233)  and  a8081a );
 a8085a <=( (not A266)  and  A265 );
 a8088a <=( A269  and  A267 );
 a8089a <=( a8088a  and  a8085a );
 a8090a <=( a8089a  and  a8082a );
 a8094a <=( A167  and  A169 );
 a8095a <=( (not A170)  and  a8094a );
 a8098a <=( A199  and  A166 );
 a8101a <=( A232  and  (not A201) );
 a8102a <=( a8101a  and  a8098a );
 a8103a <=( a8102a  and  a8095a );
 a8107a <=( A236  and  A234 );
 a8108a <=( (not A233)  and  a8107a );
 a8111a <=( (not A299)  and  A298 );
 a8114a <=( A301  and  A300 );
 a8115a <=( a8114a  and  a8111a );
 a8116a <=( a8115a  and  a8108a );
 a8120a <=( A167  and  A169 );
 a8121a <=( (not A170)  and  a8120a );
 a8124a <=( A199  and  A166 );
 a8127a <=( A232  and  (not A201) );
 a8128a <=( a8127a  and  a8124a );
 a8129a <=( a8128a  and  a8121a );
 a8133a <=( A236  and  A234 );
 a8134a <=( (not A233)  and  a8133a );
 a8137a <=( (not A299)  and  A298 );
 a8140a <=( A302  and  A300 );
 a8141a <=( a8140a  and  a8137a );
 a8142a <=( a8141a  and  a8134a );
 a8146a <=( A167  and  A169 );
 a8147a <=( (not A170)  and  a8146a );
 a8150a <=( A199  and  A166 );
 a8153a <=( A232  and  (not A201) );
 a8154a <=( a8153a  and  a8150a );
 a8155a <=( a8154a  and  a8147a );
 a8159a <=( A236  and  A234 );
 a8160a <=( (not A233)  and  a8159a );
 a8163a <=( (not A266)  and  A265 );
 a8166a <=( A268  and  A267 );
 a8167a <=( a8166a  and  a8163a );
 a8168a <=( a8167a  and  a8160a );
 a8172a <=( A167  and  A169 );
 a8173a <=( (not A170)  and  a8172a );
 a8176a <=( A199  and  A166 );
 a8179a <=( A232  and  (not A201) );
 a8180a <=( a8179a  and  a8176a );
 a8181a <=( a8180a  and  a8173a );
 a8185a <=( A236  and  A234 );
 a8186a <=( (not A233)  and  a8185a );
 a8189a <=( (not A266)  and  A265 );
 a8192a <=( A269  and  A267 );
 a8193a <=( a8192a  and  a8189a );
 a8194a <=( a8193a  and  a8186a );
 a8198a <=( A167  and  A169 );
 a8199a <=( (not A170)  and  a8198a );
 a8202a <=( A199  and  A166 );
 a8205a <=( A232  and  A200 );
 a8206a <=( a8205a  and  a8202a );
 a8207a <=( a8206a  and  a8199a );
 a8211a <=( A235  and  A234 );
 a8212a <=( (not A233)  and  a8211a );
 a8215a <=( (not A299)  and  A298 );
 a8218a <=( A301  and  A300 );
 a8219a <=( a8218a  and  a8215a );
 a8220a <=( a8219a  and  a8212a );
 a8224a <=( A167  and  A169 );
 a8225a <=( (not A170)  and  a8224a );
 a8228a <=( A199  and  A166 );
 a8231a <=( A232  and  A200 );
 a8232a <=( a8231a  and  a8228a );
 a8233a <=( a8232a  and  a8225a );
 a8237a <=( A235  and  A234 );
 a8238a <=( (not A233)  and  a8237a );
 a8241a <=( (not A299)  and  A298 );
 a8244a <=( A302  and  A300 );
 a8245a <=( a8244a  and  a8241a );
 a8246a <=( a8245a  and  a8238a );
 a8250a <=( A167  and  A169 );
 a8251a <=( (not A170)  and  a8250a );
 a8254a <=( A199  and  A166 );
 a8257a <=( A232  and  A200 );
 a8258a <=( a8257a  and  a8254a );
 a8259a <=( a8258a  and  a8251a );
 a8263a <=( A235  and  A234 );
 a8264a <=( (not A233)  and  a8263a );
 a8267a <=( (not A266)  and  A265 );
 a8270a <=( A268  and  A267 );
 a8271a <=( a8270a  and  a8267a );
 a8272a <=( a8271a  and  a8264a );
 a8276a <=( A167  and  A169 );
 a8277a <=( (not A170)  and  a8276a );
 a8280a <=( A199  and  A166 );
 a8283a <=( A232  and  A200 );
 a8284a <=( a8283a  and  a8280a );
 a8285a <=( a8284a  and  a8277a );
 a8289a <=( A235  and  A234 );
 a8290a <=( (not A233)  and  a8289a );
 a8293a <=( (not A266)  and  A265 );
 a8296a <=( A269  and  A267 );
 a8297a <=( a8296a  and  a8293a );
 a8298a <=( a8297a  and  a8290a );
 a8302a <=( A167  and  A169 );
 a8303a <=( (not A170)  and  a8302a );
 a8306a <=( A199  and  A166 );
 a8309a <=( A232  and  A200 );
 a8310a <=( a8309a  and  a8306a );
 a8311a <=( a8310a  and  a8303a );
 a8315a <=( A236  and  A234 );
 a8316a <=( (not A233)  and  a8315a );
 a8319a <=( (not A299)  and  A298 );
 a8322a <=( A301  and  A300 );
 a8323a <=( a8322a  and  a8319a );
 a8324a <=( a8323a  and  a8316a );
 a8328a <=( A167  and  A169 );
 a8329a <=( (not A170)  and  a8328a );
 a8332a <=( A199  and  A166 );
 a8335a <=( A232  and  A200 );
 a8336a <=( a8335a  and  a8332a );
 a8337a <=( a8336a  and  a8329a );
 a8341a <=( A236  and  A234 );
 a8342a <=( (not A233)  and  a8341a );
 a8345a <=( (not A299)  and  A298 );
 a8348a <=( A302  and  A300 );
 a8349a <=( a8348a  and  a8345a );
 a8350a <=( a8349a  and  a8342a );
 a8354a <=( A167  and  A169 );
 a8355a <=( (not A170)  and  a8354a );
 a8358a <=( A199  and  A166 );
 a8361a <=( A232  and  A200 );
 a8362a <=( a8361a  and  a8358a );
 a8363a <=( a8362a  and  a8355a );
 a8367a <=( A236  and  A234 );
 a8368a <=( (not A233)  and  a8367a );
 a8371a <=( (not A266)  and  A265 );
 a8374a <=( A268  and  A267 );
 a8375a <=( a8374a  and  a8371a );
 a8376a <=( a8375a  and  a8368a );
 a8380a <=( A167  and  A169 );
 a8381a <=( (not A170)  and  a8380a );
 a8384a <=( A199  and  A166 );
 a8387a <=( A232  and  A200 );
 a8388a <=( a8387a  and  a8384a );
 a8389a <=( a8388a  and  a8381a );
 a8393a <=( A236  and  A234 );
 a8394a <=( (not A233)  and  a8393a );
 a8397a <=( (not A266)  and  A265 );
 a8400a <=( A269  and  A267 );
 a8401a <=( a8400a  and  a8397a );
 a8402a <=( a8401a  and  a8394a );
 a8406a <=( A167  and  A169 );
 a8407a <=( (not A170)  and  a8406a );
 a8410a <=( (not A199)  and  A166 );
 a8413a <=( A232  and  (not A200) );
 a8414a <=( a8413a  and  a8410a );
 a8415a <=( a8414a  and  a8407a );
 a8419a <=( A235  and  A234 );
 a8420a <=( (not A233)  and  a8419a );
 a8423a <=( (not A299)  and  A298 );
 a8426a <=( A301  and  A300 );
 a8427a <=( a8426a  and  a8423a );
 a8428a <=( a8427a  and  a8420a );
 a8432a <=( A167  and  A169 );
 a8433a <=( (not A170)  and  a8432a );
 a8436a <=( (not A199)  and  A166 );
 a8439a <=( A232  and  (not A200) );
 a8440a <=( a8439a  and  a8436a );
 a8441a <=( a8440a  and  a8433a );
 a8445a <=( A235  and  A234 );
 a8446a <=( (not A233)  and  a8445a );
 a8449a <=( (not A299)  and  A298 );
 a8452a <=( A302  and  A300 );
 a8453a <=( a8452a  and  a8449a );
 a8454a <=( a8453a  and  a8446a );
 a8458a <=( A167  and  A169 );
 a8459a <=( (not A170)  and  a8458a );
 a8462a <=( (not A199)  and  A166 );
 a8465a <=( A232  and  (not A200) );
 a8466a <=( a8465a  and  a8462a );
 a8467a <=( a8466a  and  a8459a );
 a8471a <=( A235  and  A234 );
 a8472a <=( (not A233)  and  a8471a );
 a8475a <=( (not A266)  and  A265 );
 a8478a <=( A268  and  A267 );
 a8479a <=( a8478a  and  a8475a );
 a8480a <=( a8479a  and  a8472a );
 a8484a <=( A167  and  A169 );
 a8485a <=( (not A170)  and  a8484a );
 a8488a <=( (not A199)  and  A166 );
 a8491a <=( A232  and  (not A200) );
 a8492a <=( a8491a  and  a8488a );
 a8493a <=( a8492a  and  a8485a );
 a8497a <=( A235  and  A234 );
 a8498a <=( (not A233)  and  a8497a );
 a8501a <=( (not A266)  and  A265 );
 a8504a <=( A269  and  A267 );
 a8505a <=( a8504a  and  a8501a );
 a8506a <=( a8505a  and  a8498a );
 a8510a <=( A167  and  A169 );
 a8511a <=( (not A170)  and  a8510a );
 a8514a <=( (not A199)  and  A166 );
 a8517a <=( A232  and  (not A200) );
 a8518a <=( a8517a  and  a8514a );
 a8519a <=( a8518a  and  a8511a );
 a8523a <=( A236  and  A234 );
 a8524a <=( (not A233)  and  a8523a );
 a8527a <=( (not A299)  and  A298 );
 a8530a <=( A301  and  A300 );
 a8531a <=( a8530a  and  a8527a );
 a8532a <=( a8531a  and  a8524a );
 a8536a <=( A167  and  A169 );
 a8537a <=( (not A170)  and  a8536a );
 a8540a <=( (not A199)  and  A166 );
 a8543a <=( A232  and  (not A200) );
 a8544a <=( a8543a  and  a8540a );
 a8545a <=( a8544a  and  a8537a );
 a8549a <=( A236  and  A234 );
 a8550a <=( (not A233)  and  a8549a );
 a8553a <=( (not A299)  and  A298 );
 a8556a <=( A302  and  A300 );
 a8557a <=( a8556a  and  a8553a );
 a8558a <=( a8557a  and  a8550a );
 a8562a <=( A167  and  A169 );
 a8563a <=( (not A170)  and  a8562a );
 a8566a <=( (not A199)  and  A166 );
 a8569a <=( A232  and  (not A200) );
 a8570a <=( a8569a  and  a8566a );
 a8571a <=( a8570a  and  a8563a );
 a8575a <=( A236  and  A234 );
 a8576a <=( (not A233)  and  a8575a );
 a8579a <=( (not A266)  and  A265 );
 a8582a <=( A268  and  A267 );
 a8583a <=( a8582a  and  a8579a );
 a8584a <=( a8583a  and  a8576a );
 a8588a <=( A167  and  A169 );
 a8589a <=( (not A170)  and  a8588a );
 a8592a <=( (not A199)  and  A166 );
 a8595a <=( A232  and  (not A200) );
 a8596a <=( a8595a  and  a8592a );
 a8597a <=( a8596a  and  a8589a );
 a8601a <=( A236  and  A234 );
 a8602a <=( (not A233)  and  a8601a );
 a8605a <=( (not A266)  and  A265 );
 a8608a <=( A269  and  A267 );
 a8609a <=( a8608a  and  a8605a );
 a8610a <=( a8609a  and  a8602a );
 a8614a <=( (not A167)  and  A169 );
 a8615a <=( (not A170)  and  a8614a );
 a8618a <=( A199  and  (not A166) );
 a8621a <=( A232  and  (not A201) );
 a8622a <=( a8621a  and  a8618a );
 a8623a <=( a8622a  and  a8615a );
 a8627a <=( A235  and  A234 );
 a8628a <=( (not A233)  and  a8627a );
 a8631a <=( (not A299)  and  A298 );
 a8634a <=( A301  and  A300 );
 a8635a <=( a8634a  and  a8631a );
 a8636a <=( a8635a  and  a8628a );
 a8640a <=( (not A167)  and  A169 );
 a8641a <=( (not A170)  and  a8640a );
 a8644a <=( A199  and  (not A166) );
 a8647a <=( A232  and  (not A201) );
 a8648a <=( a8647a  and  a8644a );
 a8649a <=( a8648a  and  a8641a );
 a8653a <=( A235  and  A234 );
 a8654a <=( (not A233)  and  a8653a );
 a8657a <=( (not A299)  and  A298 );
 a8660a <=( A302  and  A300 );
 a8661a <=( a8660a  and  a8657a );
 a8662a <=( a8661a  and  a8654a );
 a8666a <=( (not A167)  and  A169 );
 a8667a <=( (not A170)  and  a8666a );
 a8670a <=( A199  and  (not A166) );
 a8673a <=( A232  and  (not A201) );
 a8674a <=( a8673a  and  a8670a );
 a8675a <=( a8674a  and  a8667a );
 a8679a <=( A235  and  A234 );
 a8680a <=( (not A233)  and  a8679a );
 a8683a <=( (not A266)  and  A265 );
 a8686a <=( A268  and  A267 );
 a8687a <=( a8686a  and  a8683a );
 a8688a <=( a8687a  and  a8680a );
 a8692a <=( (not A167)  and  A169 );
 a8693a <=( (not A170)  and  a8692a );
 a8696a <=( A199  and  (not A166) );
 a8699a <=( A232  and  (not A201) );
 a8700a <=( a8699a  and  a8696a );
 a8701a <=( a8700a  and  a8693a );
 a8705a <=( A235  and  A234 );
 a8706a <=( (not A233)  and  a8705a );
 a8709a <=( (not A266)  and  A265 );
 a8712a <=( A269  and  A267 );
 a8713a <=( a8712a  and  a8709a );
 a8714a <=( a8713a  and  a8706a );
 a8718a <=( (not A167)  and  A169 );
 a8719a <=( (not A170)  and  a8718a );
 a8722a <=( A199  and  (not A166) );
 a8725a <=( A232  and  (not A201) );
 a8726a <=( a8725a  and  a8722a );
 a8727a <=( a8726a  and  a8719a );
 a8731a <=( A236  and  A234 );
 a8732a <=( (not A233)  and  a8731a );
 a8735a <=( (not A299)  and  A298 );
 a8738a <=( A301  and  A300 );
 a8739a <=( a8738a  and  a8735a );
 a8740a <=( a8739a  and  a8732a );
 a8744a <=( (not A167)  and  A169 );
 a8745a <=( (not A170)  and  a8744a );
 a8748a <=( A199  and  (not A166) );
 a8751a <=( A232  and  (not A201) );
 a8752a <=( a8751a  and  a8748a );
 a8753a <=( a8752a  and  a8745a );
 a8757a <=( A236  and  A234 );
 a8758a <=( (not A233)  and  a8757a );
 a8761a <=( (not A299)  and  A298 );
 a8764a <=( A302  and  A300 );
 a8765a <=( a8764a  and  a8761a );
 a8766a <=( a8765a  and  a8758a );
 a8770a <=( (not A167)  and  A169 );
 a8771a <=( (not A170)  and  a8770a );
 a8774a <=( A199  and  (not A166) );
 a8777a <=( A232  and  (not A201) );
 a8778a <=( a8777a  and  a8774a );
 a8779a <=( a8778a  and  a8771a );
 a8783a <=( A236  and  A234 );
 a8784a <=( (not A233)  and  a8783a );
 a8787a <=( (not A266)  and  A265 );
 a8790a <=( A268  and  A267 );
 a8791a <=( a8790a  and  a8787a );
 a8792a <=( a8791a  and  a8784a );
 a8796a <=( (not A167)  and  A169 );
 a8797a <=( (not A170)  and  a8796a );
 a8800a <=( A199  and  (not A166) );
 a8803a <=( A232  and  (not A201) );
 a8804a <=( a8803a  and  a8800a );
 a8805a <=( a8804a  and  a8797a );
 a8809a <=( A236  and  A234 );
 a8810a <=( (not A233)  and  a8809a );
 a8813a <=( (not A266)  and  A265 );
 a8816a <=( A269  and  A267 );
 a8817a <=( a8816a  and  a8813a );
 a8818a <=( a8817a  and  a8810a );
 a8822a <=( (not A167)  and  A169 );
 a8823a <=( (not A170)  and  a8822a );
 a8826a <=( A199  and  (not A166) );
 a8829a <=( A232  and  A200 );
 a8830a <=( a8829a  and  a8826a );
 a8831a <=( a8830a  and  a8823a );
 a8835a <=( A235  and  A234 );
 a8836a <=( (not A233)  and  a8835a );
 a8839a <=( (not A299)  and  A298 );
 a8842a <=( A301  and  A300 );
 a8843a <=( a8842a  and  a8839a );
 a8844a <=( a8843a  and  a8836a );
 a8848a <=( (not A167)  and  A169 );
 a8849a <=( (not A170)  and  a8848a );
 a8852a <=( A199  and  (not A166) );
 a8855a <=( A232  and  A200 );
 a8856a <=( a8855a  and  a8852a );
 a8857a <=( a8856a  and  a8849a );
 a8861a <=( A235  and  A234 );
 a8862a <=( (not A233)  and  a8861a );
 a8865a <=( (not A299)  and  A298 );
 a8868a <=( A302  and  A300 );
 a8869a <=( a8868a  and  a8865a );
 a8870a <=( a8869a  and  a8862a );
 a8874a <=( (not A167)  and  A169 );
 a8875a <=( (not A170)  and  a8874a );
 a8878a <=( A199  and  (not A166) );
 a8881a <=( A232  and  A200 );
 a8882a <=( a8881a  and  a8878a );
 a8883a <=( a8882a  and  a8875a );
 a8887a <=( A235  and  A234 );
 a8888a <=( (not A233)  and  a8887a );
 a8891a <=( (not A266)  and  A265 );
 a8894a <=( A268  and  A267 );
 a8895a <=( a8894a  and  a8891a );
 a8896a <=( a8895a  and  a8888a );
 a8900a <=( (not A167)  and  A169 );
 a8901a <=( (not A170)  and  a8900a );
 a8904a <=( A199  and  (not A166) );
 a8907a <=( A232  and  A200 );
 a8908a <=( a8907a  and  a8904a );
 a8909a <=( a8908a  and  a8901a );
 a8913a <=( A235  and  A234 );
 a8914a <=( (not A233)  and  a8913a );
 a8917a <=( (not A266)  and  A265 );
 a8920a <=( A269  and  A267 );
 a8921a <=( a8920a  and  a8917a );
 a8922a <=( a8921a  and  a8914a );
 a8926a <=( (not A167)  and  A169 );
 a8927a <=( (not A170)  and  a8926a );
 a8930a <=( A199  and  (not A166) );
 a8933a <=( A232  and  A200 );
 a8934a <=( a8933a  and  a8930a );
 a8935a <=( a8934a  and  a8927a );
 a8939a <=( A236  and  A234 );
 a8940a <=( (not A233)  and  a8939a );
 a8943a <=( (not A299)  and  A298 );
 a8946a <=( A301  and  A300 );
 a8947a <=( a8946a  and  a8943a );
 a8948a <=( a8947a  and  a8940a );
 a8952a <=( (not A167)  and  A169 );
 a8953a <=( (not A170)  and  a8952a );
 a8956a <=( A199  and  (not A166) );
 a8959a <=( A232  and  A200 );
 a8960a <=( a8959a  and  a8956a );
 a8961a <=( a8960a  and  a8953a );
 a8965a <=( A236  and  A234 );
 a8966a <=( (not A233)  and  a8965a );
 a8969a <=( (not A299)  and  A298 );
 a8972a <=( A302  and  A300 );
 a8973a <=( a8972a  and  a8969a );
 a8974a <=( a8973a  and  a8966a );
 a8978a <=( (not A167)  and  A169 );
 a8979a <=( (not A170)  and  a8978a );
 a8982a <=( A199  and  (not A166) );
 a8985a <=( A232  and  A200 );
 a8986a <=( a8985a  and  a8982a );
 a8987a <=( a8986a  and  a8979a );
 a8991a <=( A236  and  A234 );
 a8992a <=( (not A233)  and  a8991a );
 a8995a <=( (not A266)  and  A265 );
 a8998a <=( A268  and  A267 );
 a8999a <=( a8998a  and  a8995a );
 a9000a <=( a8999a  and  a8992a );
 a9004a <=( (not A167)  and  A169 );
 a9005a <=( (not A170)  and  a9004a );
 a9008a <=( A199  and  (not A166) );
 a9011a <=( A232  and  A200 );
 a9012a <=( a9011a  and  a9008a );
 a9013a <=( a9012a  and  a9005a );
 a9017a <=( A236  and  A234 );
 a9018a <=( (not A233)  and  a9017a );
 a9021a <=( (not A266)  and  A265 );
 a9024a <=( A269  and  A267 );
 a9025a <=( a9024a  and  a9021a );
 a9026a <=( a9025a  and  a9018a );
 a9030a <=( (not A167)  and  A169 );
 a9031a <=( (not A170)  and  a9030a );
 a9034a <=( (not A199)  and  (not A166) );
 a9037a <=( A232  and  (not A200) );
 a9038a <=( a9037a  and  a9034a );
 a9039a <=( a9038a  and  a9031a );
 a9043a <=( A235  and  A234 );
 a9044a <=( (not A233)  and  a9043a );
 a9047a <=( (not A299)  and  A298 );
 a9050a <=( A301  and  A300 );
 a9051a <=( a9050a  and  a9047a );
 a9052a <=( a9051a  and  a9044a );
 a9056a <=( (not A167)  and  A169 );
 a9057a <=( (not A170)  and  a9056a );
 a9060a <=( (not A199)  and  (not A166) );
 a9063a <=( A232  and  (not A200) );
 a9064a <=( a9063a  and  a9060a );
 a9065a <=( a9064a  and  a9057a );
 a9069a <=( A235  and  A234 );
 a9070a <=( (not A233)  and  a9069a );
 a9073a <=( (not A299)  and  A298 );
 a9076a <=( A302  and  A300 );
 a9077a <=( a9076a  and  a9073a );
 a9078a <=( a9077a  and  a9070a );
 a9082a <=( (not A167)  and  A169 );
 a9083a <=( (not A170)  and  a9082a );
 a9086a <=( (not A199)  and  (not A166) );
 a9089a <=( A232  and  (not A200) );
 a9090a <=( a9089a  and  a9086a );
 a9091a <=( a9090a  and  a9083a );
 a9095a <=( A235  and  A234 );
 a9096a <=( (not A233)  and  a9095a );
 a9099a <=( (not A266)  and  A265 );
 a9102a <=( A268  and  A267 );
 a9103a <=( a9102a  and  a9099a );
 a9104a <=( a9103a  and  a9096a );
 a9108a <=( (not A167)  and  A169 );
 a9109a <=( (not A170)  and  a9108a );
 a9112a <=( (not A199)  and  (not A166) );
 a9115a <=( A232  and  (not A200) );
 a9116a <=( a9115a  and  a9112a );
 a9117a <=( a9116a  and  a9109a );
 a9121a <=( A235  and  A234 );
 a9122a <=( (not A233)  and  a9121a );
 a9125a <=( (not A266)  and  A265 );
 a9128a <=( A269  and  A267 );
 a9129a <=( a9128a  and  a9125a );
 a9130a <=( a9129a  and  a9122a );
 a9134a <=( (not A167)  and  A169 );
 a9135a <=( (not A170)  and  a9134a );
 a9138a <=( (not A199)  and  (not A166) );
 a9141a <=( A232  and  (not A200) );
 a9142a <=( a9141a  and  a9138a );
 a9143a <=( a9142a  and  a9135a );
 a9147a <=( A236  and  A234 );
 a9148a <=( (not A233)  and  a9147a );
 a9151a <=( (not A299)  and  A298 );
 a9154a <=( A301  and  A300 );
 a9155a <=( a9154a  and  a9151a );
 a9156a <=( a9155a  and  a9148a );
 a9160a <=( (not A167)  and  A169 );
 a9161a <=( (not A170)  and  a9160a );
 a9164a <=( (not A199)  and  (not A166) );
 a9167a <=( A232  and  (not A200) );
 a9168a <=( a9167a  and  a9164a );
 a9169a <=( a9168a  and  a9161a );
 a9173a <=( A236  and  A234 );
 a9174a <=( (not A233)  and  a9173a );
 a9177a <=( (not A299)  and  A298 );
 a9180a <=( A302  and  A300 );
 a9181a <=( a9180a  and  a9177a );
 a9182a <=( a9181a  and  a9174a );
 a9186a <=( (not A167)  and  A169 );
 a9187a <=( (not A170)  and  a9186a );
 a9190a <=( (not A199)  and  (not A166) );
 a9193a <=( A232  and  (not A200) );
 a9194a <=( a9193a  and  a9190a );
 a9195a <=( a9194a  and  a9187a );
 a9199a <=( A236  and  A234 );
 a9200a <=( (not A233)  and  a9199a );
 a9203a <=( (not A266)  and  A265 );
 a9206a <=( A268  and  A267 );
 a9207a <=( a9206a  and  a9203a );
 a9208a <=( a9207a  and  a9200a );
 a9212a <=( (not A167)  and  A169 );
 a9213a <=( (not A170)  and  a9212a );
 a9216a <=( (not A199)  and  (not A166) );
 a9219a <=( A232  and  (not A200) );
 a9220a <=( a9219a  and  a9216a );
 a9221a <=( a9220a  and  a9213a );
 a9225a <=( A236  and  A234 );
 a9226a <=( (not A233)  and  a9225a );
 a9229a <=( (not A266)  and  A265 );
 a9232a <=( A269  and  A267 );
 a9233a <=( a9232a  and  a9229a );
 a9234a <=( a9233a  and  a9226a );
 a9238a <=( A167  and  (not A169) );
 a9239a <=( A170  and  a9238a );
 a9242a <=( A199  and  (not A166) );
 a9245a <=( A232  and  (not A201) );
 a9246a <=( a9245a  and  a9242a );
 a9247a <=( a9246a  and  a9239a );
 a9251a <=( A235  and  A234 );
 a9252a <=( (not A233)  and  a9251a );
 a9255a <=( (not A299)  and  A298 );
 a9258a <=( A301  and  A300 );
 a9259a <=( a9258a  and  a9255a );
 a9260a <=( a9259a  and  a9252a );
 a9264a <=( A167  and  (not A169) );
 a9265a <=( A170  and  a9264a );
 a9268a <=( A199  and  (not A166) );
 a9271a <=( A232  and  (not A201) );
 a9272a <=( a9271a  and  a9268a );
 a9273a <=( a9272a  and  a9265a );
 a9277a <=( A235  and  A234 );
 a9278a <=( (not A233)  and  a9277a );
 a9281a <=( (not A299)  and  A298 );
 a9284a <=( A302  and  A300 );
 a9285a <=( a9284a  and  a9281a );
 a9286a <=( a9285a  and  a9278a );
 a9290a <=( A167  and  (not A169) );
 a9291a <=( A170  and  a9290a );
 a9294a <=( A199  and  (not A166) );
 a9297a <=( A232  and  (not A201) );
 a9298a <=( a9297a  and  a9294a );
 a9299a <=( a9298a  and  a9291a );
 a9303a <=( A235  and  A234 );
 a9304a <=( (not A233)  and  a9303a );
 a9307a <=( (not A266)  and  A265 );
 a9310a <=( A268  and  A267 );
 a9311a <=( a9310a  and  a9307a );
 a9312a <=( a9311a  and  a9304a );
 a9316a <=( A167  and  (not A169) );
 a9317a <=( A170  and  a9316a );
 a9320a <=( A199  and  (not A166) );
 a9323a <=( A232  and  (not A201) );
 a9324a <=( a9323a  and  a9320a );
 a9325a <=( a9324a  and  a9317a );
 a9329a <=( A235  and  A234 );
 a9330a <=( (not A233)  and  a9329a );
 a9333a <=( (not A266)  and  A265 );
 a9336a <=( A269  and  A267 );
 a9337a <=( a9336a  and  a9333a );
 a9338a <=( a9337a  and  a9330a );
 a9342a <=( A167  and  (not A169) );
 a9343a <=( A170  and  a9342a );
 a9346a <=( A199  and  (not A166) );
 a9349a <=( A232  and  (not A201) );
 a9350a <=( a9349a  and  a9346a );
 a9351a <=( a9350a  and  a9343a );
 a9355a <=( A236  and  A234 );
 a9356a <=( (not A233)  and  a9355a );
 a9359a <=( (not A299)  and  A298 );
 a9362a <=( A301  and  A300 );
 a9363a <=( a9362a  and  a9359a );
 a9364a <=( a9363a  and  a9356a );
 a9368a <=( A167  and  (not A169) );
 a9369a <=( A170  and  a9368a );
 a9372a <=( A199  and  (not A166) );
 a9375a <=( A232  and  (not A201) );
 a9376a <=( a9375a  and  a9372a );
 a9377a <=( a9376a  and  a9369a );
 a9381a <=( A236  and  A234 );
 a9382a <=( (not A233)  and  a9381a );
 a9385a <=( (not A299)  and  A298 );
 a9388a <=( A302  and  A300 );
 a9389a <=( a9388a  and  a9385a );
 a9390a <=( a9389a  and  a9382a );
 a9394a <=( A167  and  (not A169) );
 a9395a <=( A170  and  a9394a );
 a9398a <=( A199  and  (not A166) );
 a9401a <=( A232  and  (not A201) );
 a9402a <=( a9401a  and  a9398a );
 a9403a <=( a9402a  and  a9395a );
 a9407a <=( A236  and  A234 );
 a9408a <=( (not A233)  and  a9407a );
 a9411a <=( (not A266)  and  A265 );
 a9414a <=( A268  and  A267 );
 a9415a <=( a9414a  and  a9411a );
 a9416a <=( a9415a  and  a9408a );
 a9420a <=( A167  and  (not A169) );
 a9421a <=( A170  and  a9420a );
 a9424a <=( A199  and  (not A166) );
 a9427a <=( A232  and  (not A201) );
 a9428a <=( a9427a  and  a9424a );
 a9429a <=( a9428a  and  a9421a );
 a9433a <=( A236  and  A234 );
 a9434a <=( (not A233)  and  a9433a );
 a9437a <=( (not A266)  and  A265 );
 a9440a <=( A269  and  A267 );
 a9441a <=( a9440a  and  a9437a );
 a9442a <=( a9441a  and  a9434a );
 a9446a <=( A167  and  (not A169) );
 a9447a <=( A170  and  a9446a );
 a9450a <=( A199  and  (not A166) );
 a9453a <=( A232  and  A200 );
 a9454a <=( a9453a  and  a9450a );
 a9455a <=( a9454a  and  a9447a );
 a9459a <=( A235  and  A234 );
 a9460a <=( (not A233)  and  a9459a );
 a9463a <=( (not A299)  and  A298 );
 a9466a <=( A301  and  A300 );
 a9467a <=( a9466a  and  a9463a );
 a9468a <=( a9467a  and  a9460a );
 a9472a <=( A167  and  (not A169) );
 a9473a <=( A170  and  a9472a );
 a9476a <=( A199  and  (not A166) );
 a9479a <=( A232  and  A200 );
 a9480a <=( a9479a  and  a9476a );
 a9481a <=( a9480a  and  a9473a );
 a9485a <=( A235  and  A234 );
 a9486a <=( (not A233)  and  a9485a );
 a9489a <=( (not A299)  and  A298 );
 a9492a <=( A302  and  A300 );
 a9493a <=( a9492a  and  a9489a );
 a9494a <=( a9493a  and  a9486a );
 a9498a <=( A167  and  (not A169) );
 a9499a <=( A170  and  a9498a );
 a9502a <=( A199  and  (not A166) );
 a9505a <=( A232  and  A200 );
 a9506a <=( a9505a  and  a9502a );
 a9507a <=( a9506a  and  a9499a );
 a9511a <=( A235  and  A234 );
 a9512a <=( (not A233)  and  a9511a );
 a9515a <=( (not A266)  and  A265 );
 a9518a <=( A268  and  A267 );
 a9519a <=( a9518a  and  a9515a );
 a9520a <=( a9519a  and  a9512a );
 a9524a <=( A167  and  (not A169) );
 a9525a <=( A170  and  a9524a );
 a9528a <=( A199  and  (not A166) );
 a9531a <=( A232  and  A200 );
 a9532a <=( a9531a  and  a9528a );
 a9533a <=( a9532a  and  a9525a );
 a9537a <=( A235  and  A234 );
 a9538a <=( (not A233)  and  a9537a );
 a9541a <=( (not A266)  and  A265 );
 a9544a <=( A269  and  A267 );
 a9545a <=( a9544a  and  a9541a );
 a9546a <=( a9545a  and  a9538a );
 a9550a <=( A167  and  (not A169) );
 a9551a <=( A170  and  a9550a );
 a9554a <=( A199  and  (not A166) );
 a9557a <=( A232  and  A200 );
 a9558a <=( a9557a  and  a9554a );
 a9559a <=( a9558a  and  a9551a );
 a9563a <=( A236  and  A234 );
 a9564a <=( (not A233)  and  a9563a );
 a9567a <=( (not A299)  and  A298 );
 a9570a <=( A301  and  A300 );
 a9571a <=( a9570a  and  a9567a );
 a9572a <=( a9571a  and  a9564a );
 a9576a <=( A167  and  (not A169) );
 a9577a <=( A170  and  a9576a );
 a9580a <=( A199  and  (not A166) );
 a9583a <=( A232  and  A200 );
 a9584a <=( a9583a  and  a9580a );
 a9585a <=( a9584a  and  a9577a );
 a9589a <=( A236  and  A234 );
 a9590a <=( (not A233)  and  a9589a );
 a9593a <=( (not A299)  and  A298 );
 a9596a <=( A302  and  A300 );
 a9597a <=( a9596a  and  a9593a );
 a9598a <=( a9597a  and  a9590a );
 a9602a <=( A167  and  (not A169) );
 a9603a <=( A170  and  a9602a );
 a9606a <=( A199  and  (not A166) );
 a9609a <=( A232  and  A200 );
 a9610a <=( a9609a  and  a9606a );
 a9611a <=( a9610a  and  a9603a );
 a9615a <=( A236  and  A234 );
 a9616a <=( (not A233)  and  a9615a );
 a9619a <=( (not A266)  and  A265 );
 a9622a <=( A268  and  A267 );
 a9623a <=( a9622a  and  a9619a );
 a9624a <=( a9623a  and  a9616a );
 a9628a <=( A167  and  (not A169) );
 a9629a <=( A170  and  a9628a );
 a9632a <=( A199  and  (not A166) );
 a9635a <=( A232  and  A200 );
 a9636a <=( a9635a  and  a9632a );
 a9637a <=( a9636a  and  a9629a );
 a9641a <=( A236  and  A234 );
 a9642a <=( (not A233)  and  a9641a );
 a9645a <=( (not A266)  and  A265 );
 a9648a <=( A269  and  A267 );
 a9649a <=( a9648a  and  a9645a );
 a9650a <=( a9649a  and  a9642a );
 a9654a <=( A167  and  (not A169) );
 a9655a <=( A170  and  a9654a );
 a9658a <=( (not A199)  and  (not A166) );
 a9661a <=( A232  and  (not A200) );
 a9662a <=( a9661a  and  a9658a );
 a9663a <=( a9662a  and  a9655a );
 a9667a <=( A235  and  A234 );
 a9668a <=( (not A233)  and  a9667a );
 a9671a <=( (not A299)  and  A298 );
 a9674a <=( A301  and  A300 );
 a9675a <=( a9674a  and  a9671a );
 a9676a <=( a9675a  and  a9668a );
 a9680a <=( A167  and  (not A169) );
 a9681a <=( A170  and  a9680a );
 a9684a <=( (not A199)  and  (not A166) );
 a9687a <=( A232  and  (not A200) );
 a9688a <=( a9687a  and  a9684a );
 a9689a <=( a9688a  and  a9681a );
 a9693a <=( A235  and  A234 );
 a9694a <=( (not A233)  and  a9693a );
 a9697a <=( (not A299)  and  A298 );
 a9700a <=( A302  and  A300 );
 a9701a <=( a9700a  and  a9697a );
 a9702a <=( a9701a  and  a9694a );
 a9706a <=( A167  and  (not A169) );
 a9707a <=( A170  and  a9706a );
 a9710a <=( (not A199)  and  (not A166) );
 a9713a <=( A232  and  (not A200) );
 a9714a <=( a9713a  and  a9710a );
 a9715a <=( a9714a  and  a9707a );
 a9719a <=( A235  and  A234 );
 a9720a <=( (not A233)  and  a9719a );
 a9723a <=( (not A266)  and  A265 );
 a9726a <=( A268  and  A267 );
 a9727a <=( a9726a  and  a9723a );
 a9728a <=( a9727a  and  a9720a );
 a9732a <=( A167  and  (not A169) );
 a9733a <=( A170  and  a9732a );
 a9736a <=( (not A199)  and  (not A166) );
 a9739a <=( A232  and  (not A200) );
 a9740a <=( a9739a  and  a9736a );
 a9741a <=( a9740a  and  a9733a );
 a9745a <=( A235  and  A234 );
 a9746a <=( (not A233)  and  a9745a );
 a9749a <=( (not A266)  and  A265 );
 a9752a <=( A269  and  A267 );
 a9753a <=( a9752a  and  a9749a );
 a9754a <=( a9753a  and  a9746a );
 a9758a <=( A167  and  (not A169) );
 a9759a <=( A170  and  a9758a );
 a9762a <=( (not A199)  and  (not A166) );
 a9765a <=( A232  and  (not A200) );
 a9766a <=( a9765a  and  a9762a );
 a9767a <=( a9766a  and  a9759a );
 a9771a <=( A236  and  A234 );
 a9772a <=( (not A233)  and  a9771a );
 a9775a <=( (not A299)  and  A298 );
 a9778a <=( A301  and  A300 );
 a9779a <=( a9778a  and  a9775a );
 a9780a <=( a9779a  and  a9772a );
 a9784a <=( A167  and  (not A169) );
 a9785a <=( A170  and  a9784a );
 a9788a <=( (not A199)  and  (not A166) );
 a9791a <=( A232  and  (not A200) );
 a9792a <=( a9791a  and  a9788a );
 a9793a <=( a9792a  and  a9785a );
 a9797a <=( A236  and  A234 );
 a9798a <=( (not A233)  and  a9797a );
 a9801a <=( (not A299)  and  A298 );
 a9804a <=( A302  and  A300 );
 a9805a <=( a9804a  and  a9801a );
 a9806a <=( a9805a  and  a9798a );
 a9810a <=( A167  and  (not A169) );
 a9811a <=( A170  and  a9810a );
 a9814a <=( (not A199)  and  (not A166) );
 a9817a <=( A232  and  (not A200) );
 a9818a <=( a9817a  and  a9814a );
 a9819a <=( a9818a  and  a9811a );
 a9823a <=( A236  and  A234 );
 a9824a <=( (not A233)  and  a9823a );
 a9827a <=( (not A266)  and  A265 );
 a9830a <=( A268  and  A267 );
 a9831a <=( a9830a  and  a9827a );
 a9832a <=( a9831a  and  a9824a );
 a9836a <=( A167  and  (not A169) );
 a9837a <=( A170  and  a9836a );
 a9840a <=( (not A199)  and  (not A166) );
 a9843a <=( A232  and  (not A200) );
 a9844a <=( a9843a  and  a9840a );
 a9845a <=( a9844a  and  a9837a );
 a9849a <=( A236  and  A234 );
 a9850a <=( (not A233)  and  a9849a );
 a9853a <=( (not A266)  and  A265 );
 a9856a <=( A269  and  A267 );
 a9857a <=( a9856a  and  a9853a );
 a9858a <=( a9857a  and  a9850a );
 a9862a <=( (not A167)  and  (not A169) );
 a9863a <=( A170  and  a9862a );
 a9866a <=( A199  and  A166 );
 a9869a <=( A232  and  (not A201) );
 a9870a <=( a9869a  and  a9866a );
 a9871a <=( a9870a  and  a9863a );
 a9875a <=( A235  and  A234 );
 a9876a <=( (not A233)  and  a9875a );
 a9879a <=( (not A299)  and  A298 );
 a9882a <=( A301  and  A300 );
 a9883a <=( a9882a  and  a9879a );
 a9884a <=( a9883a  and  a9876a );
 a9888a <=( (not A167)  and  (not A169) );
 a9889a <=( A170  and  a9888a );
 a9892a <=( A199  and  A166 );
 a9895a <=( A232  and  (not A201) );
 a9896a <=( a9895a  and  a9892a );
 a9897a <=( a9896a  and  a9889a );
 a9901a <=( A235  and  A234 );
 a9902a <=( (not A233)  and  a9901a );
 a9905a <=( (not A299)  and  A298 );
 a9908a <=( A302  and  A300 );
 a9909a <=( a9908a  and  a9905a );
 a9910a <=( a9909a  and  a9902a );
 a9914a <=( (not A167)  and  (not A169) );
 a9915a <=( A170  and  a9914a );
 a9918a <=( A199  and  A166 );
 a9921a <=( A232  and  (not A201) );
 a9922a <=( a9921a  and  a9918a );
 a9923a <=( a9922a  and  a9915a );
 a9927a <=( A235  and  A234 );
 a9928a <=( (not A233)  and  a9927a );
 a9931a <=( (not A266)  and  A265 );
 a9934a <=( A268  and  A267 );
 a9935a <=( a9934a  and  a9931a );
 a9936a <=( a9935a  and  a9928a );
 a9940a <=( (not A167)  and  (not A169) );
 a9941a <=( A170  and  a9940a );
 a9944a <=( A199  and  A166 );
 a9947a <=( A232  and  (not A201) );
 a9948a <=( a9947a  and  a9944a );
 a9949a <=( a9948a  and  a9941a );
 a9953a <=( A235  and  A234 );
 a9954a <=( (not A233)  and  a9953a );
 a9957a <=( (not A266)  and  A265 );
 a9960a <=( A269  and  A267 );
 a9961a <=( a9960a  and  a9957a );
 a9962a <=( a9961a  and  a9954a );
 a9966a <=( (not A167)  and  (not A169) );
 a9967a <=( A170  and  a9966a );
 a9970a <=( A199  and  A166 );
 a9973a <=( A232  and  (not A201) );
 a9974a <=( a9973a  and  a9970a );
 a9975a <=( a9974a  and  a9967a );
 a9979a <=( A236  and  A234 );
 a9980a <=( (not A233)  and  a9979a );
 a9983a <=( (not A299)  and  A298 );
 a9986a <=( A301  and  A300 );
 a9987a <=( a9986a  and  a9983a );
 a9988a <=( a9987a  and  a9980a );
 a9992a <=( (not A167)  and  (not A169) );
 a9993a <=( A170  and  a9992a );
 a9996a <=( A199  and  A166 );
 a9999a <=( A232  and  (not A201) );
 a10000a <=( a9999a  and  a9996a );
 a10001a <=( a10000a  and  a9993a );
 a10005a <=( A236  and  A234 );
 a10006a <=( (not A233)  and  a10005a );
 a10009a <=( (not A299)  and  A298 );
 a10012a <=( A302  and  A300 );
 a10013a <=( a10012a  and  a10009a );
 a10014a <=( a10013a  and  a10006a );
 a10018a <=( (not A167)  and  (not A169) );
 a10019a <=( A170  and  a10018a );
 a10022a <=( A199  and  A166 );
 a10025a <=( A232  and  (not A201) );
 a10026a <=( a10025a  and  a10022a );
 a10027a <=( a10026a  and  a10019a );
 a10031a <=( A236  and  A234 );
 a10032a <=( (not A233)  and  a10031a );
 a10035a <=( (not A266)  and  A265 );
 a10038a <=( A268  and  A267 );
 a10039a <=( a10038a  and  a10035a );
 a10040a <=( a10039a  and  a10032a );
 a10044a <=( (not A167)  and  (not A169) );
 a10045a <=( A170  and  a10044a );
 a10048a <=( A199  and  A166 );
 a10051a <=( A232  and  (not A201) );
 a10052a <=( a10051a  and  a10048a );
 a10053a <=( a10052a  and  a10045a );
 a10057a <=( A236  and  A234 );
 a10058a <=( (not A233)  and  a10057a );
 a10061a <=( (not A266)  and  A265 );
 a10064a <=( A269  and  A267 );
 a10065a <=( a10064a  and  a10061a );
 a10066a <=( a10065a  and  a10058a );
 a10070a <=( (not A167)  and  (not A169) );
 a10071a <=( A170  and  a10070a );
 a10074a <=( A199  and  A166 );
 a10077a <=( A232  and  A200 );
 a10078a <=( a10077a  and  a10074a );
 a10079a <=( a10078a  and  a10071a );
 a10083a <=( A235  and  A234 );
 a10084a <=( (not A233)  and  a10083a );
 a10087a <=( (not A299)  and  A298 );
 a10090a <=( A301  and  A300 );
 a10091a <=( a10090a  and  a10087a );
 a10092a <=( a10091a  and  a10084a );
 a10096a <=( (not A167)  and  (not A169) );
 a10097a <=( A170  and  a10096a );
 a10100a <=( A199  and  A166 );
 a10103a <=( A232  and  A200 );
 a10104a <=( a10103a  and  a10100a );
 a10105a <=( a10104a  and  a10097a );
 a10109a <=( A235  and  A234 );
 a10110a <=( (not A233)  and  a10109a );
 a10113a <=( (not A299)  and  A298 );
 a10116a <=( A302  and  A300 );
 a10117a <=( a10116a  and  a10113a );
 a10118a <=( a10117a  and  a10110a );
 a10122a <=( (not A167)  and  (not A169) );
 a10123a <=( A170  and  a10122a );
 a10126a <=( A199  and  A166 );
 a10129a <=( A232  and  A200 );
 a10130a <=( a10129a  and  a10126a );
 a10131a <=( a10130a  and  a10123a );
 a10135a <=( A235  and  A234 );
 a10136a <=( (not A233)  and  a10135a );
 a10139a <=( (not A266)  and  A265 );
 a10142a <=( A268  and  A267 );
 a10143a <=( a10142a  and  a10139a );
 a10144a <=( a10143a  and  a10136a );
 a10148a <=( (not A167)  and  (not A169) );
 a10149a <=( A170  and  a10148a );
 a10152a <=( A199  and  A166 );
 a10155a <=( A232  and  A200 );
 a10156a <=( a10155a  and  a10152a );
 a10157a <=( a10156a  and  a10149a );
 a10161a <=( A235  and  A234 );
 a10162a <=( (not A233)  and  a10161a );
 a10165a <=( (not A266)  and  A265 );
 a10168a <=( A269  and  A267 );
 a10169a <=( a10168a  and  a10165a );
 a10170a <=( a10169a  and  a10162a );
 a10174a <=( (not A167)  and  (not A169) );
 a10175a <=( A170  and  a10174a );
 a10178a <=( A199  and  A166 );
 a10181a <=( A232  and  A200 );
 a10182a <=( a10181a  and  a10178a );
 a10183a <=( a10182a  and  a10175a );
 a10187a <=( A236  and  A234 );
 a10188a <=( (not A233)  and  a10187a );
 a10191a <=( (not A299)  and  A298 );
 a10194a <=( A301  and  A300 );
 a10195a <=( a10194a  and  a10191a );
 a10196a <=( a10195a  and  a10188a );
 a10200a <=( (not A167)  and  (not A169) );
 a10201a <=( A170  and  a10200a );
 a10204a <=( A199  and  A166 );
 a10207a <=( A232  and  A200 );
 a10208a <=( a10207a  and  a10204a );
 a10209a <=( a10208a  and  a10201a );
 a10213a <=( A236  and  A234 );
 a10214a <=( (not A233)  and  a10213a );
 a10217a <=( (not A299)  and  A298 );
 a10220a <=( A302  and  A300 );
 a10221a <=( a10220a  and  a10217a );
 a10222a <=( a10221a  and  a10214a );
 a10226a <=( (not A167)  and  (not A169) );
 a10227a <=( A170  and  a10226a );
 a10230a <=( A199  and  A166 );
 a10233a <=( A232  and  A200 );
 a10234a <=( a10233a  and  a10230a );
 a10235a <=( a10234a  and  a10227a );
 a10239a <=( A236  and  A234 );
 a10240a <=( (not A233)  and  a10239a );
 a10243a <=( (not A266)  and  A265 );
 a10246a <=( A268  and  A267 );
 a10247a <=( a10246a  and  a10243a );
 a10248a <=( a10247a  and  a10240a );
 a10252a <=( (not A167)  and  (not A169) );
 a10253a <=( A170  and  a10252a );
 a10256a <=( A199  and  A166 );
 a10259a <=( A232  and  A200 );
 a10260a <=( a10259a  and  a10256a );
 a10261a <=( a10260a  and  a10253a );
 a10265a <=( A236  and  A234 );
 a10266a <=( (not A233)  and  a10265a );
 a10269a <=( (not A266)  and  A265 );
 a10272a <=( A269  and  A267 );
 a10273a <=( a10272a  and  a10269a );
 a10274a <=( a10273a  and  a10266a );
 a10278a <=( (not A167)  and  (not A169) );
 a10279a <=( A170  and  a10278a );
 a10282a <=( (not A199)  and  A166 );
 a10285a <=( A232  and  (not A200) );
 a10286a <=( a10285a  and  a10282a );
 a10287a <=( a10286a  and  a10279a );
 a10291a <=( A235  and  A234 );
 a10292a <=( (not A233)  and  a10291a );
 a10295a <=( (not A299)  and  A298 );
 a10298a <=( A301  and  A300 );
 a10299a <=( a10298a  and  a10295a );
 a10300a <=( a10299a  and  a10292a );
 a10304a <=( (not A167)  and  (not A169) );
 a10305a <=( A170  and  a10304a );
 a10308a <=( (not A199)  and  A166 );
 a10311a <=( A232  and  (not A200) );
 a10312a <=( a10311a  and  a10308a );
 a10313a <=( a10312a  and  a10305a );
 a10317a <=( A235  and  A234 );
 a10318a <=( (not A233)  and  a10317a );
 a10321a <=( (not A299)  and  A298 );
 a10324a <=( A302  and  A300 );
 a10325a <=( a10324a  and  a10321a );
 a10326a <=( a10325a  and  a10318a );
 a10330a <=( (not A167)  and  (not A169) );
 a10331a <=( A170  and  a10330a );
 a10334a <=( (not A199)  and  A166 );
 a10337a <=( A232  and  (not A200) );
 a10338a <=( a10337a  and  a10334a );
 a10339a <=( a10338a  and  a10331a );
 a10343a <=( A235  and  A234 );
 a10344a <=( (not A233)  and  a10343a );
 a10347a <=( (not A266)  and  A265 );
 a10350a <=( A268  and  A267 );
 a10351a <=( a10350a  and  a10347a );
 a10352a <=( a10351a  and  a10344a );
 a10356a <=( (not A167)  and  (not A169) );
 a10357a <=( A170  and  a10356a );
 a10360a <=( (not A199)  and  A166 );
 a10363a <=( A232  and  (not A200) );
 a10364a <=( a10363a  and  a10360a );
 a10365a <=( a10364a  and  a10357a );
 a10369a <=( A235  and  A234 );
 a10370a <=( (not A233)  and  a10369a );
 a10373a <=( (not A266)  and  A265 );
 a10376a <=( A269  and  A267 );
 a10377a <=( a10376a  and  a10373a );
 a10378a <=( a10377a  and  a10370a );
 a10382a <=( (not A167)  and  (not A169) );
 a10383a <=( A170  and  a10382a );
 a10386a <=( (not A199)  and  A166 );
 a10389a <=( A232  and  (not A200) );
 a10390a <=( a10389a  and  a10386a );
 a10391a <=( a10390a  and  a10383a );
 a10395a <=( A236  and  A234 );
 a10396a <=( (not A233)  and  a10395a );
 a10399a <=( (not A299)  and  A298 );
 a10402a <=( A301  and  A300 );
 a10403a <=( a10402a  and  a10399a );
 a10404a <=( a10403a  and  a10396a );
 a10408a <=( (not A167)  and  (not A169) );
 a10409a <=( A170  and  a10408a );
 a10412a <=( (not A199)  and  A166 );
 a10415a <=( A232  and  (not A200) );
 a10416a <=( a10415a  and  a10412a );
 a10417a <=( a10416a  and  a10409a );
 a10421a <=( A236  and  A234 );
 a10422a <=( (not A233)  and  a10421a );
 a10425a <=( (not A299)  and  A298 );
 a10428a <=( A302  and  A300 );
 a10429a <=( a10428a  and  a10425a );
 a10430a <=( a10429a  and  a10422a );
 a10434a <=( (not A167)  and  (not A169) );
 a10435a <=( A170  and  a10434a );
 a10438a <=( (not A199)  and  A166 );
 a10441a <=( A232  and  (not A200) );
 a10442a <=( a10441a  and  a10438a );
 a10443a <=( a10442a  and  a10435a );
 a10447a <=( A236  and  A234 );
 a10448a <=( (not A233)  and  a10447a );
 a10451a <=( (not A266)  and  A265 );
 a10454a <=( A268  and  A267 );
 a10455a <=( a10454a  and  a10451a );
 a10456a <=( a10455a  and  a10448a );
 a10460a <=( (not A167)  and  (not A169) );
 a10461a <=( A170  and  a10460a );
 a10464a <=( (not A199)  and  A166 );
 a10467a <=( A232  and  (not A200) );
 a10468a <=( a10467a  and  a10464a );
 a10469a <=( a10468a  and  a10461a );
 a10473a <=( A236  and  A234 );
 a10474a <=( (not A233)  and  a10473a );
 a10477a <=( (not A266)  and  A265 );
 a10480a <=( A269  and  A267 );
 a10481a <=( a10480a  and  a10477a );
 a10482a <=( a10481a  and  a10474a );
 a10486a <=( A167  and  A169 );
 a10487a <=( (not A170)  and  a10486a );
 a10490a <=( A199  and  A166 );
 a10493a <=( (not A203)  and  (not A202) );
 a10494a <=( a10493a  and  a10490a );
 a10495a <=( a10494a  and  a10487a );
 a10498a <=( (not A233)  and  A232 );
 a10501a <=( A235  and  A234 );
 a10502a <=( a10501a  and  a10498a );
 a10505a <=( (not A299)  and  A298 );
 a10508a <=( A301  and  A300 );
 a10509a <=( a10508a  and  a10505a );
 a10510a <=( a10509a  and  a10502a );
 a10514a <=( A167  and  A169 );
 a10515a <=( (not A170)  and  a10514a );
 a10518a <=( A199  and  A166 );
 a10521a <=( (not A203)  and  (not A202) );
 a10522a <=( a10521a  and  a10518a );
 a10523a <=( a10522a  and  a10515a );
 a10526a <=( (not A233)  and  A232 );
 a10529a <=( A235  and  A234 );
 a10530a <=( a10529a  and  a10526a );
 a10533a <=( (not A299)  and  A298 );
 a10536a <=( A302  and  A300 );
 a10537a <=( a10536a  and  a10533a );
 a10538a <=( a10537a  and  a10530a );
 a10542a <=( A167  and  A169 );
 a10543a <=( (not A170)  and  a10542a );
 a10546a <=( A199  and  A166 );
 a10549a <=( (not A203)  and  (not A202) );
 a10550a <=( a10549a  and  a10546a );
 a10551a <=( a10550a  and  a10543a );
 a10554a <=( (not A233)  and  A232 );
 a10557a <=( A235  and  A234 );
 a10558a <=( a10557a  and  a10554a );
 a10561a <=( (not A266)  and  A265 );
 a10564a <=( A268  and  A267 );
 a10565a <=( a10564a  and  a10561a );
 a10566a <=( a10565a  and  a10558a );
 a10570a <=( A167  and  A169 );
 a10571a <=( (not A170)  and  a10570a );
 a10574a <=( A199  and  A166 );
 a10577a <=( (not A203)  and  (not A202) );
 a10578a <=( a10577a  and  a10574a );
 a10579a <=( a10578a  and  a10571a );
 a10582a <=( (not A233)  and  A232 );
 a10585a <=( A235  and  A234 );
 a10586a <=( a10585a  and  a10582a );
 a10589a <=( (not A266)  and  A265 );
 a10592a <=( A269  and  A267 );
 a10593a <=( a10592a  and  a10589a );
 a10594a <=( a10593a  and  a10586a );
 a10598a <=( A167  and  A169 );
 a10599a <=( (not A170)  and  a10598a );
 a10602a <=( A199  and  A166 );
 a10605a <=( (not A203)  and  (not A202) );
 a10606a <=( a10605a  and  a10602a );
 a10607a <=( a10606a  and  a10599a );
 a10610a <=( (not A233)  and  A232 );
 a10613a <=( A236  and  A234 );
 a10614a <=( a10613a  and  a10610a );
 a10617a <=( (not A299)  and  A298 );
 a10620a <=( A301  and  A300 );
 a10621a <=( a10620a  and  a10617a );
 a10622a <=( a10621a  and  a10614a );
 a10626a <=( A167  and  A169 );
 a10627a <=( (not A170)  and  a10626a );
 a10630a <=( A199  and  A166 );
 a10633a <=( (not A203)  and  (not A202) );
 a10634a <=( a10633a  and  a10630a );
 a10635a <=( a10634a  and  a10627a );
 a10638a <=( (not A233)  and  A232 );
 a10641a <=( A236  and  A234 );
 a10642a <=( a10641a  and  a10638a );
 a10645a <=( (not A299)  and  A298 );
 a10648a <=( A302  and  A300 );
 a10649a <=( a10648a  and  a10645a );
 a10650a <=( a10649a  and  a10642a );
 a10654a <=( A167  and  A169 );
 a10655a <=( (not A170)  and  a10654a );
 a10658a <=( A199  and  A166 );
 a10661a <=( (not A203)  and  (not A202) );
 a10662a <=( a10661a  and  a10658a );
 a10663a <=( a10662a  and  a10655a );
 a10666a <=( (not A233)  and  A232 );
 a10669a <=( A236  and  A234 );
 a10670a <=( a10669a  and  a10666a );
 a10673a <=( (not A266)  and  A265 );
 a10676a <=( A268  and  A267 );
 a10677a <=( a10676a  and  a10673a );
 a10678a <=( a10677a  and  a10670a );
 a10682a <=( A167  and  A169 );
 a10683a <=( (not A170)  and  a10682a );
 a10686a <=( A199  and  A166 );
 a10689a <=( (not A203)  and  (not A202) );
 a10690a <=( a10689a  and  a10686a );
 a10691a <=( a10690a  and  a10683a );
 a10694a <=( (not A233)  and  A232 );
 a10697a <=( A236  and  A234 );
 a10698a <=( a10697a  and  a10694a );
 a10701a <=( (not A266)  and  A265 );
 a10704a <=( A269  and  A267 );
 a10705a <=( a10704a  and  a10701a );
 a10706a <=( a10705a  and  a10698a );
 a10710a <=( (not A167)  and  A169 );
 a10711a <=( (not A170)  and  a10710a );
 a10714a <=( A199  and  (not A166) );
 a10717a <=( (not A203)  and  (not A202) );
 a10718a <=( a10717a  and  a10714a );
 a10719a <=( a10718a  and  a10711a );
 a10722a <=( (not A233)  and  A232 );
 a10725a <=( A235  and  A234 );
 a10726a <=( a10725a  and  a10722a );
 a10729a <=( (not A299)  and  A298 );
 a10732a <=( A301  and  A300 );
 a10733a <=( a10732a  and  a10729a );
 a10734a <=( a10733a  and  a10726a );
 a10738a <=( (not A167)  and  A169 );
 a10739a <=( (not A170)  and  a10738a );
 a10742a <=( A199  and  (not A166) );
 a10745a <=( (not A203)  and  (not A202) );
 a10746a <=( a10745a  and  a10742a );
 a10747a <=( a10746a  and  a10739a );
 a10750a <=( (not A233)  and  A232 );
 a10753a <=( A235  and  A234 );
 a10754a <=( a10753a  and  a10750a );
 a10757a <=( (not A299)  and  A298 );
 a10760a <=( A302  and  A300 );
 a10761a <=( a10760a  and  a10757a );
 a10762a <=( a10761a  and  a10754a );
 a10766a <=( (not A167)  and  A169 );
 a10767a <=( (not A170)  and  a10766a );
 a10770a <=( A199  and  (not A166) );
 a10773a <=( (not A203)  and  (not A202) );
 a10774a <=( a10773a  and  a10770a );
 a10775a <=( a10774a  and  a10767a );
 a10778a <=( (not A233)  and  A232 );
 a10781a <=( A235  and  A234 );
 a10782a <=( a10781a  and  a10778a );
 a10785a <=( (not A266)  and  A265 );
 a10788a <=( A268  and  A267 );
 a10789a <=( a10788a  and  a10785a );
 a10790a <=( a10789a  and  a10782a );
 a10794a <=( (not A167)  and  A169 );
 a10795a <=( (not A170)  and  a10794a );
 a10798a <=( A199  and  (not A166) );
 a10801a <=( (not A203)  and  (not A202) );
 a10802a <=( a10801a  and  a10798a );
 a10803a <=( a10802a  and  a10795a );
 a10806a <=( (not A233)  and  A232 );
 a10809a <=( A235  and  A234 );
 a10810a <=( a10809a  and  a10806a );
 a10813a <=( (not A266)  and  A265 );
 a10816a <=( A269  and  A267 );
 a10817a <=( a10816a  and  a10813a );
 a10818a <=( a10817a  and  a10810a );
 a10822a <=( (not A167)  and  A169 );
 a10823a <=( (not A170)  and  a10822a );
 a10826a <=( A199  and  (not A166) );
 a10829a <=( (not A203)  and  (not A202) );
 a10830a <=( a10829a  and  a10826a );
 a10831a <=( a10830a  and  a10823a );
 a10834a <=( (not A233)  and  A232 );
 a10837a <=( A236  and  A234 );
 a10838a <=( a10837a  and  a10834a );
 a10841a <=( (not A299)  and  A298 );
 a10844a <=( A301  and  A300 );
 a10845a <=( a10844a  and  a10841a );
 a10846a <=( a10845a  and  a10838a );
 a10850a <=( (not A167)  and  A169 );
 a10851a <=( (not A170)  and  a10850a );
 a10854a <=( A199  and  (not A166) );
 a10857a <=( (not A203)  and  (not A202) );
 a10858a <=( a10857a  and  a10854a );
 a10859a <=( a10858a  and  a10851a );
 a10862a <=( (not A233)  and  A232 );
 a10865a <=( A236  and  A234 );
 a10866a <=( a10865a  and  a10862a );
 a10869a <=( (not A299)  and  A298 );
 a10872a <=( A302  and  A300 );
 a10873a <=( a10872a  and  a10869a );
 a10874a <=( a10873a  and  a10866a );
 a10878a <=( (not A167)  and  A169 );
 a10879a <=( (not A170)  and  a10878a );
 a10882a <=( A199  and  (not A166) );
 a10885a <=( (not A203)  and  (not A202) );
 a10886a <=( a10885a  and  a10882a );
 a10887a <=( a10886a  and  a10879a );
 a10890a <=( (not A233)  and  A232 );
 a10893a <=( A236  and  A234 );
 a10894a <=( a10893a  and  a10890a );
 a10897a <=( (not A266)  and  A265 );
 a10900a <=( A268  and  A267 );
 a10901a <=( a10900a  and  a10897a );
 a10902a <=( a10901a  and  a10894a );
 a10906a <=( (not A167)  and  A169 );
 a10907a <=( (not A170)  and  a10906a );
 a10910a <=( A199  and  (not A166) );
 a10913a <=( (not A203)  and  (not A202) );
 a10914a <=( a10913a  and  a10910a );
 a10915a <=( a10914a  and  a10907a );
 a10918a <=( (not A233)  and  A232 );
 a10921a <=( A236  and  A234 );
 a10922a <=( a10921a  and  a10918a );
 a10925a <=( (not A266)  and  A265 );
 a10928a <=( A269  and  A267 );
 a10929a <=( a10928a  and  a10925a );
 a10930a <=( a10929a  and  a10922a );
 a10934a <=( A167  and  (not A169) );
 a10935a <=( A170  and  a10934a );
 a10938a <=( A199  and  (not A166) );
 a10941a <=( (not A203)  and  (not A202) );
 a10942a <=( a10941a  and  a10938a );
 a10943a <=( a10942a  and  a10935a );
 a10946a <=( (not A233)  and  A232 );
 a10949a <=( A235  and  A234 );
 a10950a <=( a10949a  and  a10946a );
 a10953a <=( (not A299)  and  A298 );
 a10956a <=( A301  and  A300 );
 a10957a <=( a10956a  and  a10953a );
 a10958a <=( a10957a  and  a10950a );
 a10962a <=( A167  and  (not A169) );
 a10963a <=( A170  and  a10962a );
 a10966a <=( A199  and  (not A166) );
 a10969a <=( (not A203)  and  (not A202) );
 a10970a <=( a10969a  and  a10966a );
 a10971a <=( a10970a  and  a10963a );
 a10974a <=( (not A233)  and  A232 );
 a10977a <=( A235  and  A234 );
 a10978a <=( a10977a  and  a10974a );
 a10981a <=( (not A299)  and  A298 );
 a10984a <=( A302  and  A300 );
 a10985a <=( a10984a  and  a10981a );
 a10986a <=( a10985a  and  a10978a );
 a10990a <=( A167  and  (not A169) );
 a10991a <=( A170  and  a10990a );
 a10994a <=( A199  and  (not A166) );
 a10997a <=( (not A203)  and  (not A202) );
 a10998a <=( a10997a  and  a10994a );
 a10999a <=( a10998a  and  a10991a );
 a11002a <=( (not A233)  and  A232 );
 a11005a <=( A235  and  A234 );
 a11006a <=( a11005a  and  a11002a );
 a11009a <=( (not A266)  and  A265 );
 a11012a <=( A268  and  A267 );
 a11013a <=( a11012a  and  a11009a );
 a11014a <=( a11013a  and  a11006a );
 a11018a <=( A167  and  (not A169) );
 a11019a <=( A170  and  a11018a );
 a11022a <=( A199  and  (not A166) );
 a11025a <=( (not A203)  and  (not A202) );
 a11026a <=( a11025a  and  a11022a );
 a11027a <=( a11026a  and  a11019a );
 a11030a <=( (not A233)  and  A232 );
 a11033a <=( A235  and  A234 );
 a11034a <=( a11033a  and  a11030a );
 a11037a <=( (not A266)  and  A265 );
 a11040a <=( A269  and  A267 );
 a11041a <=( a11040a  and  a11037a );
 a11042a <=( a11041a  and  a11034a );
 a11046a <=( A167  and  (not A169) );
 a11047a <=( A170  and  a11046a );
 a11050a <=( A199  and  (not A166) );
 a11053a <=( (not A203)  and  (not A202) );
 a11054a <=( a11053a  and  a11050a );
 a11055a <=( a11054a  and  a11047a );
 a11058a <=( (not A233)  and  A232 );
 a11061a <=( A236  and  A234 );
 a11062a <=( a11061a  and  a11058a );
 a11065a <=( (not A299)  and  A298 );
 a11068a <=( A301  and  A300 );
 a11069a <=( a11068a  and  a11065a );
 a11070a <=( a11069a  and  a11062a );
 a11074a <=( A167  and  (not A169) );
 a11075a <=( A170  and  a11074a );
 a11078a <=( A199  and  (not A166) );
 a11081a <=( (not A203)  and  (not A202) );
 a11082a <=( a11081a  and  a11078a );
 a11083a <=( a11082a  and  a11075a );
 a11086a <=( (not A233)  and  A232 );
 a11089a <=( A236  and  A234 );
 a11090a <=( a11089a  and  a11086a );
 a11093a <=( (not A299)  and  A298 );
 a11096a <=( A302  and  A300 );
 a11097a <=( a11096a  and  a11093a );
 a11098a <=( a11097a  and  a11090a );
 a11102a <=( A167  and  (not A169) );
 a11103a <=( A170  and  a11102a );
 a11106a <=( A199  and  (not A166) );
 a11109a <=( (not A203)  and  (not A202) );
 a11110a <=( a11109a  and  a11106a );
 a11111a <=( a11110a  and  a11103a );
 a11114a <=( (not A233)  and  A232 );
 a11117a <=( A236  and  A234 );
 a11118a <=( a11117a  and  a11114a );
 a11121a <=( (not A266)  and  A265 );
 a11124a <=( A268  and  A267 );
 a11125a <=( a11124a  and  a11121a );
 a11126a <=( a11125a  and  a11118a );
 a11130a <=( A167  and  (not A169) );
 a11131a <=( A170  and  a11130a );
 a11134a <=( A199  and  (not A166) );
 a11137a <=( (not A203)  and  (not A202) );
 a11138a <=( a11137a  and  a11134a );
 a11139a <=( a11138a  and  a11131a );
 a11142a <=( (not A233)  and  A232 );
 a11145a <=( A236  and  A234 );
 a11146a <=( a11145a  and  a11142a );
 a11149a <=( (not A266)  and  A265 );
 a11152a <=( A269  and  A267 );
 a11153a <=( a11152a  and  a11149a );
 a11154a <=( a11153a  and  a11146a );
 a11158a <=( (not A167)  and  (not A169) );
 a11159a <=( A170  and  a11158a );
 a11162a <=( A199  and  A166 );
 a11165a <=( (not A203)  and  (not A202) );
 a11166a <=( a11165a  and  a11162a );
 a11167a <=( a11166a  and  a11159a );
 a11170a <=( (not A233)  and  A232 );
 a11173a <=( A235  and  A234 );
 a11174a <=( a11173a  and  a11170a );
 a11177a <=( (not A299)  and  A298 );
 a11180a <=( A301  and  A300 );
 a11181a <=( a11180a  and  a11177a );
 a11182a <=( a11181a  and  a11174a );
 a11186a <=( (not A167)  and  (not A169) );
 a11187a <=( A170  and  a11186a );
 a11190a <=( A199  and  A166 );
 a11193a <=( (not A203)  and  (not A202) );
 a11194a <=( a11193a  and  a11190a );
 a11195a <=( a11194a  and  a11187a );
 a11198a <=( (not A233)  and  A232 );
 a11201a <=( A235  and  A234 );
 a11202a <=( a11201a  and  a11198a );
 a11205a <=( (not A299)  and  A298 );
 a11208a <=( A302  and  A300 );
 a11209a <=( a11208a  and  a11205a );
 a11210a <=( a11209a  and  a11202a );
 a11214a <=( (not A167)  and  (not A169) );
 a11215a <=( A170  and  a11214a );
 a11218a <=( A199  and  A166 );
 a11221a <=( (not A203)  and  (not A202) );
 a11222a <=( a11221a  and  a11218a );
 a11223a <=( a11222a  and  a11215a );
 a11226a <=( (not A233)  and  A232 );
 a11229a <=( A235  and  A234 );
 a11230a <=( a11229a  and  a11226a );
 a11233a <=( (not A266)  and  A265 );
 a11236a <=( A268  and  A267 );
 a11237a <=( a11236a  and  a11233a );
 a11238a <=( a11237a  and  a11230a );
 a11242a <=( (not A167)  and  (not A169) );
 a11243a <=( A170  and  a11242a );
 a11246a <=( A199  and  A166 );
 a11249a <=( (not A203)  and  (not A202) );
 a11250a <=( a11249a  and  a11246a );
 a11251a <=( a11250a  and  a11243a );
 a11254a <=( (not A233)  and  A232 );
 a11257a <=( A235  and  A234 );
 a11258a <=( a11257a  and  a11254a );
 a11261a <=( (not A266)  and  A265 );
 a11264a <=( A269  and  A267 );
 a11265a <=( a11264a  and  a11261a );
 a11266a <=( a11265a  and  a11258a );
 a11270a <=( (not A167)  and  (not A169) );
 a11271a <=( A170  and  a11270a );
 a11274a <=( A199  and  A166 );
 a11277a <=( (not A203)  and  (not A202) );
 a11278a <=( a11277a  and  a11274a );
 a11279a <=( a11278a  and  a11271a );
 a11282a <=( (not A233)  and  A232 );
 a11285a <=( A236  and  A234 );
 a11286a <=( a11285a  and  a11282a );
 a11289a <=( (not A299)  and  A298 );
 a11292a <=( A301  and  A300 );
 a11293a <=( a11292a  and  a11289a );
 a11294a <=( a11293a  and  a11286a );
 a11298a <=( (not A167)  and  (not A169) );
 a11299a <=( A170  and  a11298a );
 a11302a <=( A199  and  A166 );
 a11305a <=( (not A203)  and  (not A202) );
 a11306a <=( a11305a  and  a11302a );
 a11307a <=( a11306a  and  a11299a );
 a11310a <=( (not A233)  and  A232 );
 a11313a <=( A236  and  A234 );
 a11314a <=( a11313a  and  a11310a );
 a11317a <=( (not A299)  and  A298 );
 a11320a <=( A302  and  A300 );
 a11321a <=( a11320a  and  a11317a );
 a11322a <=( a11321a  and  a11314a );
 a11326a <=( (not A167)  and  (not A169) );
 a11327a <=( A170  and  a11326a );
 a11330a <=( A199  and  A166 );
 a11333a <=( (not A203)  and  (not A202) );
 a11334a <=( a11333a  and  a11330a );
 a11335a <=( a11334a  and  a11327a );
 a11338a <=( (not A233)  and  A232 );
 a11341a <=( A236  and  A234 );
 a11342a <=( a11341a  and  a11338a );
 a11345a <=( (not A266)  and  A265 );
 a11348a <=( A268  and  A267 );
 a11349a <=( a11348a  and  a11345a );
 a11350a <=( a11349a  and  a11342a );
 a11354a <=( (not A167)  and  (not A169) );
 a11355a <=( A170  and  a11354a );
 a11358a <=( A199  and  A166 );
 a11361a <=( (not A203)  and  (not A202) );
 a11362a <=( a11361a  and  a11358a );
 a11363a <=( a11362a  and  a11355a );
 a11366a <=( (not A233)  and  A232 );
 a11369a <=( A236  and  A234 );
 a11370a <=( a11369a  and  a11366a );
 a11373a <=( (not A266)  and  A265 );
 a11376a <=( A269  and  A267 );
 a11377a <=( a11376a  and  a11373a );
 a11378a <=( a11377a  and  a11370a );


end x25_7x_behav;
