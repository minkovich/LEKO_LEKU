Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_8x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A107: buffer std_logic
);
end x25_8x;

architecture x25_8x_behav of x25_8x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a168a,a172a,a173a,a174a,a177a,a181a,a182a,a183a,a184a,a187a,a191a,a192a,a193a,a196a,a200a,a201a,a202a,a203a,a204a,a207a,a211a,a212a,a213a,a216a,a220a,a221a,a222a,a223a,a226a,a230a,a231a,a232a,a236a,a237a,a241a,a242a,a243a,a244a,a245a,a246a,a249a,a253a,a254a,a255a,a258a,a262a,a263a,a264a,a265a,a268a,a272a,a273a,a274a,a277a,a281a,a282a,a283a,a284a,a285a,a288a,a292a,a293a,a294a,a297a,a301a,a302a,a303a,a304a,a307a,a311a,a312a,a313a,a317a,a318a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a331a,a335a,a336a,a337a,a340a,a344a,a345a,a346a,a347a,a350a,a354a,a355a,a356a,a359a,a363a,a364a,a365a,a366a,a367a,a370a,a374a,a375a,a376a,a379a,a383a,a384a,a385a,a386a,a389a,a393a,a394a,a395a,a399a,a400a,a404a,a405a,a406a,a407a,a408a,a409a,a412a,a416a,a417a,a418a,a421a,a425a,a426a,a427a,a428a,a431a,a435a,a436a,a437a,a441a,a442a,a446a,a447a,a448a,a449a,a450a,a453a,a457a,a458a,a459a,a462a,a466a,a467a,a468a,a469a,a472a,a476a,a477a,a478a,a482a,a483a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a498a,a501a,a504a,a507a,a510a,a513a,a516a,a519a,a522a,a525a,a529a,a530a,a534a,a535a,a539a,a540a,a544a,a545a,a549a,a550a,a554a,a555a,a559a,a560a,a564a,a565a,a569a,a570a,a574a,a575a,a579a,a580a,a584a,a585a,a589a,a590a,a594a,a595a,a599a,a600a,a604a,a605a,a609a,a610a,a614a,a615a,a619a,a620a,a624a,a625a,a629a,a630a,a634a,a635a,a639a,a640a,a644a,a645a,a649a,a650a,a654a,a655a,a659a,a660a,a664a,a665a,a669a,a670a,a674a,a675a,a679a,a680a,a684a,a685a,a689a,a690a,a694a,a695a,a699a,a700a,a704a,a705a,a709a,a710a,a713a,a716a,a717a,a721a,a722a,a725a,a728a,a729a,a733a,a734a,a737a,a740a,a741a,a745a,a746a,a749a,a752a,a753a,a757a,a758a,a761a,a764a,a765a,a769a,a770a,a773a,a776a,a777a,a780a,a783a,a784a,a787a,a790a,a791a,a794a,a797a,a798a,a801a,a804a,a805a,a808a,a811a,a812a,a815a,a818a,a819a,a822a,a825a,a826a,a829a,a832a,a833a,a836a,a839a,a840a,a843a,a846a,a847a,a850a,a853a,a854a,a857a,a860a,a861a,a864a,a867a,a868a,a871a,a874a,a875a,a878a,a881a,a882a,a885a,a888a,a889a,a892a,a895a,a896a,a899a,a902a,a903a,a906a,a909a,a910a,a913a,a916a,a917a,a920a,a923a,a924a,a927a,a930a,a931a,a934a,a937a,a938a,a941a,a944a,a945a,a948a,a951a,a952a,a955a,a958a,a959a,a962a,a965a,a966a,a969a,a972a,a973a,a976a,a979a,a980a,a983a,a986a,a987a,a990a,a993a,a994a,a997a,a1000a,a1001a,a1004a,a1007a,a1008a,a1011a,a1014a,a1015a,a1018a,a1021a,a1022a,a1025a,a1028a,a1029a,a1032a,a1035a,a1036a,a1039a,a1042a,a1043a,a1046a,a1049a,a1050a,a1053a,a1056a,a1057a,a1060a,a1063a,a1064a,a1067a,a1070a,a1071a,a1074a,a1077a,a1078a,a1081a,a1084a,a1085a,a1088a,a1091a,a1092a,a1095a,a1098a,a1099a,a1102a,a1105a,a1106a,a1109a,a1112a,a1113a,a1116a,a1119a,a1120a,a1123a,a1126a,a1127a,a1130a,a1133a,a1134a,a1137a,a1140a,a1141a,a1144a,a1147a,a1148a,a1151a,a1154a,a1155a,a1158a,a1161a,a1162a,a1165a,a1168a,a1169a,a1172a,a1175a,a1176a,a1179a,a1182a,a1183a,a1186a,a1189a,a1190a,a1193a,a1196a,a1197a,a1200a,a1203a,a1204a,a1207a,a1210a,a1211a,a1214a,a1217a,a1218a,a1221a,a1224a,a1225a,a1228a,a1231a,a1232a,a1235a,a1238a,a1239a,a1242a,a1245a,a1246a,a1249a,a1252a,a1253a,a1256a,a1259a,a1260a,a1263a,a1266a,a1267a,a1270a,a1273a,a1274a,a1277a,a1280a,a1281a,a1284a,a1287a,a1288a,a1291a,a1294a,a1295a,a1298a,a1301a,a1302a,a1305a,a1308a,a1309a,a1312a,a1315a,a1316a,a1319a,a1322a,a1323a,a1326a,a1329a,a1330a,a1333a,a1337a,a1338a,a1339a,a1342a,a1345a,a1346a,a1349a,a1353a,a1354a,a1355a,a1358a,a1361a,a1362a,a1365a,a1369a,a1370a,a1371a,a1374a,a1377a,a1378a,a1381a,a1385a,a1386a,a1387a,a1390a,a1393a,a1394a,a1397a,a1401a,a1402a,a1403a,a1406a,a1409a,a1410a,a1413a,a1417a,a1418a,a1419a,a1422a,a1425a,a1426a,a1429a,a1433a,a1434a,a1435a,a1438a,a1441a,a1442a,a1445a,a1449a,a1450a,a1451a,a1454a,a1457a,a1458a,a1461a,a1465a,a1466a,a1467a,a1470a,a1473a,a1474a,a1477a,a1481a,a1482a,a1483a,a1486a,a1489a,a1490a,a1493a,a1497a,a1498a,a1499a,a1502a,a1505a,a1506a,a1509a,a1513a,a1514a,a1515a,a1518a,a1521a,a1522a,a1525a,a1529a,a1530a,a1531a,a1534a,a1537a,a1538a,a1541a,a1545a,a1546a,a1547a,a1550a,a1553a,a1554a,a1557a,a1561a,a1562a,a1563a,a1566a,a1569a,a1570a,a1573a,a1577a,a1578a,a1579a,a1582a,a1585a,a1586a,a1589a,a1593a,a1594a,a1595a,a1598a,a1601a,a1602a,a1605a,a1609a,a1610a,a1611a,a1614a,a1617a,a1618a,a1621a,a1625a,a1626a,a1627a,a1630a,a1633a,a1634a,a1637a,a1641a,a1642a,a1643a,a1646a,a1649a,a1650a,a1653a,a1657a,a1658a,a1659a,a1662a,a1665a,a1666a,a1669a,a1673a,a1674a,a1675a,a1678a,a1681a,a1682a,a1685a,a1689a,a1690a,a1691a,a1694a,a1697a,a1698a,a1701a,a1705a,a1706a,a1707a,a1710a,a1714a,a1715a,a1716a,a1719a,a1723a,a1724a,a1725a,a1728a,a1732a,a1733a,a1734a,a1737a,a1741a,a1742a,a1743a,a1746a,a1750a,a1751a,a1752a,a1755a,a1759a,a1760a,a1761a,a1764a,a1768a,a1769a,a1770a,a1773a,a1777a,a1778a,a1779a,a1782a,a1786a,a1787a,a1788a,a1791a,a1795a,a1796a,a1797a,a1800a,a1804a,a1805a,a1806a,a1809a,a1813a,a1814a,a1815a,a1818a,a1822a,a1823a,a1824a,a1827a,a1831a,a1832a,a1833a,a1836a,a1840a,a1841a,a1842a,a1845a,a1849a,a1850a,a1851a,a1854a,a1858a,a1859a,a1860a,a1863a,a1867a,a1868a,a1869a,a1872a,a1876a,a1877a,a1878a,a1881a,a1885a,a1886a,a1887a,a1890a,a1894a,a1895a,a1896a,a1899a,a1903a,a1904a,a1905a,a1908a,a1912a,a1913a,a1914a,a1917a,a1921a,a1922a,a1923a,a1926a,a1930a,a1931a,a1932a,a1935a,a1939a,a1940a,a1941a,a1944a,a1948a,a1949a,a1950a,a1953a,a1957a,a1958a,a1959a,a1962a,a1966a,a1967a,a1968a,a1971a,a1975a,a1976a,a1977a,a1980a,a1984a,a1985a,a1986a,a1989a,a1993a,a1994a,a1995a,a1998a,a2002a,a2003a,a2004a,a2007a,a2011a,a2012a,a2013a,a2016a,a2020a,a2021a,a2022a,a2025a,a2029a,a2030a,a2031a,a2034a,a2038a,a2039a,a2040a,a2043a,a2047a,a2048a,a2049a,a2052a,a2056a,a2057a,a2058a,a2061a,a2065a,a2066a,a2067a,a2070a,a2074a,a2075a,a2076a,a2079a,a2083a,a2084a,a2085a,a2088a,a2092a,a2093a,a2094a,a2097a,a2101a,a2102a,a2103a,a2106a,a2110a,a2111a,a2112a,a2115a,a2119a,a2120a,a2121a,a2124a,a2128a,a2129a,a2130a,a2133a,a2137a,a2138a,a2139a,a2142a,a2146a,a2147a,a2148a,a2151a,a2155a,a2156a,a2157a,a2160a,a2164a,a2165a,a2166a,a2169a,a2173a,a2174a,a2175a,a2178a,a2182a,a2183a,a2184a,a2187a,a2191a,a2192a,a2193a,a2196a,a2200a,a2201a,a2202a,a2205a,a2209a,a2210a,a2211a,a2214a,a2218a,a2219a,a2220a,a2223a,a2227a,a2228a,a2229a,a2232a,a2236a,a2237a,a2238a,a2241a,a2245a,a2246a,a2247a,a2250a,a2254a,a2255a,a2256a,a2259a,a2263a,a2264a,a2265a,a2268a,a2272a,a2273a,a2274a,a2277a,a2281a,a2282a,a2283a,a2286a,a2290a,a2291a,a2292a,a2295a,a2299a,a2300a,a2301a,a2304a,a2308a,a2309a,a2310a,a2313a,a2317a,a2318a,a2319a,a2322a,a2326a,a2327a,a2328a,a2331a,a2335a,a2336a,a2337a,a2340a,a2344a,a2345a,a2346a,a2349a,a2353a,a2354a,a2355a,a2358a,a2362a,a2363a,a2364a,a2368a,a2369a,a2373a,a2374a,a2375a,a2378a,a2382a,a2383a,a2384a,a2388a,a2389a,a2393a,a2394a,a2395a,a2398a,a2402a,a2403a,a2404a,a2408a,a2409a,a2413a,a2414a,a2415a,a2418a,a2422a,a2423a,a2424a,a2428a,a2429a,a2433a,a2434a,a2435a,a2438a,a2442a,a2443a,a2444a,a2448a,a2449a,a2453a,a2454a,a2455a,a2458a,a2462a,a2463a,a2464a,a2468a,a2469a,a2473a,a2474a,a2475a,a2478a,a2482a,a2483a,a2484a,a2488a,a2489a,a2493a,a2494a,a2495a,a2498a,a2502a,a2503a,a2504a,a2508a,a2509a,a2513a,a2514a,a2515a,a2518a,a2522a,a2523a,a2524a,a2528a,a2529a,a2533a,a2534a,a2535a,a2538a,a2542a,a2543a,a2544a,a2548a,a2549a,a2553a,a2554a,a2555a,a2558a,a2562a,a2563a,a2564a,a2568a,a2569a,a2573a,a2574a,a2575a,a2578a,a2582a,a2583a,a2584a,a2588a,a2589a,a2593a,a2594a,a2595a,a2598a,a2602a,a2603a,a2604a,a2608a,a2609a,a2613a,a2614a,a2615a,a2618a,a2622a,a2623a,a2624a,a2628a,a2629a,a2633a,a2634a,a2635a,a2638a,a2642a,a2643a,a2644a,a2648a,a2649a,a2653a,a2654a,a2655a,a2658a,a2662a,a2663a,a2664a,a2668a,a2669a,a2673a,a2674a,a2675a,a2678a,a2682a,a2683a,a2684a,a2688a,a2689a,a2693a,a2694a,a2695a,a2698a,a2702a,a2703a,a2704a,a2708a,a2709a,a2713a,a2714a,a2715a,a2718a,a2722a,a2723a,a2724a,a2728a,a2729a,a2733a,a2734a,a2735a,a2738a,a2742a,a2743a,a2744a,a2748a,a2749a,a2753a,a2754a,a2755a,a2758a,a2762a,a2763a,a2764a,a2768a,a2769a,a2773a,a2774a,a2775a,a2778a,a2782a,a2783a,a2784a,a2788a,a2789a,a2793a,a2794a,a2795a,a2798a,a2802a,a2803a,a2804a,a2808a,a2809a,a2813a,a2814a,a2815a,a2818a,a2822a,a2823a,a2824a,a2828a,a2829a,a2833a,a2834a,a2835a,a2839a,a2840a,a2844a,a2845a,a2846a,a2850a,a2851a,a2855a,a2856a,a2857a,a2861a,a2862a,a2866a,a2867a,a2868a,a2872a,a2873a,a2877a,a2878a,a2879a,a2883a,a2884a,a2888a,a2889a,a2890a,a2894a,a2895a,a2899a,a2900a,a2901a,a2905a,a2906a,a2910a,a2911a,a2912a,a2916a,a2917a,a2921a,a2922a,a2923a,a2927a,a2928a,a2932a,a2933a,a2934a,a2938a,a2939a,a2943a,a2944a,a2945a,a2949a,a2950a,a2954a,a2955a,a2956a,a2960a,a2961a,a2965a,a2966a,a2967a,a2971a,a2972a,a2976a,a2977a,a2978a,a2982a,a2983a,a2987a,a2988a,a2989a,a2993a,a2994a,a2998a,a2999a,a3000a,a3004a,a3005a,a3009a,a3010a,a3011a,a3015a,a3016a,a3020a,a3021a,a3022a,a3026a,a3027a,a3031a,a3032a,a3033a,a3037a,a3038a,a3042a,a3043a,a3044a,a3048a,a3049a,a3053a,a3054a,a3055a,a3059a,a3060a,a3064a,a3065a,a3066a,a3070a,a3071a,a3075a,a3076a,a3077a,a3081a,a3082a,a3086a,a3087a,a3088a,a3092a,a3093a,a3097a,a3098a,a3099a: std_logic;
begin

A107 <=( a493a ) or ( a328a );
 a1a <=( a3099a  and  a3088a );
 a2a <=( a3077a  and  a3066a );
 a3a <=( a3055a  and  a3044a );
 a4a <=( a3033a  and  a3022a );
 a5a <=( a3011a  and  a3000a );
 a6a <=( a2989a  and  a2978a );
 a7a <=( a2967a  and  a2956a );
 a8a <=( a2945a  and  a2934a );
 a9a <=( a2923a  and  a2912a );
 a10a <=( a2901a  and  a2890a );
 a11a <=( a2879a  and  a2868a );
 a12a <=( a2857a  and  a2846a );
 a13a <=( a2835a  and  a2824a );
 a14a <=( a2815a  and  a2804a );
 a15a <=( a2795a  and  a2784a );
 a16a <=( a2775a  and  a2764a );
 a17a <=( a2755a  and  a2744a );
 a18a <=( a2735a  and  a2724a );
 a19a <=( a2715a  and  a2704a );
 a20a <=( a2695a  and  a2684a );
 a21a <=( a2675a  and  a2664a );
 a22a <=( a2655a  and  a2644a );
 a23a <=( a2635a  and  a2624a );
 a24a <=( a2615a  and  a2604a );
 a25a <=( a2595a  and  a2584a );
 a26a <=( a2575a  and  a2564a );
 a27a <=( a2555a  and  a2544a );
 a28a <=( a2535a  and  a2524a );
 a29a <=( a2515a  and  a2504a );
 a30a <=( a2495a  and  a2484a );
 a31a <=( a2475a  and  a2464a );
 a32a <=( a2455a  and  a2444a );
 a33a <=( a2435a  and  a2424a );
 a34a <=( a2415a  and  a2404a );
 a35a <=( a2395a  and  a2384a );
 a36a <=( a2375a  and  a2364a );
 a37a <=( a2355a  and  a2346a );
 a38a <=( a2337a  and  a2328a );
 a39a <=( a2319a  and  a2310a );
 a40a <=( a2301a  and  a2292a );
 a41a <=( a2283a  and  a2274a );
 a42a <=( a2265a  and  a2256a );
 a43a <=( a2247a  and  a2238a );
 a44a <=( a2229a  and  a2220a );
 a45a <=( a2211a  and  a2202a );
 a46a <=( a2193a  and  a2184a );
 a47a <=( a2175a  and  a2166a );
 a48a <=( a2157a  and  a2148a );
 a49a <=( a2139a  and  a2130a );
 a50a <=( a2121a  and  a2112a );
 a51a <=( a2103a  and  a2094a );
 a52a <=( a2085a  and  a2076a );
 a53a <=( a2067a  and  a2058a );
 a54a <=( a2049a  and  a2040a );
 a55a <=( a2031a  and  a2022a );
 a56a <=( a2013a  and  a2004a );
 a57a <=( a1995a  and  a1986a );
 a58a <=( a1977a  and  a1968a );
 a59a <=( a1959a  and  a1950a );
 a60a <=( a1941a  and  a1932a );
 a61a <=( a1923a  and  a1914a );
 a62a <=( a1905a  and  a1896a );
 a63a <=( a1887a  and  a1878a );
 a64a <=( a1869a  and  a1860a );
 a65a <=( a1851a  and  a1842a );
 a66a <=( a1833a  and  a1824a );
 a67a <=( a1815a  and  a1806a );
 a68a <=( a1797a  and  a1788a );
 a69a <=( a1779a  and  a1770a );
 a70a <=( a1761a  and  a1752a );
 a71a <=( a1743a  and  a1734a );
 a72a <=( a1725a  and  a1716a );
 a73a <=( a1707a  and  a1698a );
 a74a <=( a1691a  and  a1682a );
 a75a <=( a1675a  and  a1666a );
 a76a <=( a1659a  and  a1650a );
 a77a <=( a1643a  and  a1634a );
 a78a <=( a1627a  and  a1618a );
 a79a <=( a1611a  and  a1602a );
 a80a <=( a1595a  and  a1586a );
 a81a <=( a1579a  and  a1570a );
 a82a <=( a1563a  and  a1554a );
 a83a <=( a1547a  and  a1538a );
 a84a <=( a1531a  and  a1522a );
 a85a <=( a1515a  and  a1506a );
 a86a <=( a1499a  and  a1490a );
 a87a <=( a1483a  and  a1474a );
 a88a <=( a1467a  and  a1458a );
 a89a <=( a1451a  and  a1442a );
 a90a <=( a1435a  and  a1426a );
 a91a <=( a1419a  and  a1410a );
 a92a <=( a1403a  and  a1394a );
 a93a <=( a1387a  and  a1378a );
 a94a <=( a1371a  and  a1362a );
 a95a <=( a1355a  and  a1346a );
 a96a <=( a1339a  and  a1330a );
 a97a <=( a1323a  and  a1316a );
 a98a <=( a1309a  and  a1302a );
 a99a <=( a1295a  and  a1288a );
 a100a <=( a1281a  and  a1274a );
 a101a <=( a1267a  and  a1260a );
 a102a <=( a1253a  and  a1246a );
 a103a <=( a1239a  and  a1232a );
 a104a <=( a1225a  and  a1218a );
 a105a <=( a1211a  and  a1204a );
 a106a <=( a1197a  and  a1190a );
 a107a <=( a1183a  and  a1176a );
 a108a <=( a1169a  and  a1162a );
 a109a <=( a1155a  and  a1148a );
 a110a <=( a1141a  and  a1134a );
 a111a <=( a1127a  and  a1120a );
 a112a <=( a1113a  and  a1106a );
 a113a <=( a1099a  and  a1092a );
 a114a <=( a1085a  and  a1078a );
 a115a <=( a1071a  and  a1064a );
 a116a <=( a1057a  and  a1050a );
 a117a <=( a1043a  and  a1036a );
 a118a <=( a1029a  and  a1022a );
 a119a <=( a1015a  and  a1008a );
 a120a <=( a1001a  and  a994a );
 a121a <=( a987a  and  a980a );
 a122a <=( a973a  and  a966a );
 a123a <=( a959a  and  a952a );
 a124a <=( a945a  and  a938a );
 a125a <=( a931a  and  a924a );
 a126a <=( a917a  and  a910a );
 a127a <=( a903a  and  a896a );
 a128a <=( a889a  and  a882a );
 a129a <=( a875a  and  a868a );
 a130a <=( a861a  and  a854a );
 a131a <=( a847a  and  a840a );
 a132a <=( a833a  and  a826a );
 a133a <=( a819a  and  a812a );
 a134a <=( a805a  and  a798a );
 a135a <=( a791a  and  a784a );
 a136a <=( a777a  and  a770a );
 a137a <=( a765a  and  a758a );
 a138a <=( a753a  and  a746a );
 a139a <=( a741a  and  a734a );
 a140a <=( a729a  and  a722a );
 a141a <=( a717a  and  a710a );
 a142a <=( a705a  and  a700a );
 a143a <=( a695a  and  a690a );
 a144a <=( a685a  and  a680a );
 a145a <=( a675a  and  a670a );
 a146a <=( a665a  and  a660a );
 a147a <=( a655a  and  a650a );
 a148a <=( a645a  and  a640a );
 a149a <=( a635a  and  a630a );
 a150a <=( a625a  and  a620a );
 a151a <=( a615a  and  a610a );
 a152a <=( a605a  and  a600a );
 a153a <=( a595a  and  a590a );
 a154a <=( a585a  and  a580a );
 a155a <=( a575a  and  a570a );
 a156a <=( a565a  and  a560a );
 a157a <=( a555a  and  a550a );
 a158a <=( a545a  and  a540a );
 a159a <=( a535a  and  a530a );
 a160a <=( a525a  and  a522a );
 a161a <=( a519a  and  a516a );
 a162a <=( a513a  and  a510a );
 a163a <=( a507a  and  a504a );
 a164a <=( a501a  and  a498a );
 a165a <=( A266  and  (not A265) );
 a168a <=( a164a ) or ( a165a );
 a172a <=( a161a ) or ( a162a );
 a173a <=( a163a ) or ( a172a );
 a174a <=( a173a ) or ( a168a );
 a177a <=( a159a ) or ( a160a );
 a181a <=( a156a ) or ( a157a );
 a182a <=( a158a ) or ( a181a );
 a183a <=( a182a ) or ( a177a );
 a184a <=( a183a ) or ( a174a );
 a187a <=( a154a ) or ( a155a );
 a191a <=( a151a ) or ( a152a );
 a192a <=( a153a ) or ( a191a );
 a193a <=( a192a ) or ( a187a );
 a196a <=( a149a ) or ( a150a );
 a200a <=( a146a ) or ( a147a );
 a201a <=( a148a ) or ( a200a );
 a202a <=( a201a ) or ( a196a );
 a203a <=( a202a ) or ( a193a );
 a204a <=( a203a ) or ( a184a );
 a207a <=( a144a ) or ( a145a );
 a211a <=( a141a ) or ( a142a );
 a212a <=( a143a ) or ( a211a );
 a213a <=( a212a ) or ( a207a );
 a216a <=( a139a ) or ( a140a );
 a220a <=( a136a ) or ( a137a );
 a221a <=( a138a ) or ( a220a );
 a222a <=( a221a ) or ( a216a );
 a223a <=( a222a ) or ( a213a );
 a226a <=( a134a ) or ( a135a );
 a230a <=( a131a ) or ( a132a );
 a231a <=( a133a ) or ( a230a );
 a232a <=( a231a ) or ( a226a );
 a236a <=( a128a ) or ( a129a );
 a237a <=( a130a ) or ( a236a );
 a241a <=( a125a ) or ( a126a );
 a242a <=( a127a ) or ( a241a );
 a243a <=( a242a ) or ( a237a );
 a244a <=( a243a ) or ( a232a );
 a245a <=( a244a ) or ( a223a );
 a246a <=( a245a ) or ( a204a );
 a249a <=( a123a ) or ( a124a );
 a253a <=( a120a ) or ( a121a );
 a254a <=( a122a ) or ( a253a );
 a255a <=( a254a ) or ( a249a );
 a258a <=( a118a ) or ( a119a );
 a262a <=( a115a ) or ( a116a );
 a263a <=( a117a ) or ( a262a );
 a264a <=( a263a ) or ( a258a );
 a265a <=( a264a ) or ( a255a );
 a268a <=( a113a ) or ( a114a );
 a272a <=( a110a ) or ( a111a );
 a273a <=( a112a ) or ( a272a );
 a274a <=( a273a ) or ( a268a );
 a277a <=( a108a ) or ( a109a );
 a281a <=( a105a ) or ( a106a );
 a282a <=( a107a ) or ( a281a );
 a283a <=( a282a ) or ( a277a );
 a284a <=( a283a ) or ( a274a );
 a285a <=( a284a ) or ( a265a );
 a288a <=( a103a ) or ( a104a );
 a292a <=( a100a ) or ( a101a );
 a293a <=( a102a ) or ( a292a );
 a294a <=( a293a ) or ( a288a );
 a297a <=( a98a ) or ( a99a );
 a301a <=( a95a ) or ( a96a );
 a302a <=( a97a ) or ( a301a );
 a303a <=( a302a ) or ( a297a );
 a304a <=( a303a ) or ( a294a );
 a307a <=( a93a ) or ( a94a );
 a311a <=( a90a ) or ( a91a );
 a312a <=( a92a ) or ( a311a );
 a313a <=( a312a ) or ( a307a );
 a317a <=( a87a ) or ( a88a );
 a318a <=( a89a ) or ( a317a );
 a322a <=( a84a ) or ( a85a );
 a323a <=( a86a ) or ( a322a );
 a324a <=( a323a ) or ( a318a );
 a325a <=( a324a ) or ( a313a );
 a326a <=( a325a ) or ( a304a );
 a327a <=( a326a ) or ( a285a );
 a328a <=( a327a ) or ( a246a );
 a331a <=( a82a ) or ( a83a );
 a335a <=( a79a ) or ( a80a );
 a336a <=( a81a ) or ( a335a );
 a337a <=( a336a ) or ( a331a );
 a340a <=( a77a ) or ( a78a );
 a344a <=( a74a ) or ( a75a );
 a345a <=( a76a ) or ( a344a );
 a346a <=( a345a ) or ( a340a );
 a347a <=( a346a ) or ( a337a );
 a350a <=( a72a ) or ( a73a );
 a354a <=( a69a ) or ( a70a );
 a355a <=( a71a ) or ( a354a );
 a356a <=( a355a ) or ( a350a );
 a359a <=( a67a ) or ( a68a );
 a363a <=( a64a ) or ( a65a );
 a364a <=( a66a ) or ( a363a );
 a365a <=( a364a ) or ( a359a );
 a366a <=( a365a ) or ( a356a );
 a367a <=( a366a ) or ( a347a );
 a370a <=( a62a ) or ( a63a );
 a374a <=( a59a ) or ( a60a );
 a375a <=( a61a ) or ( a374a );
 a376a <=( a375a ) or ( a370a );
 a379a <=( a57a ) or ( a58a );
 a383a <=( a54a ) or ( a55a );
 a384a <=( a56a ) or ( a383a );
 a385a <=( a384a ) or ( a379a );
 a386a <=( a385a ) or ( a376a );
 a389a <=( a52a ) or ( a53a );
 a393a <=( a49a ) or ( a50a );
 a394a <=( a51a ) or ( a393a );
 a395a <=( a394a ) or ( a389a );
 a399a <=( a46a ) or ( a47a );
 a400a <=( a48a ) or ( a399a );
 a404a <=( a43a ) or ( a44a );
 a405a <=( a45a ) or ( a404a );
 a406a <=( a405a ) or ( a400a );
 a407a <=( a406a ) or ( a395a );
 a408a <=( a407a ) or ( a386a );
 a409a <=( a408a ) or ( a367a );
 a412a <=( a41a ) or ( a42a );
 a416a <=( a38a ) or ( a39a );
 a417a <=( a40a ) or ( a416a );
 a418a <=( a417a ) or ( a412a );
 a421a <=( a36a ) or ( a37a );
 a425a <=( a33a ) or ( a34a );
 a426a <=( a35a ) or ( a425a );
 a427a <=( a426a ) or ( a421a );
 a428a <=( a427a ) or ( a418a );
 a431a <=( a31a ) or ( a32a );
 a435a <=( a28a ) or ( a29a );
 a436a <=( a30a ) or ( a435a );
 a437a <=( a436a ) or ( a431a );
 a441a <=( a25a ) or ( a26a );
 a442a <=( a27a ) or ( a441a );
 a446a <=( a22a ) or ( a23a );
 a447a <=( a24a ) or ( a446a );
 a448a <=( a447a ) or ( a442a );
 a449a <=( a448a ) or ( a437a );
 a450a <=( a449a ) or ( a428a );
 a453a <=( a20a ) or ( a21a );
 a457a <=( a17a ) or ( a18a );
 a458a <=( a19a ) or ( a457a );
 a459a <=( a458a ) or ( a453a );
 a462a <=( a15a ) or ( a16a );
 a466a <=( a12a ) or ( a13a );
 a467a <=( a14a ) or ( a466a );
 a468a <=( a467a ) or ( a462a );
 a469a <=( a468a ) or ( a459a );
 a472a <=( a10a ) or ( a11a );
 a476a <=( a7a ) or ( a8a );
 a477a <=( a9a ) or ( a476a );
 a478a <=( a477a ) or ( a472a );
 a482a <=( a4a ) or ( a5a );
 a483a <=( a6a ) or ( a482a );
 a487a <=( a1a ) or ( a2a );
 a488a <=( a3a ) or ( a487a );
 a489a <=( a488a ) or ( a483a );
 a490a <=( a489a ) or ( a478a );
 a491a <=( a490a ) or ( a469a );
 a492a <=( a491a ) or ( a450a );
 a493a <=( a492a ) or ( a409a );
 a498a <=( (not A266)  and  A265 );
 a501a <=( A268  and  A267 );
 a504a <=( (not A266)  and  A265 );
 a507a <=( A269  and  A267 );
 a510a <=( A200  and  (not A199) );
 a513a <=( A233  and  (not A232) );
 a516a <=( A166  and  A168 );
 a519a <=( A233  and  (not A232) );
 a522a <=( A167  and  A168 );
 a525a <=( A233  and  (not A232) );
 a529a <=( A232  and  A200 );
 a530a <=( (not A199)  and  a529a );
 a534a <=( A235  and  A234 );
 a535a <=( (not A233)  and  a534a );
 a539a <=( A232  and  A200 );
 a540a <=( (not A199)  and  a539a );
 a544a <=( A236  and  A234 );
 a545a <=( (not A233)  and  a544a );
 a549a <=( A201  and  (not A200) );
 a550a <=( A199  and  a549a );
 a554a <=( A233  and  (not A232) );
 a555a <=( A202  and  a554a );
 a559a <=( A201  and  (not A200) );
 a560a <=( A199  and  a559a );
 a564a <=( A233  and  (not A232) );
 a565a <=( A203  and  a564a );
 a569a <=( A232  and  A166 );
 a570a <=( A168  and  a569a );
 a574a <=( A235  and  A234 );
 a575a <=( (not A233)  and  a574a );
 a579a <=( A232  and  A166 );
 a580a <=( A168  and  a579a );
 a584a <=( A236  and  A234 );
 a585a <=( (not A233)  and  a584a );
 a589a <=( A199  and  A166 );
 a590a <=( A168  and  a589a );
 a594a <=( A299  and  (not A298) );
 a595a <=( A200  and  a594a );
 a599a <=( (not A200)  and  A166 );
 a600a <=( A168  and  a599a );
 a604a <=( A299  and  (not A298) );
 a605a <=( (not A201)  and  a604a );
 a609a <=( (not A199)  and  A166 );
 a610a <=( A168  and  a609a );
 a614a <=( A299  and  (not A298) );
 a615a <=( (not A200)  and  a614a );
 a619a <=( A232  and  A167 );
 a620a <=( A168  and  a619a );
 a624a <=( A235  and  A234 );
 a625a <=( (not A233)  and  a624a );
 a629a <=( A232  and  A167 );
 a630a <=( A168  and  a629a );
 a634a <=( A236  and  A234 );
 a635a <=( (not A233)  and  a634a );
 a639a <=( A199  and  A167 );
 a640a <=( A168  and  a639a );
 a644a <=( A299  and  (not A298) );
 a645a <=( A200  and  a644a );
 a649a <=( (not A200)  and  A167 );
 a650a <=( A168  and  a649a );
 a654a <=( A299  and  (not A298) );
 a655a <=( (not A201)  and  a654a );
 a659a <=( (not A199)  and  A167 );
 a660a <=( A168  and  a659a );
 a664a <=( A299  and  (not A298) );
 a665a <=( (not A200)  and  a664a );
 a669a <=( A167  and  A169 );
 a670a <=( (not A170)  and  a669a );
 a674a <=( A233  and  (not A232) );
 a675a <=( A166  and  a674a );
 a679a <=( (not A167)  and  A169 );
 a680a <=( (not A170)  and  a679a );
 a684a <=( A233  and  (not A232) );
 a685a <=( (not A166)  and  a684a );
 a689a <=( A167  and  (not A169) );
 a690a <=( A170  and  a689a );
 a694a <=( A233  and  (not A232) );
 a695a <=( (not A166)  and  a694a );
 a699a <=( (not A167)  and  (not A169) );
 a700a <=( A170  and  a699a );
 a704a <=( A233  and  (not A232) );
 a705a <=( A166  and  a704a );
 a709a <=( (not A200)  and  A166 );
 a710a <=( A168  and  a709a );
 a713a <=( (not A203)  and  (not A202) );
 a716a <=( A299  and  (not A298) );
 a717a <=( a716a  and  a713a );
 a721a <=( (not A200)  and  A167 );
 a722a <=( A168  and  a721a );
 a725a <=( (not A203)  and  (not A202) );
 a728a <=( A299  and  (not A298) );
 a729a <=( a728a  and  a725a );
 a733a <=( (not A166)  and  (not A167) );
 a734a <=( A170  and  a733a );
 a737a <=( A200  and  (not A199) );
 a740a <=( A299  and  (not A298) );
 a741a <=( a740a  and  a737a );
 a745a <=( (not A168)  and  A169 );
 a746a <=( A170  and  a745a );
 a749a <=( A200  and  (not A199) );
 a752a <=( A299  and  (not A298) );
 a753a <=( a752a  and  a749a );
 a757a <=( (not A166)  and  (not A167) );
 a758a <=( (not A169)  and  a757a );
 a761a <=( A200  and  (not A199) );
 a764a <=( A299  and  (not A298) );
 a765a <=( a764a  and  a761a );
 a769a <=( (not A168)  and  (not A169) );
 a770a <=( (not A170)  and  a769a );
 a773a <=( A200  and  (not A199) );
 a776a <=( A299  and  (not A298) );
 a777a <=( a776a  and  a773a );
 a780a <=( (not A200)  and  A199 );
 a783a <=( A202  and  A201 );
 a784a <=( a783a  and  a780a );
 a787a <=( (not A233)  and  A232 );
 a790a <=( A235  and  A234 );
 a791a <=( a790a  and  a787a );
 a794a <=( (not A200)  and  A199 );
 a797a <=( A202  and  A201 );
 a798a <=( a797a  and  a794a );
 a801a <=( (not A233)  and  A232 );
 a804a <=( A236  and  A234 );
 a805a <=( a804a  and  a801a );
 a808a <=( (not A200)  and  A199 );
 a811a <=( A203  and  A201 );
 a812a <=( a811a  and  a808a );
 a815a <=( (not A233)  and  A232 );
 a818a <=( A235  and  A234 );
 a819a <=( a818a  and  a815a );
 a822a <=( (not A200)  and  A199 );
 a825a <=( A203  and  A201 );
 a826a <=( a825a  and  a822a );
 a829a <=( (not A233)  and  A232 );
 a832a <=( A236  and  A234 );
 a833a <=( a832a  and  a829a );
 a836a <=( A166  and  A168 );
 a839a <=( A200  and  A199 );
 a840a <=( a839a  and  a836a );
 a843a <=( (not A299)  and  A298 );
 a846a <=( A301  and  A300 );
 a847a <=( a846a  and  a843a );
 a850a <=( A166  and  A168 );
 a853a <=( A200  and  A199 );
 a854a <=( a853a  and  a850a );
 a857a <=( (not A299)  and  A298 );
 a860a <=( A302  and  A300 );
 a861a <=( a860a  and  a857a );
 a864a <=( A166  and  A168 );
 a867a <=( (not A201)  and  (not A200) );
 a868a <=( a867a  and  a864a );
 a871a <=( (not A299)  and  A298 );
 a874a <=( A301  and  A300 );
 a875a <=( a874a  and  a871a );
 a878a <=( A166  and  A168 );
 a881a <=( (not A201)  and  (not A200) );
 a882a <=( a881a  and  a878a );
 a885a <=( (not A299)  and  A298 );
 a888a <=( A302  and  A300 );
 a889a <=( a888a  and  a885a );
 a892a <=( A166  and  A168 );
 a895a <=( (not A200)  and  (not A199) );
 a896a <=( a895a  and  a892a );
 a899a <=( (not A299)  and  A298 );
 a902a <=( A301  and  A300 );
 a903a <=( a902a  and  a899a );
 a906a <=( A166  and  A168 );
 a909a <=( (not A200)  and  (not A199) );
 a910a <=( a909a  and  a906a );
 a913a <=( (not A299)  and  A298 );
 a916a <=( A302  and  A300 );
 a917a <=( a916a  and  a913a );
 a920a <=( A167  and  A168 );
 a923a <=( A200  and  A199 );
 a924a <=( a923a  and  a920a );
 a927a <=( (not A299)  and  A298 );
 a930a <=( A301  and  A300 );
 a931a <=( a930a  and  a927a );
 a934a <=( A167  and  A168 );
 a937a <=( A200  and  A199 );
 a938a <=( a937a  and  a934a );
 a941a <=( (not A299)  and  A298 );
 a944a <=( A302  and  A300 );
 a945a <=( a944a  and  a941a );
 a948a <=( A167  and  A168 );
 a951a <=( (not A201)  and  (not A200) );
 a952a <=( a951a  and  a948a );
 a955a <=( (not A299)  and  A298 );
 a958a <=( A301  and  A300 );
 a959a <=( a958a  and  a955a );
 a962a <=( A167  and  A168 );
 a965a <=( (not A201)  and  (not A200) );
 a966a <=( a965a  and  a962a );
 a969a <=( (not A299)  and  A298 );
 a972a <=( A302  and  A300 );
 a973a <=( a972a  and  a969a );
 a976a <=( A167  and  A168 );
 a979a <=( (not A200)  and  (not A199) );
 a980a <=( a979a  and  a976a );
 a983a <=( (not A299)  and  A298 );
 a986a <=( A301  and  A300 );
 a987a <=( a986a  and  a983a );
 a990a <=( A167  and  A168 );
 a993a <=( (not A200)  and  (not A199) );
 a994a <=( a993a  and  a990a );
 a997a <=( (not A299)  and  A298 );
 a1000a <=( A302  and  A300 );
 a1001a <=( a1000a  and  a997a );
 a1004a <=( (not A168)  and  A169 );
 a1007a <=( (not A166)  and  A167 );
 a1008a <=( a1007a  and  a1004a );
 a1011a <=( A200  and  (not A199) );
 a1014a <=( A299  and  (not A298) );
 a1015a <=( a1014a  and  a1011a );
 a1018a <=( (not A168)  and  A169 );
 a1021a <=( A166  and  (not A167) );
 a1022a <=( a1021a  and  a1018a );
 a1025a <=( A200  and  (not A199) );
 a1028a <=( A299  and  (not A298) );
 a1029a <=( a1028a  and  a1025a );
 a1032a <=( A169  and  (not A170) );
 a1035a <=( A166  and  A167 );
 a1036a <=( a1035a  and  a1032a );
 a1039a <=( (not A233)  and  A232 );
 a1042a <=( A235  and  A234 );
 a1043a <=( a1042a  and  a1039a );
 a1046a <=( A169  and  (not A170) );
 a1049a <=( A166  and  A167 );
 a1050a <=( a1049a  and  a1046a );
 a1053a <=( (not A233)  and  A232 );
 a1056a <=( A236  and  A234 );
 a1057a <=( a1056a  and  a1053a );
 a1060a <=( A169  and  (not A170) );
 a1063a <=( A166  and  A167 );
 a1064a <=( a1063a  and  a1060a );
 a1067a <=( A200  and  A199 );
 a1070a <=( A299  and  (not A298) );
 a1071a <=( a1070a  and  a1067a );
 a1074a <=( A169  and  (not A170) );
 a1077a <=( A166  and  A167 );
 a1078a <=( a1077a  and  a1074a );
 a1081a <=( (not A201)  and  (not A200) );
 a1084a <=( A299  and  (not A298) );
 a1085a <=( a1084a  and  a1081a );
 a1088a <=( A169  and  (not A170) );
 a1091a <=( A166  and  A167 );
 a1092a <=( a1091a  and  a1088a );
 a1095a <=( (not A200)  and  (not A199) );
 a1098a <=( A299  and  (not A298) );
 a1099a <=( a1098a  and  a1095a );
 a1102a <=( A169  and  (not A170) );
 a1105a <=( (not A166)  and  (not A167) );
 a1106a <=( a1105a  and  a1102a );
 a1109a <=( (not A233)  and  A232 );
 a1112a <=( A235  and  A234 );
 a1113a <=( a1112a  and  a1109a );
 a1116a <=( A169  and  (not A170) );
 a1119a <=( (not A166)  and  (not A167) );
 a1120a <=( a1119a  and  a1116a );
 a1123a <=( (not A233)  and  A232 );
 a1126a <=( A236  and  A234 );
 a1127a <=( a1126a  and  a1123a );
 a1130a <=( A169  and  (not A170) );
 a1133a <=( (not A166)  and  (not A167) );
 a1134a <=( a1133a  and  a1130a );
 a1137a <=( A200  and  A199 );
 a1140a <=( A299  and  (not A298) );
 a1141a <=( a1140a  and  a1137a );
 a1144a <=( A169  and  (not A170) );
 a1147a <=( (not A166)  and  (not A167) );
 a1148a <=( a1147a  and  a1144a );
 a1151a <=( (not A201)  and  (not A200) );
 a1154a <=( A299  and  (not A298) );
 a1155a <=( a1154a  and  a1151a );
 a1158a <=( A169  and  (not A170) );
 a1161a <=( (not A166)  and  (not A167) );
 a1162a <=( a1161a  and  a1158a );
 a1165a <=( (not A200)  and  (not A199) );
 a1168a <=( A299  and  (not A298) );
 a1169a <=( a1168a  and  a1165a );
 a1172a <=( (not A168)  and  (not A169) );
 a1175a <=( A166  and  A167 );
 a1176a <=( a1175a  and  a1172a );
 a1179a <=( A200  and  (not A199) );
 a1182a <=( A299  and  (not A298) );
 a1183a <=( a1182a  and  a1179a );
 a1186a <=( (not A169)  and  A170 );
 a1189a <=( (not A166)  and  A167 );
 a1190a <=( a1189a  and  a1186a );
 a1193a <=( (not A233)  and  A232 );
 a1196a <=( A235  and  A234 );
 a1197a <=( a1196a  and  a1193a );
 a1200a <=( (not A169)  and  A170 );
 a1203a <=( (not A166)  and  A167 );
 a1204a <=( a1203a  and  a1200a );
 a1207a <=( (not A233)  and  A232 );
 a1210a <=( A236  and  A234 );
 a1211a <=( a1210a  and  a1207a );
 a1214a <=( (not A169)  and  A170 );
 a1217a <=( (not A166)  and  A167 );
 a1218a <=( a1217a  and  a1214a );
 a1221a <=( A200  and  A199 );
 a1224a <=( A299  and  (not A298) );
 a1225a <=( a1224a  and  a1221a );
 a1228a <=( (not A169)  and  A170 );
 a1231a <=( (not A166)  and  A167 );
 a1232a <=( a1231a  and  a1228a );
 a1235a <=( (not A201)  and  (not A200) );
 a1238a <=( A299  and  (not A298) );
 a1239a <=( a1238a  and  a1235a );
 a1242a <=( (not A169)  and  A170 );
 a1245a <=( (not A166)  and  A167 );
 a1246a <=( a1245a  and  a1242a );
 a1249a <=( (not A200)  and  (not A199) );
 a1252a <=( A299  and  (not A298) );
 a1253a <=( a1252a  and  a1249a );
 a1256a <=( (not A169)  and  A170 );
 a1259a <=( A166  and  (not A167) );
 a1260a <=( a1259a  and  a1256a );
 a1263a <=( (not A233)  and  A232 );
 a1266a <=( A235  and  A234 );
 a1267a <=( a1266a  and  a1263a );
 a1270a <=( (not A169)  and  A170 );
 a1273a <=( A166  and  (not A167) );
 a1274a <=( a1273a  and  a1270a );
 a1277a <=( (not A233)  and  A232 );
 a1280a <=( A236  and  A234 );
 a1281a <=( a1280a  and  a1277a );
 a1284a <=( (not A169)  and  A170 );
 a1287a <=( A166  and  (not A167) );
 a1288a <=( a1287a  and  a1284a );
 a1291a <=( A200  and  A199 );
 a1294a <=( A299  and  (not A298) );
 a1295a <=( a1294a  and  a1291a );
 a1298a <=( (not A169)  and  A170 );
 a1301a <=( A166  and  (not A167) );
 a1302a <=( a1301a  and  a1298a );
 a1305a <=( (not A201)  and  (not A200) );
 a1308a <=( A299  and  (not A298) );
 a1309a <=( a1308a  and  a1305a );
 a1312a <=( (not A169)  and  A170 );
 a1315a <=( A166  and  (not A167) );
 a1316a <=( a1315a  and  a1312a );
 a1319a <=( (not A200)  and  (not A199) );
 a1322a <=( A299  and  (not A298) );
 a1323a <=( a1322a  and  a1319a );
 a1326a <=( A166  and  A168 );
 a1329a <=( (not A202)  and  (not A200) );
 a1330a <=( a1329a  and  a1326a );
 a1333a <=( A298  and  (not A203) );
 a1337a <=( A301  and  A300 );
 a1338a <=( (not A299)  and  a1337a );
 a1339a <=( a1338a  and  a1333a );
 a1342a <=( A166  and  A168 );
 a1345a <=( (not A202)  and  (not A200) );
 a1346a <=( a1345a  and  a1342a );
 a1349a <=( A298  and  (not A203) );
 a1353a <=( A302  and  A300 );
 a1354a <=( (not A299)  and  a1353a );
 a1355a <=( a1354a  and  a1349a );
 a1358a <=( A167  and  A168 );
 a1361a <=( (not A202)  and  (not A200) );
 a1362a <=( a1361a  and  a1358a );
 a1365a <=( A298  and  (not A203) );
 a1369a <=( A301  and  A300 );
 a1370a <=( (not A299)  and  a1369a );
 a1371a <=( a1370a  and  a1365a );
 a1374a <=( A167  and  A168 );
 a1377a <=( (not A202)  and  (not A200) );
 a1378a <=( a1377a  and  a1374a );
 a1381a <=( A298  and  (not A203) );
 a1385a <=( A302  and  A300 );
 a1386a <=( (not A299)  and  a1385a );
 a1387a <=( a1386a  and  a1381a );
 a1390a <=( (not A167)  and  A170 );
 a1393a <=( (not A199)  and  (not A166) );
 a1394a <=( a1393a  and  a1390a );
 a1397a <=( A298  and  A200 );
 a1401a <=( A301  and  A300 );
 a1402a <=( (not A299)  and  a1401a );
 a1403a <=( a1402a  and  a1397a );
 a1406a <=( (not A167)  and  A170 );
 a1409a <=( (not A199)  and  (not A166) );
 a1410a <=( a1409a  and  a1406a );
 a1413a <=( A298  and  A200 );
 a1417a <=( A302  and  A300 );
 a1418a <=( (not A299)  and  a1417a );
 a1419a <=( a1418a  and  a1413a );
 a1422a <=( (not A167)  and  A170 );
 a1425a <=( A199  and  (not A166) );
 a1426a <=( a1425a  and  a1422a );
 a1429a <=( A201  and  (not A200) );
 a1433a <=( A299  and  (not A298) );
 a1434a <=( A202  and  a1433a );
 a1435a <=( a1434a  and  a1429a );
 a1438a <=( (not A167)  and  A170 );
 a1441a <=( A199  and  (not A166) );
 a1442a <=( a1441a  and  a1438a );
 a1445a <=( A201  and  (not A200) );
 a1449a <=( A299  and  (not A298) );
 a1450a <=( A203  and  a1449a );
 a1451a <=( a1450a  and  a1445a );
 a1454a <=( A169  and  A170 );
 a1457a <=( (not A199)  and  (not A168) );
 a1458a <=( a1457a  and  a1454a );
 a1461a <=( A298  and  A200 );
 a1465a <=( A301  and  A300 );
 a1466a <=( (not A299)  and  a1465a );
 a1467a <=( a1466a  and  a1461a );
 a1470a <=( A169  and  A170 );
 a1473a <=( (not A199)  and  (not A168) );
 a1474a <=( a1473a  and  a1470a );
 a1477a <=( A298  and  A200 );
 a1481a <=( A302  and  A300 );
 a1482a <=( (not A299)  and  a1481a );
 a1483a <=( a1482a  and  a1477a );
 a1486a <=( A169  and  A170 );
 a1489a <=( A199  and  (not A168) );
 a1490a <=( a1489a  and  a1486a );
 a1493a <=( A201  and  (not A200) );
 a1497a <=( A299  and  (not A298) );
 a1498a <=( A202  and  a1497a );
 a1499a <=( a1498a  and  a1493a );
 a1502a <=( A169  and  A170 );
 a1505a <=( A199  and  (not A168) );
 a1506a <=( a1505a  and  a1502a );
 a1509a <=( A201  and  (not A200) );
 a1513a <=( A299  and  (not A298) );
 a1514a <=( A203  and  a1513a );
 a1515a <=( a1514a  and  a1509a );
 a1518a <=( A169  and  (not A170) );
 a1521a <=( A166  and  A167 );
 a1522a <=( a1521a  and  a1518a );
 a1525a <=( (not A202)  and  (not A200) );
 a1529a <=( A299  and  (not A298) );
 a1530a <=( (not A203)  and  a1529a );
 a1531a <=( a1530a  and  a1525a );
 a1534a <=( A169  and  (not A170) );
 a1537a <=( (not A166)  and  (not A167) );
 a1538a <=( a1537a  and  a1534a );
 a1541a <=( (not A202)  and  (not A200) );
 a1545a <=( A299  and  (not A298) );
 a1546a <=( (not A203)  and  a1545a );
 a1547a <=( a1546a  and  a1541a );
 a1550a <=( (not A167)  and  (not A169) );
 a1553a <=( (not A199)  and  (not A166) );
 a1554a <=( a1553a  and  a1550a );
 a1557a <=( A298  and  A200 );
 a1561a <=( A301  and  A300 );
 a1562a <=( (not A299)  and  a1561a );
 a1563a <=( a1562a  and  a1557a );
 a1566a <=( (not A167)  and  (not A169) );
 a1569a <=( (not A199)  and  (not A166) );
 a1570a <=( a1569a  and  a1566a );
 a1573a <=( A298  and  A200 );
 a1577a <=( A302  and  A300 );
 a1578a <=( (not A299)  and  a1577a );
 a1579a <=( a1578a  and  a1573a );
 a1582a <=( (not A167)  and  (not A169) );
 a1585a <=( A199  and  (not A166) );
 a1586a <=( a1585a  and  a1582a );
 a1589a <=( A201  and  (not A200) );
 a1593a <=( A299  and  (not A298) );
 a1594a <=( A202  and  a1593a );
 a1595a <=( a1594a  and  a1589a );
 a1598a <=( (not A167)  and  (not A169) );
 a1601a <=( A199  and  (not A166) );
 a1602a <=( a1601a  and  a1598a );
 a1605a <=( A201  and  (not A200) );
 a1609a <=( A299  and  (not A298) );
 a1610a <=( A203  and  a1609a );
 a1611a <=( a1610a  and  a1605a );
 a1614a <=( (not A169)  and  A170 );
 a1617a <=( (not A166)  and  A167 );
 a1618a <=( a1617a  and  a1614a );
 a1621a <=( (not A202)  and  (not A200) );
 a1625a <=( A299  and  (not A298) );
 a1626a <=( (not A203)  and  a1625a );
 a1627a <=( a1626a  and  a1621a );
 a1630a <=( (not A169)  and  A170 );
 a1633a <=( A166  and  (not A167) );
 a1634a <=( a1633a  and  a1630a );
 a1637a <=( (not A202)  and  (not A200) );
 a1641a <=( A299  and  (not A298) );
 a1642a <=( (not A203)  and  a1641a );
 a1643a <=( a1642a  and  a1637a );
 a1646a <=( (not A169)  and  (not A170) );
 a1649a <=( (not A199)  and  (not A168) );
 a1650a <=( a1649a  and  a1646a );
 a1653a <=( A298  and  A200 );
 a1657a <=( A301  and  A300 );
 a1658a <=( (not A299)  and  a1657a );
 a1659a <=( a1658a  and  a1653a );
 a1662a <=( (not A169)  and  (not A170) );
 a1665a <=( (not A199)  and  (not A168) );
 a1666a <=( a1665a  and  a1662a );
 a1669a <=( A298  and  A200 );
 a1673a <=( A302  and  A300 );
 a1674a <=( (not A299)  and  a1673a );
 a1675a <=( a1674a  and  a1669a );
 a1678a <=( (not A169)  and  (not A170) );
 a1681a <=( A199  and  (not A168) );
 a1682a <=( a1681a  and  a1678a );
 a1685a <=( A201  and  (not A200) );
 a1689a <=( A299  and  (not A298) );
 a1690a <=( A202  and  a1689a );
 a1691a <=( a1690a  and  a1685a );
 a1694a <=( (not A169)  and  (not A170) );
 a1697a <=( A199  and  (not A168) );
 a1698a <=( a1697a  and  a1694a );
 a1701a <=( A201  and  (not A200) );
 a1705a <=( A299  and  (not A298) );
 a1706a <=( A203  and  a1705a );
 a1707a <=( a1706a  and  a1701a );
 a1710a <=( (not A168)  and  A169 );
 a1714a <=( (not A199)  and  (not A166) );
 a1715a <=( A167  and  a1714a );
 a1716a <=( a1715a  and  a1710a );
 a1719a <=( A298  and  A200 );
 a1723a <=( A301  and  A300 );
 a1724a <=( (not A299)  and  a1723a );
 a1725a <=( a1724a  and  a1719a );
 a1728a <=( (not A168)  and  A169 );
 a1732a <=( (not A199)  and  (not A166) );
 a1733a <=( A167  and  a1732a );
 a1734a <=( a1733a  and  a1728a );
 a1737a <=( A298  and  A200 );
 a1741a <=( A302  and  A300 );
 a1742a <=( (not A299)  and  a1741a );
 a1743a <=( a1742a  and  a1737a );
 a1746a <=( (not A168)  and  A169 );
 a1750a <=( A199  and  (not A166) );
 a1751a <=( A167  and  a1750a );
 a1752a <=( a1751a  and  a1746a );
 a1755a <=( A201  and  (not A200) );
 a1759a <=( A299  and  (not A298) );
 a1760a <=( A202  and  a1759a );
 a1761a <=( a1760a  and  a1755a );
 a1764a <=( (not A168)  and  A169 );
 a1768a <=( A199  and  (not A166) );
 a1769a <=( A167  and  a1768a );
 a1770a <=( a1769a  and  a1764a );
 a1773a <=( A201  and  (not A200) );
 a1777a <=( A299  and  (not A298) );
 a1778a <=( A203  and  a1777a );
 a1779a <=( a1778a  and  a1773a );
 a1782a <=( (not A168)  and  A169 );
 a1786a <=( (not A199)  and  A166 );
 a1787a <=( (not A167)  and  a1786a );
 a1788a <=( a1787a  and  a1782a );
 a1791a <=( A298  and  A200 );
 a1795a <=( A301  and  A300 );
 a1796a <=( (not A299)  and  a1795a );
 a1797a <=( a1796a  and  a1791a );
 a1800a <=( (not A168)  and  A169 );
 a1804a <=( (not A199)  and  A166 );
 a1805a <=( (not A167)  and  a1804a );
 a1806a <=( a1805a  and  a1800a );
 a1809a <=( A298  and  A200 );
 a1813a <=( A302  and  A300 );
 a1814a <=( (not A299)  and  a1813a );
 a1815a <=( a1814a  and  a1809a );
 a1818a <=( (not A168)  and  A169 );
 a1822a <=( A199  and  A166 );
 a1823a <=( (not A167)  and  a1822a );
 a1824a <=( a1823a  and  a1818a );
 a1827a <=( A201  and  (not A200) );
 a1831a <=( A299  and  (not A298) );
 a1832a <=( A202  and  a1831a );
 a1833a <=( a1832a  and  a1827a );
 a1836a <=( (not A168)  and  A169 );
 a1840a <=( A199  and  A166 );
 a1841a <=( (not A167)  and  a1840a );
 a1842a <=( a1841a  and  a1836a );
 a1845a <=( A201  and  (not A200) );
 a1849a <=( A299  and  (not A298) );
 a1850a <=( A203  and  a1849a );
 a1851a <=( a1850a  and  a1845a );
 a1854a <=( A169  and  (not A170) );
 a1858a <=( A199  and  A166 );
 a1859a <=( A167  and  a1858a );
 a1860a <=( a1859a  and  a1854a );
 a1863a <=( A298  and  A200 );
 a1867a <=( A301  and  A300 );
 a1868a <=( (not A299)  and  a1867a );
 a1869a <=( a1868a  and  a1863a );
 a1872a <=( A169  and  (not A170) );
 a1876a <=( A199  and  A166 );
 a1877a <=( A167  and  a1876a );
 a1878a <=( a1877a  and  a1872a );
 a1881a <=( A298  and  A200 );
 a1885a <=( A302  and  A300 );
 a1886a <=( (not A299)  and  a1885a );
 a1887a <=( a1886a  and  a1881a );
 a1890a <=( A169  and  (not A170) );
 a1894a <=( (not A200)  and  A166 );
 a1895a <=( A167  and  a1894a );
 a1896a <=( a1895a  and  a1890a );
 a1899a <=( A298  and  (not A201) );
 a1903a <=( A301  and  A300 );
 a1904a <=( (not A299)  and  a1903a );
 a1905a <=( a1904a  and  a1899a );
 a1908a <=( A169  and  (not A170) );
 a1912a <=( (not A200)  and  A166 );
 a1913a <=( A167  and  a1912a );
 a1914a <=( a1913a  and  a1908a );
 a1917a <=( A298  and  (not A201) );
 a1921a <=( A302  and  A300 );
 a1922a <=( (not A299)  and  a1921a );
 a1923a <=( a1922a  and  a1917a );
 a1926a <=( A169  and  (not A170) );
 a1930a <=( (not A199)  and  A166 );
 a1931a <=( A167  and  a1930a );
 a1932a <=( a1931a  and  a1926a );
 a1935a <=( A298  and  (not A200) );
 a1939a <=( A301  and  A300 );
 a1940a <=( (not A299)  and  a1939a );
 a1941a <=( a1940a  and  a1935a );
 a1944a <=( A169  and  (not A170) );
 a1948a <=( (not A199)  and  A166 );
 a1949a <=( A167  and  a1948a );
 a1950a <=( a1949a  and  a1944a );
 a1953a <=( A298  and  (not A200) );
 a1957a <=( A302  and  A300 );
 a1958a <=( (not A299)  and  a1957a );
 a1959a <=( a1958a  and  a1953a );
 a1962a <=( A169  and  (not A170) );
 a1966a <=( A199  and  (not A166) );
 a1967a <=( (not A167)  and  a1966a );
 a1968a <=( a1967a  and  a1962a );
 a1971a <=( A298  and  A200 );
 a1975a <=( A301  and  A300 );
 a1976a <=( (not A299)  and  a1975a );
 a1977a <=( a1976a  and  a1971a );
 a1980a <=( A169  and  (not A170) );
 a1984a <=( A199  and  (not A166) );
 a1985a <=( (not A167)  and  a1984a );
 a1986a <=( a1985a  and  a1980a );
 a1989a <=( A298  and  A200 );
 a1993a <=( A302  and  A300 );
 a1994a <=( (not A299)  and  a1993a );
 a1995a <=( a1994a  and  a1989a );
 a1998a <=( A169  and  (not A170) );
 a2002a <=( (not A200)  and  (not A166) );
 a2003a <=( (not A167)  and  a2002a );
 a2004a <=( a2003a  and  a1998a );
 a2007a <=( A298  and  (not A201) );
 a2011a <=( A301  and  A300 );
 a2012a <=( (not A299)  and  a2011a );
 a2013a <=( a2012a  and  a2007a );
 a2016a <=( A169  and  (not A170) );
 a2020a <=( (not A200)  and  (not A166) );
 a2021a <=( (not A167)  and  a2020a );
 a2022a <=( a2021a  and  a2016a );
 a2025a <=( A298  and  (not A201) );
 a2029a <=( A302  and  A300 );
 a2030a <=( (not A299)  and  a2029a );
 a2031a <=( a2030a  and  a2025a );
 a2034a <=( A169  and  (not A170) );
 a2038a <=( (not A199)  and  (not A166) );
 a2039a <=( (not A167)  and  a2038a );
 a2040a <=( a2039a  and  a2034a );
 a2043a <=( A298  and  (not A200) );
 a2047a <=( A301  and  A300 );
 a2048a <=( (not A299)  and  a2047a );
 a2049a <=( a2048a  and  a2043a );
 a2052a <=( A169  and  (not A170) );
 a2056a <=( (not A199)  and  (not A166) );
 a2057a <=( (not A167)  and  a2056a );
 a2058a <=( a2057a  and  a2052a );
 a2061a <=( A298  and  (not A200) );
 a2065a <=( A302  and  A300 );
 a2066a <=( (not A299)  and  a2065a );
 a2067a <=( a2066a  and  a2061a );
 a2070a <=( (not A168)  and  (not A169) );
 a2074a <=( (not A199)  and  A166 );
 a2075a <=( A167  and  a2074a );
 a2076a <=( a2075a  and  a2070a );
 a2079a <=( A298  and  A200 );
 a2083a <=( A301  and  A300 );
 a2084a <=( (not A299)  and  a2083a );
 a2085a <=( a2084a  and  a2079a );
 a2088a <=( (not A168)  and  (not A169) );
 a2092a <=( (not A199)  and  A166 );
 a2093a <=( A167  and  a2092a );
 a2094a <=( a2093a  and  a2088a );
 a2097a <=( A298  and  A200 );
 a2101a <=( A302  and  A300 );
 a2102a <=( (not A299)  and  a2101a );
 a2103a <=( a2102a  and  a2097a );
 a2106a <=( (not A168)  and  (not A169) );
 a2110a <=( A199  and  A166 );
 a2111a <=( A167  and  a2110a );
 a2112a <=( a2111a  and  a2106a );
 a2115a <=( A201  and  (not A200) );
 a2119a <=( A299  and  (not A298) );
 a2120a <=( A202  and  a2119a );
 a2121a <=( a2120a  and  a2115a );
 a2124a <=( (not A168)  and  (not A169) );
 a2128a <=( A199  and  A166 );
 a2129a <=( A167  and  a2128a );
 a2130a <=( a2129a  and  a2124a );
 a2133a <=( A201  and  (not A200) );
 a2137a <=( A299  and  (not A298) );
 a2138a <=( A203  and  a2137a );
 a2139a <=( a2138a  and  a2133a );
 a2142a <=( (not A169)  and  A170 );
 a2146a <=( A199  and  (not A166) );
 a2147a <=( A167  and  a2146a );
 a2148a <=( a2147a  and  a2142a );
 a2151a <=( A298  and  A200 );
 a2155a <=( A301  and  A300 );
 a2156a <=( (not A299)  and  a2155a );
 a2157a <=( a2156a  and  a2151a );
 a2160a <=( (not A169)  and  A170 );
 a2164a <=( A199  and  (not A166) );
 a2165a <=( A167  and  a2164a );
 a2166a <=( a2165a  and  a2160a );
 a2169a <=( A298  and  A200 );
 a2173a <=( A302  and  A300 );
 a2174a <=( (not A299)  and  a2173a );
 a2175a <=( a2174a  and  a2169a );
 a2178a <=( (not A169)  and  A170 );
 a2182a <=( (not A200)  and  (not A166) );
 a2183a <=( A167  and  a2182a );
 a2184a <=( a2183a  and  a2178a );
 a2187a <=( A298  and  (not A201) );
 a2191a <=( A301  and  A300 );
 a2192a <=( (not A299)  and  a2191a );
 a2193a <=( a2192a  and  a2187a );
 a2196a <=( (not A169)  and  A170 );
 a2200a <=( (not A200)  and  (not A166) );
 a2201a <=( A167  and  a2200a );
 a2202a <=( a2201a  and  a2196a );
 a2205a <=( A298  and  (not A201) );
 a2209a <=( A302  and  A300 );
 a2210a <=( (not A299)  and  a2209a );
 a2211a <=( a2210a  and  a2205a );
 a2214a <=( (not A169)  and  A170 );
 a2218a <=( (not A199)  and  (not A166) );
 a2219a <=( A167  and  a2218a );
 a2220a <=( a2219a  and  a2214a );
 a2223a <=( A298  and  (not A200) );
 a2227a <=( A301  and  A300 );
 a2228a <=( (not A299)  and  a2227a );
 a2229a <=( a2228a  and  a2223a );
 a2232a <=( (not A169)  and  A170 );
 a2236a <=( (not A199)  and  (not A166) );
 a2237a <=( A167  and  a2236a );
 a2238a <=( a2237a  and  a2232a );
 a2241a <=( A298  and  (not A200) );
 a2245a <=( A302  and  A300 );
 a2246a <=( (not A299)  and  a2245a );
 a2247a <=( a2246a  and  a2241a );
 a2250a <=( (not A169)  and  A170 );
 a2254a <=( A199  and  A166 );
 a2255a <=( (not A167)  and  a2254a );
 a2256a <=( a2255a  and  a2250a );
 a2259a <=( A298  and  A200 );
 a2263a <=( A301  and  A300 );
 a2264a <=( (not A299)  and  a2263a );
 a2265a <=( a2264a  and  a2259a );
 a2268a <=( (not A169)  and  A170 );
 a2272a <=( A199  and  A166 );
 a2273a <=( (not A167)  and  a2272a );
 a2274a <=( a2273a  and  a2268a );
 a2277a <=( A298  and  A200 );
 a2281a <=( A302  and  A300 );
 a2282a <=( (not A299)  and  a2281a );
 a2283a <=( a2282a  and  a2277a );
 a2286a <=( (not A169)  and  A170 );
 a2290a <=( (not A200)  and  A166 );
 a2291a <=( (not A167)  and  a2290a );
 a2292a <=( a2291a  and  a2286a );
 a2295a <=( A298  and  (not A201) );
 a2299a <=( A301  and  A300 );
 a2300a <=( (not A299)  and  a2299a );
 a2301a <=( a2300a  and  a2295a );
 a2304a <=( (not A169)  and  A170 );
 a2308a <=( (not A200)  and  A166 );
 a2309a <=( (not A167)  and  a2308a );
 a2310a <=( a2309a  and  a2304a );
 a2313a <=( A298  and  (not A201) );
 a2317a <=( A302  and  A300 );
 a2318a <=( (not A299)  and  a2317a );
 a2319a <=( a2318a  and  a2313a );
 a2322a <=( (not A169)  and  A170 );
 a2326a <=( (not A199)  and  A166 );
 a2327a <=( (not A167)  and  a2326a );
 a2328a <=( a2327a  and  a2322a );
 a2331a <=( A298  and  (not A200) );
 a2335a <=( A301  and  A300 );
 a2336a <=( (not A299)  and  a2335a );
 a2337a <=( a2336a  and  a2331a );
 a2340a <=( (not A169)  and  A170 );
 a2344a <=( (not A199)  and  A166 );
 a2345a <=( (not A167)  and  a2344a );
 a2346a <=( a2345a  and  a2340a );
 a2349a <=( A298  and  (not A200) );
 a2353a <=( A302  and  A300 );
 a2354a <=( (not A299)  and  a2353a );
 a2355a <=( a2354a  and  a2349a );
 a2358a <=( (not A167)  and  A170 );
 a2362a <=( (not A200)  and  A199 );
 a2363a <=( (not A166)  and  a2362a );
 a2364a <=( a2363a  and  a2358a );
 a2368a <=( A298  and  A202 );
 a2369a <=( A201  and  a2368a );
 a2373a <=( A301  and  A300 );
 a2374a <=( (not A299)  and  a2373a );
 a2375a <=( a2374a  and  a2369a );
 a2378a <=( (not A167)  and  A170 );
 a2382a <=( (not A200)  and  A199 );
 a2383a <=( (not A166)  and  a2382a );
 a2384a <=( a2383a  and  a2378a );
 a2388a <=( A298  and  A202 );
 a2389a <=( A201  and  a2388a );
 a2393a <=( A302  and  A300 );
 a2394a <=( (not A299)  and  a2393a );
 a2395a <=( a2394a  and  a2389a );
 a2398a <=( (not A167)  and  A170 );
 a2402a <=( (not A200)  and  A199 );
 a2403a <=( (not A166)  and  a2402a );
 a2404a <=( a2403a  and  a2398a );
 a2408a <=( A298  and  A203 );
 a2409a <=( A201  and  a2408a );
 a2413a <=( A301  and  A300 );
 a2414a <=( (not A299)  and  a2413a );
 a2415a <=( a2414a  and  a2409a );
 a2418a <=( (not A167)  and  A170 );
 a2422a <=( (not A200)  and  A199 );
 a2423a <=( (not A166)  and  a2422a );
 a2424a <=( a2423a  and  a2418a );
 a2428a <=( A298  and  A203 );
 a2429a <=( A201  and  a2428a );
 a2433a <=( A302  and  A300 );
 a2434a <=( (not A299)  and  a2433a );
 a2435a <=( a2434a  and  a2429a );
 a2438a <=( A169  and  A170 );
 a2442a <=( (not A200)  and  A199 );
 a2443a <=( (not A168)  and  a2442a );
 a2444a <=( a2443a  and  a2438a );
 a2448a <=( A298  and  A202 );
 a2449a <=( A201  and  a2448a );
 a2453a <=( A301  and  A300 );
 a2454a <=( (not A299)  and  a2453a );
 a2455a <=( a2454a  and  a2449a );
 a2458a <=( A169  and  A170 );
 a2462a <=( (not A200)  and  A199 );
 a2463a <=( (not A168)  and  a2462a );
 a2464a <=( a2463a  and  a2458a );
 a2468a <=( A298  and  A202 );
 a2469a <=( A201  and  a2468a );
 a2473a <=( A302  and  A300 );
 a2474a <=( (not A299)  and  a2473a );
 a2475a <=( a2474a  and  a2469a );
 a2478a <=( A169  and  A170 );
 a2482a <=( (not A200)  and  A199 );
 a2483a <=( (not A168)  and  a2482a );
 a2484a <=( a2483a  and  a2478a );
 a2488a <=( A298  and  A203 );
 a2489a <=( A201  and  a2488a );
 a2493a <=( A301  and  A300 );
 a2494a <=( (not A299)  and  a2493a );
 a2495a <=( a2494a  and  a2489a );
 a2498a <=( A169  and  A170 );
 a2502a <=( (not A200)  and  A199 );
 a2503a <=( (not A168)  and  a2502a );
 a2504a <=( a2503a  and  a2498a );
 a2508a <=( A298  and  A203 );
 a2509a <=( A201  and  a2508a );
 a2513a <=( A302  and  A300 );
 a2514a <=( (not A299)  and  a2513a );
 a2515a <=( a2514a  and  a2509a );
 a2518a <=( A169  and  (not A170) );
 a2522a <=( (not A200)  and  A166 );
 a2523a <=( A167  and  a2522a );
 a2524a <=( a2523a  and  a2518a );
 a2528a <=( A298  and  (not A203) );
 a2529a <=( (not A202)  and  a2528a );
 a2533a <=( A301  and  A300 );
 a2534a <=( (not A299)  and  a2533a );
 a2535a <=( a2534a  and  a2529a );
 a2538a <=( A169  and  (not A170) );
 a2542a <=( (not A200)  and  A166 );
 a2543a <=( A167  and  a2542a );
 a2544a <=( a2543a  and  a2538a );
 a2548a <=( A298  and  (not A203) );
 a2549a <=( (not A202)  and  a2548a );
 a2553a <=( A302  and  A300 );
 a2554a <=( (not A299)  and  a2553a );
 a2555a <=( a2554a  and  a2549a );
 a2558a <=( A169  and  (not A170) );
 a2562a <=( (not A200)  and  (not A166) );
 a2563a <=( (not A167)  and  a2562a );
 a2564a <=( a2563a  and  a2558a );
 a2568a <=( A298  and  (not A203) );
 a2569a <=( (not A202)  and  a2568a );
 a2573a <=( A301  and  A300 );
 a2574a <=( (not A299)  and  a2573a );
 a2575a <=( a2574a  and  a2569a );
 a2578a <=( A169  and  (not A170) );
 a2582a <=( (not A200)  and  (not A166) );
 a2583a <=( (not A167)  and  a2582a );
 a2584a <=( a2583a  and  a2578a );
 a2588a <=( A298  and  (not A203) );
 a2589a <=( (not A202)  and  a2588a );
 a2593a <=( A302  and  A300 );
 a2594a <=( (not A299)  and  a2593a );
 a2595a <=( a2594a  and  a2589a );
 a2598a <=( (not A167)  and  (not A169) );
 a2602a <=( (not A200)  and  A199 );
 a2603a <=( (not A166)  and  a2602a );
 a2604a <=( a2603a  and  a2598a );
 a2608a <=( A298  and  A202 );
 a2609a <=( A201  and  a2608a );
 a2613a <=( A301  and  A300 );
 a2614a <=( (not A299)  and  a2613a );
 a2615a <=( a2614a  and  a2609a );
 a2618a <=( (not A167)  and  (not A169) );
 a2622a <=( (not A200)  and  A199 );
 a2623a <=( (not A166)  and  a2622a );
 a2624a <=( a2623a  and  a2618a );
 a2628a <=( A298  and  A202 );
 a2629a <=( A201  and  a2628a );
 a2633a <=( A302  and  A300 );
 a2634a <=( (not A299)  and  a2633a );
 a2635a <=( a2634a  and  a2629a );
 a2638a <=( (not A167)  and  (not A169) );
 a2642a <=( (not A200)  and  A199 );
 a2643a <=( (not A166)  and  a2642a );
 a2644a <=( a2643a  and  a2638a );
 a2648a <=( A298  and  A203 );
 a2649a <=( A201  and  a2648a );
 a2653a <=( A301  and  A300 );
 a2654a <=( (not A299)  and  a2653a );
 a2655a <=( a2654a  and  a2649a );
 a2658a <=( (not A167)  and  (not A169) );
 a2662a <=( (not A200)  and  A199 );
 a2663a <=( (not A166)  and  a2662a );
 a2664a <=( a2663a  and  a2658a );
 a2668a <=( A298  and  A203 );
 a2669a <=( A201  and  a2668a );
 a2673a <=( A302  and  A300 );
 a2674a <=( (not A299)  and  a2673a );
 a2675a <=( a2674a  and  a2669a );
 a2678a <=( (not A169)  and  A170 );
 a2682a <=( (not A200)  and  (not A166) );
 a2683a <=( A167  and  a2682a );
 a2684a <=( a2683a  and  a2678a );
 a2688a <=( A298  and  (not A203) );
 a2689a <=( (not A202)  and  a2688a );
 a2693a <=( A301  and  A300 );
 a2694a <=( (not A299)  and  a2693a );
 a2695a <=( a2694a  and  a2689a );
 a2698a <=( (not A169)  and  A170 );
 a2702a <=( (not A200)  and  (not A166) );
 a2703a <=( A167  and  a2702a );
 a2704a <=( a2703a  and  a2698a );
 a2708a <=( A298  and  (not A203) );
 a2709a <=( (not A202)  and  a2708a );
 a2713a <=( A302  and  A300 );
 a2714a <=( (not A299)  and  a2713a );
 a2715a <=( a2714a  and  a2709a );
 a2718a <=( (not A169)  and  A170 );
 a2722a <=( (not A200)  and  A166 );
 a2723a <=( (not A167)  and  a2722a );
 a2724a <=( a2723a  and  a2718a );
 a2728a <=( A298  and  (not A203) );
 a2729a <=( (not A202)  and  a2728a );
 a2733a <=( A301  and  A300 );
 a2734a <=( (not A299)  and  a2733a );
 a2735a <=( a2734a  and  a2729a );
 a2738a <=( (not A169)  and  A170 );
 a2742a <=( (not A200)  and  A166 );
 a2743a <=( (not A167)  and  a2742a );
 a2744a <=( a2743a  and  a2738a );
 a2748a <=( A298  and  (not A203) );
 a2749a <=( (not A202)  and  a2748a );
 a2753a <=( A302  and  A300 );
 a2754a <=( (not A299)  and  a2753a );
 a2755a <=( a2754a  and  a2749a );
 a2758a <=( (not A169)  and  (not A170) );
 a2762a <=( (not A200)  and  A199 );
 a2763a <=( (not A168)  and  a2762a );
 a2764a <=( a2763a  and  a2758a );
 a2768a <=( A298  and  A202 );
 a2769a <=( A201  and  a2768a );
 a2773a <=( A301  and  A300 );
 a2774a <=( (not A299)  and  a2773a );
 a2775a <=( a2774a  and  a2769a );
 a2778a <=( (not A169)  and  (not A170) );
 a2782a <=( (not A200)  and  A199 );
 a2783a <=( (not A168)  and  a2782a );
 a2784a <=( a2783a  and  a2778a );
 a2788a <=( A298  and  A202 );
 a2789a <=( A201  and  a2788a );
 a2793a <=( A302  and  A300 );
 a2794a <=( (not A299)  and  a2793a );
 a2795a <=( a2794a  and  a2789a );
 a2798a <=( (not A169)  and  (not A170) );
 a2802a <=( (not A200)  and  A199 );
 a2803a <=( (not A168)  and  a2802a );
 a2804a <=( a2803a  and  a2798a );
 a2808a <=( A298  and  A203 );
 a2809a <=( A201  and  a2808a );
 a2813a <=( A301  and  A300 );
 a2814a <=( (not A299)  and  a2813a );
 a2815a <=( a2814a  and  a2809a );
 a2818a <=( (not A169)  and  (not A170) );
 a2822a <=( (not A200)  and  A199 );
 a2823a <=( (not A168)  and  a2822a );
 a2824a <=( a2823a  and  a2818a );
 a2828a <=( A298  and  A203 );
 a2829a <=( A201  and  a2828a );
 a2833a <=( A302  and  A300 );
 a2834a <=( (not A299)  and  a2833a );
 a2835a <=( a2834a  and  a2829a );
 a2839a <=( A167  and  (not A168) );
 a2840a <=( A169  and  a2839a );
 a2844a <=( (not A200)  and  A199 );
 a2845a <=( (not A166)  and  a2844a );
 a2846a <=( a2845a  and  a2840a );
 a2850a <=( A298  and  A202 );
 a2851a <=( A201  and  a2850a );
 a2855a <=( A301  and  A300 );
 a2856a <=( (not A299)  and  a2855a );
 a2857a <=( a2856a  and  a2851a );
 a2861a <=( A167  and  (not A168) );
 a2862a <=( A169  and  a2861a );
 a2866a <=( (not A200)  and  A199 );
 a2867a <=( (not A166)  and  a2866a );
 a2868a <=( a2867a  and  a2862a );
 a2872a <=( A298  and  A202 );
 a2873a <=( A201  and  a2872a );
 a2877a <=( A302  and  A300 );
 a2878a <=( (not A299)  and  a2877a );
 a2879a <=( a2878a  and  a2873a );
 a2883a <=( A167  and  (not A168) );
 a2884a <=( A169  and  a2883a );
 a2888a <=( (not A200)  and  A199 );
 a2889a <=( (not A166)  and  a2888a );
 a2890a <=( a2889a  and  a2884a );
 a2894a <=( A298  and  A203 );
 a2895a <=( A201  and  a2894a );
 a2899a <=( A301  and  A300 );
 a2900a <=( (not A299)  and  a2899a );
 a2901a <=( a2900a  and  a2895a );
 a2905a <=( A167  and  (not A168) );
 a2906a <=( A169  and  a2905a );
 a2910a <=( (not A200)  and  A199 );
 a2911a <=( (not A166)  and  a2910a );
 a2912a <=( a2911a  and  a2906a );
 a2916a <=( A298  and  A203 );
 a2917a <=( A201  and  a2916a );
 a2921a <=( A302  and  A300 );
 a2922a <=( (not A299)  and  a2921a );
 a2923a <=( a2922a  and  a2917a );
 a2927a <=( (not A167)  and  (not A168) );
 a2928a <=( A169  and  a2927a );
 a2932a <=( (not A200)  and  A199 );
 a2933a <=( A166  and  a2932a );
 a2934a <=( a2933a  and  a2928a );
 a2938a <=( A298  and  A202 );
 a2939a <=( A201  and  a2938a );
 a2943a <=( A301  and  A300 );
 a2944a <=( (not A299)  and  a2943a );
 a2945a <=( a2944a  and  a2939a );
 a2949a <=( (not A167)  and  (not A168) );
 a2950a <=( A169  and  a2949a );
 a2954a <=( (not A200)  and  A199 );
 a2955a <=( A166  and  a2954a );
 a2956a <=( a2955a  and  a2950a );
 a2960a <=( A298  and  A202 );
 a2961a <=( A201  and  a2960a );
 a2965a <=( A302  and  A300 );
 a2966a <=( (not A299)  and  a2965a );
 a2967a <=( a2966a  and  a2961a );
 a2971a <=( (not A167)  and  (not A168) );
 a2972a <=( A169  and  a2971a );
 a2976a <=( (not A200)  and  A199 );
 a2977a <=( A166  and  a2976a );
 a2978a <=( a2977a  and  a2972a );
 a2982a <=( A298  and  A203 );
 a2983a <=( A201  and  a2982a );
 a2987a <=( A301  and  A300 );
 a2988a <=( (not A299)  and  a2987a );
 a2989a <=( a2988a  and  a2983a );
 a2993a <=( (not A167)  and  (not A168) );
 a2994a <=( A169  and  a2993a );
 a2998a <=( (not A200)  and  A199 );
 a2999a <=( A166  and  a2998a );
 a3000a <=( a2999a  and  a2994a );
 a3004a <=( A298  and  A203 );
 a3005a <=( A201  and  a3004a );
 a3009a <=( A302  and  A300 );
 a3010a <=( (not A299)  and  a3009a );
 a3011a <=( a3010a  and  a3005a );
 a3015a <=( A167  and  (not A168) );
 a3016a <=( (not A169)  and  a3015a );
 a3020a <=( (not A200)  and  A199 );
 a3021a <=( A166  and  a3020a );
 a3022a <=( a3021a  and  a3016a );
 a3026a <=( A298  and  A202 );
 a3027a <=( A201  and  a3026a );
 a3031a <=( A301  and  A300 );
 a3032a <=( (not A299)  and  a3031a );
 a3033a <=( a3032a  and  a3027a );
 a3037a <=( A167  and  (not A168) );
 a3038a <=( (not A169)  and  a3037a );
 a3042a <=( (not A200)  and  A199 );
 a3043a <=( A166  and  a3042a );
 a3044a <=( a3043a  and  a3038a );
 a3048a <=( A298  and  A202 );
 a3049a <=( A201  and  a3048a );
 a3053a <=( A302  and  A300 );
 a3054a <=( (not A299)  and  a3053a );
 a3055a <=( a3054a  and  a3049a );
 a3059a <=( A167  and  (not A168) );
 a3060a <=( (not A169)  and  a3059a );
 a3064a <=( (not A200)  and  A199 );
 a3065a <=( A166  and  a3064a );
 a3066a <=( a3065a  and  a3060a );
 a3070a <=( A298  and  A203 );
 a3071a <=( A201  and  a3070a );
 a3075a <=( A301  and  A300 );
 a3076a <=( (not A299)  and  a3075a );
 a3077a <=( a3076a  and  a3071a );
 a3081a <=( A167  and  (not A168) );
 a3082a <=( (not A169)  and  a3081a );
 a3086a <=( (not A200)  and  A199 );
 a3087a <=( A166  and  a3086a );
 a3088a <=( a3087a  and  a3082a );
 a3092a <=( A298  and  A203 );
 a3093a <=( A201  and  a3092a );
 a3097a <=( A302  and  A300 );
 a3098a <=( (not A299)  and  a3097a );
 a3099a <=( a3098a  and  a3093a );


end x25_8x_behav;
