Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_19x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A40: buffer std_logic
);
end x25_19x;

architecture x25_19x_behav of x25_19x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1753a,a1754a,a1755a,a1756a,a1757a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1765a,a1766a,a1767a,a1768a,a1769a,a1770a,a1771a,a1772a,a1773a,a1774a,a1775a,a1776a,a1777a,a1778a,a1779a,a1780a,a1781a,a1782a,a1783a,a1784a,a1785a,a1786a,a1787a,a1788a,a1789a,a1790a,a1791a,a1792a,a1793a,a1794a,a1795a,a1796a,a1797a,a1798a,a1799a,a1800a,a1801a,a1802a,a1803a,a1804a,a1805a,a1806a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1816a,a1817a,a1818a,a1819a,a1820a,a1821a,a1822a,a1823a,a1824a,a1825a,a1826a,a1827a,a1828a,a1829a,a1830a,a1831a,a1832a,a1833a,a1834a,a1835a,a1836a,a1837a,a1838a,a1839a,a1840a,a1841a,a1842a,a1843a,a1844a,a1845a,a1846a,a1847a,a1848a,a1849a,a1850a,a1851a,a1852a,a1853a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1860a,a1861a,a1862a,a1863a,a1864a,a1865a,a1866a,a1867a,a1868a,a1869a,a1870a,a1871a,a1872a,a1873a,a1874a,a1875a,a1876a,a1877a,a1878a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1890a,a1891a,a1892a,a1893a,a1894a,a1895a,a1896a,a1897a,a1898a,a1899a,a1900a,a1901a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1910a,a1911a,a1912a,a1913a,a1914a,a1915a,a1916a,a1917a,a1918a,a1919a,a1920a,a1921a,a1922a,a1923a,a1924a,a1925a,a1926a,a1927a,a1928a,a1929a,a1930a,a1931a,a1932a,a1933a,a1934a,a1935a,a1936a,a1937a,a1938a,a1939a,a1940a,a1941a,a1942a,a1943a,a1944a,a1945a,a1946a,a1947a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1956a,a1957a,a1958a,a1959a,a1960a,a1961a,a1962a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1970a,a1971a,a1972a,a1973a,a1974a,a1975a,a1976a,a1977a,a1978a,a1979a,a1980a,a1981a,a1982a,a1983a,a1984a,a1985a,a1986a,a1987a,a1988a,a1989a,a1990a,a1991a,a1992a,a1993a,a1994a,a1995a,a1996a,a1997a,a1998a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2005a,a2006a,a2007a,a2008a,a2009a,a2010a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2025a,a2026a,a2027a,a2028a,a2029a,a2030a,a2031a,a2032a,a2033a,a2034a,a2035a,a2036a,a2037a,a2038a,a2039a,a2040a,a2041a,a2042a,a2043a,a2044a,a2045a,a2046a,a2047a,a2048a,a2049a,a2050a,a2051a,a2052a,a2053a,a2054a,a2055a,a2056a,a2057a,a2058a,a2059a,a2060a,a2061a,a2062a,a2063a,a2064a,a2065a,a2066a,a2067a,a2068a,a2069a,a2070a,a2071a,a2072a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2079a,a2080a,a2081a,a2082a,a2083a,a2084a,a2085a,a2086a,a2087a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2101a,a2102a,a2103a,a2104a,a2105a,a2106a,a2107a,a2108a,a2109a,a2110a,a2111a,a2112a,a2113a,a2114a,a2115a,a2116a,a2117a,a2118a,a2119a,a2120a,a2121a,a2122a,a2123a,a2124a,a2125a,a2126a,a2127a,a2128a,a2129a,a2130a,a2131a,a2132a,a2133a,a2134a,a2135a,a2136a,a2137a,a2138a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2145a,a2146a,a2147a,a2148a,a2149a,a2150a,a2151a,a2152a,a2153a,a2154a,a2155a,a2156a,a2157a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2164a,a2165a,a2166a,a2167a,a2168a,a2169a,a2170a,a2171a,a2172a,a2173a,a2174a,a2175a,a2176a,a2177a,a2178a,a2179a,a2180a,a2181a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2190a,a2191a,a2192a,a2193a,a2194a,a2195a,a2196a,a2197a,a2198a,a2199a,a2200a,a2201a,a2202a,a2203a,a2204a,a2205a,a2206a,a2207a,a2208a,a2209a,a2210a,a2211a,a2212a,a2213a,a2214a,a2215a,a2216a,a2217a,a2218a,a2219a,a2220a,a2221a,a2222a,a2223a,a2224a,a2225a,a2226a,a2227a,a2228a,a2229a,a2230a,a2231a,a2232a,a2233a,a2234a,a2235a,a2236a,a2237a,a2238a,a2239a,a2240a,a2241a,a2242a,a2243a,a2244a,a2245a,a2246a,a2247a,a2248a,a2249a,a2250a,a2251a,a2252a,a2253a,a2254a,a2255a,a2256a,a2257a,a2258a,a2259a,a2260a,a2261a,a2262a,a2263a,a2264a,a2265a,a2266a,a2267a,a2268a,a2269a,a2270a,a2271a,a2272a,a2273a,a2274a,a2275a,a2276a,a2277a,a2278a,a2279a,a2280a,a2281a,a2282a,a2283a,a2284a,a2285a,a2286a,a2287a,a2288a,a2289a,a2290a,a2291a,a2292a,a2293a,a2294a,a2295a,a2296a,a2297a,a2298a,a2299a,a2300a,a2301a,a2302a,a2303a,a2304a,a2305a,a2306a,a2307a,a2308a,a2309a,a2310a,a2311a,a2312a,a2313a,a2314a,a2315a,a2316a,a2317a,a2318a,a2319a,a2320a,a2321a,a2322a,a2323a,a2324a,a2325a,a2326a,a2327a,a2328a,a2329a,a2330a,a2331a,a2332a,a2333a,a2334a,a2335a,a2336a,a2337a,a2338a,a2339a,a2340a,a2341a,a2342a,a2343a,a2344a,a2345a,a2346a,a2347a,a2348a,a2349a,a2350a,a2351a,a2352a,a2353a,a2354a,a2355a,a2356a,a2357a,a2358a,a2359a,a2360a,a2361a,a2362a,a2363a,a2364a,a2365a,a2366a,a2367a,a2368a,a2369a,a2370a,a2371a,a2372a,a2373a,a2374a,a2375a,a2376a,a2377a,a2378a,a2379a,a2380a,a2381a,a2382a,a2383a,a2384a,a2385a,a2386a,a2387a,a2388a,a2389a,a2390a,a2391a,a2392a,a2393a,a2394a,a2395a,a2396a,a2397a,a2398a,a2399a,a2400a,a2401a,a2402a,a2403a,a2404a,a2405a,a2406a,a2407a,a2408a,a2409a,a2410a,a2411a,a2412a,a2413a,a2414a,a2415a,a2416a,a2417a,a2418a,a2419a,a2420a,a2421a,a2422a,a2423a,a2424a,a2425a,a2426a,a2427a,a2428a,a2429a,a2430a,a2431a,a2432a,a2433a,a2434a,a2435a,a2436a,a2437a,a2438a,a2439a,a2440a,a2441a,a2442a,a2443a,a2444a,a2445a,a2446a,a2447a,a2448a,a2449a,a2450a,a2451a,a2452a,a2453a,a2454a,a2455a,a2456a,a2457a,a2458a,a2459a,a2460a,a2461a,a2462a,a2463a,a2464a,a2465a,a2466a,a2467a,a2468a,a2469a,a2470a,a2471a,a2472a,a2473a,a2474a,a2475a,a2476a,a2477a,a2478a,a2479a,a2480a,a2481a,a2482a,a2483a,a2484a,a2485a,a2486a,a2487a,a2488a,a2489a,a2490a,a2491a,a2492a,a2493a,a2494a,a2495a,a2496a,a2497a,a2498a,a2499a,a2500a,a2501a,a2502a,a2503a,a2504a,a2505a,a2506a,a2507a,a2508a,a2509a,a2510a,a2511a,a2512a,a2513a,a2514a,a2515a,a2516a,a2517a,a2518a,a2519a,a2520a,a2521a,a2522a,a2523a,a2524a,a2525a,a2526a,a2527a,a2528a,a2529a,a2530a,a2531a,a2532a,a2533a,a2534a,a2535a,a2536a,a2537a,a2538a,a2539a,a2540a,a2541a,a2542a,a2543a,a2544a,a2545a,a2546a,a2547a,a2548a,a2549a,a2550a,a2551a,a2552a,a2553a,a2554a,a2555a,a2556a,a2557a,a2558a,a2559a,a2560a,a2561a,a2562a,a2563a,a2564a,a2565a,a2566a,a2567a,a2568a,a2569a,a2570a,a2571a,a2572a,a2573a,a2574a,a2575a,a2576a,a2577a,a2578a,a2579a,a2580a,a2581a,a2582a,a2583a,a2584a,a2585a,a2586a,a2587a,a2588a,a2589a,a2590a,a2591a,a2592a,a2593a,a2594a,a2595a,a2596a,a2597a,a2598a,a2599a,a2600a,a2601a,a2602a,a2603a,a2604a,a2605a,a2606a,a2607a,a2608a,a2609a,a2610a,a2611a,a2612a,a2613a,a2614a,a2615a,a2616a,a2617a,a2618a,a2619a,a2620a,a2621a,a2622a,a2623a,a2624a,a2625a,a2626a,a2627a,a2628a,a2629a,a2630a,a2631a,a2632a,a2633a,a2634a,a2635a,a2636a,a2637a,a2638a,a2639a,a2640a,a2641a,a2642a,a2643a,a2644a,a2645a,a2646a,a2647a,a2648a,a2649a,a2650a,a2651a,a2652a,a2653a,a2654a,a2655a,a2656a,a2657a,a2658a,a2659a,a2660a,a2661a,a2662a,a2663a,a2664a,a2665a,a2666a,a2667a,a2668a,a2669a,a2670a,a2671a,a2672a,a2673a,a2674a,a2675a,a2676a,a2677a,a2678a,a2679a,a2680a,a2681a,a2682a,a2683a,a2684a,a2685a,a2686a,a2687a,a2688a,a2689a,a2690a,a2691a,a2692a,a2693a,a2694a,a2695a,a2696a,a2697a,a2698a,a2699a,a2700a,a2701a,a2702a,a2703a,a2704a,a2705a,a2706a,a2707a,a2708a,a2709a,a2710a,a2711a,a2712a,a2713a,a2714a,a2715a,a2716a,a2717a,a2718a,a2719a,a2720a,a2721a,a2722a,a2723a,a2724a,a2725a,a2726a,a2727a,a2728a,a2729a,a2730a,a2731a,a2732a,a2733a,a2734a,a2735a,a2736a,a2737a,a2738a,a2739a,a2740a,a2741a,a2742a,a2743a,a2744a,a2745a,a2746a,a2747a,a2748a,a2749a,a2750a,a2751a,a2752a,a2753a,a2754a,a2755a,a2756a,a2757a,a2758a,a2759a,a2760a,a2761a,a2762a,a2763a,a2764a,a2765a,a2766a,a2767a,a2768a,a2769a,a2770a,a2771a,a2772a,a2773a,a2774a,a2775a,a2776a,a2777a,a2778a,a2779a,a2780a,a2781a,a2782a,a2783a,a2784a,a2785a,a2786a,a2787a,a2788a,a2789a,a2790a,a2791a,a2792a,a2793a,a2794a,a2795a,a2796a,a2797a,a2798a,a2799a,a2800a,a2801a,a2802a,a2803a,a2804a,a2805a,a2806a,a2807a,a2808a,a2809a,a2810a,a2811a,a2812a,a2813a,a2814a,a2815a,a2816a,a2817a,a2818a,a2819a,a2820a,a2821a,a2822a,a2823a,a2824a,a2825a,a2826a,a2827a,a2828a,a2829a,a2830a,a2831a,a2832a,a2833a,a2834a,a2835a,a2836a,a2837a,a2838a,a2839a,a2840a,a2841a,a2842a,a2843a,a2844a,a2845a,a2846a,a2847a,a2848a,a2849a,a2850a,a2851a,a2852a,a2853a,a2854a,a2855a,a2856a,a2857a,a2858a,a2859a,a2860a,a2861a,a2862a,a2863a,a2864a,a2865a,a2866a,a2867a,a2868a,a2869a,a2870a,a2871a,a2872a,a2873a,a2874a,a2875a,a2876a,a2877a,a2878a,a2879a,a2880a,a2881a,a2882a,a2883a,a2884a,a2885a,a2886a,a2887a,a2888a,a2889a,a2890a,a2891a,a2892a,a2893a,a2894a,a2895a,a2896a,a2897a,a2898a,a2899a,a2900a,a2901a,a2902a,a2903a,a2904a,a2905a,a2906a,a2907a,a2908a,a2909a,a2910a,a2911a,a2912a,a2913a,a2914a,a2915a,a2916a,a2917a,a2918a,a2919a,a2920a,a2921a,a2922a,a2923a,a2924a,a2925a,a2926a,a2927a,a2928a,a2929a,a2930a,a2931a,a2932a,a2933a,a2934a,a2935a,a2936a,a2937a,a2938a,a2939a,a2940a,a2941a,a2942a,a2943a,a2944a,a2945a,a2946a,a2947a,a2948a,a2949a,a2950a,a2951a,a2952a,a2953a,a2954a,a2955a,a2956a,a2957a,a2958a,a2959a,a2960a,a2961a,a2962a,a2963a,a2964a,a2965a,a2966a,a2967a,a2968a,a2969a,a2970a,a2971a,a2972a,a2973a,a2974a,a2975a,a2976a,a2977a,a2978a,a2979a,a2980a,a2981a,a2982a,a2983a,a2984a,a2985a,a2986a,a2987a,a2988a,a2989a,a2990a,a2991a,a2992a,a2993a,a2994a,a2995a,a2996a,a2997a,a2998a,a2999a,a3000a,a3001a,a3002a,a3003a,a3004a,a3005a,a3006a,a3007a,a3008a,a3009a,a3010a,a3011a,a3012a,a3013a,a3014a,a3015a,a3016a,a3017a,a3018a,a3019a,a3020a,a3021a,a3022a,a3023a,a3024a,a3025a,a3026a,a3027a,a3028a,a3029a,a3030a,a3031a,a3032a,a3033a,a3034a,a3035a,a3036a,a3037a,a3038a,a3039a,a3040a,a3041a,a3042a,a3043a,a3044a,a3045a,a3046a,a3047a,a3048a,a3049a,a3050a,a3051a,a3052a,a3053a,a3054a,a3055a,a3056a,a3057a,a3058a,a3059a,a3060a,a3061a,a3062a,a3063a,a3064a,a3065a,a3066a,a3067a,a3068a,a3069a,a3070a,a3071a,a3072a,a3073a,a3074a,a3075a,a3076a,a3077a,a3078a,a3079a,a3080a,a3081a,a3082a,a3083a,a3084a,a3085a,a3086a,a3087a,a3088a,a3089a,a3090a,a3091a,a3092a,a3093a,a3094a,a3095a,a3096a,a3097a,a3098a,a3099a,a3100a,a3101a,a3102a,a3103a,a3104a,a3105a,a3106a,a3107a,a3108a,a3109a,a3110a,a3111a,a3112a,a3113a,a3114a,a3115a,a3116a,a3117a,a3118a,a3119a,a3120a,a3121a,a3122a,a3123a,a3124a,a3125a,a3126a,a3127a,a3128a,a3129a,a3130a,a3131a,a3132a,a3133a,a3134a,a3135a,a3136a,a3137a,a3138a,a3139a,a3140a,a3141a,a3142a,a3143a,a3144a,a3145a,a3146a,a3147a,a3148a,a3149a,a3150a,a3151a,a3152a,a3153a,a3154a,a3155a,a3156a,a3157a,a3158a,a3159a,a3160a,a3161a,a3162a,a3163a,a3164a,a3165a,a3166a,a3167a,a3168a,a3169a,a3170a,a3171a,a3172a,a3173a,a3174a,a3175a,a3176a,a3177a,a3178a,a3179a,a3180a,a3181a,a3182a,a3183a,a3184a,a3185a,a3186a,a3187a,a3188a,a3189a,a3190a,a3191a,a3192a,a3193a,a3194a,a3195a,a3196a,a3197a,a3198a,a3199a,a3200a,a3201a,a3202a,a3203a,a3204a,a3205a,a3206a,a3207a,a3208a,a3209a,a3210a,a3211a,a3212a,a3213a,a3214a,a3215a,a3216a,a3217a,a3218a,a3219a,a3220a,a3221a,a3222a,a3223a,a3224a,a3225a,a3226a,a3227a,a3228a,a3229a,a3230a,a3231a,a3232a,a3233a,a3234a,a3235a,a3236a,a3237a,a3238a,a3239a,a3240a,a3241a,a3242a,a3243a,a3244a,a3245a,a3246a,a3247a,a3248a,a3249a,a3250a,a3251a,a3252a,a3253a,a3254a,a3255a,a3256a,a3257a,a3258a,a3259a,a3260a,a3261a,a3262a,a3263a,a3264a,a3265a,a3266a,a3267a,a3268a,a3269a,a3270a,a3271a,a3272a,a3273a,a3274a,a3275a,a3276a,a3277a,a3278a,a3279a,a3280a,a3281a,a3282a,a3283a,a3284a,a3285a,a3286a,a3287a,a3288a,a3289a,a3290a,a3291a,a3292a,a3293a,a3294a,a3295a,a3296a,a3297a,a3298a,a3299a,a3300a,a3301a,a3302a,a3303a,a3304a,a3305a,a3306a,a3307a,a3308a,a3309a,a3310a,a3311a,a3312a,a3313a,a3314a,a3315a,a3316a,a3317a,a3318a,a3319a,a3320a,a3321a,a3322a,a3323a,a3324a,a3325a,a3326a,a3327a,a3328a,a3329a,a3330a,a3331a,a3332a,a3333a,a3334a,a3335a,a3336a,a3337a,a3338a,a3339a,a3340a,a3341a,a3342a,a3343a,a3344a,a3345a,a3346a,a3347a,a3348a,a3349a,a3350a,a3351a,a3352a,a3353a,a3354a,a3355a,a3356a,a3357a,a3358a,a3359a,a3360a,a3361a,a3362a,a3363a,a3364a,a3365a,a3366a,a3367a,a3368a,a3369a,a3370a,a3371a,a3372a,a3373a,a3374a,a3375a,a3376a,a3377a,a3378a,a3379a,a3380a,a3381a,a3382a,a3383a,a3384a,a3385a,a3386a,a3387a,a3388a,a3389a,a3390a,a3391a,a3392a,a3393a,a3394a,a3395a,a3396a,a3397a,a3398a,a3399a,a3400a,a3401a,a3402a,a3403a,a3404a,a3405a,a3406a,a3407a,a3408a,a3409a,a3410a,a3411a,a3412a,a3413a,a3414a,a3415a,a3416a,a3417a,a3418a,a3419a,a3420a,a3421a,a3422a,a3423a,a3424a,a3425a,a3426a,a3427a,a3428a,a3429a,a3430a,a3431a,a3432a,a3433a,a3434a,a3435a,a3436a,a3437a,a3438a,a3439a,a3440a,a3441a,a3442a,a3443a,a3444a,a3445a,a3446a,a3447a,a3448a,a3449a,a3450a,a3451a,a3452a,a3453a,a3454a,a3455a,a3456a,a3457a,a3458a,a3459a,a3460a,a3461a,a3462a,a3463a,a3464a,a3465a,a3466a,a3467a,a3468a,a3469a,a3470a,a3471a,a3472a,a3473a,a3474a,a3475a,a3476a,a3477a,a3478a,a3479a,a3480a,a3481a,a3482a,a3483a,a3484a,a3485a,a3486a,a3487a,a3488a,a3489a,a3490a,a3491a,a3492a,a3493a,a3494a,a3495a,a3496a,a3497a,a3498a,a3499a,a3500a,a3501a,a3502a,a3503a,a3504a,a3505a,a3506a,a3507a,a3508a,a3509a,a3510a,a3511a,a3512a,a3513a,a3514a,a3515a,a3516a,a3517a,a3518a,a3519a,a3520a,a3521a,a3522a,a3523a,a3524a,a3525a,a3526a,a3527a,a3528a,a3529a,a3530a,a3531a,a3532a,a3533a,a3534a,a3535a,a3536a,a3537a,a3538a,a3539a,a3540a,a3541a,a3542a,a3543a,a3544a,a3545a,a3546a,a3547a,a3548a,a3549a,a3550a,a3551a,a3552a,a3553a,a3554a,a3555a,a3556a,a3557a,a3558a,a3559a,a3560a,a3561a,a3562a,a3563a,a3564a,a3565a,a3566a,a3567a,a3568a,a3569a,a3570a,a3571a,a3572a,a3573a,a3574a,a3575a,a3576a,a3577a,a3578a,a3579a,a3580a,a3581a,a3582a,a3583a,a3584a,a3585a,a3586a,a3587a,a3588a,a3589a,a3590a,a3591a,a3592a,a3593a,a3594a,a3595a,a3596a,a3597a,a3598a,a3599a,a3600a,a3601a,a3602a,a3603a,a3604a,a3605a,a3606a,a3607a,a3608a,a3609a,a3610a,a3611a,a3612a,a3613a,a3614a,a3615a,a3616a,a3617a,a3618a,a3619a,a3620a,a3621a,a3622a,a3623a,a3624a,a3625a,a3626a,a3627a,a3628a,a3629a,a3630a,a3631a,a3632a,a3633a,a3634a,a3635a,a3636a,a3637a,a3638a,a3639a,a3640a,a3641a,a3642a,a3643a,a3644a,a3645a,a3646a,a3647a,a3648a,a3649a,a3650a,a3651a,a3652a,a3653a,a3654a,a3655a,a3656a,a3657a,a3658a,a3659a,a3660a,a3661a,a3662a,a3663a,a3664a,a3665a,a3666a,a3667a,a3668a,a3669a,a3670a,a3671a,a3672a,a3673a,a3674a,a3675a,a3676a,a3677a,a3678a,a3679a,a3680a,a3681a,a3682a,a3683a,a3684a,a3685a,a3686a,a3687a,a3688a,a3689a,a3690a,a3691a,a3692a,a3693a,a3694a,a3695a,a3696a,a3697a,a3698a,a3699a,a3700a,a3701a,a3702a,a3703a,a3704a,a3705a,a3706a,a3707a,a3708a,a3709a,a3710a,a3711a,a3712a,a3713a,a3714a,a3715a,a3716a,a3717a,a3718a,a3719a,a3720a,a3721a,a3722a,a3723a,a3724a,a3725a,a3726a,a3727a,a3728a,a3729a,a3730a,a3731a,a3732a,a3733a,a3734a,a3735a,a3736a,a3737a,a3738a,a3739a,a3740a,a3741a,a3742a,a3743a,a3744a,a3745a,a3746a,a3747a,a3748a,a3749a,a3750a,a3751a,a3752a,a3753a,a3754a,a3755a,a3756a,a3757a,a3758a,a3759a,a3760a,a3761a,a3762a,a3763a,a3764a,a3765a,a3766a,a3767a,a3768a,a3769a,a3770a,a3771a,a3772a,a3773a,a3774a,a3775a,a3776a,a3777a,a3778a,a3779a,a3780a,a3781a,a3782a,a3783a,a3784a,a3785a,a3786a,a3787a,a3788a,a3789a,a3790a,a3791a,a3792a,a3793a,a3794a,a3795a,a3796a,a3797a,a3798a,a3799a,a3800a,a3801a,a3802a,a3803a,a3804a,a3805a,a3806a,a3807a,a3808a,a3809a,a3810a,a3811a,a3812a,a3813a,a3814a,a3815a,a3816a,a3817a,a3818a,a3819a,a3820a,a3821a,a3822a,a3823a,a3824a,a3825a,a3826a,a3827a,a3828a,a3829a,a3830a,a3831a,a3832a,a3833a,a3834a,a3835a,a3836a,a3837a,a3838a,a3839a,a3840a,a3841a,a3842a,a3843a,a3844a,a3845a,a3846a,a3847a,a3848a,a3849a,a3850a,a3851a,a3852a,a3853a,a3854a,a3855a,a3856a,a3857a,a3858a,a3859a,a3860a,a3861a,a3862a,a3863a,a3864a,a3865a,a3866a,a3867a,a3868a,a3869a,a3870a,a3871a,a3872a,a3873a,a3874a,a3875a,a3876a,a3877a,a3878a,a3879a,a3880a,a3881a,a3882a,a3883a,a3884a,a3885a,a3886a,a3887a,a3888a,a3889a,a3890a,a3891a,a3892a,a3893a,a3894a,a3895a,a3896a,a3897a,a3898a,a3899a,a3900a,a3901a,a3902a,a3903a,a3904a,a3905a,a3906a,a3907a,a3908a,a3909a,a3910a,a3911a,a3912a,a3913a,a3914a,a3915a,a3916a,a3917a,a3918a,a3919a,a3920a,a3921a,a3922a,a3923a,a3924a,a3925a,a3926a,a3927a,a3928a,a3929a,a3930a,a3931a,a3932a,a3933a,a3934a,a3935a,a3936a,a3937a,a3938a,a3939a,a3940a,a3941a,a3942a,a3943a,a3944a,a3945a,a3946a,a3947a,a3948a,a3949a,a3950a,a3951a,a3952a,a3953a,a3954a,a3955a,a3956a,a3957a,a3958a,a3959a,a3960a,a3961a,a3962a,a3963a,a3964a,a3965a,a3966a,a3967a,a3968a,a3969a,a3970a,a3971a,a3972a,a3973a,a3974a,a3975a,a3976a,a3977a,a3978a,a3979a,a3980a,a3981a,a3982a,a3983a,a3984a,a3985a,a3986a,a3987a,a3988a,a3989a,a3990a,a3991a,a3992a,a3993a,a3994a,a3995a,a3996a,a3997a,a3998a,a3999a,a4000a,a4001a,a4002a,a4003a,a4004a,a4005a,a4006a,a4007a,a4008a,a4009a,a4010a,a4011a,a4012a,a4013a,a4014a,a4015a,a4016a,a4017a,a4018a,a4019a,a4020a,a4021a,a4022a,a4023a,a4024a,a4025a,a4026a,a4027a,a4028a,a4029a,a4030a,a4031a,a4032a,a4033a,a4034a,a4035a,a4036a,a4037a,a4038a,a4039a,a4040a,a4041a,a4042a,a4043a,a4044a,a4045a,a4046a,a4047a,a4048a,a4049a,a4050a,a4051a,a4052a,a4053a,a4054a,a4055a,a4056a,a4057a,a4058a,a4059a,a4060a,a4061a,a4062a,a4063a,a4064a,a4065a,a4066a,a4067a,a4068a,a4069a,a4070a,a4071a,a4072a,a4073a,a4074a,a4075a,a4076a,a4077a,a4078a,a4079a,a4080a,a4081a,a4082a,a4083a,a4084a,a4085a,a4086a,a4087a,a4088a,a4089a,a4090a,a4091a,a4092a,a4093a,a4094a,a4095a,a4096a,a4097a,a4098a,a4099a,a4100a,a4101a,a4102a,a4103a,a4104a,a4105a,a4106a,a4107a,a4108a,a4109a,a4110a,a4111a,a4112a,a4113a,a4114a,a4115a,a4116a,a4117a,a4118a,a4119a,a4120a,a4121a,a4122a,a4123a,a4124a,a4125a,a4126a,a4127a,a4128a,a4129a,a4130a,a4131a,a4132a,a4133a,a4134a,a4135a,a4136a,a4137a,a4138a,a4139a,a4140a,a4141a,a4142a,a4143a,a4144a,a4145a,a4146a,a4147a,a4148a,a4149a,a4150a,a4151a,a4152a,a4153a,a4154a,a4155a,a4156a,a4157a,a4158a,a4159a,a4160a,a4161a,a4162a,a4163a,a4164a,a4165a,a4166a,a4167a,a4168a,a4169a,a4170a,a4171a,a4172a,a4173a,a4174a,a4175a,a4176a,a4177a,a4178a,a4179a,a4180a,a4181a,a4182a,a4183a,a4184a,a4185a,a4186a,a4187a,a4188a,a4189a,a4190a,a4191a,a4192a,a4193a,a4194a,a4195a,a4196a,a4197a,a4198a,a4199a,a4200a,a4201a,a4202a,a4203a,a4204a,a4205a,a4206a,a4207a,a4208a,a4209a,a4210a,a4211a,a4212a,a4213a,a4214a,a4215a,a4216a,a4217a,a4218a,a4219a,a4220a,a4221a,a4222a,a4223a,a4224a,a4225a,a4226a,a4227a,a4228a,a4229a,a4230a,a4231a,a4232a,a4233a,a4234a,a4235a,a4236a,a4237a,a4238a,a4239a,a4240a,a4241a,a4242a,a4243a,a4244a,a4245a,a4246a,a4247a,a4248a,a4249a,a4250a,a4251a,a4252a,a4253a,a4254a,a4255a,a4256a,a4257a,a4258a,a4259a,a4260a,a4261a,a4262a,a4263a,a4264a,a4265a,a4266a,a4267a,a4268a,a4269a,a4270a,a4271a,a4272a,a4273a,a4274a,a4275a,a4276a,a4277a,a4278a,a4279a,a4280a,a4281a,a4282a,a4283a,a4284a,a4285a,a4286a,a4287a,a4288a,a4289a,a4290a,a4291a,a4292a,a4293a,a4294a,a4295a,a4296a,a4297a,a4298a,a4299a,a4300a,a4301a,a4302a,a4303a,a4304a,a4305a,a4306a,a4307a,a4308a,a4309a,a4310a,a4311a,a4312a,a4313a,a4314a,a4315a,a4316a,a4317a,a4318a,a4319a,a4320a,a4321a,a4322a,a4323a,a4324a,a4325a,a4326a,a4327a,a4328a,a4329a,a4330a,a4331a,a4332a,a4333a,a4334a,a4335a,a4336a,a4337a,a4338a,a4339a,a4340a,a4341a,a4342a,a4343a,a4344a,a4345a,a4346a,a4347a,a4348a,a4349a,a4350a,a4351a,a4352a,a4353a,a4354a,a4355a,a4356a,a4357a,a4358a,a4359a,a4360a,a4361a,a4362a,a4363a,a4364a,a4365a,a4366a,a4367a,a4368a,a4369a,a4370a,a4371a,a4372a,a4373a,a4374a,a4375a,a4376a,a4377a,a4378a,a4379a,a4380a,a4381a,a4382a,a4383a,a4384a,a4385a,a4386a,a4387a,a4388a,a4389a,a4390a,a4391a,a4392a,a4393a,a4394a,a4395a,a4396a,a4397a,a4398a,a4399a,a4400a,a4401a,a4402a,a4403a,a4404a,a4405a,a4406a,a4407a,a4408a,a4409a,a4410a,a4411a,a4412a,a4413a,a4414a,a4415a,a4416a,a4417a,a4418a,a4419a,a4420a,a4421a,a4422a,a4423a,a4424a,a4425a,a4426a,a4427a,a4428a,a4429a,a4430a,a4431a,a4432a,a4433a,a4434a,a4435a,a4436a,a4437a,a4438a,a4439a,a4440a,a4441a,a4442a,a4443a,a4444a,a4445a,a4446a,a4447a,a4448a,a4449a,a4450a,a4451a,a4452a,a4453a,a4454a,a4455a,a4456a,a4457a,a4458a,a4459a,a4460a,a4461a,a4462a,a4463a,a4464a,a4465a,a4466a,a4467a,a4468a,a4469a,a4470a,a4471a,a4472a,a4473a,a4474a,a4475a,a4476a,a4477a,a4478a,a4479a,a4480a,a4481a,a4482a,a4483a,a4484a,a4485a,a4486a,a4487a,a4488a,a4489a,a4490a,a4491a,a4492a,a4493a,a4494a,a4495a,a4496a,a4497a,a4498a,a4499a,a4500a,a4501a,a4502a,a4503a,a4504a,a4505a,a4506a,a4507a,a4508a,a4509a,a4510a,a4511a,a4512a,a4513a,a4514a,a4515a,a4516a,a4517a,a4518a,a4519a,a4520a,a4521a,a4522a,a4523a,a4524a,a4525a,a4526a,a4527a,a4528a,a4529a,a4530a,a4531a,a4532a,a4533a,a4534a,a4535a,a4536a,a4537a,a4538a,a4539a,a4540a,a4541a,a4542a,a4543a,a4544a,a4545a,a4546a,a4547a,a4548a,a4549a,a4550a,a4551a,a4552a,a4553a,a4554a,a4555a,a4556a,a4557a,a4558a,a4559a,a4560a,a4561a,a4562a,a4563a,a4564a,a4565a,a4566a,a4567a,a4568a,a4569a,a4570a,a4571a,a4572a,a4573a,a4574a,a4575a,a4576a,a4577a,a4578a,a4579a,a4580a,a4581a,a4582a,a4583a,a4584a,a4585a,a4586a,a4587a,a4588a,a4589a,a4590a,a4591a,a4592a,a4593a,a4594a,a4595a,a4596a,a4597a,a4598a,a4599a,a4600a,a4601a,a4602a,a4603a,a4604a,a4605a,a4606a,a4607a,a4608a,a4609a,a4610a,a4611a,a4612a,a4613a,a4614a,a4615a,a4616a,a4617a,a4618a,a4619a,a4620a,a4621a,a4622a,a4623a,a4624a,a4625a,a4626a,a4627a,a4628a,a4629a,a4630a,a4631a,a4632a,a4633a,a4634a,a4635a,a4636a,a4637a,a4638a,a4639a,a4640a,a4641a,a4642a,a4643a,a4644a,a4645a,a4646a,a4647a,a4648a,a4649a,a4650a,a4651a,a4652a,a4653a,a4654a,a4655a,a4656a,a4657a,a4658a,a4659a,a4660a,a4661a,a4662a,a4663a,a4664a,a4665a,a4666a,a4667a,a4668a,a4669a,a4670a,a4671a,a4672a,a4673a,a4674a,a4675a,a4676a,a4677a,a4678a,a4679a,a4680a,a4681a,a4682a,a4683a,a4684a,a4685a,a4686a,a4687a,a4688a,a4689a,a4690a,a4691a,a4692a,a4693a,a4694a,a4695a,a4696a,a4697a,a4698a,a4699a,a4700a,a4701a,a4702a,a4703a,a4704a,a4705a,a4706a,a4707a,a4708a,a4709a,a4710a,a4711a,a4712a,a4713a,a4714a,a4715a,a4716a,a4717a,a4718a,a4719a,a4720a,a4721a,a4722a,a4723a,a4724a,a4725a,a4726a,a4727a,a4728a,a4729a,a4730a,a4731a,a4732a,a4733a,a4734a,a4735a,a4736a,a4737a,a4738a,a4739a,a4740a,a4741a,a4742a,a4743a,a4744a,a4745a,a4746a,a4747a,a4748a,a4749a,a4750a,a4751a,a4752a,a4753a,a4754a,a4755a,a4756a,a4757a,a4758a,a4761a,a4764a,a4765a,a4768a,a4772a,a4773a,a4774a,a4775a,a4778a,a4781a,a4782a,a4785a,a4789a,a4790a,a4791a,a4792a,a4793a,a4796a,a4799a,a4800a,a4803a,a4807a,a4808a,a4809a,a4810a,a4813a,a4817a,a4818a,a4819a,a4822a,a4826a,a4827a,a4828a,a4829a,a4830a,a4831a,a4834a,a4837a,a4838a,a4841a,a4845a,a4846a,a4847a,a4848a,a4851a,a4854a,a4855a,a4858a,a4862a,a4863a,a4864a,a4865a,a4866a,a4869a,a4872a,a4873a,a4876a,a4880a,a4881a,a4882a,a4883a,a4886a,a4890a,a4891a,a4892a,a4895a,a4899a,a4900a,a4901a,a4902a,a4903a,a4904a,a4905a,a4908a,a4911a,a4912a,a4915a,a4919a,a4920a,a4921a,a4922a,a4925a,a4928a,a4929a,a4932a,a4936a,a4937a,a4938a,a4939a,a4940a,a4943a,a4946a,a4947a,a4950a,a4954a,a4955a,a4956a,a4957a,a4960a,a4964a,a4965a,a4966a,a4969a,a4973a,a4974a,a4975a,a4976a,a4977a,a4978a,a4981a,a4984a,a4985a,a4988a,a4992a,a4993a,a4994a,a4995a,a4998a,a5001a,a5002a,a5005a,a5009a,a5010a,a5011a,a5012a,a5013a,a5016a,a5019a,a5020a,a5023a,a5027a,a5028a,a5029a,a5030a,a5033a,a5037a,a5038a,a5039a,a5042a,a5046a,a5047a,a5048a,a5049a,a5050a,a5051a,a5052a,a5053a,a5056a,a5059a,a5060a,a5063a,a5067a,a5068a,a5069a,a5070a,a5073a,a5076a,a5077a,a5080a,a5084a,a5085a,a5086a,a5087a,a5088a,a5091a,a5094a,a5095a,a5098a,a5102a,a5103a,a5104a,a5105a,a5108a,a5112a,a5113a,a5114a,a5117a,a5121a,a5122a,a5123a,a5124a,a5125a,a5126a,a5129a,a5132a,a5133a,a5136a,a5140a,a5141a,a5142a,a5143a,a5146a,a5149a,a5150a,a5153a,a5157a,a5158a,a5159a,a5160a,a5161a,a5164a,a5167a,a5168a,a5171a,a5175a,a5176a,a5177a,a5178a,a5181a,a5185a,a5186a,a5187a,a5190a,a5194a,a5195a,a5196a,a5197a,a5198a,a5199a,a5200a,a5203a,a5206a,a5207a,a5210a,a5214a,a5215a,a5216a,a5217a,a5220a,a5223a,a5224a,a5227a,a5231a,a5232a,a5233a,a5234a,a5235a,a5238a,a5241a,a5242a,a5245a,a5249a,a5250a,a5251a,a5252a,a5255a,a5259a,a5260a,a5261a,a5264a,a5268a,a5269a,a5270a,a5271a,a5272a,a5273a,a5276a,a5279a,a5280a,a5283a,a5287a,a5288a,a5289a,a5290a,a5293a,a5297a,a5298a,a5299a,a5302a,a5306a,a5307a,a5308a,a5309a,a5310a,a5313a,a5316a,a5317a,a5320a,a5324a,a5325a,a5326a,a5327a,a5330a,a5334a,a5335a,a5336a,a5339a,a5343a,a5344a,a5345a,a5346a,a5347a,a5348a,a5349a,a5350a,a5351a,a5354a,a5357a,a5358a,a5361a,a5365a,a5366a,a5367a,a5368a,a5371a,a5374a,a5375a,a5378a,a5382a,a5383a,a5384a,a5385a,a5386a,a5389a,a5392a,a5393a,a5396a,a5400a,a5401a,a5402a,a5403a,a5406a,a5410a,a5411a,a5412a,a5415a,a5419a,a5420a,a5421a,a5422a,a5423a,a5424a,a5427a,a5430a,a5431a,a5434a,a5438a,a5439a,a5440a,a5441a,a5444a,a5447a,a5448a,a5451a,a5455a,a5456a,a5457a,a5458a,a5459a,a5462a,a5465a,a5466a,a5469a,a5473a,a5474a,a5475a,a5476a,a5479a,a5483a,a5484a,a5485a,a5488a,a5492a,a5493a,a5494a,a5495a,a5496a,a5497a,a5498a,a5501a,a5504a,a5505a,a5508a,a5512a,a5513a,a5514a,a5515a,a5518a,a5521a,a5522a,a5525a,a5529a,a5530a,a5531a,a5532a,a5533a,a5536a,a5539a,a5540a,a5543a,a5547a,a5548a,a5549a,a5550a,a5553a,a5557a,a5558a,a5559a,a5562a,a5566a,a5567a,a5568a,a5569a,a5570a,a5571a,a5574a,a5577a,a5578a,a5581a,a5585a,a5586a,a5587a,a5588a,a5591a,a5594a,a5595a,a5598a,a5602a,a5603a,a5604a,a5605a,a5606a,a5609a,a5612a,a5613a,a5616a,a5620a,a5621a,a5622a,a5623a,a5626a,a5630a,a5631a,a5632a,a5635a,a5639a,a5640a,a5641a,a5642a,a5643a,a5644a,a5645a,a5646a,a5649a,a5652a,a5653a,a5656a,a5660a,a5661a,a5662a,a5663a,a5666a,a5669a,a5670a,a5673a,a5677a,a5678a,a5679a,a5680a,a5681a,a5684a,a5687a,a5688a,a5691a,a5695a,a5696a,a5697a,a5698a,a5701a,a5705a,a5706a,a5707a,a5710a,a5714a,a5715a,a5716a,a5717a,a5718a,a5719a,a5722a,a5725a,a5726a,a5729a,a5733a,a5734a,a5735a,a5736a,a5739a,a5742a,a5743a,a5746a,a5750a,a5751a,a5752a,a5753a,a5754a,a5757a,a5760a,a5761a,a5764a,a5768a,a5769a,a5770a,a5771a,a5774a,a5778a,a5779a,a5780a,a5783a,a5787a,a5788a,a5789a,a5790a,a5791a,a5792a,a5793a,a5796a,a5799a,a5800a,a5803a,a5807a,a5808a,a5809a,a5810a,a5813a,a5816a,a5817a,a5820a,a5824a,a5825a,a5826a,a5827a,a5828a,a5831a,a5834a,a5835a,a5838a,a5842a,a5843a,a5844a,a5845a,a5848a,a5852a,a5853a,a5854a,a5857a,a5861a,a5862a,a5863a,a5864a,a5865a,a5866a,a5869a,a5872a,a5873a,a5876a,a5880a,a5881a,a5882a,a5883a,a5886a,a5890a,a5891a,a5892a,a5895a,a5899a,a5900a,a5901a,a5902a,a5903a,a5906a,a5909a,a5910a,a5913a,a5917a,a5918a,a5919a,a5920a,a5923a,a5927a,a5928a,a5929a,a5932a,a5936a,a5937a,a5938a,a5939a,a5940a,a5941a,a5942a,a5943a,a5944a,a5945a,a5948a,a5951a,a5952a,a5955a,a5959a,a5960a,a5961a,a5962a,a5965a,a5968a,a5969a,a5972a,a5976a,a5977a,a5978a,a5979a,a5980a,a5983a,a5986a,a5987a,a5990a,a5994a,a5995a,a5996a,a5997a,a6000a,a6004a,a6005a,a6006a,a6009a,a6013a,a6014a,a6015a,a6016a,a6017a,a6018a,a6021a,a6024a,a6025a,a6028a,a6032a,a6033a,a6034a,a6035a,a6038a,a6041a,a6042a,a6045a,a6049a,a6050a,a6051a,a6052a,a6053a,a6056a,a6059a,a6060a,a6063a,a6067a,a6068a,a6069a,a6070a,a6073a,a6077a,a6078a,a6079a,a6082a,a6086a,a6087a,a6088a,a6089a,a6090a,a6091a,a6092a,a6095a,a6098a,a6099a,a6102a,a6106a,a6107a,a6108a,a6109a,a6112a,a6115a,a6116a,a6119a,a6123a,a6124a,a6125a,a6126a,a6127a,a6130a,a6133a,a6134a,a6137a,a6141a,a6142a,a6143a,a6144a,a6147a,a6151a,a6152a,a6153a,a6156a,a6160a,a6161a,a6162a,a6163a,a6164a,a6165a,a6168a,a6171a,a6172a,a6175a,a6179a,a6180a,a6181a,a6182a,a6185a,a6188a,a6189a,a6192a,a6196a,a6197a,a6198a,a6199a,a6200a,a6203a,a6206a,a6207a,a6210a,a6214a,a6215a,a6216a,a6217a,a6220a,a6224a,a6225a,a6226a,a6229a,a6233a,a6234a,a6235a,a6236a,a6237a,a6238a,a6239a,a6240a,a6243a,a6246a,a6247a,a6250a,a6254a,a6255a,a6256a,a6257a,a6260a,a6263a,a6264a,a6267a,a6271a,a6272a,a6273a,a6274a,a6275a,a6278a,a6281a,a6282a,a6285a,a6289a,a6290a,a6291a,a6292a,a6295a,a6299a,a6300a,a6301a,a6304a,a6308a,a6309a,a6310a,a6311a,a6312a,a6313a,a6316a,a6319a,a6320a,a6323a,a6327a,a6328a,a6329a,a6330a,a6333a,a6336a,a6337a,a6340a,a6344a,a6345a,a6346a,a6347a,a6348a,a6351a,a6354a,a6355a,a6358a,a6362a,a6363a,a6364a,a6365a,a6368a,a6372a,a6373a,a6374a,a6377a,a6381a,a6382a,a6383a,a6384a,a6385a,a6386a,a6387a,a6390a,a6393a,a6394a,a6397a,a6401a,a6402a,a6403a,a6404a,a6407a,a6410a,a6411a,a6414a,a6418a,a6419a,a6420a,a6421a,a6422a,a6425a,a6428a,a6429a,a6432a,a6436a,a6437a,a6438a,a6439a,a6442a,a6446a,a6447a,a6448a,a6451a,a6455a,a6456a,a6457a,a6458a,a6459a,a6460a,a6463a,a6466a,a6467a,a6470a,a6474a,a6475a,a6476a,a6477a,a6480a,a6484a,a6485a,a6486a,a6489a,a6493a,a6494a,a6495a,a6496a,a6497a,a6500a,a6503a,a6504a,a6507a,a6511a,a6512a,a6513a,a6514a,a6517a,a6521a,a6522a,a6523a,a6526a,a6530a,a6531a,a6532a,a6533a,a6534a,a6535a,a6536a,a6537a,a6538a,a6541a,a6544a,a6545a,a6548a,a6552a,a6553a,a6554a,a6555a,a6558a,a6561a,a6562a,a6565a,a6569a,a6570a,a6571a,a6572a,a6573a,a6576a,a6579a,a6580a,a6583a,a6587a,a6588a,a6589a,a6590a,a6593a,a6597a,a6598a,a6599a,a6602a,a6606a,a6607a,a6608a,a6609a,a6610a,a6611a,a6614a,a6617a,a6618a,a6621a,a6625a,a6626a,a6627a,a6628a,a6631a,a6634a,a6635a,a6638a,a6642a,a6643a,a6644a,a6645a,a6646a,a6649a,a6652a,a6653a,a6656a,a6660a,a6661a,a6662a,a6663a,a6666a,a6670a,a6671a,a6672a,a6675a,a6679a,a6680a,a6681a,a6682a,a6683a,a6684a,a6685a,a6688a,a6691a,a6692a,a6695a,a6699a,a6700a,a6701a,a6702a,a6705a,a6708a,a6709a,a6712a,a6716a,a6717a,a6718a,a6719a,a6720a,a6723a,a6726a,a6727a,a6730a,a6734a,a6735a,a6736a,a6737a,a6740a,a6744a,a6745a,a6746a,a6749a,a6753a,a6754a,a6755a,a6756a,a6757a,a6758a,a6761a,a6764a,a6765a,a6768a,a6772a,a6773a,a6774a,a6775a,a6778a,a6782a,a6783a,a6784a,a6787a,a6791a,a6792a,a6793a,a6794a,a6795a,a6798a,a6801a,a6802a,a6805a,a6809a,a6810a,a6811a,a6812a,a6815a,a6819a,a6820a,a6821a,a6824a,a6828a,a6829a,a6830a,a6831a,a6832a,a6833a,a6834a,a6835a,a6838a,a6841a,a6842a,a6845a,a6849a,a6850a,a6851a,a6852a,a6855a,a6858a,a6859a,a6862a,a6866a,a6867a,a6868a,a6869a,a6870a,a6873a,a6876a,a6877a,a6880a,a6884a,a6885a,a6886a,a6887a,a6890a,a6894a,a6895a,a6896a,a6899a,a6903a,a6904a,a6905a,a6906a,a6907a,a6908a,a6911a,a6914a,a6915a,a6918a,a6922a,a6923a,a6924a,a6925a,a6928a,a6931a,a6932a,a6935a,a6939a,a6940a,a6941a,a6942a,a6943a,a6946a,a6949a,a6950a,a6953a,a6957a,a6958a,a6959a,a6960a,a6963a,a6967a,a6968a,a6969a,a6972a,a6976a,a6977a,a6978a,a6979a,a6980a,a6981a,a6982a,a6985a,a6988a,a6989a,a6992a,a6996a,a6997a,a6998a,a6999a,a7002a,a7005a,a7006a,a7009a,a7013a,a7014a,a7015a,a7016a,a7017a,a7020a,a7023a,a7024a,a7027a,a7031a,a7032a,a7033a,a7034a,a7037a,a7041a,a7042a,a7043a,a7046a,a7050a,a7051a,a7052a,a7053a,a7054a,a7055a,a7058a,a7061a,a7062a,a7065a,a7069a,a7070a,a7071a,a7072a,a7075a,a7079a,a7080a,a7081a,a7084a,a7088a,a7089a,a7090a,a7091a,a7092a,a7095a,a7098a,a7099a,a7102a,a7106a,a7107a,a7108a,a7109a,a7112a,a7116a,a7117a,a7118a,a7121a,a7125a,a7126a,a7127a,a7128a,a7129a,a7130a,a7131a,a7132a,a7133a,a7134a,a7135a,a7138a,a7141a,a7142a,a7145a,a7149a,a7150a,a7151a,a7152a,a7155a,a7158a,a7159a,a7162a,a7166a,a7167a,a7168a,a7169a,a7170a,a7173a,a7176a,a7177a,a7180a,a7184a,a7185a,a7186a,a7187a,a7190a,a7194a,a7195a,a7196a,a7199a,a7203a,a7204a,a7205a,a7206a,a7207a,a7208a,a7211a,a7214a,a7215a,a7218a,a7222a,a7223a,a7224a,a7225a,a7228a,a7231a,a7232a,a7235a,a7239a,a7240a,a7241a,a7242a,a7243a,a7246a,a7249a,a7250a,a7253a,a7257a,a7258a,a7259a,a7260a,a7263a,a7267a,a7268a,a7269a,a7272a,a7276a,a7277a,a7278a,a7279a,a7280a,a7281a,a7282a,a7285a,a7288a,a7289a,a7292a,a7296a,a7297a,a7298a,a7299a,a7302a,a7305a,a7306a,a7309a,a7313a,a7314a,a7315a,a7316a,a7317a,a7320a,a7323a,a7324a,a7327a,a7331a,a7332a,a7333a,a7334a,a7337a,a7341a,a7342a,a7343a,a7346a,a7350a,a7351a,a7352a,a7353a,a7354a,a7355a,a7358a,a7361a,a7362a,a7365a,a7369a,a7370a,a7371a,a7372a,a7375a,a7378a,a7379a,a7382a,a7386a,a7387a,a7388a,a7389a,a7390a,a7393a,a7396a,a7397a,a7400a,a7404a,a7405a,a7406a,a7407a,a7410a,a7414a,a7415a,a7416a,a7419a,a7423a,a7424a,a7425a,a7426a,a7427a,a7428a,a7429a,a7430a,a7433a,a7436a,a7437a,a7440a,a7444a,a7445a,a7446a,a7447a,a7450a,a7453a,a7454a,a7457a,a7461a,a7462a,a7463a,a7464a,a7465a,a7468a,a7471a,a7472a,a7475a,a7479a,a7480a,a7481a,a7482a,a7485a,a7489a,a7490a,a7491a,a7494a,a7498a,a7499a,a7500a,a7501a,a7502a,a7503a,a7506a,a7509a,a7510a,a7513a,a7517a,a7518a,a7519a,a7520a,a7523a,a7526a,a7527a,a7530a,a7534a,a7535a,a7536a,a7537a,a7538a,a7541a,a7544a,a7545a,a7548a,a7552a,a7553a,a7554a,a7555a,a7558a,a7562a,a7563a,a7564a,a7567a,a7571a,a7572a,a7573a,a7574a,a7575a,a7576a,a7577a,a7580a,a7583a,a7584a,a7587a,a7591a,a7592a,a7593a,a7594a,a7597a,a7600a,a7601a,a7604a,a7608a,a7609a,a7610a,a7611a,a7612a,a7615a,a7618a,a7619a,a7622a,a7626a,a7627a,a7628a,a7629a,a7632a,a7636a,a7637a,a7638a,a7641a,a7645a,a7646a,a7647a,a7648a,a7649a,a7650a,a7653a,a7656a,a7657a,a7660a,a7664a,a7665a,a7666a,a7667a,a7670a,a7674a,a7675a,a7676a,a7679a,a7683a,a7684a,a7685a,a7686a,a7687a,a7690a,a7693a,a7694a,a7697a,a7701a,a7702a,a7703a,a7704a,a7707a,a7711a,a7712a,a7713a,a7716a,a7720a,a7721a,a7722a,a7723a,a7724a,a7725a,a7726a,a7727a,a7728a,a7731a,a7734a,a7735a,a7738a,a7742a,a7743a,a7744a,a7745a,a7748a,a7751a,a7752a,a7755a,a7759a,a7760a,a7761a,a7762a,a7763a,a7766a,a7769a,a7770a,a7773a,a7777a,a7778a,a7779a,a7780a,a7783a,a7787a,a7788a,a7789a,a7792a,a7796a,a7797a,a7798a,a7799a,a7800a,a7801a,a7804a,a7807a,a7808a,a7811a,a7815a,a7816a,a7817a,a7818a,a7821a,a7824a,a7825a,a7828a,a7832a,a7833a,a7834a,a7835a,a7836a,a7839a,a7842a,a7843a,a7846a,a7850a,a7851a,a7852a,a7853a,a7856a,a7860a,a7861a,a7862a,a7865a,a7869a,a7870a,a7871a,a7872a,a7873a,a7874a,a7875a,a7878a,a7881a,a7882a,a7885a,a7889a,a7890a,a7891a,a7892a,a7895a,a7898a,a7899a,a7902a,a7906a,a7907a,a7908a,a7909a,a7910a,a7913a,a7916a,a7917a,a7920a,a7924a,a7925a,a7926a,a7927a,a7930a,a7934a,a7935a,a7936a,a7939a,a7943a,a7944a,a7945a,a7946a,a7947a,a7948a,a7951a,a7954a,a7955a,a7958a,a7962a,a7963a,a7964a,a7965a,a7968a,a7972a,a7973a,a7974a,a7977a,a7981a,a7982a,a7983a,a7984a,a7985a,a7988a,a7991a,a7992a,a7995a,a7999a,a8000a,a8001a,a8002a,a8005a,a8009a,a8010a,a8011a,a8014a,a8018a,a8019a,a8020a,a8021a,a8022a,a8023a,a8024a,a8025a,a8028a,a8031a,a8032a,a8035a,a8039a,a8040a,a8041a,a8042a,a8045a,a8048a,a8049a,a8052a,a8056a,a8057a,a8058a,a8059a,a8060a,a8063a,a8066a,a8067a,a8070a,a8074a,a8075a,a8076a,a8077a,a8080a,a8084a,a8085a,a8086a,a8089a,a8093a,a8094a,a8095a,a8096a,a8097a,a8098a,a8101a,a8104a,a8105a,a8108a,a8112a,a8113a,a8114a,a8115a,a8118a,a8121a,a8122a,a8125a,a8129a,a8130a,a8131a,a8132a,a8133a,a8136a,a8139a,a8140a,a8143a,a8147a,a8148a,a8149a,a8150a,a8153a,a8157a,a8158a,a8159a,a8162a,a8166a,a8167a,a8168a,a8169a,a8170a,a8171a,a8172a,a8175a,a8178a,a8179a,a8182a,a8186a,a8187a,a8188a,a8189a,a8192a,a8195a,a8196a,a8199a,a8203a,a8204a,a8205a,a8206a,a8207a,a8210a,a8213a,a8214a,a8217a,a8221a,a8222a,a8223a,a8224a,a8227a,a8231a,a8232a,a8233a,a8236a,a8240a,a8241a,a8242a,a8243a,a8244a,a8245a,a8248a,a8251a,a8252a,a8255a,a8259a,a8260a,a8261a,a8262a,a8265a,a8269a,a8270a,a8271a,a8274a,a8278a,a8279a,a8280a,a8281a,a8282a,a8285a,a8288a,a8289a,a8292a,a8296a,a8297a,a8298a,a8299a,a8302a,a8306a,a8307a,a8308a,a8311a,a8315a,a8316a,a8317a,a8318a,a8319a,a8320a,a8321a,a8322a,a8323a,a8324a,a8327a,a8330a,a8331a,a8334a,a8338a,a8339a,a8340a,a8341a,a8344a,a8347a,a8348a,a8351a,a8355a,a8356a,a8357a,a8358a,a8359a,a8362a,a8365a,a8366a,a8369a,a8373a,a8374a,a8375a,a8376a,a8379a,a8383a,a8384a,a8385a,a8388a,a8392a,a8393a,a8394a,a8395a,a8396a,a8397a,a8400a,a8403a,a8404a,a8407a,a8411a,a8412a,a8413a,a8414a,a8417a,a8420a,a8421a,a8424a,a8428a,a8429a,a8430a,a8431a,a8432a,a8435a,a8438a,a8439a,a8442a,a8446a,a8447a,a8448a,a8449a,a8452a,a8456a,a8457a,a8458a,a8461a,a8465a,a8466a,a8467a,a8468a,a8469a,a8470a,a8471a,a8474a,a8477a,a8478a,a8481a,a8485a,a8486a,a8487a,a8488a,a8491a,a8494a,a8495a,a8498a,a8502a,a8503a,a8504a,a8505a,a8506a,a8509a,a8512a,a8513a,a8516a,a8520a,a8521a,a8522a,a8523a,a8526a,a8530a,a8531a,a8532a,a8535a,a8539a,a8540a,a8541a,a8542a,a8543a,a8544a,a8547a,a8550a,a8551a,a8554a,a8558a,a8559a,a8560a,a8561a,a8564a,a8567a,a8568a,a8571a,a8575a,a8576a,a8577a,a8578a,a8579a,a8582a,a8585a,a8586a,a8589a,a8593a,a8594a,a8595a,a8596a,a8599a,a8603a,a8604a,a8605a,a8608a,a8612a,a8613a,a8614a,a8615a,a8616a,a8617a,a8618a,a8619a,a8622a,a8625a,a8626a,a8629a,a8633a,a8634a,a8635a,a8636a,a8639a,a8642a,a8643a,a8646a,a8650a,a8651a,a8652a,a8653a,a8654a,a8657a,a8660a,a8661a,a8664a,a8668a,a8669a,a8670a,a8671a,a8674a,a8678a,a8679a,a8680a,a8683a,a8687a,a8688a,a8689a,a8690a,a8691a,a8692a,a8695a,a8698a,a8699a,a8702a,a8706a,a8707a,a8708a,a8709a,a8712a,a8715a,a8716a,a8719a,a8723a,a8724a,a8725a,a8726a,a8727a,a8730a,a8733a,a8734a,a8737a,a8741a,a8742a,a8743a,a8744a,a8747a,a8751a,a8752a,a8753a,a8756a,a8760a,a8761a,a8762a,a8763a,a8764a,a8765a,a8766a,a8769a,a8772a,a8773a,a8776a,a8780a,a8781a,a8782a,a8783a,a8786a,a8789a,a8790a,a8793a,a8797a,a8798a,a8799a,a8800a,a8801a,a8804a,a8807a,a8808a,a8811a,a8815a,a8816a,a8817a,a8818a,a8821a,a8825a,a8826a,a8827a,a8830a,a8834a,a8835a,a8836a,a8837a,a8838a,a8839a,a8842a,a8845a,a8846a,a8849a,a8853a,a8854a,a8855a,a8856a,a8859a,a8863a,a8864a,a8865a,a8868a,a8872a,a8873a,a8874a,a8875a,a8876a,a8879a,a8882a,a8883a,a8886a,a8890a,a8891a,a8892a,a8893a,a8896a,a8900a,a8901a,a8902a,a8905a,a8909a,a8910a,a8911a,a8912a,a8913a,a8914a,a8915a,a8916a,a8917a,a8920a,a8923a,a8924a,a8927a,a8931a,a8932a,a8933a,a8934a,a8937a,a8940a,a8941a,a8944a,a8948a,a8949a,a8950a,a8951a,a8952a,a8955a,a8958a,a8959a,a8962a,a8966a,a8967a,a8968a,a8969a,a8972a,a8976a,a8977a,a8978a,a8981a,a8985a,a8986a,a8987a,a8988a,a8989a,a8990a,a8993a,a8996a,a8997a,a9000a,a9004a,a9005a,a9006a,a9007a,a9010a,a9013a,a9014a,a9017a,a9021a,a9022a,a9023a,a9024a,a9025a,a9028a,a9031a,a9032a,a9035a,a9039a,a9040a,a9041a,a9042a,a9045a,a9049a,a9050a,a9051a,a9054a,a9058a,a9059a,a9060a,a9061a,a9062a,a9063a,a9064a,a9067a,a9070a,a9071a,a9074a,a9078a,a9079a,a9080a,a9081a,a9084a,a9087a,a9088a,a9091a,a9095a,a9096a,a9097a,a9098a,a9099a,a9102a,a9105a,a9106a,a9109a,a9113a,a9114a,a9115a,a9116a,a9119a,a9123a,a9124a,a9125a,a9128a,a9132a,a9133a,a9134a,a9135a,a9136a,a9137a,a9140a,a9143a,a9144a,a9147a,a9151a,a9152a,a9153a,a9154a,a9157a,a9161a,a9162a,a9163a,a9166a,a9170a,a9171a,a9172a,a9173a,a9174a,a9177a,a9180a,a9181a,a9184a,a9188a,a9189a,a9190a,a9191a,a9194a,a9198a,a9199a,a9200a,a9203a,a9207a,a9208a,a9209a,a9210a,a9211a,a9212a,a9213a,a9214a,a9217a,a9220a,a9221a,a9224a,a9228a,a9229a,a9230a,a9231a,a9234a,a9237a,a9238a,a9241a,a9245a,a9246a,a9247a,a9248a,a9249a,a9252a,a9255a,a9256a,a9259a,a9263a,a9264a,a9265a,a9266a,a9269a,a9273a,a9274a,a9275a,a9278a,a9282a,a9283a,a9284a,a9285a,a9286a,a9287a,a9290a,a9293a,a9294a,a9297a,a9301a,a9302a,a9303a,a9304a,a9307a,a9310a,a9311a,a9314a,a9318a,a9319a,a9320a,a9321a,a9322a,a9325a,a9328a,a9329a,a9332a,a9336a,a9337a,a9338a,a9339a,a9342a,a9346a,a9347a,a9348a,a9351a,a9355a,a9356a,a9357a,a9358a,a9359a,a9360a,a9361a,a9364a,a9367a,a9368a,a9371a,a9375a,a9376a,a9377a,a9378a,a9381a,a9384a,a9385a,a9388a,a9392a,a9393a,a9394a,a9395a,a9396a,a9399a,a9402a,a9403a,a9406a,a9410a,a9411a,a9412a,a9413a,a9416a,a9420a,a9421a,a9422a,a9425a,a9429a,a9430a,a9431a,a9432a,a9433a,a9434a,a9437a,a9440a,a9441a,a9444a,a9448a,a9449a,a9450a,a9451a,a9454a,a9458a,a9459a,a9460a,a9463a,a9467a,a9468a,a9469a,a9470a,a9471a,a9474a,a9477a,a9478a,a9481a,a9485a,a9486a,a9487a,a9488a,a9491a,a9495a,a9496a,a9497a,a9500a,a9504a,a9505a,a9506a,a9507a,a9508a,a9509a,a9510a,a9511a,a9512a,a9513a,a9514a,a9515a,a9518a,a9521a,a9522a,a9525a,a9529a,a9530a,a9531a,a9532a,a9535a,a9538a,a9539a,a9542a,a9546a,a9547a,a9548a,a9549a,a9550a,a9553a,a9556a,a9557a,a9560a,a9564a,a9565a,a9566a,a9567a,a9570a,a9574a,a9575a,a9576a,a9579a,a9583a,a9584a,a9585a,a9586a,a9587a,a9588a,a9591a,a9594a,a9595a,a9598a,a9602a,a9603a,a9604a,a9605a,a9608a,a9611a,a9612a,a9615a,a9619a,a9620a,a9621a,a9622a,a9623a,a9626a,a9629a,a9630a,a9633a,a9637a,a9638a,a9639a,a9640a,a9643a,a9647a,a9648a,a9649a,a9652a,a9656a,a9657a,a9658a,a9659a,a9660a,a9661a,a9662a,a9665a,a9668a,a9669a,a9672a,a9676a,a9677a,a9678a,a9679a,a9682a,a9685a,a9686a,a9689a,a9693a,a9694a,a9695a,a9696a,a9697a,a9700a,a9703a,a9704a,a9707a,a9711a,a9712a,a9713a,a9714a,a9717a,a9721a,a9722a,a9723a,a9726a,a9730a,a9731a,a9732a,a9733a,a9734a,a9735a,a9738a,a9741a,a9742a,a9745a,a9749a,a9750a,a9751a,a9752a,a9755a,a9758a,a9759a,a9762a,a9766a,a9767a,a9768a,a9769a,a9770a,a9773a,a9776a,a9777a,a9780a,a9784a,a9785a,a9786a,a9787a,a9790a,a9794a,a9795a,a9796a,a9799a,a9803a,a9804a,a9805a,a9806a,a9807a,a9808a,a9809a,a9810a,a9813a,a9816a,a9817a,a9820a,a9824a,a9825a,a9826a,a9827a,a9830a,a9833a,a9834a,a9837a,a9841a,a9842a,a9843a,a9844a,a9845a,a9848a,a9851a,a9852a,a9855a,a9859a,a9860a,a9861a,a9862a,a9865a,a9869a,a9870a,a9871a,a9874a,a9878a,a9879a,a9880a,a9881a,a9882a,a9883a,a9886a,a9889a,a9890a,a9893a,a9897a,a9898a,a9899a,a9900a,a9903a,a9906a,a9907a,a9910a,a9914a,a9915a,a9916a,a9917a,a9918a,a9921a,a9924a,a9925a,a9928a,a9932a,a9933a,a9934a,a9935a,a9938a,a9942a,a9943a,a9944a,a9947a,a9951a,a9952a,a9953a,a9954a,a9955a,a9956a,a9957a,a9960a,a9963a,a9964a,a9967a,a9971a,a9972a,a9973a,a9974a,a9977a,a9980a,a9981a,a9984a,a9988a,a9989a,a9990a,a9991a,a9992a,a9995a,a9998a,a9999a,a10002a,a10006a,a10007a,a10008a,a10009a,a10012a,a10016a,a10017a,a10018a,a10021a,a10025a,a10026a,a10027a,a10028a,a10029a,a10030a,a10033a,a10036a,a10037a,a10040a,a10044a,a10045a,a10046a,a10047a,a10050a,a10054a,a10055a,a10056a,a10059a,a10063a,a10064a,a10065a,a10066a,a10067a,a10070a,a10073a,a10074a,a10077a,a10081a,a10082a,a10083a,a10084a,a10087a,a10091a,a10092a,a10093a,a10096a,a10100a,a10101a,a10102a,a10103a,a10104a,a10105a,a10106a,a10107a,a10108a,a10111a,a10114a,a10115a,a10118a,a10122a,a10123a,a10124a,a10125a,a10128a,a10131a,a10132a,a10135a,a10139a,a10140a,a10141a,a10142a,a10143a,a10146a,a10149a,a10150a,a10153a,a10157a,a10158a,a10159a,a10160a,a10163a,a10167a,a10168a,a10169a,a10172a,a10176a,a10177a,a10178a,a10179a,a10180a,a10181a,a10184a,a10187a,a10188a,a10191a,a10195a,a10196a,a10197a,a10198a,a10201a,a10204a,a10205a,a10208a,a10212a,a10213a,a10214a,a10215a,a10216a,a10219a,a10222a,a10223a,a10226a,a10230a,a10231a,a10232a,a10233a,a10236a,a10240a,a10241a,a10242a,a10245a,a10249a,a10250a,a10251a,a10252a,a10253a,a10254a,a10255a,a10258a,a10261a,a10262a,a10265a,a10269a,a10270a,a10271a,a10272a,a10275a,a10278a,a10279a,a10282a,a10286a,a10287a,a10288a,a10289a,a10290a,a10293a,a10296a,a10297a,a10300a,a10304a,a10305a,a10306a,a10307a,a10310a,a10314a,a10315a,a10316a,a10319a,a10323a,a10324a,a10325a,a10326a,a10327a,a10328a,a10331a,a10334a,a10335a,a10338a,a10342a,a10343a,a10344a,a10345a,a10348a,a10351a,a10352a,a10355a,a10359a,a10360a,a10361a,a10362a,a10363a,a10366a,a10369a,a10370a,a10373a,a10377a,a10378a,a10379a,a10380a,a10383a,a10387a,a10388a,a10389a,a10392a,a10396a,a10397a,a10398a,a10399a,a10400a,a10401a,a10402a,a10403a,a10406a,a10409a,a10410a,a10413a,a10417a,a10418a,a10419a,a10420a,a10423a,a10426a,a10427a,a10430a,a10434a,a10435a,a10436a,a10437a,a10438a,a10441a,a10444a,a10445a,a10448a,a10452a,a10453a,a10454a,a10455a,a10458a,a10462a,a10463a,a10464a,a10467a,a10471a,a10472a,a10473a,a10474a,a10475a,a10476a,a10479a,a10482a,a10483a,a10486a,a10490a,a10491a,a10492a,a10493a,a10496a,a10499a,a10500a,a10503a,a10507a,a10508a,a10509a,a10510a,a10511a,a10514a,a10517a,a10518a,a10521a,a10525a,a10526a,a10527a,a10528a,a10531a,a10535a,a10536a,a10537a,a10540a,a10544a,a10545a,a10546a,a10547a,a10548a,a10549a,a10550a,a10553a,a10556a,a10557a,a10560a,a10564a,a10565a,a10566a,a10567a,a10570a,a10573a,a10574a,a10577a,a10581a,a10582a,a10583a,a10584a,a10585a,a10588a,a10591a,a10592a,a10595a,a10599a,a10600a,a10601a,a10602a,a10605a,a10609a,a10610a,a10611a,a10614a,a10618a,a10619a,a10620a,a10621a,a10622a,a10623a,a10626a,a10629a,a10630a,a10633a,a10637a,a10638a,a10639a,a10640a,a10643a,a10647a,a10648a,a10649a,a10652a,a10656a,a10657a,a10658a,a10659a,a10660a,a10663a,a10666a,a10667a,a10670a,a10674a,a10675a,a10676a,a10677a,a10680a,a10684a,a10685a,a10686a,a10689a,a10693a,a10694a,a10695a,a10696a,a10697a,a10698a,a10699a,a10700a,a10701a,a10702a,a10705a,a10708a,a10709a,a10712a,a10716a,a10717a,a10718a,a10719a,a10722a,a10725a,a10726a,a10729a,a10733a,a10734a,a10735a,a10736a,a10737a,a10740a,a10743a,a10744a,a10747a,a10751a,a10752a,a10753a,a10754a,a10757a,a10761a,a10762a,a10763a,a10766a,a10770a,a10771a,a10772a,a10773a,a10774a,a10775a,a10778a,a10781a,a10782a,a10785a,a10789a,a10790a,a10791a,a10792a,a10795a,a10798a,a10799a,a10802a,a10806a,a10807a,a10808a,a10809a,a10810a,a10813a,a10816a,a10817a,a10820a,a10824a,a10825a,a10826a,a10827a,a10830a,a10834a,a10835a,a10836a,a10839a,a10843a,a10844a,a10845a,a10846a,a10847a,a10848a,a10849a,a10852a,a10855a,a10856a,a10859a,a10863a,a10864a,a10865a,a10866a,a10869a,a10872a,a10873a,a10876a,a10880a,a10881a,a10882a,a10883a,a10884a,a10887a,a10890a,a10891a,a10894a,a10898a,a10899a,a10900a,a10901a,a10904a,a10908a,a10909a,a10910a,a10913a,a10917a,a10918a,a10919a,a10920a,a10921a,a10922a,a10925a,a10928a,a10929a,a10932a,a10936a,a10937a,a10938a,a10939a,a10942a,a10945a,a10946a,a10949a,a10953a,a10954a,a10955a,a10956a,a10957a,a10960a,a10963a,a10964a,a10967a,a10971a,a10972a,a10973a,a10974a,a10977a,a10981a,a10982a,a10983a,a10986a,a10990a,a10991a,a10992a,a10993a,a10994a,a10995a,a10996a,a10997a,a11000a,a11003a,a11004a,a11007a,a11011a,a11012a,a11013a,a11014a,a11017a,a11020a,a11021a,a11024a,a11028a,a11029a,a11030a,a11031a,a11032a,a11035a,a11038a,a11039a,a11042a,a11046a,a11047a,a11048a,a11049a,a11052a,a11056a,a11057a,a11058a,a11061a,a11065a,a11066a,a11067a,a11068a,a11069a,a11070a,a11073a,a11076a,a11077a,a11080a,a11084a,a11085a,a11086a,a11087a,a11090a,a11093a,a11094a,a11097a,a11101a,a11102a,a11103a,a11104a,a11105a,a11108a,a11111a,a11112a,a11115a,a11119a,a11120a,a11121a,a11122a,a11125a,a11129a,a11130a,a11131a,a11134a,a11138a,a11139a,a11140a,a11141a,a11142a,a11143a,a11144a,a11147a,a11150a,a11151a,a11154a,a11158a,a11159a,a11160a,a11161a,a11164a,a11167a,a11168a,a11171a,a11175a,a11176a,a11177a,a11178a,a11179a,a11182a,a11185a,a11186a,a11189a,a11193a,a11194a,a11195a,a11196a,a11199a,a11203a,a11204a,a11205a,a11208a,a11212a,a11213a,a11214a,a11215a,a11216a,a11217a,a11220a,a11223a,a11224a,a11227a,a11231a,a11232a,a11233a,a11234a,a11237a,a11241a,a11242a,a11243a,a11246a,a11250a,a11251a,a11252a,a11253a,a11254a,a11257a,a11260a,a11261a,a11264a,a11268a,a11269a,a11270a,a11271a,a11274a,a11278a,a11279a,a11280a,a11283a,a11287a,a11288a,a11289a,a11290a,a11291a,a11292a,a11293a,a11294a,a11295a,a11298a,a11301a,a11302a,a11305a,a11309a,a11310a,a11311a,a11312a,a11315a,a11318a,a11319a,a11322a,a11326a,a11327a,a11328a,a11329a,a11330a,a11333a,a11336a,a11337a,a11340a,a11344a,a11345a,a11346a,a11347a,a11350a,a11354a,a11355a,a11356a,a11359a,a11363a,a11364a,a11365a,a11366a,a11367a,a11368a,a11371a,a11374a,a11375a,a11378a,a11382a,a11383a,a11384a,a11385a,a11388a,a11391a,a11392a,a11395a,a11399a,a11400a,a11401a,a11402a,a11403a,a11406a,a11409a,a11410a,a11413a,a11417a,a11418a,a11419a,a11420a,a11423a,a11427a,a11428a,a11429a,a11432a,a11436a,a11437a,a11438a,a11439a,a11440a,a11441a,a11442a,a11445a,a11448a,a11449a,a11452a,a11456a,a11457a,a11458a,a11459a,a11462a,a11465a,a11466a,a11469a,a11473a,a11474a,a11475a,a11476a,a11477a,a11480a,a11483a,a11484a,a11487a,a11491a,a11492a,a11493a,a11494a,a11497a,a11501a,a11502a,a11503a,a11506a,a11510a,a11511a,a11512a,a11513a,a11514a,a11515a,a11518a,a11521a,a11522a,a11525a,a11529a,a11530a,a11531a,a11532a,a11535a,a11539a,a11540a,a11541a,a11544a,a11548a,a11549a,a11550a,a11551a,a11552a,a11555a,a11558a,a11559a,a11562a,a11566a,a11567a,a11568a,a11569a,a11572a,a11576a,a11577a,a11578a,a11581a,a11585a,a11586a,a11587a,a11588a,a11589a,a11590a,a11591a,a11592a,a11595a,a11598a,a11599a,a11602a,a11606a,a11607a,a11608a,a11609a,a11612a,a11615a,a11616a,a11619a,a11623a,a11624a,a11625a,a11626a,a11627a,a11630a,a11633a,a11634a,a11637a,a11641a,a11642a,a11643a,a11644a,a11647a,a11651a,a11652a,a11653a,a11656a,a11660a,a11661a,a11662a,a11663a,a11664a,a11665a,a11668a,a11671a,a11672a,a11675a,a11679a,a11680a,a11681a,a11682a,a11685a,a11688a,a11689a,a11692a,a11696a,a11697a,a11698a,a11699a,a11700a,a11703a,a11706a,a11707a,a11710a,a11714a,a11715a,a11716a,a11717a,a11720a,a11724a,a11725a,a11726a,a11729a,a11733a,a11734a,a11735a,a11736a,a11737a,a11738a,a11739a,a11742a,a11745a,a11746a,a11749a,a11753a,a11754a,a11755a,a11756a,a11759a,a11762a,a11763a,a11766a,a11770a,a11771a,a11772a,a11773a,a11774a,a11777a,a11780a,a11781a,a11784a,a11788a,a11789a,a11790a,a11791a,a11794a,a11798a,a11799a,a11800a,a11803a,a11807a,a11808a,a11809a,a11810a,a11811a,a11812a,a11815a,a11818a,a11819a,a11822a,a11826a,a11827a,a11828a,a11829a,a11832a,a11836a,a11837a,a11838a,a11841a,a11845a,a11846a,a11847a,a11848a,a11849a,a11852a,a11855a,a11856a,a11859a,a11863a,a11864a,a11865a,a11866a,a11869a,a11873a,a11874a,a11875a,a11878a,a11882a,a11883a,a11884a,a11885a,a11886a,a11887a,a11888a,a11889a,a11890a,a11891a,a11892a,a11895a,a11898a,a11899a,a11902a,a11906a,a11907a,a11908a,a11909a,a11912a,a11915a,a11916a,a11919a,a11923a,a11924a,a11925a,a11926a,a11927a,a11930a,a11933a,a11934a,a11937a,a11941a,a11942a,a11943a,a11944a,a11947a,a11951a,a11952a,a11953a,a11956a,a11960a,a11961a,a11962a,a11963a,a11964a,a11965a,a11968a,a11971a,a11972a,a11975a,a11979a,a11980a,a11981a,a11982a,a11985a,a11988a,a11989a,a11992a,a11996a,a11997a,a11998a,a11999a,a12000a,a12003a,a12006a,a12007a,a12010a,a12014a,a12015a,a12016a,a12017a,a12020a,a12024a,a12025a,a12026a,a12029a,a12033a,a12034a,a12035a,a12036a,a12037a,a12038a,a12039a,a12042a,a12045a,a12046a,a12049a,a12053a,a12054a,a12055a,a12056a,a12059a,a12062a,a12063a,a12066a,a12070a,a12071a,a12072a,a12073a,a12074a,a12077a,a12080a,a12081a,a12084a,a12088a,a12089a,a12090a,a12091a,a12094a,a12098a,a12099a,a12100a,a12103a,a12107a,a12108a,a12109a,a12110a,a12111a,a12112a,a12115a,a12118a,a12119a,a12122a,a12126a,a12127a,a12128a,a12129a,a12132a,a12135a,a12136a,a12139a,a12143a,a12144a,a12145a,a12146a,a12147a,a12150a,a12153a,a12154a,a12157a,a12161a,a12162a,a12163a,a12164a,a12167a,a12171a,a12172a,a12173a,a12176a,a12180a,a12181a,a12182a,a12183a,a12184a,a12185a,a12186a,a12187a,a12190a,a12193a,a12194a,a12197a,a12201a,a12202a,a12203a,a12204a,a12207a,a12210a,a12211a,a12214a,a12218a,a12219a,a12220a,a12221a,a12222a,a12225a,a12228a,a12229a,a12232a,a12236a,a12237a,a12238a,a12239a,a12242a,a12246a,a12247a,a12248a,a12251a,a12255a,a12256a,a12257a,a12258a,a12259a,a12260a,a12263a,a12266a,a12267a,a12270a,a12274a,a12275a,a12276a,a12277a,a12280a,a12283a,a12284a,a12287a,a12291a,a12292a,a12293a,a12294a,a12295a,a12298a,a12301a,a12302a,a12305a,a12309a,a12310a,a12311a,a12312a,a12315a,a12319a,a12320a,a12321a,a12324a,a12328a,a12329a,a12330a,a12331a,a12332a,a12333a,a12334a,a12337a,a12340a,a12341a,a12344a,a12348a,a12349a,a12350a,a12351a,a12354a,a12357a,a12358a,a12361a,a12365a,a12366a,a12367a,a12368a,a12369a,a12372a,a12375a,a12376a,a12379a,a12383a,a12384a,a12385a,a12386a,a12389a,a12393a,a12394a,a12395a,a12398a,a12402a,a12403a,a12404a,a12405a,a12406a,a12407a,a12410a,a12413a,a12414a,a12417a,a12421a,a12422a,a12423a,a12424a,a12427a,a12431a,a12432a,a12433a,a12436a,a12440a,a12441a,a12442a,a12443a,a12444a,a12447a,a12450a,a12451a,a12454a,a12458a,a12459a,a12460a,a12461a,a12464a,a12468a,a12469a,a12470a,a12473a,a12477a,a12478a,a12479a,a12480a,a12481a,a12482a,a12483a,a12484a,a12485a,a12488a,a12491a,a12492a,a12495a,a12499a,a12500a,a12501a,a12502a,a12505a,a12508a,a12509a,a12512a,a12516a,a12517a,a12518a,a12519a,a12520a,a12523a,a12526a,a12527a,a12530a,a12534a,a12535a,a12536a,a12537a,a12540a,a12544a,a12545a,a12546a,a12549a,a12553a,a12554a,a12555a,a12556a,a12557a,a12558a,a12561a,a12564a,a12565a,a12568a,a12572a,a12573a,a12574a,a12575a,a12578a,a12581a,a12582a,a12585a,a12589a,a12590a,a12591a,a12592a,a12593a,a12596a,a12599a,a12600a,a12603a,a12607a,a12608a,a12609a,a12610a,a12613a,a12617a,a12618a,a12619a,a12622a,a12626a,a12627a,a12628a,a12629a,a12630a,a12631a,a12632a,a12635a,a12638a,a12639a,a12642a,a12646a,a12647a,a12648a,a12649a,a12652a,a12655a,a12656a,a12659a,a12663a,a12664a,a12665a,a12666a,a12667a,a12670a,a12673a,a12674a,a12677a,a12681a,a12682a,a12683a,a12684a,a12687a,a12691a,a12692a,a12693a,a12696a,a12700a,a12701a,a12702a,a12703a,a12704a,a12705a,a12708a,a12711a,a12712a,a12715a,a12719a,a12720a,a12721a,a12722a,a12725a,a12729a,a12730a,a12731a,a12734a,a12738a,a12739a,a12740a,a12741a,a12742a,a12745a,a12748a,a12749a,a12752a,a12756a,a12757a,a12758a,a12759a,a12762a,a12766a,a12767a,a12768a,a12771a,a12775a,a12776a,a12777a,a12778a,a12779a,a12780a,a12781a,a12782a,a12785a,a12788a,a12789a,a12792a,a12796a,a12797a,a12798a,a12799a,a12802a,a12805a,a12806a,a12809a,a12813a,a12814a,a12815a,a12816a,a12817a,a12820a,a12823a,a12824a,a12827a,a12831a,a12832a,a12833a,a12834a,a12837a,a12841a,a12842a,a12843a,a12846a,a12850a,a12851a,a12852a,a12853a,a12854a,a12855a,a12858a,a12861a,a12862a,a12865a,a12869a,a12870a,a12871a,a12872a,a12875a,a12878a,a12879a,a12882a,a12886a,a12887a,a12888a,a12889a,a12890a,a12893a,a12896a,a12897a,a12900a,a12904a,a12905a,a12906a,a12907a,a12910a,a12914a,a12915a,a12916a,a12919a,a12923a,a12924a,a12925a,a12926a,a12927a,a12928a,a12929a,a12932a,a12935a,a12936a,a12939a,a12943a,a12944a,a12945a,a12946a,a12949a,a12952a,a12953a,a12956a,a12960a,a12961a,a12962a,a12963a,a12964a,a12967a,a12970a,a12971a,a12974a,a12978a,a12979a,a12980a,a12981a,a12984a,a12988a,a12989a,a12990a,a12993a,a12997a,a12998a,a12999a,a13000a,a13001a,a13002a,a13005a,a13008a,a13009a,a13012a,a13016a,a13017a,a13018a,a13019a,a13022a,a13026a,a13027a,a13028a,a13031a,a13035a,a13036a,a13037a,a13038a,a13039a,a13042a,a13045a,a13046a,a13049a,a13053a,a13054a,a13055a,a13056a,a13059a,a13063a,a13064a,a13065a,a13068a,a13072a,a13073a,a13074a,a13075a,a13076a,a13077a,a13078a,a13079a,a13080a,a13081a,a13084a,a13087a,a13088a,a13091a,a13095a,a13096a,a13097a,a13098a,a13101a,a13104a,a13105a,a13108a,a13112a,a13113a,a13114a,a13115a,a13116a,a13119a,a13122a,a13123a,a13126a,a13130a,a13131a,a13132a,a13133a,a13136a,a13140a,a13141a,a13142a,a13145a,a13149a,a13150a,a13151a,a13152a,a13153a,a13154a,a13157a,a13160a,a13161a,a13164a,a13168a,a13169a,a13170a,a13171a,a13174a,a13177a,a13178a,a13181a,a13185a,a13186a,a13187a,a13188a,a13189a,a13192a,a13195a,a13196a,a13199a,a13203a,a13204a,a13205a,a13206a,a13209a,a13213a,a13214a,a13215a,a13218a,a13222a,a13223a,a13224a,a13225a,a13226a,a13227a,a13228a,a13231a,a13234a,a13235a,a13238a,a13242a,a13243a,a13244a,a13245a,a13248a,a13251a,a13252a,a13255a,a13259a,a13260a,a13261a,a13262a,a13263a,a13266a,a13269a,a13270a,a13273a,a13277a,a13278a,a13279a,a13280a,a13283a,a13287a,a13288a,a13289a,a13292a,a13296a,a13297a,a13298a,a13299a,a13300a,a13301a,a13304a,a13307a,a13308a,a13311a,a13315a,a13316a,a13317a,a13318a,a13321a,a13324a,a13325a,a13328a,a13332a,a13333a,a13334a,a13335a,a13336a,a13339a,a13342a,a13343a,a13346a,a13350a,a13351a,a13352a,a13353a,a13356a,a13360a,a13361a,a13362a,a13365a,a13369a,a13370a,a13371a,a13372a,a13373a,a13374a,a13375a,a13376a,a13379a,a13382a,a13383a,a13386a,a13390a,a13391a,a13392a,a13393a,a13396a,a13399a,a13400a,a13403a,a13407a,a13408a,a13409a,a13410a,a13411a,a13414a,a13417a,a13418a,a13421a,a13425a,a13426a,a13427a,a13428a,a13431a,a13435a,a13436a,a13437a,a13440a,a13444a,a13445a,a13446a,a13447a,a13448a,a13449a,a13452a,a13455a,a13456a,a13459a,a13463a,a13464a,a13465a,a13466a,a13469a,a13472a,a13473a,a13476a,a13480a,a13481a,a13482a,a13483a,a13484a,a13487a,a13490a,a13491a,a13494a,a13498a,a13499a,a13500a,a13501a,a13504a,a13508a,a13509a,a13510a,a13513a,a13517a,a13518a,a13519a,a13520a,a13521a,a13522a,a13523a,a13526a,a13529a,a13530a,a13533a,a13537a,a13538a,a13539a,a13540a,a13543a,a13546a,a13547a,a13550a,a13554a,a13555a,a13556a,a13557a,a13558a,a13561a,a13564a,a13565a,a13568a,a13572a,a13573a,a13574a,a13575a,a13578a,a13582a,a13583a,a13584a,a13587a,a13591a,a13592a,a13593a,a13594a,a13595a,a13596a,a13599a,a13602a,a13603a,a13606a,a13610a,a13611a,a13612a,a13613a,a13616a,a13620a,a13621a,a13622a,a13625a,a13629a,a13630a,a13631a,a13632a,a13633a,a13636a,a13639a,a13640a,a13643a,a13647a,a13648a,a13649a,a13650a,a13653a,a13657a,a13658a,a13659a,a13662a,a13666a,a13667a,a13668a,a13669a,a13670a,a13671a,a13672a,a13673a,a13674a,a13677a,a13680a,a13681a,a13684a,a13688a,a13689a,a13690a,a13691a,a13694a,a13697a,a13698a,a13701a,a13705a,a13706a,a13707a,a13708a,a13709a,a13712a,a13715a,a13716a,a13719a,a13723a,a13724a,a13725a,a13726a,a13729a,a13733a,a13734a,a13735a,a13738a,a13742a,a13743a,a13744a,a13745a,a13746a,a13747a,a13750a,a13753a,a13754a,a13757a,a13761a,a13762a,a13763a,a13764a,a13767a,a13770a,a13771a,a13774a,a13778a,a13779a,a13780a,a13781a,a13782a,a13785a,a13788a,a13789a,a13792a,a13796a,a13797a,a13798a,a13799a,a13802a,a13806a,a13807a,a13808a,a13811a,a13815a,a13816a,a13817a,a13818a,a13819a,a13820a,a13821a,a13824a,a13827a,a13828a,a13831a,a13835a,a13836a,a13837a,a13838a,a13841a,a13844a,a13845a,a13848a,a13852a,a13853a,a13854a,a13855a,a13856a,a13859a,a13862a,a13863a,a13866a,a13870a,a13871a,a13872a,a13873a,a13876a,a13880a,a13881a,a13882a,a13885a,a13889a,a13890a,a13891a,a13892a,a13893a,a13894a,a13897a,a13900a,a13901a,a13904a,a13908a,a13909a,a13910a,a13911a,a13914a,a13918a,a13919a,a13920a,a13923a,a13927a,a13928a,a13929a,a13930a,a13931a,a13934a,a13937a,a13938a,a13941a,a13945a,a13946a,a13947a,a13948a,a13951a,a13955a,a13956a,a13957a,a13960a,a13964a,a13965a,a13966a,a13967a,a13968a,a13969a,a13970a,a13971a,a13974a,a13977a,a13978a,a13981a,a13985a,a13986a,a13987a,a13988a,a13991a,a13994a,a13995a,a13998a,a14002a,a14003a,a14004a,a14005a,a14006a,a14009a,a14012a,a14013a,a14016a,a14020a,a14021a,a14022a,a14023a,a14026a,a14030a,a14031a,a14032a,a14035a,a14039a,a14040a,a14041a,a14042a,a14043a,a14044a,a14047a,a14050a,a14051a,a14054a,a14058a,a14059a,a14060a,a14061a,a14064a,a14067a,a14068a,a14071a,a14075a,a14076a,a14077a,a14078a,a14079a,a14082a,a14085a,a14086a,a14089a,a14093a,a14094a,a14095a,a14096a,a14099a,a14103a,a14104a,a14105a,a14108a,a14112a,a14113a,a14114a,a14115a,a14116a,a14117a,a14118a,a14121a,a14124a,a14125a,a14128a,a14132a,a14133a,a14134a,a14135a,a14138a,a14141a,a14142a,a14145a,a14149a,a14150a,a14151a,a14152a,a14153a,a14156a,a14159a,a14160a,a14163a,a14167a,a14168a,a14169a,a14170a,a14173a,a14177a,a14178a,a14179a,a14182a,a14186a,a14187a,a14188a,a14189a,a14190a,a14191a,a14194a,a14197a,a14198a,a14201a,a14205a,a14206a,a14207a,a14208a,a14211a,a14215a,a14216a,a14217a,a14220a,a14224a,a14225a,a14226a,a14227a,a14228a,a14231a,a14234a,a14235a,a14238a,a14242a,a14243a,a14244a,a14245a,a14248a,a14252a,a14253a,a14254a,a14257a,a14261a,a14262a,a14263a,a14264a,a14265a,a14266a,a14267a,a14268a,a14269a,a14270a,a14271a,a14272a,a14275a,a14278a,a14281a,a14284a,a14287a,a14290a,a14293a,a14296a,a14299a,a14302a,a14305a,a14308a,a14312a,a14313a,a14317a,a14318a,a14322a,a14323a,a14327a,a14328a,a14332a,a14333a,a14337a,a14338a,a14342a,a14343a,a14347a,a14348a,a14352a,a14353a,a14357a,a14358a,a14362a,a14363a,a14367a,a14368a,a14372a,a14373a,a14377a,a14378a,a14382a,a14383a,a14387a,a14388a,a14392a,a14393a,a14397a,a14398a,a14402a,a14403a,a14407a,a14408a,a14412a,a14413a,a14417a,a14418a,a14422a,a14423a,a14427a,a14428a,a14432a,a14433a,a14437a,a14438a,a14442a,a14443a,a14447a,a14448a,a14452a,a14453a,a14457a,a14458a,a14462a,a14463a,a14467a,a14468a,a14472a,a14473a,a14477a,a14478a,a14482a,a14483a,a14487a,a14488a,a14492a,a14493a,a14497a,a14498a,a14502a,a14503a,a14507a,a14508a,a14512a,a14513a,a14517a,a14518a,a14522a,a14523a,a14527a,a14528a,a14532a,a14533a,a14537a,a14538a,a14542a,a14543a,a14547a,a14548a,a14551a,a14554a,a14555a,a14558a,a14561a,a14562a,a14565a,a14568a,a14569a,a14572a,a14575a,a14576a,a14579a,a14582a,a14583a,a14586a,a14589a,a14590a,a14593a,a14596a,a14597a,a14600a,a14603a,a14604a,a14607a,a14610a,a14611a,a14614a,a14617a,a14618a,a14621a,a14624a,a14625a,a14628a,a14631a,a14632a,a14635a,a14638a,a14639a,a14642a,a14645a,a14646a,a14649a,a14652a,a14653a,a14656a,a14659a,a14660a,a14663a,a14666a,a14667a,a14670a,a14673a,a14674a,a14677a,a14680a,a14681a,a14684a,a14687a,a14688a,a14691a,a14694a,a14695a,a14698a,a14701a,a14702a,a14705a,a14708a,a14709a,a14712a,a14715a,a14716a,a14719a,a14722a,a14723a,a14726a,a14729a,a14730a,a14733a,a14736a,a14737a,a14740a,a14743a,a14744a,a14747a,a14750a,a14751a,a14754a,a14757a,a14758a,a14761a,a14764a,a14765a,a14768a,a14771a,a14772a,a14775a,a14778a,a14779a,a14782a,a14785a,a14786a,a14789a,a14792a,a14793a,a14796a,a14799a,a14800a,a14803a,a14806a,a14807a,a14810a,a14813a,a14814a,a14817a,a14820a,a14821a,a14824a,a14827a,a14828a,a14831a,a14834a,a14835a,a14838a,a14841a,a14842a,a14845a,a14848a,a14849a,a14852a,a14855a,a14856a,a14859a,a14862a,a14863a,a14866a,a14869a,a14870a,a14873a,a14876a,a14877a,a14880a,a14883a,a14884a,a14887a,a14890a,a14891a,a14894a,a14898a,a14899a,a14900a,a14903a,a14906a,a14907a,a14910a,a14914a,a14915a,a14916a,a14919a,a14922a,a14923a,a14926a,a14930a,a14931a,a14932a,a14935a,a14938a,a14939a,a14942a,a14946a,a14947a,a14948a,a14951a,a14954a,a14955a,a14958a,a14962a,a14963a,a14964a,a14967a,a14970a,a14971a,a14974a,a14978a,a14979a,a14980a,a14983a,a14986a,a14987a,a14990a,a14994a,a14995a,a14996a,a14999a,a15002a,a15003a,a15006a,a15010a,a15011a,a15012a,a15015a,a15018a,a15019a,a15022a,a15026a,a15027a,a15028a,a15031a,a15034a,a15035a,a15038a,a15042a,a15043a,a15044a,a15047a,a15050a,a15051a,a15054a,a15058a,a15059a,a15060a,a15063a,a15066a,a15067a,a15070a,a15074a,a15075a,a15076a,a15079a,a15082a,a15083a,a15086a,a15090a,a15091a,a15092a,a15095a,a15098a,a15099a,a15102a,a15106a,a15107a,a15108a,a15111a,a15114a,a15115a,a15118a,a15122a,a15123a,a15124a,a15127a,a15130a,a15131a,a15134a,a15138a,a15139a,a15140a,a15143a,a15146a,a15147a,a15150a,a15154a,a15155a,a15156a,a15159a,a15162a,a15163a,a15166a,a15170a,a15171a,a15172a,a15175a,a15178a,a15179a,a15182a,a15186a,a15187a,a15188a,a15191a,a15194a,a15195a,a15198a,a15202a,a15203a,a15204a,a15207a,a15210a,a15211a,a15214a,a15218a,a15219a,a15220a,a15223a,a15226a,a15227a,a15230a,a15234a,a15235a,a15236a,a15239a,a15242a,a15243a,a15246a,a15250a,a15251a,a15252a,a15255a,a15258a,a15259a,a15262a,a15266a,a15267a,a15268a,a15271a,a15274a,a15275a,a15278a,a15282a,a15283a,a15284a,a15287a,a15290a,a15291a,a15294a,a15298a,a15299a,a15300a,a15303a,a15306a,a15307a,a15310a,a15314a,a15315a,a15316a,a15319a,a15322a,a15323a,a15326a,a15330a,a15331a,a15332a,a15335a,a15338a,a15339a,a15342a,a15346a,a15347a,a15348a,a15351a,a15354a,a15355a,a15358a,a15362a,a15363a,a15364a,a15367a,a15370a,a15371a,a15374a,a15378a,a15379a,a15380a,a15383a,a15386a,a15387a,a15390a,a15394a,a15395a,a15396a,a15399a,a15403a,a15404a,a15405a,a15408a,a15412a,a15413a,a15414a,a15417a,a15421a,a15422a,a15423a,a15426a,a15430a,a15431a,a15432a,a15435a,a15439a,a15440a,a15441a,a15444a,a15448a,a15449a,a15450a,a15453a,a15457a,a15458a,a15459a,a15462a,a15466a,a15467a,a15468a,a15471a,a15475a,a15476a,a15477a,a15480a,a15484a,a15485a,a15486a,a15489a,a15493a,a15494a,a15495a,a15498a,a15502a,a15503a,a15504a,a15507a,a15511a,a15512a,a15513a,a15516a,a15520a,a15521a,a15522a,a15525a,a15529a,a15530a,a15531a,a15534a,a15538a,a15539a,a15540a,a15543a,a15547a,a15548a,a15549a,a15552a,a15556a,a15557a,a15558a,a15561a,a15565a,a15566a,a15567a,a15570a,a15574a,a15575a,a15576a,a15579a,a15583a,a15584a,a15585a,a15588a,a15592a,a15593a,a15594a,a15597a,a15601a,a15602a,a15603a,a15606a,a15610a,a15611a,a15612a,a15615a,a15619a,a15620a,a15621a,a15624a,a15628a,a15629a,a15630a,a15633a,a15637a,a15638a,a15639a,a15642a,a15646a,a15647a,a15648a,a15651a,a15655a,a15656a,a15657a,a15660a,a15664a,a15665a,a15666a,a15669a,a15673a,a15674a,a15675a,a15678a,a15682a,a15683a,a15684a,a15687a,a15691a,a15692a,a15693a,a15696a,a15700a,a15701a,a15702a,a15705a,a15709a,a15710a,a15711a,a15714a,a15718a,a15719a,a15720a,a15723a,a15727a,a15728a,a15729a,a15732a,a15736a,a15737a,a15738a,a15741a,a15745a,a15746a,a15747a,a15750a,a15754a,a15755a,a15756a,a15759a,a15763a,a15764a,a15765a,a15768a,a15772a,a15773a,a15774a,a15777a,a15781a,a15782a,a15783a,a15786a,a15790a,a15791a,a15792a,a15795a,a15799a,a15800a,a15801a,a15804a,a15808a,a15809a,a15810a,a15813a,a15817a,a15818a,a15819a,a15822a,a15826a,a15827a,a15828a,a15831a,a15835a,a15836a,a15837a,a15840a,a15844a,a15845a,a15846a,a15849a,a15853a,a15854a,a15855a,a15858a,a15862a,a15863a,a15864a,a15867a,a15871a,a15872a,a15873a,a15876a,a15880a,a15881a,a15882a,a15885a,a15889a,a15890a,a15891a,a15894a,a15898a,a15899a,a15900a,a15903a,a15907a,a15908a,a15909a,a15912a,a15916a,a15917a,a15918a,a15921a,a15925a,a15926a,a15927a,a15930a,a15934a,a15935a,a15936a,a15939a,a15943a,a15944a,a15945a,a15948a,a15952a,a15953a,a15954a,a15957a,a15961a,a15962a,a15963a,a15966a,a15970a,a15971a,a15972a,a15975a,a15979a,a15980a,a15981a,a15984a,a15988a,a15989a,a15990a,a15993a,a15997a,a15998a,a15999a,a16002a,a16006a,a16007a,a16008a,a16011a,a16015a,a16016a,a16017a,a16020a,a16024a,a16025a,a16026a,a16029a,a16033a,a16034a,a16035a,a16038a,a16042a,a16043a,a16044a,a16047a,a16051a,a16052a,a16053a,a16056a,a16060a,a16061a,a16062a,a16065a,a16069a,a16070a,a16071a,a16074a,a16078a,a16079a,a16080a,a16083a,a16087a,a16088a,a16089a,a16092a,a16096a,a16097a,a16098a,a16101a,a16105a,a16106a,a16107a,a16110a,a16114a,a16115a,a16116a,a16119a,a16123a,a16124a,a16125a,a16128a,a16132a,a16133a,a16134a,a16137a,a16141a,a16142a,a16143a,a16146a,a16150a,a16151a,a16152a,a16155a,a16159a,a16160a,a16161a,a16164a,a16168a,a16169a,a16170a,a16173a,a16177a,a16178a,a16179a,a16182a,a16186a,a16187a,a16188a,a16191a,a16195a,a16196a,a16197a,a16200a,a16204a,a16205a,a16206a,a16209a,a16213a,a16214a,a16215a,a16218a,a16222a,a16223a,a16224a,a16227a,a16231a,a16232a,a16233a,a16236a,a16240a,a16241a,a16242a,a16245a,a16249a,a16250a,a16251a,a16254a,a16258a,a16259a,a16260a,a16263a,a16267a,a16268a,a16269a,a16272a,a16276a,a16277a,a16278a,a16281a,a16285a,a16286a,a16287a,a16290a,a16294a,a16295a,a16296a,a16299a,a16303a,a16304a,a16305a,a16308a,a16312a,a16313a,a16314a,a16317a,a16321a,a16322a,a16323a,a16326a,a16330a,a16331a,a16332a,a16335a,a16339a,a16340a,a16341a,a16344a,a16348a,a16349a,a16350a,a16353a,a16357a,a16358a,a16359a,a16362a,a16366a,a16367a,a16368a,a16371a,a16375a,a16376a,a16377a,a16380a,a16384a,a16385a,a16386a,a16389a,a16393a,a16394a,a16395a,a16398a,a16402a,a16403a,a16404a,a16407a,a16411a,a16412a,a16413a,a16416a,a16420a,a16421a,a16422a,a16425a,a16429a,a16430a,a16431a,a16434a,a16438a,a16439a,a16440a,a16443a,a16447a,a16448a,a16449a,a16452a,a16456a,a16457a,a16458a,a16461a,a16465a,a16466a,a16467a,a16470a,a16474a,a16475a,a16476a,a16479a,a16483a,a16484a,a16485a,a16488a,a16492a,a16493a,a16494a,a16497a,a16501a,a16502a,a16503a,a16506a,a16510a,a16511a,a16512a,a16515a,a16519a,a16520a,a16521a,a16524a,a16528a,a16529a,a16530a,a16533a,a16537a,a16538a,a16539a,a16542a,a16546a,a16547a,a16548a,a16551a,a16555a,a16556a,a16557a,a16560a,a16564a,a16565a,a16566a,a16569a,a16573a,a16574a,a16575a,a16578a,a16582a,a16583a,a16584a,a16587a,a16591a,a16592a,a16593a,a16596a,a16600a,a16601a,a16602a,a16605a,a16609a,a16610a,a16611a,a16614a,a16618a,a16619a,a16620a,a16623a,a16627a,a16628a,a16629a,a16632a,a16636a,a16637a,a16638a,a16641a,a16645a,a16646a,a16647a,a16650a,a16654a,a16655a,a16656a,a16659a,a16663a,a16664a,a16665a,a16668a,a16672a,a16673a,a16674a,a16677a,a16681a,a16682a,a16683a,a16686a,a16690a,a16691a,a16692a,a16695a,a16699a,a16700a,a16701a,a16704a,a16708a,a16709a,a16710a,a16713a,a16717a,a16718a,a16719a,a16722a,a16726a,a16727a,a16728a,a16731a,a16735a,a16736a,a16737a,a16740a,a16744a,a16745a,a16746a,a16749a,a16753a,a16754a,a16755a,a16758a,a16762a,a16763a,a16764a,a16767a,a16771a,a16772a,a16773a,a16776a,a16780a,a16781a,a16782a,a16785a,a16789a,a16790a,a16791a,a16794a,a16798a,a16799a,a16800a,a16803a,a16807a,a16808a,a16809a,a16812a,a16816a,a16817a,a16818a,a16821a,a16825a,a16826a,a16827a,a16830a,a16834a,a16835a,a16836a,a16839a,a16843a,a16844a,a16845a,a16848a,a16852a,a16853a,a16854a,a16857a,a16861a,a16862a,a16863a,a16866a,a16870a,a16871a,a16872a,a16875a,a16879a,a16880a,a16881a,a16884a,a16888a,a16889a,a16890a,a16893a,a16897a,a16898a,a16899a,a16902a,a16906a,a16907a,a16908a,a16911a,a16915a,a16916a,a16917a,a16920a,a16924a,a16925a,a16926a,a16929a,a16933a,a16934a,a16935a,a16938a,a16942a,a16943a,a16944a,a16947a,a16951a,a16952a,a16953a,a16956a,a16960a,a16961a,a16962a,a16965a,a16969a,a16970a,a16971a,a16974a,a16978a,a16979a,a16980a,a16983a,a16987a,a16988a,a16989a,a16992a,a16996a,a16997a,a16998a,a17001a,a17005a,a17006a,a17007a,a17010a,a17014a,a17015a,a17016a,a17019a,a17023a,a17024a,a17025a,a17028a,a17032a,a17033a,a17034a,a17037a,a17041a,a17042a,a17043a,a17046a,a17050a,a17051a,a17052a,a17055a,a17059a,a17060a,a17061a,a17064a,a17068a,a17069a,a17070a,a17073a,a17077a,a17078a,a17079a,a17082a,a17086a,a17087a,a17088a,a17091a,a17095a,a17096a,a17097a,a17100a,a17104a,a17105a,a17106a,a17109a,a17113a,a17114a,a17115a,a17118a,a17122a,a17123a,a17124a,a17127a,a17131a,a17132a,a17133a,a17136a,a17140a,a17141a,a17142a,a17145a,a17149a,a17150a,a17151a,a17154a,a17158a,a17159a,a17160a,a17163a,a17167a,a17168a,a17169a,a17172a,a17176a,a17177a,a17178a,a17181a,a17185a,a17186a,a17187a,a17190a,a17194a,a17195a,a17196a,a17199a,a17203a,a17204a,a17205a,a17208a,a17212a,a17213a,a17214a,a17217a,a17221a,a17222a,a17223a,a17226a,a17230a,a17231a,a17232a,a17235a,a17239a,a17240a,a17241a,a17244a,a17248a,a17249a,a17250a,a17253a,a17257a,a17258a,a17259a,a17262a,a17266a,a17267a,a17268a,a17271a,a17275a,a17276a,a17277a,a17280a,a17284a,a17285a,a17286a,a17289a,a17293a,a17294a,a17295a,a17298a,a17302a,a17303a,a17304a,a17307a,a17311a,a17312a,a17313a,a17316a,a17320a,a17321a,a17322a,a17325a,a17329a,a17330a,a17331a,a17334a,a17338a,a17339a,a17340a,a17343a,a17347a,a17348a,a17349a,a17352a,a17356a,a17357a,a17358a,a17361a,a17365a,a17366a,a17367a,a17370a,a17374a,a17375a,a17376a,a17379a,a17383a,a17384a,a17385a,a17388a,a17392a,a17393a,a17394a,a17397a,a17401a,a17402a,a17403a,a17406a,a17410a,a17411a,a17412a,a17415a,a17419a,a17420a,a17421a,a17424a,a17428a,a17429a,a17430a,a17433a,a17437a,a17438a,a17439a,a17442a,a17446a,a17447a,a17448a,a17451a,a17455a,a17456a,a17457a,a17460a,a17464a,a17465a,a17466a,a17469a,a17473a,a17474a,a17475a,a17478a,a17482a,a17483a,a17484a,a17487a,a17491a,a17492a,a17493a,a17496a,a17500a,a17501a,a17502a,a17505a,a17509a,a17510a,a17511a,a17514a,a17518a,a17519a,a17520a,a17523a,a17527a,a17528a,a17529a,a17532a,a17536a,a17537a,a17538a,a17541a,a17545a,a17546a,a17547a,a17550a,a17554a,a17555a,a17556a,a17559a,a17563a,a17564a,a17565a,a17568a,a17572a,a17573a,a17574a,a17577a,a17581a,a17582a,a17583a,a17586a,a17590a,a17591a,a17592a,a17595a,a17599a,a17600a,a17601a,a17604a,a17608a,a17609a,a17610a,a17613a,a17617a,a17618a,a17619a,a17622a,a17626a,a17627a,a17628a,a17631a,a17635a,a17636a,a17637a,a17640a,a17644a,a17645a,a17646a,a17649a,a17653a,a17654a,a17655a,a17658a,a17662a,a17663a,a17664a,a17667a,a17671a,a17672a,a17673a,a17676a,a17680a,a17681a,a17682a,a17685a,a17689a,a17690a,a17691a,a17694a,a17698a,a17699a,a17700a,a17703a,a17707a,a17708a,a17709a,a17712a,a17716a,a17717a,a17718a,a17721a,a17725a,a17726a,a17727a,a17730a,a17734a,a17735a,a17736a,a17739a,a17743a,a17744a,a17745a,a17748a,a17752a,a17753a,a17754a,a17757a,a17761a,a17762a,a17763a,a17766a,a17770a,a17771a,a17772a,a17775a,a17779a,a17780a,a17781a,a17784a,a17788a,a17789a,a17790a,a17793a,a17797a,a17798a,a17799a,a17802a,a17806a,a17807a,a17808a,a17811a,a17815a,a17816a,a17817a,a17820a,a17824a,a17825a,a17826a,a17829a,a17833a,a17834a,a17835a,a17838a,a17842a,a17843a,a17844a,a17847a,a17851a,a17852a,a17853a,a17857a,a17858a,a17862a,a17863a,a17864a,a17867a,a17871a,a17872a,a17873a,a17877a,a17878a,a17882a,a17883a,a17884a,a17887a,a17891a,a17892a,a17893a,a17897a,a17898a,a17902a,a17903a,a17904a,a17907a,a17911a,a17912a,a17913a,a17917a,a17918a,a17922a,a17923a,a17924a,a17927a,a17931a,a17932a,a17933a,a17937a,a17938a,a17942a,a17943a,a17944a,a17947a,a17951a,a17952a,a17953a,a17957a,a17958a,a17962a,a17963a,a17964a,a17967a,a17971a,a17972a,a17973a,a17977a,a17978a,a17982a,a17983a,a17984a,a17987a,a17991a,a17992a,a17993a,a17997a,a17998a,a18002a,a18003a,a18004a,a18007a,a18011a,a18012a,a18013a,a18017a,a18018a,a18022a,a18023a,a18024a,a18027a,a18031a,a18032a,a18033a,a18037a,a18038a,a18042a,a18043a,a18044a,a18047a,a18051a,a18052a,a18053a,a18057a,a18058a,a18062a,a18063a,a18064a,a18067a,a18071a,a18072a,a18073a,a18077a,a18078a,a18082a,a18083a,a18084a,a18087a,a18091a,a18092a,a18093a,a18097a,a18098a,a18102a,a18103a,a18104a,a18107a,a18111a,a18112a,a18113a,a18117a,a18118a,a18122a,a18123a,a18124a,a18127a,a18131a,a18132a,a18133a,a18137a,a18138a,a18142a,a18143a,a18144a,a18147a,a18151a,a18152a,a18153a,a18157a,a18158a,a18162a,a18163a,a18164a,a18167a,a18171a,a18172a,a18173a,a18177a,a18178a,a18182a,a18183a,a18184a,a18187a,a18191a,a18192a,a18193a,a18197a,a18198a,a18202a,a18203a,a18204a,a18207a,a18211a,a18212a,a18213a,a18217a,a18218a,a18222a,a18223a,a18224a,a18227a,a18231a,a18232a,a18233a,a18237a,a18238a,a18242a,a18243a,a18244a,a18247a,a18251a,a18252a,a18253a,a18257a,a18258a,a18262a,a18263a,a18264a,a18267a,a18271a,a18272a,a18273a,a18277a,a18278a,a18282a,a18283a,a18284a,a18287a,a18291a,a18292a,a18293a,a18297a,a18298a,a18302a,a18303a,a18304a,a18307a,a18311a,a18312a,a18313a,a18317a,a18318a,a18322a,a18323a,a18324a,a18327a,a18331a,a18332a,a18333a,a18337a,a18338a,a18342a,a18343a,a18344a,a18347a,a18351a,a18352a,a18353a,a18357a,a18358a,a18362a,a18363a,a18364a,a18367a,a18371a,a18372a,a18373a,a18377a,a18378a,a18382a,a18383a,a18384a,a18387a,a18391a,a18392a,a18393a,a18397a,a18398a,a18402a,a18403a,a18404a,a18407a,a18411a,a18412a,a18413a,a18417a,a18418a,a18422a,a18423a,a18424a,a18427a,a18431a,a18432a,a18433a,a18437a,a18438a,a18442a,a18443a,a18444a,a18447a,a18451a,a18452a,a18453a,a18457a,a18458a,a18462a,a18463a,a18464a,a18467a,a18471a,a18472a,a18473a,a18477a,a18478a,a18482a,a18483a,a18484a,a18487a,a18491a,a18492a,a18493a,a18497a,a18498a,a18502a,a18503a,a18504a,a18507a,a18511a,a18512a,a18513a,a18517a,a18518a,a18522a,a18523a,a18524a,a18527a,a18531a,a18532a,a18533a,a18537a,a18538a,a18542a,a18543a,a18544a,a18547a,a18551a,a18552a,a18553a,a18557a,a18558a,a18562a,a18563a,a18564a,a18567a,a18571a,a18572a,a18573a,a18577a,a18578a,a18582a,a18583a,a18584a,a18587a,a18591a,a18592a,a18593a,a18597a,a18598a,a18602a,a18603a,a18604a,a18607a,a18611a,a18612a,a18613a,a18617a,a18618a,a18622a,a18623a,a18624a,a18627a,a18631a,a18632a,a18633a,a18637a,a18638a,a18642a,a18643a,a18644a,a18647a,a18651a,a18652a,a18653a,a18657a,a18658a,a18662a,a18663a,a18664a,a18667a,a18671a,a18672a,a18673a,a18677a,a18678a,a18682a,a18683a,a18684a,a18687a,a18691a,a18692a,a18693a,a18697a,a18698a,a18702a,a18703a,a18704a,a18707a,a18711a,a18712a,a18713a,a18717a,a18718a,a18722a,a18723a,a18724a,a18727a,a18731a,a18732a,a18733a,a18737a,a18738a,a18742a,a18743a,a18744a,a18747a,a18751a,a18752a,a18753a,a18757a,a18758a,a18762a,a18763a,a18764a,a18767a,a18771a,a18772a,a18773a,a18777a,a18778a,a18782a,a18783a,a18784a,a18787a,a18791a,a18792a,a18793a,a18797a,a18798a,a18802a,a18803a,a18804a,a18807a,a18811a,a18812a,a18813a,a18817a,a18818a,a18822a,a18823a,a18824a,a18827a,a18831a,a18832a,a18833a,a18837a,a18838a,a18842a,a18843a,a18844a,a18847a,a18851a,a18852a,a18853a,a18857a,a18858a,a18862a,a18863a,a18864a,a18867a,a18871a,a18872a,a18873a,a18877a,a18878a,a18882a,a18883a,a18884a,a18887a,a18891a,a18892a,a18893a,a18897a,a18898a,a18902a,a18903a,a18904a,a18907a,a18911a,a18912a,a18913a,a18917a,a18918a,a18922a,a18923a,a18924a,a18927a,a18931a,a18932a,a18933a,a18937a,a18938a,a18942a,a18943a,a18944a,a18947a,a18951a,a18952a,a18953a,a18957a,a18958a,a18962a,a18963a,a18964a,a18967a,a18971a,a18972a,a18973a,a18977a,a18978a,a18982a,a18983a,a18984a,a18987a,a18991a,a18992a,a18993a,a18997a,a18998a,a19002a,a19003a,a19004a,a19007a,a19011a,a19012a,a19013a,a19017a,a19018a,a19022a,a19023a,a19024a,a19027a,a19031a,a19032a,a19033a,a19037a,a19038a,a19042a,a19043a,a19044a,a19047a,a19051a,a19052a,a19053a,a19057a,a19058a,a19062a,a19063a,a19064a,a19067a,a19071a,a19072a,a19073a,a19077a,a19078a,a19082a,a19083a,a19084a,a19087a,a19091a,a19092a,a19093a,a19097a,a19098a,a19102a,a19103a,a19104a,a19107a,a19111a,a19112a,a19113a,a19117a,a19118a,a19122a,a19123a,a19124a,a19127a,a19131a,a19132a,a19133a,a19137a,a19138a,a19142a,a19143a,a19144a,a19147a,a19151a,a19152a,a19153a,a19157a,a19158a,a19162a,a19163a,a19164a,a19167a,a19171a,a19172a,a19173a,a19177a,a19178a,a19182a,a19183a,a19184a,a19187a,a19191a,a19192a,a19193a,a19197a,a19198a,a19202a,a19203a,a19204a,a19207a,a19211a,a19212a,a19213a,a19217a,a19218a,a19222a,a19223a,a19224a,a19227a,a19231a,a19232a,a19233a,a19237a,a19238a,a19242a,a19243a,a19244a,a19247a,a19251a,a19252a,a19253a,a19257a,a19258a,a19262a,a19263a,a19264a,a19267a,a19271a,a19272a,a19273a,a19277a,a19278a,a19282a,a19283a,a19284a,a19287a,a19291a,a19292a,a19293a,a19297a,a19298a,a19302a,a19303a,a19304a,a19307a,a19311a,a19312a,a19313a,a19317a,a19318a,a19322a,a19323a,a19324a,a19327a,a19331a,a19332a,a19333a,a19337a,a19338a,a19342a,a19343a,a19344a,a19347a,a19351a,a19352a,a19353a,a19357a,a19358a,a19362a,a19363a,a19364a,a19367a,a19371a,a19372a,a19373a,a19377a,a19378a,a19382a,a19383a,a19384a,a19387a,a19391a,a19392a,a19393a,a19397a,a19398a,a19402a,a19403a,a19404a,a19407a,a19411a,a19412a,a19413a,a19417a,a19418a,a19422a,a19423a,a19424a,a19427a,a19431a,a19432a,a19433a,a19437a,a19438a,a19442a,a19443a,a19444a,a19447a,a19451a,a19452a,a19453a,a19457a,a19458a,a19462a,a19463a,a19464a,a19467a,a19471a,a19472a,a19473a,a19477a,a19478a,a19482a,a19483a,a19484a,a19487a,a19491a,a19492a,a19493a,a19497a,a19498a,a19502a,a19503a,a19504a,a19507a,a19511a,a19512a,a19513a,a19517a,a19518a,a19522a,a19523a,a19524a,a19527a,a19531a,a19532a,a19533a,a19537a,a19538a,a19542a,a19543a,a19544a,a19547a,a19551a,a19552a,a19553a,a19557a,a19558a,a19562a,a19563a,a19564a,a19567a,a19571a,a19572a,a19573a,a19577a,a19578a,a19582a,a19583a,a19584a,a19587a,a19591a,a19592a,a19593a,a19597a,a19598a,a19602a,a19603a,a19604a,a19607a,a19611a,a19612a,a19613a,a19617a,a19618a,a19622a,a19623a,a19624a,a19627a,a19631a,a19632a,a19633a,a19637a,a19638a,a19642a,a19643a,a19644a,a19647a,a19651a,a19652a,a19653a,a19657a,a19658a,a19662a,a19663a,a19664a,a19667a,a19671a,a19672a,a19673a,a19677a,a19678a,a19682a,a19683a,a19684a,a19687a,a19691a,a19692a,a19693a,a19697a,a19698a,a19702a,a19703a,a19704a,a19707a,a19711a,a19712a,a19713a,a19717a,a19718a,a19722a,a19723a,a19724a,a19727a,a19731a,a19732a,a19733a,a19737a,a19738a,a19742a,a19743a,a19744a,a19747a,a19751a,a19752a,a19753a,a19757a,a19758a,a19762a,a19763a,a19764a,a19767a,a19771a,a19772a,a19773a,a19777a,a19778a,a19782a,a19783a,a19784a,a19787a,a19791a,a19792a,a19793a,a19797a,a19798a,a19802a,a19803a,a19804a,a19807a,a19811a,a19812a,a19813a,a19817a,a19818a,a19822a,a19823a,a19824a,a19827a,a19831a,a19832a,a19833a,a19837a,a19838a,a19842a,a19843a,a19844a,a19847a,a19851a,a19852a,a19853a,a19857a,a19858a,a19862a,a19863a,a19864a,a19867a,a19871a,a19872a,a19873a,a19877a,a19878a,a19882a,a19883a,a19884a,a19887a,a19891a,a19892a,a19893a,a19897a,a19898a,a19902a,a19903a,a19904a,a19907a,a19911a,a19912a,a19913a,a19917a,a19918a,a19922a,a19923a,a19924a,a19927a,a19931a,a19932a,a19933a,a19937a,a19938a,a19942a,a19943a,a19944a,a19947a,a19951a,a19952a,a19953a,a19957a,a19958a,a19962a,a19963a,a19964a,a19967a,a19971a,a19972a,a19973a,a19977a,a19978a,a19982a,a19983a,a19984a,a19987a,a19991a,a19992a,a19993a,a19997a,a19998a,a20002a,a20003a,a20004a,a20007a,a20011a,a20012a,a20013a,a20017a,a20018a,a20022a,a20023a,a20024a,a20027a,a20031a,a20032a,a20033a,a20037a,a20038a,a20042a,a20043a,a20044a,a20047a,a20051a,a20052a,a20053a,a20057a,a20058a,a20062a,a20063a,a20064a,a20067a,a20071a,a20072a,a20073a,a20077a,a20078a,a20082a,a20083a,a20084a,a20087a,a20091a,a20092a,a20093a,a20097a,a20098a,a20102a,a20103a,a20104a,a20107a,a20111a,a20112a,a20113a,a20117a,a20118a,a20122a,a20123a,a20124a,a20127a,a20131a,a20132a,a20133a,a20137a,a20138a,a20142a,a20143a,a20144a,a20147a,a20151a,a20152a,a20153a,a20157a,a20158a,a20162a,a20163a,a20164a,a20167a,a20171a,a20172a,a20173a,a20177a,a20178a,a20182a,a20183a,a20184a,a20187a,a20191a,a20192a,a20193a,a20197a,a20198a,a20202a,a20203a,a20204a,a20207a,a20211a,a20212a,a20213a,a20217a,a20218a,a20222a,a20223a,a20224a,a20227a,a20231a,a20232a,a20233a,a20237a,a20238a,a20242a,a20243a,a20244a,a20247a,a20251a,a20252a,a20253a,a20257a,a20258a,a20262a,a20263a,a20264a,a20267a,a20271a,a20272a,a20273a,a20277a,a20278a,a20282a,a20283a,a20284a,a20287a,a20291a,a20292a,a20293a,a20297a,a20298a,a20302a,a20303a,a20304a,a20307a,a20311a,a20312a,a20313a,a20317a,a20318a,a20322a,a20323a,a20324a,a20327a,a20331a,a20332a,a20333a,a20337a,a20338a,a20342a,a20343a,a20344a,a20347a,a20351a,a20352a,a20353a,a20357a,a20358a,a20362a,a20363a,a20364a,a20367a,a20371a,a20372a,a20373a,a20377a,a20378a,a20382a,a20383a,a20384a,a20387a,a20391a,a20392a,a20393a,a20397a,a20398a,a20402a,a20403a,a20404a,a20407a,a20411a,a20412a,a20413a,a20417a,a20418a,a20422a,a20423a,a20424a,a20427a,a20431a,a20432a,a20433a,a20437a,a20438a,a20442a,a20443a,a20444a,a20447a,a20451a,a20452a,a20453a,a20457a,a20458a,a20462a,a20463a,a20464a,a20467a,a20471a,a20472a,a20473a,a20477a,a20478a,a20482a,a20483a,a20484a,a20487a,a20491a,a20492a,a20493a,a20497a,a20498a,a20502a,a20503a,a20504a,a20507a,a20511a,a20512a,a20513a,a20517a,a20518a,a20522a,a20523a,a20524a,a20527a,a20531a,a20532a,a20533a,a20537a,a20538a,a20542a,a20543a,a20544a,a20547a,a20551a,a20552a,a20553a,a20557a,a20558a,a20562a,a20563a,a20564a,a20567a,a20571a,a20572a,a20573a,a20577a,a20578a,a20582a,a20583a,a20584a,a20587a,a20591a,a20592a,a20593a,a20597a,a20598a,a20602a,a20603a,a20604a,a20607a,a20611a,a20612a,a20613a,a20617a,a20618a,a20622a,a20623a,a20624a,a20627a,a20631a,a20632a,a20633a,a20637a,a20638a,a20642a,a20643a,a20644a,a20647a,a20651a,a20652a,a20653a,a20657a,a20658a,a20662a,a20663a,a20664a,a20667a,a20671a,a20672a,a20673a,a20677a,a20678a,a20682a,a20683a,a20684a,a20687a,a20691a,a20692a,a20693a,a20697a,a20698a,a20702a,a20703a,a20704a,a20707a,a20711a,a20712a,a20713a,a20717a,a20718a,a20722a,a20723a,a20724a,a20727a,a20731a,a20732a,a20733a,a20737a,a20738a,a20742a,a20743a,a20744a,a20747a,a20751a,a20752a,a20753a,a20757a,a20758a,a20762a,a20763a,a20764a,a20767a,a20771a,a20772a,a20773a,a20777a,a20778a,a20782a,a20783a,a20784a,a20787a,a20791a,a20792a,a20793a,a20797a,a20798a,a20802a,a20803a,a20804a,a20807a,a20811a,a20812a,a20813a,a20817a,a20818a,a20822a,a20823a,a20824a,a20827a,a20831a,a20832a,a20833a,a20837a,a20838a,a20842a,a20843a,a20844a,a20847a,a20851a,a20852a,a20853a,a20857a,a20858a,a20862a,a20863a,a20864a,a20867a,a20871a,a20872a,a20873a,a20877a,a20878a,a20882a,a20883a,a20884a,a20887a,a20891a,a20892a,a20893a,a20897a,a20898a,a20902a,a20903a,a20904a,a20907a,a20911a,a20912a,a20913a,a20917a,a20918a,a20922a,a20923a,a20924a,a20927a,a20931a,a20932a,a20933a,a20937a,a20938a,a20942a,a20943a,a20944a,a20947a,a20951a,a20952a,a20953a,a20957a,a20958a,a20962a,a20963a,a20964a,a20967a,a20971a,a20972a,a20973a,a20977a,a20978a,a20982a,a20983a,a20984a,a20987a,a20991a,a20992a,a20993a,a20997a,a20998a,a21002a,a21003a,a21004a,a21007a,a21011a,a21012a,a21013a,a21017a,a21018a,a21022a,a21023a,a21024a,a21027a,a21031a,a21032a,a21033a,a21037a,a21038a,a21042a,a21043a,a21044a,a21047a,a21051a,a21052a,a21053a,a21057a,a21058a,a21062a,a21063a,a21064a,a21067a,a21071a,a21072a,a21073a,a21077a,a21078a,a21082a,a21083a,a21084a,a21087a,a21091a,a21092a,a21093a,a21097a,a21098a,a21102a,a21103a,a21104a,a21107a,a21111a,a21112a,a21113a,a21117a,a21118a,a21122a,a21123a,a21124a,a21127a,a21131a,a21132a,a21133a,a21137a,a21138a,a21142a,a21143a,a21144a,a21147a,a21151a,a21152a,a21153a,a21157a,a21158a,a21162a,a21163a,a21164a,a21167a,a21171a,a21172a,a21173a,a21177a,a21178a,a21182a,a21183a,a21184a,a21187a,a21191a,a21192a,a21193a,a21197a,a21198a,a21202a,a21203a,a21204a,a21207a,a21211a,a21212a,a21213a,a21217a,a21218a,a21222a,a21223a,a21224a,a21227a,a21231a,a21232a,a21233a,a21237a,a21238a,a21242a,a21243a,a21244a,a21247a,a21251a,a21252a,a21253a,a21257a,a21258a,a21262a,a21263a,a21264a,a21267a,a21271a,a21272a,a21273a,a21277a,a21278a,a21282a,a21283a,a21284a,a21287a,a21291a,a21292a,a21293a,a21297a,a21298a,a21302a,a21303a,a21304a,a21307a,a21311a,a21312a,a21313a,a21317a,a21318a,a21322a,a21323a,a21324a,a21327a,a21331a,a21332a,a21333a,a21337a,a21338a,a21342a,a21343a,a21344a,a21347a,a21351a,a21352a,a21353a,a21357a,a21358a,a21362a,a21363a,a21364a,a21367a,a21371a,a21372a,a21373a,a21377a,a21378a,a21382a,a21383a,a21384a,a21387a,a21391a,a21392a,a21393a,a21397a,a21398a,a21402a,a21403a,a21404a,a21407a,a21411a,a21412a,a21413a,a21417a,a21418a,a21422a,a21423a,a21424a,a21427a,a21431a,a21432a,a21433a,a21437a,a21438a,a21442a,a21443a,a21444a,a21447a,a21451a,a21452a,a21453a,a21457a,a21458a,a21462a,a21463a,a21464a,a21467a,a21471a,a21472a,a21473a,a21477a,a21478a,a21482a,a21483a,a21484a,a21487a,a21491a,a21492a,a21493a,a21497a,a21498a,a21502a,a21503a,a21504a,a21507a,a21511a,a21512a,a21513a,a21517a,a21518a,a21522a,a21523a,a21524a,a21527a,a21531a,a21532a,a21533a,a21537a,a21538a,a21542a,a21543a,a21544a,a21547a,a21551a,a21552a,a21553a,a21557a,a21558a,a21562a,a21563a,a21564a,a21567a,a21571a,a21572a,a21573a,a21577a,a21578a,a21582a,a21583a,a21584a,a21587a,a21591a,a21592a,a21593a,a21597a,a21598a,a21602a,a21603a,a21604a,a21607a,a21611a,a21612a,a21613a,a21617a,a21618a,a21622a,a21623a,a21624a,a21627a,a21631a,a21632a,a21633a,a21637a,a21638a,a21642a,a21643a,a21644a,a21647a,a21651a,a21652a,a21653a,a21657a,a21658a,a21662a,a21663a,a21664a,a21667a,a21671a,a21672a,a21673a,a21677a,a21678a,a21682a,a21683a,a21684a,a21687a,a21691a,a21692a,a21693a,a21697a,a21698a,a21702a,a21703a,a21704a,a21707a,a21711a,a21712a,a21713a,a21717a,a21718a,a21722a,a21723a,a21724a,a21727a,a21731a,a21732a,a21733a,a21737a,a21738a,a21742a,a21743a,a21744a,a21747a,a21751a,a21752a,a21753a,a21757a,a21758a,a21762a,a21763a,a21764a,a21767a,a21771a,a21772a,a21773a,a21777a,a21778a,a21782a,a21783a,a21784a,a21787a,a21791a,a21792a,a21793a,a21797a,a21798a,a21802a,a21803a,a21804a,a21807a,a21811a,a21812a,a21813a,a21817a,a21818a,a21822a,a21823a,a21824a,a21827a,a21831a,a21832a,a21833a,a21837a,a21838a,a21842a,a21843a,a21844a,a21847a,a21851a,a21852a,a21853a,a21857a,a21858a,a21862a,a21863a,a21864a,a21867a,a21871a,a21872a,a21873a,a21877a,a21878a,a21882a,a21883a,a21884a,a21887a,a21891a,a21892a,a21893a,a21897a,a21898a,a21902a,a21903a,a21904a,a21907a,a21911a,a21912a,a21913a,a21917a,a21918a,a21922a,a21923a,a21924a,a21927a,a21931a,a21932a,a21933a,a21937a,a21938a,a21942a,a21943a,a21944a,a21947a,a21951a,a21952a,a21953a,a21957a,a21958a,a21962a,a21963a,a21964a,a21967a,a21971a,a21972a,a21973a,a21977a,a21978a,a21982a,a21983a,a21984a,a21987a,a21991a,a21992a,a21993a,a21997a,a21998a,a22002a,a22003a,a22004a,a22007a,a22011a,a22012a,a22013a,a22017a,a22018a,a22022a,a22023a,a22024a,a22027a,a22031a,a22032a,a22033a,a22037a,a22038a,a22042a,a22043a,a22044a,a22047a,a22051a,a22052a,a22053a,a22057a,a22058a,a22062a,a22063a,a22064a,a22067a,a22071a,a22072a,a22073a,a22077a,a22078a,a22082a,a22083a,a22084a,a22087a,a22091a,a22092a,a22093a,a22097a,a22098a,a22102a,a22103a,a22104a,a22107a,a22111a,a22112a,a22113a,a22117a,a22118a,a22122a,a22123a,a22124a,a22127a,a22131a,a22132a,a22133a,a22137a,a22138a,a22142a,a22143a,a22144a,a22147a,a22151a,a22152a,a22153a,a22157a,a22158a,a22162a,a22163a,a22164a,a22167a,a22171a,a22172a,a22173a,a22177a,a22178a,a22182a,a22183a,a22184a,a22187a,a22191a,a22192a,a22193a,a22197a,a22198a,a22202a,a22203a,a22204a,a22207a,a22211a,a22212a,a22213a,a22217a,a22218a,a22222a,a22223a,a22224a,a22227a,a22231a,a22232a,a22233a,a22237a,a22238a,a22242a,a22243a,a22244a,a22247a,a22251a,a22252a,a22253a,a22257a,a22258a,a22262a,a22263a,a22264a,a22267a,a22271a,a22272a,a22273a,a22277a,a22278a,a22282a,a22283a,a22284a,a22287a,a22291a,a22292a,a22293a,a22297a,a22298a,a22302a,a22303a,a22304a,a22307a,a22311a,a22312a,a22313a,a22317a,a22318a,a22322a,a22323a,a22324a,a22327a,a22331a,a22332a,a22333a,a22337a,a22338a,a22342a,a22343a,a22344a,a22347a,a22351a,a22352a,a22353a,a22357a,a22358a,a22362a,a22363a,a22364a,a22367a,a22371a,a22372a,a22373a,a22377a,a22378a,a22382a,a22383a,a22384a,a22387a,a22391a,a22392a,a22393a,a22397a,a22398a,a22402a,a22403a,a22404a,a22407a,a22411a,a22412a,a22413a,a22417a,a22418a,a22422a,a22423a,a22424a,a22427a,a22431a,a22432a,a22433a,a22437a,a22438a,a22442a,a22443a,a22444a,a22447a,a22451a,a22452a,a22453a,a22457a,a22458a,a22462a,a22463a,a22464a,a22467a,a22471a,a22472a,a22473a,a22477a,a22478a,a22482a,a22483a,a22484a,a22487a,a22491a,a22492a,a22493a,a22497a,a22498a,a22502a,a22503a,a22504a,a22507a,a22511a,a22512a,a22513a,a22517a,a22518a,a22522a,a22523a,a22524a,a22527a,a22531a,a22532a,a22533a,a22537a,a22538a,a22542a,a22543a,a22544a,a22547a,a22551a,a22552a,a22553a,a22557a,a22558a,a22562a,a22563a,a22564a,a22567a,a22571a,a22572a,a22573a,a22577a,a22578a,a22582a,a22583a,a22584a,a22587a,a22591a,a22592a,a22593a,a22597a,a22598a,a22602a,a22603a,a22604a,a22607a,a22611a,a22612a,a22613a,a22617a,a22618a,a22622a,a22623a,a22624a,a22627a,a22631a,a22632a,a22633a,a22637a,a22638a,a22642a,a22643a,a22644a,a22647a,a22651a,a22652a,a22653a,a22657a,a22658a,a22662a,a22663a,a22664a,a22667a,a22671a,a22672a,a22673a,a22677a,a22678a,a22682a,a22683a,a22684a,a22687a,a22691a,a22692a,a22693a,a22697a,a22698a,a22702a,a22703a,a22704a,a22707a,a22711a,a22712a,a22713a,a22717a,a22718a,a22722a,a22723a,a22724a,a22727a,a22731a,a22732a,a22733a,a22737a,a22738a,a22742a,a22743a,a22744a,a22747a,a22751a,a22752a,a22753a,a22757a,a22758a,a22762a,a22763a,a22764a,a22767a,a22771a,a22772a,a22773a,a22777a,a22778a,a22782a,a22783a,a22784a,a22787a,a22791a,a22792a,a22793a,a22797a,a22798a,a22802a,a22803a,a22804a,a22807a,a22811a,a22812a,a22813a,a22817a,a22818a,a22822a,a22823a,a22824a,a22827a,a22831a,a22832a,a22833a,a22837a,a22838a,a22842a,a22843a,a22844a,a22847a,a22851a,a22852a,a22853a,a22857a,a22858a,a22862a,a22863a,a22864a,a22867a,a22871a,a22872a,a22873a,a22877a,a22878a,a22882a,a22883a,a22884a,a22887a,a22891a,a22892a,a22893a,a22897a,a22898a,a22902a,a22903a,a22904a,a22907a,a22911a,a22912a,a22913a,a22917a,a22918a,a22922a,a22923a,a22924a,a22927a,a22931a,a22932a,a22933a,a22937a,a22938a,a22942a,a22943a,a22944a,a22947a,a22951a,a22952a,a22953a,a22957a,a22958a,a22962a,a22963a,a22964a,a22967a,a22971a,a22972a,a22973a,a22977a,a22978a,a22982a,a22983a,a22984a,a22987a,a22991a,a22992a,a22993a,a22997a,a22998a,a23002a,a23003a,a23004a,a23007a,a23011a,a23012a,a23013a,a23017a,a23018a,a23022a,a23023a,a23024a,a23027a,a23031a,a23032a,a23033a,a23037a,a23038a,a23042a,a23043a,a23044a,a23047a,a23051a,a23052a,a23053a,a23057a,a23058a,a23062a,a23063a,a23064a,a23067a,a23071a,a23072a,a23073a,a23077a,a23078a,a23082a,a23083a,a23084a,a23087a,a23091a,a23092a,a23093a,a23097a,a23098a,a23102a,a23103a,a23104a,a23107a,a23111a,a23112a,a23113a,a23117a,a23118a,a23122a,a23123a,a23124a,a23127a,a23131a,a23132a,a23133a,a23137a,a23138a,a23142a,a23143a,a23144a,a23147a,a23151a,a23152a,a23153a,a23157a,a23158a,a23162a,a23163a,a23164a,a23167a,a23171a,a23172a,a23173a,a23177a,a23178a,a23182a,a23183a,a23184a,a23187a,a23191a,a23192a,a23193a,a23197a,a23198a,a23202a,a23203a,a23204a,a23207a,a23211a,a23212a,a23213a,a23217a,a23218a,a23222a,a23223a,a23224a,a23227a,a23231a,a23232a,a23233a,a23237a,a23238a,a23242a,a23243a,a23244a,a23247a,a23251a,a23252a,a23253a,a23257a,a23258a,a23262a,a23263a,a23264a,a23267a,a23271a,a23272a,a23273a,a23277a,a23278a,a23282a,a23283a,a23284a,a23287a,a23291a,a23292a,a23293a,a23297a,a23298a,a23302a,a23303a,a23304a,a23307a,a23311a,a23312a,a23313a,a23317a,a23318a,a23322a,a23323a,a23324a,a23327a,a23331a,a23332a,a23333a,a23337a,a23338a,a23342a,a23343a,a23344a,a23347a,a23351a,a23352a,a23353a,a23357a,a23358a,a23362a,a23363a,a23364a,a23367a,a23371a,a23372a,a23373a,a23377a,a23378a,a23382a,a23383a,a23384a,a23387a,a23391a,a23392a,a23393a,a23397a,a23398a,a23402a,a23403a,a23404a,a23407a,a23411a,a23412a,a23413a,a23417a,a23418a,a23422a,a23423a,a23424a,a23427a,a23431a,a23432a,a23433a,a23437a,a23438a,a23442a,a23443a,a23444a,a23447a,a23451a,a23452a,a23453a,a23457a,a23458a,a23462a,a23463a,a23464a,a23467a,a23471a,a23472a,a23473a,a23477a,a23478a,a23482a,a23483a,a23484a,a23487a,a23491a,a23492a,a23493a,a23497a,a23498a,a23502a,a23503a,a23504a,a23507a,a23511a,a23512a,a23513a,a23517a,a23518a,a23522a,a23523a,a23524a,a23527a,a23531a,a23532a,a23533a,a23537a,a23538a,a23542a,a23543a,a23544a,a23547a,a23551a,a23552a,a23553a,a23557a,a23558a,a23562a,a23563a,a23564a,a23567a,a23571a,a23572a,a23573a,a23577a,a23578a,a23582a,a23583a,a23584a,a23587a,a23591a,a23592a,a23593a,a23597a,a23598a,a23602a,a23603a,a23604a,a23607a,a23611a,a23612a,a23613a,a23617a,a23618a,a23622a,a23623a,a23624a,a23627a,a23631a,a23632a,a23633a,a23637a,a23638a,a23642a,a23643a,a23644a,a23647a,a23651a,a23652a,a23653a,a23657a,a23658a,a23662a,a23663a,a23664a,a23667a,a23671a,a23672a,a23673a,a23677a,a23678a,a23682a,a23683a,a23684a,a23687a,a23691a,a23692a,a23693a,a23697a,a23698a,a23702a,a23703a,a23704a,a23707a,a23711a,a23712a,a23713a,a23717a,a23718a,a23722a,a23723a,a23724a,a23727a,a23731a,a23732a,a23733a,a23737a,a23738a,a23742a,a23743a,a23744a,a23747a,a23751a,a23752a,a23753a,a23757a,a23758a,a23762a,a23763a,a23764a,a23767a,a23771a,a23772a,a23773a,a23777a,a23778a,a23782a,a23783a,a23784a,a23787a,a23791a,a23792a,a23793a,a23797a,a23798a,a23802a,a23803a,a23804a,a23807a,a23811a,a23812a,a23813a,a23817a,a23818a,a23822a,a23823a,a23824a,a23827a,a23831a,a23832a,a23833a,a23837a,a23838a,a23842a,a23843a,a23844a,a23847a,a23851a,a23852a,a23853a,a23857a,a23858a,a23862a,a23863a,a23864a,a23867a,a23871a,a23872a,a23873a,a23877a,a23878a,a23882a,a23883a,a23884a,a23887a,a23891a,a23892a,a23893a,a23897a,a23898a,a23902a,a23903a,a23904a,a23907a,a23911a,a23912a,a23913a,a23917a,a23918a,a23922a,a23923a,a23924a,a23927a,a23931a,a23932a,a23933a,a23937a,a23938a,a23942a,a23943a,a23944a,a23947a,a23951a,a23952a,a23953a,a23957a,a23958a,a23962a,a23963a,a23964a,a23967a,a23971a,a23972a,a23973a,a23977a,a23978a,a23982a,a23983a,a23984a,a23987a,a23991a,a23992a,a23993a,a23997a,a23998a,a24002a,a24003a,a24004a,a24007a,a24011a,a24012a,a24013a,a24017a,a24018a,a24022a,a24023a,a24024a,a24027a,a24031a,a24032a,a24033a,a24037a,a24038a,a24042a,a24043a,a24044a,a24047a,a24051a,a24052a,a24053a,a24057a,a24058a,a24062a,a24063a,a24064a,a24067a,a24071a,a24072a,a24073a,a24077a,a24078a,a24082a,a24083a,a24084a,a24087a,a24091a,a24092a,a24093a,a24097a,a24098a,a24102a,a24103a,a24104a,a24107a,a24111a,a24112a,a24113a,a24117a,a24118a,a24122a,a24123a,a24124a,a24127a,a24131a,a24132a,a24133a,a24137a,a24138a,a24142a,a24143a,a24144a,a24147a,a24151a,a24152a,a24153a,a24157a,a24158a,a24162a,a24163a,a24164a,a24167a,a24171a,a24172a,a24173a,a24177a,a24178a,a24182a,a24183a,a24184a,a24187a,a24191a,a24192a,a24193a,a24197a,a24198a,a24202a,a24203a,a24204a,a24207a,a24211a,a24212a,a24213a,a24217a,a24218a,a24222a,a24223a,a24224a,a24227a,a24231a,a24232a,a24233a,a24237a,a24238a,a24242a,a24243a,a24244a,a24247a,a24251a,a24252a,a24253a,a24257a,a24258a,a24262a,a24263a,a24264a,a24267a,a24271a,a24272a,a24273a,a24277a,a24278a,a24282a,a24283a,a24284a,a24287a,a24291a,a24292a,a24293a,a24297a,a24298a,a24302a,a24303a,a24304a,a24307a,a24311a,a24312a,a24313a,a24317a,a24318a,a24322a,a24323a,a24324a,a24327a,a24331a,a24332a,a24333a,a24337a,a24338a,a24342a,a24343a,a24344a,a24347a,a24351a,a24352a,a24353a,a24357a,a24358a,a24362a,a24363a,a24364a,a24367a,a24371a,a24372a,a24373a,a24377a,a24378a,a24382a,a24383a,a24384a,a24387a,a24391a,a24392a,a24393a,a24397a,a24398a,a24402a,a24403a,a24404a,a24407a,a24411a,a24412a,a24413a,a24417a,a24418a,a24422a,a24423a,a24424a,a24427a,a24431a,a24432a,a24433a,a24437a,a24438a,a24442a,a24443a,a24444a,a24447a,a24451a,a24452a,a24453a,a24457a,a24458a,a24462a,a24463a,a24464a,a24467a,a24471a,a24472a,a24473a,a24477a,a24478a,a24482a,a24483a,a24484a,a24487a,a24491a,a24492a,a24493a,a24497a,a24498a,a24502a,a24503a,a24504a,a24507a,a24511a,a24512a,a24513a,a24517a,a24518a,a24522a,a24523a,a24524a,a24527a,a24531a,a24532a,a24533a,a24537a,a24538a,a24542a,a24543a,a24544a,a24547a,a24551a,a24552a,a24553a,a24557a,a24558a,a24562a,a24563a,a24564a,a24567a,a24571a,a24572a,a24573a,a24577a,a24578a,a24582a,a24583a,a24584a,a24587a,a24591a,a24592a,a24593a,a24597a,a24598a,a24602a,a24603a,a24604a,a24607a,a24611a,a24612a,a24613a,a24617a,a24618a,a24622a,a24623a,a24624a,a24627a,a24631a,a24632a,a24633a,a24637a,a24638a,a24642a,a24643a,a24644a,a24647a,a24651a,a24652a,a24653a,a24657a,a24658a,a24662a,a24663a,a24664a,a24667a,a24671a,a24672a,a24673a,a24677a,a24678a,a24682a,a24683a,a24684a,a24687a,a24691a,a24692a,a24693a,a24697a,a24698a,a24702a,a24703a,a24704a,a24707a,a24711a,a24712a,a24713a,a24717a,a24718a,a24722a,a24723a,a24724a,a24727a,a24731a,a24732a,a24733a,a24737a,a24738a,a24742a,a24743a,a24744a,a24747a,a24751a,a24752a,a24753a,a24757a,a24758a,a24762a,a24763a,a24764a,a24767a,a24771a,a24772a,a24773a,a24777a,a24778a,a24782a,a24783a,a24784a,a24787a,a24791a,a24792a,a24793a,a24797a,a24798a,a24802a,a24803a,a24804a,a24807a,a24811a,a24812a,a24813a,a24817a,a24818a,a24822a,a24823a,a24824a,a24827a,a24831a,a24832a,a24833a,a24837a,a24838a,a24842a,a24843a,a24844a,a24847a,a24851a,a24852a,a24853a,a24857a,a24858a,a24862a,a24863a,a24864a,a24867a,a24871a,a24872a,a24873a,a24877a,a24878a,a24882a,a24883a,a24884a,a24887a,a24891a,a24892a,a24893a,a24897a,a24898a,a24902a,a24903a,a24904a,a24907a,a24911a,a24912a,a24913a,a24917a,a24918a,a24922a,a24923a,a24924a,a24927a,a24931a,a24932a,a24933a,a24937a,a24938a,a24942a,a24943a,a24944a,a24947a,a24951a,a24952a,a24953a,a24957a,a24958a,a24962a,a24963a,a24964a,a24967a,a24971a,a24972a,a24973a,a24977a,a24978a,a24982a,a24983a,a24984a,a24987a,a24991a,a24992a,a24993a,a24997a,a24998a,a25002a,a25003a,a25004a,a25007a,a25011a,a25012a,a25013a,a25017a,a25018a,a25022a,a25023a,a25024a,a25027a,a25031a,a25032a,a25033a,a25037a,a25038a,a25042a,a25043a,a25044a,a25047a,a25051a,a25052a,a25053a,a25057a,a25058a,a25062a,a25063a,a25064a,a25067a,a25071a,a25072a,a25073a,a25077a,a25078a,a25082a,a25083a,a25084a,a25087a,a25091a,a25092a,a25093a,a25097a,a25098a,a25102a,a25103a,a25104a,a25107a,a25111a,a25112a,a25113a,a25117a,a25118a,a25122a,a25123a,a25124a,a25127a,a25131a,a25132a,a25133a,a25137a,a25138a,a25142a,a25143a,a25144a,a25147a,a25151a,a25152a,a25153a,a25157a,a25158a,a25162a,a25163a,a25164a,a25167a,a25171a,a25172a,a25173a,a25177a,a25178a,a25182a,a25183a,a25184a,a25187a,a25191a,a25192a,a25193a,a25197a,a25198a,a25202a,a25203a,a25204a,a25208a,a25209a,a25213a,a25214a,a25215a,a25219a,a25220a,a25224a,a25225a,a25226a,a25230a,a25231a,a25235a,a25236a,a25237a,a25241a,a25242a,a25246a,a25247a,a25248a,a25252a,a25253a,a25257a,a25258a,a25259a,a25263a,a25264a,a25268a,a25269a,a25270a,a25274a,a25275a,a25279a,a25280a,a25281a,a25285a,a25286a,a25290a,a25291a,a25292a,a25296a,a25297a,a25301a,a25302a,a25303a,a25307a,a25308a,a25312a,a25313a,a25314a,a25318a,a25319a,a25323a,a25324a,a25325a,a25329a,a25330a,a25334a,a25335a,a25336a,a25340a,a25341a,a25345a,a25346a,a25347a,a25351a,a25352a,a25356a,a25357a,a25358a,a25362a,a25363a,a25367a,a25368a,a25369a,a25373a,a25374a,a25378a,a25379a,a25380a,a25384a,a25385a,a25389a,a25390a,a25391a,a25395a,a25396a,a25400a,a25401a,a25402a,a25406a,a25407a,a25411a,a25412a,a25413a,a25417a,a25418a,a25422a,a25423a,a25424a,a25428a,a25429a,a25433a,a25434a,a25435a,a25439a,a25440a,a25444a,a25445a,a25446a,a25450a,a25451a,a25455a,a25456a,a25457a,a25461a,a25462a,a25466a,a25467a,a25468a,a25472a,a25473a,a25477a,a25478a,a25479a,a25483a,a25484a,a25488a,a25489a,a25490a,a25494a,a25495a,a25499a,a25500a,a25501a,a25505a,a25506a,a25510a,a25511a,a25512a,a25516a,a25517a,a25521a,a25522a,a25523a,a25527a,a25528a,a25532a,a25533a,a25534a,a25538a,a25539a,a25543a,a25544a,a25545a,a25549a,a25550a,a25554a,a25555a,a25556a,a25560a,a25561a,a25565a,a25566a,a25567a,a25571a,a25572a,a25576a,a25577a,a25578a,a25582a,a25583a,a25587a,a25588a,a25589a,a25593a,a25594a,a25598a,a25599a,a25600a,a25604a,a25605a,a25609a,a25610a,a25611a,a25615a,a25616a,a25620a,a25621a,a25622a,a25626a,a25627a,a25631a,a25632a,a25633a,a25637a,a25638a,a25642a,a25643a,a25644a,a25648a,a25649a,a25653a,a25654a,a25655a,a25659a,a25660a,a25664a,a25665a,a25666a,a25670a,a25671a,a25675a,a25676a,a25677a,a25681a,a25682a,a25686a,a25687a,a25688a,a25692a,a25693a,a25697a,a25698a,a25699a,a25703a,a25704a,a25708a,a25709a,a25710a,a25714a,a25715a,a25719a,a25720a,a25721a,a25725a,a25726a,a25730a,a25731a,a25732a,a25736a,a25737a,a25741a,a25742a,a25743a,a25747a,a25748a,a25752a,a25753a,a25754a,a25758a,a25759a,a25763a,a25764a,a25765a,a25769a,a25770a,a25774a,a25775a,a25776a,a25780a,a25781a,a25785a,a25786a,a25787a,a25791a,a25792a,a25796a,a25797a,a25798a,a25802a,a25803a,a25807a,a25808a,a25809a,a25813a,a25814a,a25818a,a25819a,a25820a,a25824a,a25825a,a25829a,a25830a,a25831a,a25835a,a25836a,a25840a,a25841a,a25842a,a25846a,a25847a,a25851a,a25852a,a25853a,a25857a,a25858a,a25862a,a25863a,a25864a,a25868a,a25869a,a25873a,a25874a,a25875a,a25879a,a25880a,a25884a,a25885a,a25886a,a25890a,a25891a,a25895a,a25896a,a25897a,a25901a,a25902a,a25906a,a25907a,a25908a,a25912a,a25913a,a25917a,a25918a,a25919a,a25923a,a25924a,a25928a,a25929a,a25930a,a25934a,a25935a,a25939a,a25940a,a25941a,a25945a,a25946a,a25950a,a25951a,a25952a,a25956a,a25957a,a25961a,a25962a,a25963a,a25967a,a25968a,a25972a,a25973a,a25974a,a25978a,a25979a,a25983a,a25984a,a25985a,a25989a,a25990a,a25994a,a25995a,a25996a,a26000a,a26001a,a26005a,a26006a,a26007a,a26011a,a26012a,a26016a,a26017a,a26018a,a26022a,a26023a,a26027a,a26028a,a26029a,a26033a,a26034a,a26038a,a26039a,a26040a,a26044a,a26045a,a26049a,a26050a,a26051a,a26055a,a26056a,a26060a,a26061a,a26062a,a26066a,a26067a,a26071a,a26072a,a26073a,a26077a,a26078a,a26082a,a26083a,a26084a,a26088a,a26089a,a26093a,a26094a,a26095a,a26099a,a26100a,a26104a,a26105a,a26106a,a26110a,a26111a,a26115a,a26116a,a26117a,a26121a,a26122a,a26126a,a26127a,a26128a,a26132a,a26133a,a26137a,a26138a,a26139a,a26143a,a26144a,a26148a,a26149a,a26150a,a26154a,a26155a,a26159a,a26160a,a26161a,a26165a,a26166a,a26170a,a26171a,a26172a,a26176a,a26177a,a26181a,a26182a,a26183a,a26187a,a26188a,a26192a,a26193a,a26194a,a26198a,a26199a,a26203a,a26204a,a26205a,a26209a,a26210a,a26214a,a26215a,a26216a,a26220a,a26221a,a26225a,a26226a,a26227a,a26231a,a26232a,a26236a,a26237a,a26238a,a26242a,a26243a,a26247a,a26248a,a26249a,a26253a,a26254a,a26258a,a26259a,a26260a,a26264a,a26265a,a26269a,a26270a,a26271a,a26275a,a26276a,a26280a,a26281a,a26282a,a26286a,a26287a,a26291a,a26292a,a26293a,a26297a,a26298a,a26302a,a26303a,a26304a,a26308a,a26309a,a26313a,a26314a,a26315a,a26319a,a26320a,a26324a,a26325a,a26326a,a26330a,a26331a,a26335a,a26336a,a26337a,a26341a,a26342a,a26346a,a26347a,a26348a,a26352a,a26353a,a26357a,a26358a,a26359a,a26363a,a26364a,a26368a,a26369a,a26370a,a26374a,a26375a,a26379a,a26380a,a26381a,a26385a,a26386a,a26390a,a26391a,a26392a,a26396a,a26397a,a26401a,a26402a,a26403a,a26407a,a26408a,a26412a,a26413a,a26414a,a26418a,a26419a,a26423a,a26424a,a26425a,a26429a,a26430a,a26434a,a26435a,a26436a,a26440a,a26441a,a26445a,a26446a,a26447a,a26451a,a26452a,a26456a,a26457a,a26458a,a26462a,a26463a,a26467a,a26468a,a26469a,a26473a,a26474a,a26478a,a26479a,a26480a,a26484a,a26485a,a26489a,a26490a,a26491a,a26495a,a26496a,a26500a,a26501a,a26502a,a26506a,a26507a,a26511a,a26512a,a26513a,a26517a,a26518a,a26522a,a26523a,a26524a,a26528a,a26529a,a26533a,a26534a,a26535a,a26539a,a26540a,a26544a,a26545a,a26546a,a26550a,a26551a,a26555a,a26556a,a26557a,a26561a,a26562a,a26566a,a26567a,a26568a,a26572a,a26573a,a26577a,a26578a,a26579a,a26583a,a26584a,a26588a,a26589a,a26590a,a26594a,a26595a,a26599a,a26600a,a26601a,a26605a,a26606a,a26610a,a26611a,a26612a,a26616a,a26617a,a26621a,a26622a,a26623a,a26627a,a26628a,a26632a,a26633a,a26634a,a26638a,a26639a,a26643a,a26644a,a26645a,a26649a,a26650a,a26654a,a26655a,a26656a,a26660a,a26661a,a26665a,a26666a,a26667a,a26671a,a26672a,a26676a,a26677a,a26678a,a26682a,a26683a,a26687a,a26688a,a26689a,a26693a,a26694a,a26698a,a26699a,a26700a,a26704a,a26705a,a26709a,a26710a,a26711a,a26715a,a26716a,a26720a,a26721a,a26722a,a26726a,a26727a,a26731a,a26732a,a26733a,a26737a,a26738a,a26742a,a26743a,a26744a,a26748a,a26749a,a26753a,a26754a,a26755a,a26759a,a26760a,a26764a,a26765a,a26766a,a26770a,a26771a,a26775a,a26776a,a26777a,a26781a,a26782a,a26786a,a26787a,a26788a,a26792a,a26793a,a26797a,a26798a,a26799a,a26803a,a26804a,a26808a,a26809a,a26810a,a26814a,a26815a,a26819a,a26820a,a26821a,a26825a,a26826a,a26830a,a26831a,a26832a,a26836a,a26837a,a26841a,a26842a,a26843a,a26847a,a26848a,a26852a,a26853a,a26854a,a26858a,a26859a,a26863a,a26864a,a26865a,a26869a,a26870a,a26874a,a26875a,a26876a,a26880a,a26881a,a26885a,a26886a,a26887a,a26891a,a26892a,a26896a,a26897a,a26898a,a26902a,a26903a,a26907a,a26908a,a26909a,a26913a,a26914a,a26918a,a26919a,a26920a,a26924a,a26925a,a26929a,a26930a,a26931a,a26935a,a26936a,a26940a,a26941a,a26942a,a26946a,a26947a,a26951a,a26952a,a26953a,a26957a,a26958a,a26962a,a26963a,a26964a,a26968a,a26969a,a26973a,a26974a,a26975a,a26979a,a26980a,a26984a,a26985a,a26986a,a26990a,a26991a,a26995a,a26996a,a26997a,a27001a,a27002a,a27006a,a27007a,a27008a,a27012a,a27013a,a27017a,a27018a,a27019a,a27023a,a27024a,a27028a,a27029a,a27030a,a27034a,a27035a,a27039a,a27040a,a27041a,a27045a,a27046a,a27050a,a27051a,a27052a,a27056a,a27057a,a27061a,a27062a,a27063a,a27067a,a27068a,a27072a,a27073a,a27074a,a27078a,a27079a,a27083a,a27084a,a27085a,a27089a,a27090a,a27094a,a27095a,a27096a,a27100a,a27101a,a27105a,a27106a,a27107a,a27111a,a27112a,a27116a,a27117a,a27118a,a27122a,a27123a,a27127a,a27128a,a27129a,a27133a,a27134a,a27138a,a27139a,a27140a,a27144a,a27145a,a27149a,a27150a,a27151a,a27155a,a27156a,a27160a,a27161a,a27162a,a27166a,a27167a,a27171a,a27172a,a27173a,a27177a,a27178a,a27182a,a27183a,a27184a,a27188a,a27189a,a27193a,a27194a,a27195a,a27199a,a27200a,a27204a,a27205a,a27206a,a27210a,a27211a,a27215a,a27216a,a27217a,a27221a,a27222a,a27226a,a27227a,a27228a,a27232a,a27233a,a27237a,a27238a,a27239a,a27243a,a27244a,a27248a,a27249a,a27250a,a27254a,a27255a,a27259a,a27260a,a27261a,a27265a,a27266a,a27270a,a27271a,a27272a,a27276a,a27277a,a27281a,a27282a,a27283a,a27287a,a27288a,a27292a,a27293a,a27294a,a27298a,a27299a,a27303a,a27304a,a27305a,a27309a,a27310a,a27314a,a27315a,a27316a,a27320a,a27321a,a27325a,a27326a,a27327a,a27331a,a27332a,a27336a,a27337a,a27338a,a27342a,a27343a,a27347a,a27348a,a27349a,a27353a,a27354a,a27358a,a27359a,a27360a,a27364a,a27365a,a27369a,a27370a,a27371a,a27375a,a27376a,a27380a,a27381a,a27382a,a27386a,a27387a,a27391a,a27392a,a27393a,a27397a,a27398a,a27402a,a27403a,a27404a,a27408a,a27409a,a27413a,a27414a,a27415a,a27419a,a27420a,a27424a,a27425a,a27426a,a27430a,a27431a,a27435a,a27436a,a27437a,a27441a,a27442a,a27446a,a27447a,a27448a,a27452a,a27453a,a27457a,a27458a,a27459a,a27463a,a27464a,a27468a,a27469a,a27470a,a27474a,a27475a,a27479a,a27480a,a27481a,a27485a,a27486a,a27490a,a27491a,a27492a,a27496a,a27497a,a27501a,a27502a,a27503a,a27507a,a27508a,a27512a,a27513a,a27514a,a27518a,a27519a,a27523a,a27524a,a27525a,a27529a,a27530a,a27534a,a27535a,a27536a,a27540a,a27541a,a27545a,a27546a,a27547a,a27551a,a27552a,a27556a,a27557a,a27558a,a27562a,a27563a,a27567a,a27568a,a27569a,a27573a,a27574a,a27578a,a27579a,a27580a,a27584a,a27585a,a27589a,a27590a,a27591a,a27595a,a27596a,a27600a,a27601a,a27602a,a27606a,a27607a,a27611a,a27612a,a27613a,a27617a,a27618a,a27622a,a27623a,a27624a,a27628a,a27629a,a27633a,a27634a,a27635a,a27639a,a27640a,a27644a,a27645a,a27646a,a27650a,a27651a,a27655a,a27656a,a27657a,a27661a,a27662a,a27666a,a27667a,a27668a,a27672a,a27673a,a27677a,a27678a,a27679a,a27683a,a27684a,a27688a,a27689a,a27690a,a27694a,a27695a,a27699a,a27700a,a27701a,a27705a,a27706a,a27710a,a27711a,a27712a,a27716a,a27717a,a27721a,a27722a,a27723a,a27727a,a27728a,a27732a,a27733a,a27734a,a27738a,a27739a,a27743a,a27744a,a27745a,a27749a,a27750a,a27754a,a27755a,a27756a,a27760a,a27761a,a27765a,a27766a,a27767a,a27771a,a27772a,a27776a,a27777a,a27778a,a27782a,a27783a,a27787a,a27788a,a27789a,a27793a,a27794a,a27798a,a27799a,a27800a,a27804a,a27805a,a27809a,a27810a,a27811a,a27815a,a27816a,a27820a,a27821a,a27822a,a27826a,a27827a,a27831a,a27832a,a27833a,a27837a,a27838a,a27842a,a27843a,a27844a,a27848a,a27849a,a27853a,a27854a,a27855a,a27859a,a27860a,a27864a,a27865a,a27866a,a27870a,a27871a,a27875a,a27876a,a27877a,a27881a,a27882a,a27886a,a27887a,a27888a,a27892a,a27893a,a27897a,a27898a,a27899a,a27903a,a27904a,a27908a,a27909a,a27910a,a27914a,a27915a,a27919a,a27920a,a27921a,a27925a,a27926a,a27930a,a27931a,a27932a,a27936a,a27937a,a27941a,a27942a,a27943a,a27947a,a27948a,a27952a,a27953a,a27954a,a27958a,a27959a,a27963a,a27964a,a27965a,a27969a,a27970a,a27974a,a27975a,a27976a,a27980a,a27981a,a27985a,a27986a,a27987a,a27991a,a27992a,a27996a,a27997a,a27998a,a28002a,a28003a,a28007a,a28008a,a28009a,a28013a,a28014a,a28018a,a28019a,a28020a,a28024a,a28025a,a28029a,a28030a,a28031a,a28035a,a28036a,a28040a,a28041a,a28042a,a28046a,a28047a,a28051a,a28052a,a28053a,a28057a,a28058a,a28062a,a28063a,a28064a,a28068a,a28069a,a28073a,a28074a,a28075a,a28079a,a28080a,a28084a,a28085a,a28086a,a28090a,a28091a,a28095a,a28096a,a28097a,a28101a,a28102a,a28106a,a28107a,a28108a,a28112a,a28113a,a28117a,a28118a,a28119a,a28123a,a28124a,a28128a,a28129a,a28130a,a28134a,a28135a,a28139a,a28140a,a28141a,a28145a,a28146a,a28150a,a28151a,a28152a,a28156a,a28157a,a28161a,a28162a,a28163a,a28167a,a28168a,a28172a,a28173a,a28174a,a28178a,a28179a,a28183a,a28184a,a28185a,a28189a,a28190a,a28194a,a28195a,a28196a,a28200a,a28201a,a28205a,a28206a,a28207a,a28211a,a28212a,a28216a,a28217a,a28218a,a28222a,a28223a,a28227a,a28228a,a28229a,a28233a,a28234a,a28238a,a28239a,a28240a,a28244a,a28245a,a28249a,a28250a,a28251a,a28255a,a28256a,a28260a,a28261a,a28262a,a28266a,a28267a,a28271a,a28272a,a28273a,a28277a,a28278a,a28282a,a28283a,a28284a,a28288a,a28289a,a28293a,a28294a,a28295a,a28299a,a28300a,a28304a,a28305a,a28306a,a28310a,a28311a,a28315a,a28316a,a28317a,a28321a,a28322a,a28326a,a28327a,a28328a,a28332a,a28333a,a28337a,a28338a,a28339a,a28343a,a28344a,a28348a,a28349a,a28350a,a28354a,a28355a,a28359a,a28360a,a28361a,a28365a,a28366a,a28370a,a28371a,a28372a,a28376a,a28377a,a28381a,a28382a,a28383a,a28387a,a28388a,a28392a,a28393a,a28394a,a28398a,a28399a,a28403a,a28404a,a28405a,a28409a,a28410a,a28414a,a28415a,a28416a,a28420a,a28421a,a28425a,a28426a,a28427a,a28431a,a28432a,a28436a,a28437a,a28438a,a28442a,a28443a,a28447a,a28448a,a28449a,a28453a,a28454a,a28458a,a28459a,a28460a,a28464a,a28465a,a28469a,a28470a,a28471a,a28475a,a28476a,a28480a,a28481a,a28482a,a28486a,a28487a,a28491a,a28492a,a28493a,a28497a,a28498a,a28502a,a28503a,a28504a,a28508a,a28509a,a28513a,a28514a,a28515a,a28519a,a28520a,a28524a,a28525a,a28526a,a28530a,a28531a,a28535a,a28536a,a28537a,a28541a,a28542a,a28546a,a28547a,a28548a,a28552a,a28553a,a28557a,a28558a,a28559a,a28563a,a28564a,a28568a,a28569a,a28570a,a28574a,a28575a,a28579a,a28580a,a28581a,a28585a,a28586a,a28590a,a28591a,a28592a,a28596a,a28597a,a28601a,a28602a,a28603a,a28607a,a28608a,a28612a,a28613a,a28614a,a28618a,a28619a,a28623a,a28624a,a28625a,a28629a,a28630a,a28634a,a28635a,a28636a,a28640a,a28641a,a28645a,a28646a,a28647a,a28651a,a28652a,a28656a,a28657a,a28658a,a28662a,a28663a,a28667a,a28668a,a28669a,a28673a,a28674a,a28678a,a28679a,a28680a,a28684a,a28685a,a28689a,a28690a,a28691a,a28695a,a28696a,a28700a,a28701a,a28702a,a28706a,a28707a,a28711a,a28712a,a28713a,a28717a,a28718a,a28722a,a28723a,a28724a,a28728a,a28729a,a28733a,a28734a,a28735a,a28739a,a28740a,a28744a,a28745a,a28746a,a28750a,a28751a,a28755a,a28756a,a28757a,a28761a,a28762a,a28766a,a28767a,a28768a,a28772a,a28773a,a28777a,a28778a,a28779a,a28783a,a28784a,a28788a,a28789a,a28790a,a28794a,a28795a,a28799a,a28800a,a28801a,a28805a,a28806a,a28810a,a28811a,a28812a,a28816a,a28817a,a28821a,a28822a,a28823a,a28827a,a28828a,a28832a,a28833a,a28834a,a28838a,a28839a,a28843a,a28844a,a28845a,a28849a,a28850a,a28854a,a28855a,a28856a,a28860a,a28861a,a28865a,a28866a,a28867a,a28871a,a28872a,a28876a,a28877a,a28878a,a28882a,a28883a,a28887a,a28888a,a28889a,a28893a,a28894a,a28898a,a28899a,a28900a,a28904a,a28905a,a28909a,a28910a,a28911a,a28915a,a28916a,a28920a,a28921a,a28922a,a28926a,a28927a,a28931a,a28932a,a28933a,a28937a,a28938a,a28942a,a28943a,a28944a,a28948a,a28949a,a28953a,a28954a,a28955a,a28959a,a28960a,a28964a,a28965a,a28966a,a28970a,a28971a,a28975a,a28976a,a28977a,a28981a,a28982a,a28986a,a28987a,a28988a,a28992a,a28993a,a28997a,a28998a,a28999a,a29003a,a29004a,a29008a,a29009a,a29010a,a29014a,a29015a,a29019a,a29020a,a29021a,a29025a,a29026a,a29030a,a29031a,a29032a,a29036a,a29037a,a29041a,a29042a,a29043a,a29047a,a29048a,a29052a,a29053a,a29054a,a29058a,a29059a,a29063a,a29064a,a29065a,a29069a,a29070a,a29074a,a29075a,a29076a,a29080a,a29081a,a29085a,a29086a,a29087a,a29091a,a29092a,a29096a,a29097a,a29098a,a29102a,a29103a,a29107a,a29108a,a29109a,a29113a,a29114a,a29118a,a29119a,a29120a,a29124a,a29125a,a29129a,a29130a,a29131a,a29135a,a29136a,a29140a,a29141a,a29142a,a29146a,a29147a,a29151a,a29152a,a29153a,a29157a,a29158a,a29162a,a29163a,a29164a,a29168a,a29169a,a29173a,a29174a,a29175a,a29179a,a29180a,a29184a,a29185a,a29186a,a29190a,a29191a,a29195a,a29196a,a29197a,a29201a,a29202a,a29206a,a29207a,a29208a,a29212a,a29213a,a29217a,a29218a,a29219a,a29223a,a29224a,a29228a,a29229a,a29230a,a29234a,a29235a,a29239a,a29240a,a29241a,a29245a,a29246a,a29250a,a29251a,a29252a,a29256a,a29257a,a29261a,a29262a,a29263a,a29267a,a29268a,a29272a,a29273a,a29274a,a29278a,a29279a,a29283a,a29284a,a29285a,a29289a,a29290a,a29294a,a29295a,a29296a,a29300a,a29301a,a29305a,a29306a,a29307a,a29311a,a29312a,a29316a,a29317a,a29318a,a29322a,a29323a,a29327a,a29328a,a29329a,a29333a,a29334a,a29338a,a29339a,a29340a,a29344a,a29345a,a29349a,a29350a,a29351a,a29355a,a29356a,a29360a,a29361a,a29362a,a29366a,a29367a,a29371a,a29372a,a29373a,a29377a,a29378a,a29382a,a29383a,a29384a,a29388a,a29389a,a29393a,a29394a,a29395a,a29399a,a29400a,a29404a,a29405a,a29406a,a29410a,a29411a,a29415a,a29416a,a29417a,a29421a,a29422a,a29426a,a29427a,a29428a,a29432a,a29433a,a29437a,a29438a,a29439a,a29443a,a29444a,a29448a,a29449a,a29450a,a29454a,a29455a,a29459a,a29460a,a29461a,a29465a,a29466a,a29470a,a29471a,a29472a,a29476a,a29477a,a29481a,a29482a,a29483a,a29487a,a29488a,a29492a,a29493a,a29494a,a29498a,a29499a,a29503a,a29504a,a29505a,a29509a,a29510a,a29514a,a29515a,a29516a,a29520a,a29521a,a29525a,a29526a,a29527a,a29531a,a29532a,a29536a,a29537a,a29538a,a29542a,a29543a,a29547a,a29548a,a29549a,a29553a,a29554a,a29558a,a29559a,a29560a,a29564a,a29565a,a29569a,a29570a,a29571a,a29575a,a29576a,a29580a,a29581a,a29582a,a29586a,a29587a,a29591a,a29592a,a29593a,a29597a,a29598a,a29602a,a29603a,a29604a,a29608a,a29609a,a29613a,a29614a,a29615a,a29619a,a29620a,a29624a,a29625a,a29626a,a29630a,a29631a,a29635a,a29636a,a29637a,a29641a,a29642a,a29646a,a29647a,a29648a,a29652a,a29653a,a29657a,a29658a,a29659a,a29663a,a29664a,a29668a,a29669a,a29670a,a29674a,a29675a,a29679a,a29680a,a29681a,a29685a,a29686a,a29690a,a29691a,a29692a,a29696a,a29697a,a29701a,a29702a,a29703a,a29707a,a29708a,a29712a,a29713a,a29714a,a29718a,a29719a,a29723a,a29724a,a29725a,a29729a,a29730a,a29734a,a29735a,a29736a,a29740a,a29741a,a29745a,a29746a,a29747a,a29751a,a29752a,a29756a,a29757a,a29758a,a29762a,a29763a,a29767a,a29768a,a29769a,a29773a,a29774a,a29778a,a29779a,a29780a,a29784a,a29785a,a29789a,a29790a,a29791a,a29795a,a29796a,a29800a,a29801a,a29802a,a29806a,a29807a,a29811a,a29812a,a29813a,a29817a,a29818a,a29822a,a29823a,a29824a,a29828a,a29829a,a29833a,a29834a,a29835a,a29839a,a29840a,a29844a,a29845a,a29846a,a29850a,a29851a,a29855a,a29856a,a29857a,a29861a,a29862a,a29866a,a29867a,a29868a,a29872a,a29873a,a29877a,a29878a,a29879a,a29883a,a29884a,a29888a,a29889a,a29890a,a29894a,a29895a,a29899a,a29900a,a29901a,a29905a,a29906a,a29910a,a29911a,a29912a,a29916a,a29917a,a29921a,a29922a,a29923a,a29927a,a29928a,a29932a,a29933a,a29934a,a29938a,a29939a,a29943a,a29944a,a29945a,a29949a,a29950a,a29954a,a29955a,a29956a,a29960a,a29961a,a29965a,a29966a,a29967a,a29971a,a29972a,a29976a,a29977a,a29978a,a29982a,a29983a,a29987a,a29988a,a29989a,a29993a,a29994a,a29998a,a29999a,a30000a,a30004a,a30005a,a30009a,a30010a,a30011a,a30015a,a30016a,a30020a,a30021a,a30022a,a30026a,a30027a,a30031a,a30032a,a30033a,a30037a,a30038a,a30042a,a30043a,a30044a,a30048a,a30049a,a30053a,a30054a,a30055a,a30059a,a30060a,a30064a,a30065a,a30066a,a30070a,a30071a,a30075a,a30076a,a30077a,a30081a,a30082a,a30086a,a30087a,a30088a,a30092a,a30093a,a30097a,a30098a,a30099a,a30103a,a30104a,a30108a,a30109a,a30110a,a30114a,a30115a,a30119a,a30120a,a30121a,a30125a,a30126a,a30130a,a30131a,a30132a,a30136a,a30137a,a30141a,a30142a,a30143a,a30147a,a30148a,a30152a,a30153a,a30154a,a30158a,a30159a,a30163a,a30164a,a30165a,a30169a,a30170a,a30174a,a30175a,a30176a,a30180a,a30181a,a30185a,a30186a,a30187a,a30191a,a30192a,a30196a,a30197a,a30198a,a30202a,a30203a,a30207a,a30208a,a30209a,a30213a,a30214a,a30218a,a30219a,a30220a,a30224a,a30225a,a30229a,a30230a,a30231a,a30235a,a30236a,a30240a,a30241a,a30242a,a30246a,a30247a,a30251a,a30252a,a30253a,a30257a,a30258a,a30262a,a30263a,a30264a,a30268a,a30269a,a30273a,a30274a,a30275a,a30279a,a30280a,a30284a,a30285a,a30286a,a30290a,a30291a,a30295a,a30296a,a30297a,a30301a,a30302a,a30306a,a30307a,a30308a,a30312a,a30313a,a30317a,a30318a,a30319a,a30323a,a30324a,a30328a,a30329a,a30330a,a30334a,a30335a,a30339a,a30340a,a30341a,a30345a,a30346a,a30350a,a30351a,a30352a,a30356a,a30357a,a30361a,a30362a,a30363a,a30367a,a30368a,a30372a,a30373a,a30374a,a30378a,a30379a,a30383a,a30384a,a30385a,a30389a,a30390a,a30394a,a30395a,a30396a,a30400a,a30401a,a30405a,a30406a,a30407a,a30411a,a30412a,a30416a,a30417a,a30418a,a30422a,a30423a,a30427a,a30428a,a30429a,a30433a,a30434a,a30438a,a30439a,a30440a,a30444a,a30445a,a30449a,a30450a,a30451a,a30455a,a30456a,a30460a,a30461a,a30462a,a30466a,a30467a,a30471a,a30472a,a30473a,a30477a,a30478a,a30482a,a30483a,a30484a,a30488a,a30489a,a30493a,a30494a,a30495a,a30499a,a30500a,a30504a,a30505a,a30506a,a30510a,a30511a,a30515a,a30516a,a30517a,a30521a,a30522a,a30526a,a30527a,a30528a,a30532a,a30533a,a30537a,a30538a,a30539a,a30543a,a30544a,a30548a,a30549a,a30550a,a30554a,a30555a,a30559a,a30560a,a30561a,a30565a,a30566a,a30570a,a30571a,a30572a,a30576a,a30577a,a30581a,a30582a,a30583a,a30587a,a30588a,a30592a,a30593a,a30594a,a30598a,a30599a,a30603a,a30604a,a30605a,a30609a,a30610a,a30614a,a30615a,a30616a,a30620a,a30621a,a30625a,a30626a,a30627a,a30631a,a30632a,a30636a,a30637a,a30638a,a30642a,a30643a,a30647a,a30648a,a30649a,a30653a,a30654a,a30658a,a30659a,a30660a,a30664a,a30665a,a30669a,a30670a,a30671a,a30675a,a30676a,a30680a,a30681a,a30682a,a30686a,a30687a,a30691a,a30692a,a30693a,a30697a,a30698a,a30702a,a30703a,a30704a,a30708a,a30709a,a30713a,a30714a,a30715a,a30719a,a30720a,a30724a,a30725a,a30726a,a30730a,a30731a,a30735a,a30736a,a30737a,a30741a,a30742a,a30746a,a30747a,a30748a,a30752a,a30753a,a30757a,a30758a,a30759a,a30763a,a30764a,a30768a,a30769a,a30770a,a30774a,a30775a,a30779a,a30780a,a30781a,a30785a,a30786a,a30790a,a30791a,a30792a,a30796a,a30797a,a30801a,a30802a,a30803a,a30807a,a30808a,a30812a,a30813a,a30814a,a30818a,a30819a,a30823a,a30824a,a30825a,a30829a,a30830a,a30834a,a30835a,a30836a,a30840a,a30841a,a30845a,a30846a,a30847a,a30851a,a30852a,a30856a,a30857a,a30858a,a30862a,a30863a,a30867a,a30868a,a30869a,a30873a,a30874a,a30878a,a30879a,a30880a,a30884a,a30885a,a30889a,a30890a,a30891a,a30895a,a30896a,a30900a,a30901a,a30902a,a30906a,a30907a,a30911a,a30912a,a30913a,a30917a,a30918a,a30922a,a30923a,a30924a,a30928a,a30929a,a30933a,a30934a,a30935a,a30939a,a30940a,a30944a,a30945a,a30946a,a30950a,a30951a,a30955a,a30956a,a30957a,a30961a,a30962a,a30966a,a30967a,a30968a,a30972a,a30973a,a30977a,a30978a,a30979a,a30983a,a30984a,a30988a,a30989a,a30990a,a30994a,a30995a,a30999a,a31000a,a31001a,a31005a,a31006a,a31010a,a31011a,a31012a,a31016a,a31017a,a31021a,a31022a,a31023a,a31027a,a31028a,a31032a,a31033a,a31034a,a31038a,a31039a,a31043a,a31044a,a31045a,a31049a,a31050a,a31054a,a31055a,a31056a,a31060a,a31061a,a31065a,a31066a,a31067a,a31071a,a31072a,a31076a,a31077a,a31078a,a31082a,a31083a,a31087a,a31088a,a31089a,a31093a,a31094a,a31098a,a31099a,a31100a,a31104a,a31105a,a31109a,a31110a,a31111a,a31115a,a31116a,a31120a,a31121a,a31122a,a31126a,a31127a,a31131a,a31132a,a31133a,a31137a,a31138a,a31142a,a31143a,a31144a,a31148a,a31149a,a31153a,a31154a,a31155a,a31159a,a31160a,a31164a,a31165a,a31166a,a31170a,a31171a,a31175a,a31176a,a31177a,a31181a,a31182a,a31186a,a31187a,a31188a,a31192a,a31193a,a31197a,a31198a,a31199a,a31203a,a31204a,a31208a,a31209a,a31210a,a31214a,a31215a,a31219a,a31220a,a31221a,a31225a,a31226a,a31230a,a31231a,a31232a,a31236a,a31237a,a31241a,a31242a,a31243a,a31247a,a31248a,a31252a,a31253a,a31254a,a31258a,a31259a,a31263a,a31264a,a31265a,a31269a,a31270a,a31274a,a31275a,a31276a,a31280a,a31281a,a31285a,a31286a,a31287a,a31291a,a31292a,a31296a,a31297a,a31298a,a31302a,a31303a,a31307a,a31308a,a31309a,a31313a,a31314a,a31318a,a31319a,a31320a,a31324a,a31325a,a31329a,a31330a,a31331a,a31335a,a31336a,a31340a,a31341a,a31342a,a31346a,a31347a,a31351a,a31352a,a31353a,a31357a,a31358a,a31362a,a31363a,a31364a,a31368a,a31369a,a31373a,a31374a,a31375a,a31379a,a31380a,a31384a,a31385a,a31386a,a31390a,a31391a,a31395a,a31396a,a31397a,a31401a,a31402a,a31406a,a31407a,a31408a,a31412a,a31413a,a31417a,a31418a,a31419a,a31423a,a31424a,a31428a,a31429a,a31430a,a31434a,a31435a,a31439a,a31440a,a31441a,a31445a,a31446a,a31450a,a31451a,a31452a,a31456a,a31457a,a31461a,a31462a,a31463a,a31467a,a31468a,a31472a,a31473a,a31474a,a31478a,a31479a,a31483a,a31484a,a31485a,a31489a,a31490a,a31494a,a31495a,a31496a,a31500a,a31501a,a31505a,a31506a,a31507a,a31511a,a31512a,a31516a,a31517a,a31518a,a31522a,a31523a,a31527a,a31528a,a31529a,a31533a,a31534a,a31538a,a31539a,a31540a,a31544a,a31545a,a31549a,a31550a,a31551a,a31555a,a31556a,a31560a,a31561a,a31562a,a31566a,a31567a,a31571a,a31572a,a31573a,a31577a,a31578a,a31582a,a31583a,a31584a,a31588a,a31589a,a31593a,a31594a,a31595a,a31599a,a31600a,a31604a,a31605a,a31606a,a31610a,a31611a,a31615a,a31616a,a31617a,a31621a,a31622a,a31626a,a31627a,a31628a,a31632a,a31633a,a31637a,a31638a,a31639a,a31643a,a31644a,a31648a,a31649a,a31650a,a31654a,a31655a,a31659a,a31660a,a31661a,a31665a,a31666a,a31670a,a31671a,a31672a,a31676a,a31677a,a31681a,a31682a,a31683a,a31687a,a31688a,a31692a,a31693a,a31694a,a31698a,a31699a,a31703a,a31704a,a31705a,a31709a,a31710a,a31714a,a31715a,a31716a,a31720a,a31721a,a31725a,a31726a,a31727a,a31731a,a31732a,a31736a,a31737a,a31738a,a31742a,a31743a,a31747a,a31748a,a31749a,a31753a,a31754a,a31758a,a31759a,a31760a,a31764a,a31765a,a31769a,a31770a,a31771a,a31775a,a31776a,a31780a,a31781a,a31782a,a31786a,a31787a,a31791a,a31792a,a31793a,a31797a,a31798a,a31802a,a31803a,a31804a,a31808a,a31809a,a31813a,a31814a,a31815a,a31819a,a31820a,a31824a,a31825a,a31826a,a31830a,a31831a,a31835a,a31836a,a31837a,a31841a,a31842a,a31846a,a31847a,a31848a,a31852a,a31853a,a31857a,a31858a,a31859a,a31863a,a31864a,a31868a,a31869a,a31870a,a31874a,a31875a,a31879a,a31880a,a31881a,a31885a,a31886a,a31890a,a31891a,a31892a,a31896a,a31897a,a31901a,a31902a,a31903a,a31907a,a31908a,a31912a,a31913a,a31914a,a31918a,a31919a,a31923a,a31924a,a31925a,a31929a,a31930a,a31934a,a31935a,a31936a,a31940a,a31941a,a31945a,a31946a,a31947a,a31951a,a31952a,a31956a,a31957a,a31958a,a31962a,a31963a,a31967a,a31968a,a31969a,a31973a,a31974a,a31978a,a31979a,a31980a,a31984a,a31985a,a31989a,a31990a,a31991a,a31995a,a31996a,a32000a,a32001a,a32002a,a32006a,a32007a,a32011a,a32012a,a32013a,a32017a,a32018a,a32022a,a32023a,a32024a,a32028a,a32029a,a32033a,a32034a,a32035a,a32039a,a32040a,a32044a,a32045a,a32046a,a32050a,a32051a,a32055a,a32056a,a32057a,a32061a,a32062a,a32066a,a32067a,a32068a,a32072a,a32073a,a32077a,a32078a,a32079a,a32083a,a32084a,a32088a,a32089a,a32090a,a32094a,a32095a,a32099a,a32100a,a32101a,a32105a,a32106a,a32110a,a32111a,a32112a,a32116a,a32117a,a32121a,a32122a,a32123a,a32127a,a32128a,a32132a,a32133a,a32134a,a32138a,a32139a,a32143a,a32144a,a32145a,a32149a,a32150a,a32154a,a32155a,a32156a,a32160a,a32161a,a32165a,a32166a,a32167a,a32171a,a32172a,a32176a,a32177a,a32178a,a32182a,a32183a,a32187a,a32188a,a32189a,a32193a,a32194a,a32198a,a32199a,a32200a,a32204a,a32205a,a32209a,a32210a,a32211a,a32215a,a32216a,a32220a,a32221a,a32222a,a32226a,a32227a,a32231a,a32232a,a32233a,a32237a,a32238a,a32242a,a32243a,a32244a,a32248a,a32249a,a32253a,a32254a,a32255a,a32259a,a32260a,a32264a,a32265a,a32266a,a32270a,a32271a,a32275a,a32276a,a32277a,a32281a,a32282a,a32286a,a32287a,a32288a,a32292a,a32293a,a32297a,a32298a,a32299a,a32303a,a32304a,a32308a,a32309a,a32310a,a32314a,a32315a,a32319a,a32320a,a32321a,a32325a,a32326a,a32330a,a32331a,a32332a,a32336a,a32337a,a32341a,a32342a,a32343a,a32347a,a32348a,a32352a,a32353a,a32354a,a32358a,a32359a,a32363a,a32364a,a32365a,a32369a,a32370a,a32374a,a32375a,a32376a,a32380a,a32381a,a32385a,a32386a,a32387a,a32391a,a32392a,a32396a,a32397a,a32398a,a32402a,a32403a,a32407a,a32408a,a32409a,a32413a,a32414a,a32418a,a32419a,a32420a,a32424a,a32425a,a32429a,a32430a,a32431a,a32435a,a32436a,a32440a,a32441a,a32442a,a32446a,a32447a,a32451a,a32452a,a32453a,a32457a,a32458a,a32462a,a32463a,a32464a,a32468a,a32469a,a32473a,a32474a,a32475a,a32479a,a32480a,a32484a,a32485a,a32486a,a32490a,a32491a,a32495a,a32496a,a32497a,a32501a,a32502a,a32506a,a32507a,a32508a,a32512a,a32513a,a32517a,a32518a,a32519a,a32523a,a32524a,a32528a,a32529a,a32530a,a32534a,a32535a,a32539a,a32540a,a32541a,a32545a,a32546a,a32550a,a32551a,a32552a,a32556a,a32557a,a32561a,a32562a,a32563a,a32567a,a32568a,a32572a,a32573a,a32574a,a32578a,a32579a,a32583a,a32584a,a32585a,a32589a,a32590a,a32594a,a32595a,a32596a,a32600a,a32601a,a32605a,a32606a,a32607a,a32611a,a32612a,a32616a,a32617a,a32618a,a32622a,a32623a,a32627a,a32628a,a32629a,a32633a,a32634a,a32638a,a32639a,a32640a,a32644a,a32645a,a32649a,a32650a,a32651a,a32655a,a32656a,a32660a,a32661a,a32662a,a32666a,a32667a,a32671a,a32672a,a32673a,a32677a,a32678a,a32682a,a32683a,a32684a,a32688a,a32689a,a32693a,a32694a,a32695a,a32699a,a32700a,a32704a,a32705a,a32706a,a32710a,a32711a,a32715a,a32716a,a32717a,a32721a,a32722a,a32726a,a32727a,a32728a,a32732a,a32733a,a32737a,a32738a,a32739a,a32743a,a32744a,a32748a,a32749a,a32750a,a32754a,a32755a,a32759a,a32760a,a32761a,a32765a,a32766a,a32770a,a32771a,a32772a,a32776a,a32777a,a32781a,a32782a,a32783a,a32787a,a32788a,a32792a,a32793a,a32794a,a32798a,a32799a,a32803a,a32804a,a32805a,a32809a,a32810a,a32814a,a32815a,a32816a,a32820a,a32821a,a32825a,a32826a,a32827a,a32831a,a32832a,a32836a,a32837a,a32838a,a32842a,a32843a,a32847a,a32848a,a32849a,a32853a,a32854a,a32858a,a32859a,a32860a,a32864a,a32865a,a32869a,a32870a,a32871a,a32875a,a32876a,a32880a,a32881a,a32882a,a32886a,a32887a,a32891a,a32892a,a32893a,a32897a,a32898a,a32902a,a32903a,a32904a,a32908a,a32909a,a32913a,a32914a,a32915a,a32919a,a32920a,a32924a,a32925a,a32926a,a32930a,a32931a,a32935a,a32936a,a32937a,a32941a,a32942a,a32946a,a32947a,a32948a,a32952a,a32953a,a32957a,a32958a,a32959a,a32963a,a32964a,a32968a,a32969a,a32970a,a32974a,a32975a,a32979a,a32980a,a32981a,a32985a,a32986a,a32990a,a32991a,a32992a,a32996a,a32997a,a33001a,a33002a,a33003a,a33007a,a33008a,a33012a,a33013a,a33014a,a33018a,a33019a,a33023a,a33024a,a33025a,a33029a,a33030a,a33034a,a33035a,a33036a,a33040a,a33041a,a33045a,a33046a,a33047a,a33051a,a33052a,a33056a,a33057a,a33058a,a33062a,a33063a,a33067a,a33068a,a33069a,a33073a,a33074a,a33078a,a33079a,a33080a,a33084a,a33085a,a33089a,a33090a,a33091a,a33095a,a33096a,a33100a,a33101a,a33102a,a33106a,a33107a,a33111a,a33112a,a33113a,a33117a,a33118a,a33122a,a33123a,a33124a,a33128a,a33129a,a33133a,a33134a,a33135a,a33139a,a33140a,a33144a,a33145a,a33146a,a33150a,a33151a,a33155a,a33156a,a33157a,a33161a,a33162a,a33166a,a33167a,a33168a,a33172a,a33173a,a33177a,a33178a,a33179a,a33183a,a33184a,a33188a,a33189a,a33190a,a33194a,a33195a,a33199a,a33200a,a33201a,a33205a,a33206a,a33210a,a33211a,a33212a,a33216a,a33217a,a33221a,a33222a,a33223a,a33227a,a33228a,a33232a,a33233a,a33234a,a33238a,a33239a,a33243a,a33244a,a33245a,a33249a,a33250a,a33254a,a33255a,a33256a,a33260a,a33261a,a33265a,a33266a,a33267a,a33271a,a33272a,a33276a,a33277a,a33278a,a33282a,a33283a,a33287a,a33288a,a33289a,a33293a,a33294a,a33298a,a33299a,a33300a,a33304a,a33305a,a33309a,a33310a,a33311a,a33315a,a33316a,a33320a,a33321a,a33322a,a33326a,a33327a,a33331a,a33332a,a33333a,a33337a,a33338a,a33342a,a33343a,a33344a,a33348a,a33349a,a33353a,a33354a,a33355a,a33359a,a33360a,a33364a,a33365a,a33366a,a33370a,a33371a,a33375a,a33376a,a33377a,a33381a,a33382a,a33386a,a33387a,a33388a,a33392a,a33393a,a33397a,a33398a,a33399a,a33403a,a33404a,a33408a,a33409a,a33410a,a33414a,a33415a,a33419a,a33420a,a33421a,a33425a,a33426a,a33430a,a33431a,a33432a,a33436a,a33437a,a33441a,a33442a,a33443a,a33447a,a33448a,a33452a,a33453a,a33454a,a33458a,a33459a,a33463a,a33464a,a33465a,a33469a,a33470a,a33474a,a33475a,a33476a,a33480a,a33481a,a33485a,a33486a,a33487a,a33491a,a33492a,a33496a,a33497a,a33498a,a33502a,a33503a,a33507a,a33508a,a33509a,a33513a,a33514a,a33518a,a33519a,a33520a,a33524a,a33525a,a33529a,a33530a,a33531a,a33535a,a33536a,a33540a,a33541a,a33542a,a33546a,a33547a,a33551a,a33552a,a33553a,a33557a,a33558a,a33562a,a33563a,a33564a,a33568a,a33569a,a33573a,a33574a,a33575a,a33579a,a33580a,a33584a,a33585a,a33586a,a33590a,a33591a,a33595a,a33596a,a33597a,a33601a,a33602a,a33606a,a33607a,a33608a,a33612a,a33613a,a33617a,a33618a,a33619a,a33623a,a33624a,a33628a,a33629a,a33630a,a33634a,a33635a,a33639a,a33640a,a33641a,a33645a,a33646a,a33650a,a33651a,a33652a,a33656a,a33657a,a33661a,a33662a,a33663a,a33667a,a33668a,a33672a,a33673a,a33674a,a33678a,a33679a,a33683a,a33684a,a33685a,a33689a,a33690a,a33694a,a33695a,a33696a,a33700a,a33701a,a33705a,a33706a,a33707a,a33711a,a33712a,a33716a,a33717a,a33718a,a33722a,a33723a,a33727a,a33728a,a33729a,a33733a,a33734a,a33738a,a33739a,a33740a,a33744a,a33745a,a33749a,a33750a,a33751a,a33755a,a33756a,a33760a,a33761a,a33762a,a33766a,a33767a,a33771a,a33772a,a33773a,a33777a,a33778a,a33782a,a33783a,a33784a,a33788a,a33789a,a33793a,a33794a,a33795a,a33799a,a33800a,a33804a,a33805a,a33806a,a33810a,a33811a,a33815a,a33816a,a33817a,a33821a,a33822a,a33826a,a33827a,a33828a,a33832a,a33833a,a33837a,a33838a,a33839a,a33843a,a33844a,a33848a,a33849a,a33850a,a33854a,a33855a,a33859a,a33860a,a33861a,a33865a,a33866a,a33870a,a33871a,a33872a,a33876a,a33877a,a33881a,a33882a,a33883a,a33887a,a33888a,a33892a,a33893a,a33894a,a33898a,a33899a,a33903a,a33904a,a33905a,a33909a,a33910a,a33914a,a33915a,a33916a,a33920a,a33921a,a33925a,a33926a,a33927a,a33931a,a33932a,a33936a,a33937a,a33938a,a33942a,a33943a,a33947a,a33948a,a33949a,a33953a,a33954a,a33958a,a33959a,a33960a,a33964a,a33965a,a33969a,a33970a,a33971a,a33975a,a33976a,a33980a,a33981a,a33982a,a33986a,a33987a,a33991a,a33992a,a33993a,a33997a,a33998a,a34002a,a34003a,a34004a,a34008a,a34009a,a34013a,a34014a,a34015a,a34019a,a34020a,a34024a,a34025a,a34026a,a34030a,a34031a,a34035a,a34036a,a34037a,a34041a,a34042a,a34046a,a34047a,a34048a,a34052a,a34053a,a34057a,a34058a,a34059a,a34063a,a34064a,a34068a,a34069a,a34070a,a34074a,a34075a,a34079a,a34080a,a34081a,a34085a,a34086a,a34090a,a34091a,a34092a,a34096a,a34097a,a34101a,a34102a,a34103a,a34107a,a34108a,a34112a,a34113a,a34114a,a34118a,a34119a,a34123a,a34124a,a34125a,a34129a,a34130a,a34134a,a34135a,a34136a,a34140a,a34141a,a34145a,a34146a,a34147a,a34151a,a34152a,a34156a,a34157a,a34158a,a34162a,a34163a,a34167a,a34168a,a34169a,a34173a,a34174a,a34178a,a34179a,a34180a,a34184a,a34185a,a34189a,a34190a,a34191a,a34195a,a34196a,a34200a,a34201a,a34202a,a34206a,a34207a,a34211a,a34212a,a34213a,a34217a,a34218a,a34222a,a34223a,a34224a,a34228a,a34229a,a34233a,a34234a,a34235a,a34239a,a34240a,a34244a,a34245a,a34246a,a34250a,a34251a,a34255a,a34256a,a34257a,a34261a,a34262a,a34266a,a34267a,a34268a,a34272a,a34273a,a34277a,a34278a,a34279a,a34283a,a34284a,a34288a,a34289a,a34290a,a34294a,a34295a,a34299a,a34300a,a34301a,a34305a,a34306a,a34310a,a34311a,a34312a,a34316a,a34317a,a34321a,a34322a,a34323a,a34327a,a34328a,a34332a,a34333a,a34334a,a34338a,a34339a,a34343a,a34344a,a34345a,a34349a,a34350a,a34354a,a34355a,a34356a,a34360a,a34361a,a34365a,a34366a,a34367a,a34371a,a34372a,a34376a,a34377a,a34378a,a34382a,a34383a,a34387a,a34388a,a34389a,a34393a,a34394a,a34398a,a34399a,a34400a,a34404a,a34405a,a34409a,a34410a,a34411a,a34415a,a34416a,a34420a,a34421a,a34422a,a34426a,a34427a,a34431a,a34432a,a34433a,a34437a,a34438a,a34442a,a34443a,a34444a,a34448a,a34449a,a34453a,a34454a,a34455a,a34459a,a34460a,a34464a,a34465a,a34466a,a34470a,a34471a,a34475a,a34476a,a34477a,a34481a,a34482a,a34486a,a34487a,a34488a,a34492a,a34493a,a34497a,a34498a,a34499a,a34503a,a34504a,a34508a,a34509a,a34510a,a34514a,a34515a,a34519a,a34520a,a34521a,a34525a,a34526a,a34530a,a34531a,a34532a,a34536a,a34537a,a34541a,a34542a,a34543a,a34547a,a34548a,a34552a,a34553a,a34554a,a34558a,a34559a,a34563a,a34564a,a34565a,a34569a,a34570a,a34574a,a34575a,a34576a,a34580a,a34581a,a34585a,a34586a,a34587a,a34591a,a34592a,a34596a,a34597a,a34598a,a34602a,a34603a,a34607a,a34608a,a34609a,a34613a,a34614a,a34618a,a34619a,a34620a,a34624a,a34625a,a34629a,a34630a,a34631a,a34635a,a34636a,a34640a,a34641a,a34642a,a34646a,a34647a,a34651a,a34652a,a34653a,a34657a,a34658a,a34662a,a34663a,a34664a,a34668a,a34669a,a34673a,a34674a,a34675a,a34679a,a34680a,a34684a,a34685a,a34686a,a34690a,a34691a,a34695a,a34696a,a34697a,a34701a,a34702a,a34706a,a34707a,a34708a,a34712a,a34713a,a34717a,a34718a,a34719a,a34723a,a34724a,a34728a,a34729a,a34730a,a34734a,a34735a,a34739a,a34740a,a34741a,a34745a,a34746a,a34750a,a34751a,a34752a,a34756a,a34757a,a34761a,a34762a,a34763a,a34767a,a34768a,a34772a,a34773a,a34774a,a34778a,a34779a,a34783a,a34784a,a34785a,a34789a,a34790a,a34794a,a34795a,a34796a,a34800a,a34801a,a34805a,a34806a,a34807a,a34811a,a34812a,a34816a,a34817a,a34818a,a34822a,a34823a,a34827a,a34828a,a34829a,a34833a,a34834a,a34838a,a34839a,a34840a,a34844a,a34845a,a34849a,a34850a,a34851a,a34855a,a34856a,a34860a,a34861a,a34862a,a34866a,a34867a,a34871a,a34872a,a34873a,a34877a,a34878a,a34882a,a34883a,a34884a,a34888a,a34889a,a34893a,a34894a,a34895a,a34899a,a34900a,a34904a,a34905a,a34906a,a34910a,a34911a,a34915a,a34916a,a34917a,a34921a,a34922a,a34926a,a34927a,a34928a,a34932a,a34933a,a34937a,a34938a,a34939a,a34943a,a34944a,a34948a,a34949a,a34950a,a34954a,a34955a,a34959a,a34960a,a34961a,a34965a,a34966a,a34970a,a34971a,a34972a,a34976a,a34977a,a34981a,a34982a,a34983a,a34987a,a34988a,a34992a,a34993a,a34994a,a34998a,a34999a,a35003a,a35004a,a35005a,a35009a,a35010a,a35014a,a35015a,a35016a,a35020a,a35021a,a35025a,a35026a,a35027a,a35031a,a35032a,a35036a,a35037a,a35038a,a35042a,a35043a,a35047a,a35048a,a35049a,a35053a,a35054a,a35058a,a35059a,a35060a,a35064a,a35065a,a35069a,a35070a,a35071a,a35075a,a35076a,a35080a,a35081a,a35082a,a35086a,a35087a,a35091a,a35092a,a35093a,a35097a,a35098a,a35102a,a35103a,a35104a,a35108a,a35109a,a35113a,a35114a,a35115a,a35119a,a35120a,a35124a,a35125a,a35126a,a35130a,a35131a,a35135a,a35136a,a35137a,a35141a,a35142a,a35146a,a35147a,a35148a,a35152a,a35153a,a35157a,a35158a,a35159a,a35163a,a35164a,a35168a,a35169a,a35170a,a35174a,a35175a,a35179a,a35180a,a35181a,a35185a,a35186a,a35190a,a35191a,a35192a,a35196a,a35197a,a35201a,a35202a,a35203a,a35207a,a35208a,a35212a,a35213a,a35214a,a35218a,a35219a,a35223a,a35224a,a35225a,a35229a,a35230a,a35234a,a35235a,a35236a,a35240a,a35241a,a35245a,a35246a,a35247a,a35251a,a35252a,a35256a,a35257a,a35258a,a35262a,a35263a,a35267a,a35268a,a35269a,a35273a,a35274a,a35278a,a35279a,a35280a,a35284a,a35285a,a35289a,a35290a,a35291a,a35295a,a35296a,a35300a,a35301a,a35302a,a35306a,a35307a,a35311a,a35312a,a35313a,a35317a,a35318a,a35322a,a35323a,a35324a,a35328a,a35329a,a35333a,a35334a,a35335a,a35339a,a35340a,a35344a,a35345a,a35346a,a35350a,a35351a,a35355a,a35356a,a35357a,a35361a,a35362a,a35366a,a35367a,a35368a,a35372a,a35373a,a35377a,a35378a,a35379a,a35383a,a35384a,a35388a,a35389a,a35390a,a35394a,a35395a,a35399a,a35400a,a35401a,a35405a,a35406a,a35410a,a35411a,a35412a,a35416a,a35417a,a35421a,a35422a,a35423a,a35427a,a35428a,a35432a,a35433a,a35434a,a35438a,a35439a,a35443a,a35444a,a35445a,a35449a,a35450a,a35454a,a35455a,a35456a,a35460a,a35461a,a35465a,a35466a,a35467a,a35471a,a35472a,a35476a,a35477a,a35478a,a35482a,a35483a,a35487a,a35488a,a35489a,a35493a,a35494a,a35498a,a35499a,a35500a,a35504a,a35505a,a35509a,a35510a,a35511a,a35515a,a35516a,a35520a,a35521a,a35522a,a35526a,a35527a,a35531a,a35532a,a35533a,a35537a,a35538a,a35542a,a35543a,a35544a,a35548a,a35549a,a35553a,a35554a,a35555a,a35559a,a35560a,a35564a,a35565a,a35566a,a35570a,a35571a,a35575a,a35576a,a35577a,a35581a,a35582a,a35586a,a35587a,a35588a,a35592a,a35593a,a35597a,a35598a,a35599a,a35603a,a35604a,a35608a,a35609a,a35610a,a35614a,a35615a,a35619a,a35620a,a35621a,a35625a,a35626a,a35630a,a35631a,a35632a,a35636a,a35637a,a35641a,a35642a,a35643a,a35647a,a35648a,a35652a,a35653a,a35654a,a35658a,a35659a,a35663a,a35664a,a35665a,a35669a,a35670a,a35674a,a35675a,a35676a,a35680a,a35681a,a35685a,a35686a,a35687a,a35691a,a35692a,a35696a,a35697a,a35698a,a35702a,a35703a,a35707a,a35708a,a35709a,a35713a,a35714a,a35718a,a35719a,a35720a,a35724a,a35725a,a35729a,a35730a,a35731a,a35735a,a35736a,a35740a,a35741a,a35742a,a35746a,a35747a,a35751a,a35752a,a35753a,a35757a,a35758a,a35762a,a35763a,a35764a,a35768a,a35769a,a35773a,a35774a,a35775a,a35779a,a35780a,a35784a,a35785a,a35786a,a35790a,a35791a,a35795a,a35796a,a35797a,a35801a,a35802a,a35806a,a35807a,a35808a,a35812a,a35813a,a35817a,a35818a,a35819a,a35823a,a35824a,a35828a,a35829a,a35830a,a35834a,a35835a,a35839a,a35840a,a35841a,a35845a,a35846a,a35850a,a35851a,a35852a,a35856a,a35857a,a35861a,a35862a,a35863a,a35867a,a35868a,a35872a,a35873a,a35874a,a35878a,a35879a,a35883a,a35884a,a35885a,a35889a,a35890a,a35894a,a35895a,a35896a,a35900a,a35901a,a35905a,a35906a,a35907a,a35911a,a35912a,a35916a,a35917a,a35918a,a35922a,a35923a,a35927a,a35928a,a35929a,a35933a,a35934a,a35938a,a35939a,a35940a,a35944a,a35945a,a35949a,a35950a,a35951a,a35955a,a35956a,a35960a,a35961a,a35962a,a35966a,a35967a,a35971a,a35972a,a35973a,a35977a,a35978a,a35982a,a35983a,a35984a,a35988a,a35989a,a35993a,a35994a,a35995a,a35999a,a36000a,a36004a,a36005a,a36006a,a36010a,a36011a,a36015a,a36016a,a36017a,a36021a,a36022a,a36026a,a36027a,a36028a,a36032a,a36033a,a36037a,a36038a,a36039a,a36043a,a36044a,a36048a,a36049a,a36050a,a36054a,a36055a,a36059a,a36060a,a36061a,a36065a,a36066a,a36070a,a36071a,a36072a,a36076a,a36077a,a36081a,a36082a,a36083a,a36087a,a36088a,a36092a,a36093a,a36094a,a36098a,a36099a,a36103a,a36104a,a36105a,a36109a,a36110a,a36114a,a36115a,a36116a,a36120a,a36121a,a36125a,a36126a,a36127a,a36131a,a36132a,a36136a,a36137a,a36138a,a36142a,a36143a,a36147a,a36148a,a36149a,a36153a,a36154a,a36158a,a36159a,a36160a,a36164a,a36165a,a36169a,a36170a,a36171a,a36175a,a36176a,a36180a,a36181a,a36182a,a36186a,a36187a,a36191a,a36192a,a36193a,a36197a,a36198a,a36202a,a36203a,a36204a,a36208a,a36209a,a36213a,a36214a,a36215a,a36219a,a36220a,a36224a,a36225a,a36226a,a36230a,a36231a,a36235a,a36236a,a36237a,a36241a,a36242a,a36246a,a36247a,a36248a,a36252a,a36253a,a36257a,a36258a,a36259a,a36263a,a36264a,a36268a,a36269a,a36270a,a36274a,a36275a,a36279a,a36280a,a36281a,a36285a,a36286a,a36290a,a36291a,a36292a,a36296a,a36297a,a36301a,a36302a,a36303a,a36307a,a36308a,a36312a,a36313a,a36314a,a36318a,a36319a,a36323a,a36324a,a36325a,a36329a,a36330a,a36334a,a36335a,a36336a,a36340a,a36341a,a36345a,a36346a,a36347a,a36351a,a36352a,a36356a,a36357a,a36358a,a36362a,a36363a,a36367a,a36368a,a36369a,a36373a,a36374a,a36378a,a36379a,a36380a,a36384a,a36385a,a36389a,a36390a,a36391a,a36395a,a36396a,a36400a,a36401a,a36402a,a36406a,a36407a,a36411a,a36412a,a36413a,a36417a,a36418a,a36422a,a36423a,a36424a,a36428a,a36429a,a36433a,a36434a,a36435a,a36439a,a36440a,a36444a,a36445a,a36446a,a36450a,a36451a,a36455a,a36456a,a36457a,a36461a,a36462a,a36466a,a36467a,a36468a,a36472a,a36473a,a36477a,a36478a,a36479a,a36483a,a36484a,a36488a,a36489a,a36490a,a36494a,a36495a,a36499a,a36500a,a36501a,a36505a,a36506a,a36510a,a36511a,a36512a,a36516a,a36517a,a36521a,a36522a,a36523a,a36527a,a36528a,a36532a,a36533a,a36534a,a36538a,a36539a,a36543a,a36544a,a36545a,a36549a,a36550a,a36554a,a36555a,a36556a,a36560a,a36561a,a36565a,a36566a,a36567a,a36571a,a36572a,a36576a,a36577a,a36578a,a36582a,a36583a,a36587a,a36588a,a36589a,a36593a,a36594a,a36598a,a36599a,a36600a,a36604a,a36605a,a36609a,a36610a,a36611a,a36615a,a36616a,a36620a,a36621a,a36622a,a36626a,a36627a,a36631a,a36632a,a36633a,a36637a,a36638a,a36642a,a36643a,a36644a,a36648a,a36649a,a36653a,a36654a,a36655a,a36659a,a36660a,a36664a,a36665a,a36666a,a36670a,a36671a,a36675a,a36676a,a36677a,a36681a,a36682a,a36686a,a36687a,a36688a,a36692a,a36693a,a36697a,a36698a,a36699a,a36703a,a36704a,a36708a,a36709a,a36710a,a36714a,a36715a,a36719a,a36720a,a36721a,a36725a,a36726a,a36730a,a36731a,a36732a,a36736a,a36737a,a36741a,a36742a,a36743a,a36747a,a36748a,a36752a,a36753a,a36754a,a36758a,a36759a,a36763a,a36764a,a36765a,a36769a,a36770a,a36774a,a36775a,a36776a,a36780a,a36781a,a36785a,a36786a,a36787a,a36791a,a36792a,a36796a,a36797a,a36798a,a36802a,a36803a,a36807a,a36808a,a36809a,a36813a,a36814a,a36818a,a36819a,a36820a,a36824a,a36825a,a36829a,a36830a,a36831a,a36835a,a36836a,a36840a,a36841a,a36842a,a36846a,a36847a,a36851a,a36852a,a36853a,a36857a,a36858a,a36862a,a36863a,a36864a,a36868a,a36869a,a36873a,a36874a,a36875a,a36879a,a36880a,a36884a,a36885a,a36886a,a36890a,a36891a,a36895a,a36896a,a36897a,a36901a,a36902a,a36906a,a36907a,a36908a,a36912a,a36913a,a36917a,a36918a,a36919a,a36923a,a36924a,a36928a,a36929a,a36930a,a36934a,a36935a,a36939a,a36940a,a36941a,a36945a,a36946a,a36950a,a36951a,a36952a,a36956a,a36957a,a36961a,a36962a,a36963a,a36967a,a36968a,a36972a,a36973a,a36974a,a36978a,a36979a,a36983a,a36984a,a36985a,a36989a,a36990a,a36994a,a36995a,a36996a,a37000a,a37001a,a37005a,a37006a,a37007a,a37011a,a37012a,a37016a,a37017a,a37018a,a37022a,a37023a,a37027a,a37028a,a37029a,a37033a,a37034a,a37038a,a37039a,a37040a,a37044a,a37045a,a37049a,a37050a,a37051a,a37055a,a37056a,a37060a,a37061a,a37062a,a37066a,a37067a,a37071a,a37072a,a37073a,a37077a,a37078a,a37082a,a37083a,a37084a,a37088a,a37089a,a37093a,a37094a,a37095a,a37099a,a37100a,a37104a,a37105a,a37106a,a37110a,a37111a,a37115a,a37116a,a37117a,a37121a,a37122a,a37126a,a37127a,a37128a,a37132a,a37133a,a37137a,a37138a,a37139a,a37143a,a37144a,a37148a,a37149a,a37150a,a37154a,a37155a,a37159a,a37160a,a37161a,a37165a,a37166a,a37170a,a37171a,a37172a,a37176a,a37177a,a37181a,a37182a,a37183a,a37187a,a37188a,a37192a,a37193a,a37194a,a37198a,a37199a,a37203a,a37204a,a37205a,a37209a,a37210a,a37214a,a37215a,a37216a,a37220a,a37221a,a37225a,a37226a,a37227a,a37231a,a37232a,a37236a,a37237a,a37238a,a37242a,a37243a,a37247a,a37248a,a37249a,a37253a,a37254a,a37258a,a37259a,a37260a,a37264a,a37265a,a37269a,a37270a,a37271a,a37275a,a37276a,a37280a,a37281a,a37282a,a37286a,a37287a,a37291a,a37292a,a37293a,a37297a,a37298a,a37302a,a37303a,a37304a,a37308a,a37309a,a37313a,a37314a,a37315a,a37319a,a37320a,a37324a,a37325a,a37326a,a37330a,a37331a,a37335a,a37336a,a37337a,a37341a,a37342a,a37346a,a37347a,a37348a,a37352a,a37353a,a37357a,a37358a,a37359a,a37363a,a37364a,a37368a,a37369a,a37370a,a37374a,a37375a,a37379a,a37380a,a37381a,a37385a,a37386a,a37390a,a37391a,a37392a,a37396a,a37397a,a37401a,a37402a,a37403a,a37407a,a37408a,a37412a,a37413a,a37414a,a37418a,a37419a,a37423a,a37424a,a37425a,a37429a,a37430a,a37434a,a37435a,a37436a,a37440a,a37441a,a37445a,a37446a,a37447a,a37451a,a37452a,a37456a,a37457a,a37458a,a37462a,a37463a,a37467a,a37468a,a37469a,a37473a,a37474a,a37478a,a37479a,a37480a,a37484a,a37485a,a37489a,a37490a,a37491a,a37495a,a37496a,a37500a,a37501a,a37502a,a37506a,a37507a,a37511a,a37512a,a37513a,a37517a,a37518a,a37522a,a37523a,a37524a,a37528a,a37529a,a37533a,a37534a,a37535a,a37539a,a37540a,a37544a,a37545a,a37546a,a37550a,a37551a,a37555a,a37556a,a37557a,a37561a,a37562a,a37566a,a37567a,a37568a,a37572a,a37573a,a37577a,a37578a,a37579a,a37583a,a37584a,a37588a,a37589a,a37590a,a37594a,a37595a,a37599a,a37600a,a37601a,a37605a,a37606a,a37610a,a37611a,a37612a,a37616a,a37617a,a37621a,a37622a,a37623a,a37627a,a37628a,a37632a,a37633a,a37634a,a37638a,a37639a,a37643a,a37644a,a37645a,a37649a,a37650a,a37654a,a37655a,a37656a,a37660a,a37661a,a37665a,a37666a,a37667a,a37671a,a37672a,a37676a,a37677a,a37678a,a37682a,a37683a,a37687a,a37688a,a37689a,a37693a,a37694a,a37698a,a37699a,a37700a,a37704a,a37705a,a37709a,a37710a,a37711a,a37715a,a37716a,a37720a,a37721a,a37722a,a37726a,a37727a,a37731a,a37732a,a37733a,a37737a,a37738a,a37742a,a37743a,a37744a,a37748a,a37749a,a37753a,a37754a,a37755a,a37759a,a37760a,a37764a,a37765a,a37766a,a37770a,a37771a,a37775a,a37776a,a37777a,a37781a,a37782a,a37786a,a37787a,a37788a,a37792a,a37793a,a37797a,a37798a,a37799a,a37803a,a37804a,a37808a,a37809a,a37810a,a37814a,a37815a,a37819a,a37820a,a37821a,a37825a,a37826a,a37830a,a37831a,a37832a,a37836a,a37837a,a37841a,a37842a,a37843a,a37847a,a37848a,a37852a,a37853a,a37854a,a37858a,a37859a,a37863a,a37864a,a37865a,a37869a,a37870a,a37874a,a37875a,a37876a,a37880a,a37881a,a37885a,a37886a,a37887a,a37891a,a37892a,a37896a,a37897a,a37898a,a37902a,a37903a,a37907a,a37908a,a37909a,a37913a,a37914a,a37918a,a37919a,a37920a,a37924a,a37925a,a37929a,a37930a,a37931a,a37935a,a37936a,a37940a,a37941a,a37942a,a37946a,a37947a,a37951a,a37952a,a37953a,a37957a,a37958a,a37962a,a37963a,a37964a,a37968a,a37969a,a37973a,a37974a,a37975a,a37979a,a37980a,a37984a,a37985a,a37986a,a37990a,a37991a,a37995a,a37996a,a37997a,a38001a,a38002a,a38006a,a38007a,a38008a,a38012a,a38013a,a38017a,a38018a,a38019a,a38023a,a38024a,a38028a,a38029a,a38030a,a38034a,a38035a,a38039a,a38040a,a38041a,a38045a,a38046a,a38050a,a38051a,a38052a,a38056a,a38057a,a38061a,a38062a,a38063a,a38067a,a38068a,a38072a,a38073a,a38074a,a38078a,a38079a,a38083a,a38084a,a38085a,a38089a,a38090a,a38094a,a38095a,a38096a,a38100a,a38101a,a38105a,a38106a,a38107a,a38111a,a38112a,a38116a,a38117a,a38118a,a38122a,a38123a,a38127a,a38128a,a38129a,a38133a,a38134a,a38138a,a38139a,a38140a,a38144a,a38145a,a38149a,a38150a,a38151a,a38155a,a38156a,a38160a,a38161a,a38162a,a38166a,a38167a,a38171a,a38172a,a38173a,a38177a,a38178a,a38182a,a38183a,a38184a,a38188a,a38189a,a38193a,a38194a,a38195a,a38199a,a38200a,a38204a,a38205a,a38206a,a38210a,a38211a,a38215a,a38216a,a38217a,a38221a,a38222a,a38226a,a38227a,a38228a,a38232a,a38233a,a38237a,a38238a,a38239a,a38243a,a38244a,a38248a,a38249a,a38250a,a38254a,a38255a,a38259a,a38260a,a38261a,a38265a,a38266a,a38270a,a38271a,a38272a,a38276a,a38277a,a38281a,a38282a,a38283a,a38287a,a38288a,a38292a,a38293a,a38294a,a38298a,a38299a,a38303a,a38304a,a38305a,a38309a,a38310a,a38314a,a38315a,a38316a,a38320a,a38321a,a38325a,a38326a,a38327a,a38331a,a38332a,a38336a,a38337a,a38338a,a38342a,a38343a,a38347a,a38348a,a38349a,a38353a,a38354a,a38358a,a38359a,a38360a,a38364a,a38365a,a38369a,a38370a,a38371a,a38375a,a38376a,a38380a,a38381a,a38382a,a38386a,a38387a,a38391a,a38392a,a38393a,a38397a,a38398a,a38402a,a38403a,a38404a,a38408a,a38409a,a38413a,a38414a,a38415a,a38419a,a38420a,a38424a,a38425a,a38426a,a38430a,a38431a,a38435a,a38436a,a38437a,a38441a,a38442a,a38446a,a38447a,a38448a,a38452a,a38453a,a38457a,a38458a,a38459a,a38463a,a38464a,a38468a,a38469a,a38470a,a38474a,a38475a,a38479a,a38480a,a38481a,a38485a,a38486a,a38490a,a38491a,a38492a,a38496a,a38497a,a38501a,a38502a,a38503a,a38507a,a38508a,a38512a,a38513a,a38514a,a38518a,a38519a,a38523a,a38524a,a38525a,a38529a,a38530a,a38534a,a38535a,a38536a,a38540a,a38541a,a38545a,a38546a,a38547a,a38551a,a38552a,a38556a,a38557a,a38558a,a38562a,a38563a,a38567a,a38568a,a38569a,a38573a,a38574a,a38578a,a38579a,a38580a,a38584a,a38585a,a38589a,a38590a,a38591a,a38595a,a38596a,a38600a,a38601a,a38602a,a38606a,a38607a,a38611a,a38612a,a38613a,a38617a,a38618a,a38622a,a38623a,a38624a,a38628a,a38629a,a38633a,a38634a,a38635a,a38639a,a38640a,a38644a,a38645a,a38646a,a38650a,a38651a,a38655a,a38656a,a38657a,a38661a,a38662a,a38666a,a38667a,a38668a,a38672a,a38673a,a38677a,a38678a,a38679a,a38683a,a38684a,a38688a,a38689a,a38690a,a38694a,a38695a,a38699a,a38700a,a38701a,a38705a,a38706a,a38710a,a38711a,a38712a,a38716a,a38717a,a38721a,a38722a,a38723a,a38727a,a38728a,a38732a,a38733a,a38734a,a38738a,a38739a,a38743a,a38744a,a38745a,a38749a,a38750a,a38754a,a38755a,a38756a,a38760a,a38761a,a38765a,a38766a,a38767a,a38771a,a38772a,a38776a,a38777a,a38778a,a38782a,a38783a,a38787a,a38788a,a38789a,a38793a,a38794a,a38798a,a38799a,a38800a,a38804a,a38805a,a38809a,a38810a,a38811a,a38815a,a38816a,a38820a,a38821a,a38822a,a38826a,a38827a,a38831a,a38832a,a38833a,a38837a,a38838a,a38842a,a38843a,a38844a,a38848a,a38849a,a38853a,a38854a,a38855a,a38859a,a38860a,a38864a,a38865a,a38866a,a38870a,a38871a,a38875a,a38876a,a38877a,a38881a,a38882a,a38886a,a38887a,a38888a,a38892a,a38893a,a38897a,a38898a,a38899a,a38903a,a38904a,a38908a,a38909a,a38910a,a38914a,a38915a,a38919a,a38920a,a38921a,a38925a,a38926a,a38930a,a38931a,a38932a,a38936a,a38937a,a38941a,a38942a,a38943a,a38947a,a38948a,a38952a,a38953a,a38954a,a38958a,a38959a,a38963a,a38964a,a38965a,a38969a,a38970a,a38974a,a38975a,a38976a,a38980a,a38981a,a38985a,a38986a,a38987a,a38991a,a38992a,a38996a,a38997a,a38998a,a39002a,a39003a,a39007a,a39008a,a39009a,a39013a,a39014a,a39018a,a39019a,a39020a,a39024a,a39025a,a39029a,a39030a,a39031a,a39035a,a39036a,a39040a,a39041a,a39042a,a39046a,a39047a,a39051a,a39052a,a39053a,a39057a,a39058a,a39062a,a39063a,a39064a,a39068a,a39069a,a39073a,a39074a,a39075a,a39079a,a39080a,a39084a,a39085a,a39086a,a39090a,a39091a,a39095a,a39096a,a39097a,a39101a,a39102a,a39106a,a39107a,a39108a,a39112a,a39113a,a39117a,a39118a,a39119a,a39123a,a39124a,a39128a,a39129a,a39130a,a39134a,a39135a,a39139a,a39140a,a39141a,a39145a,a39146a,a39150a,a39151a,a39152a,a39156a,a39157a,a39161a,a39162a,a39163a,a39167a,a39168a,a39172a,a39173a,a39174a,a39178a,a39179a,a39183a,a39184a,a39185a,a39189a,a39190a,a39194a,a39195a,a39196a,a39200a,a39201a,a39205a,a39206a,a39207a,a39211a,a39212a,a39216a,a39217a,a39218a,a39222a,a39223a,a39227a,a39228a,a39229a,a39233a,a39234a,a39238a,a39239a,a39240a,a39244a,a39245a,a39249a,a39250a,a39251a,a39255a,a39256a,a39260a,a39261a,a39262a,a39266a,a39267a,a39271a,a39272a,a39273a,a39277a,a39278a,a39282a,a39283a,a39284a,a39288a,a39289a,a39293a,a39294a,a39295a,a39299a,a39300a,a39304a,a39305a,a39306a,a39310a,a39311a,a39315a,a39316a,a39317a,a39321a,a39322a,a39326a,a39327a,a39328a,a39332a,a39333a,a39337a,a39338a,a39339a,a39343a,a39344a,a39348a,a39349a,a39350a,a39354a,a39355a,a39359a,a39360a,a39361a,a39365a,a39366a,a39370a,a39371a,a39372a,a39376a,a39377a,a39381a,a39382a,a39383a,a39387a,a39388a,a39392a,a39393a,a39394a,a39398a,a39399a,a39403a,a39404a,a39405a,a39409a,a39410a,a39414a,a39415a,a39416a,a39420a,a39421a,a39425a,a39426a,a39427a,a39431a,a39432a,a39436a,a39437a,a39438a,a39442a,a39443a,a39447a,a39448a,a39449a,a39453a,a39454a,a39458a,a39459a,a39460a,a39464a,a39465a,a39469a,a39470a,a39471a,a39475a,a39476a,a39480a,a39481a,a39482a,a39486a,a39487a,a39491a,a39492a,a39493a,a39497a,a39498a,a39502a,a39503a,a39504a,a39508a,a39509a,a39513a,a39514a,a39515a,a39519a,a39520a,a39524a,a39525a,a39526a,a39530a,a39531a,a39535a,a39536a,a39537a,a39541a,a39542a,a39546a,a39547a,a39548a,a39552a,a39553a,a39557a,a39558a,a39559a,a39563a,a39564a,a39568a,a39569a,a39570a,a39574a,a39575a,a39579a,a39580a,a39581a,a39585a,a39586a,a39590a,a39591a,a39592a,a39596a,a39597a,a39601a,a39602a,a39603a,a39607a,a39608a,a39612a,a39613a,a39614a,a39618a,a39619a,a39623a,a39624a,a39625a,a39629a,a39630a,a39634a,a39635a,a39636a,a39640a,a39641a,a39645a,a39646a,a39647a,a39651a,a39652a,a39656a,a39657a,a39658a,a39662a,a39663a,a39667a,a39668a,a39669a,a39673a,a39674a,a39678a,a39679a,a39680a,a39684a,a39685a,a39689a,a39690a,a39691a,a39695a,a39696a,a39700a,a39701a,a39702a,a39706a,a39707a,a39711a,a39712a,a39713a,a39717a,a39718a,a39722a,a39723a,a39724a,a39728a,a39729a,a39733a,a39734a,a39735a,a39739a,a39740a,a39744a,a39745a,a39746a,a39750a,a39751a,a39755a,a39756a,a39757a,a39761a,a39762a,a39766a,a39767a,a39768a,a39772a,a39773a,a39777a,a39778a,a39779a,a39783a,a39784a,a39788a,a39789a,a39790a,a39794a,a39795a,a39799a,a39800a,a39801a,a39805a,a39806a,a39810a,a39811a,a39812a,a39816a,a39817a,a39821a,a39822a,a39823a,a39827a,a39828a,a39832a,a39833a,a39834a,a39838a,a39839a,a39843a,a39844a,a39845a,a39849a,a39850a,a39854a,a39855a,a39856a,a39860a,a39861a,a39865a,a39866a,a39867a,a39871a,a39872a,a39876a,a39877a,a39878a,a39882a,a39883a,a39887a,a39888a,a39889a,a39893a,a39894a,a39898a,a39899a,a39900a,a39904a,a39905a,a39909a,a39910a,a39911a,a39915a,a39916a,a39920a,a39921a,a39922a,a39926a,a39927a,a39931a,a39932a,a39933a,a39937a,a39938a,a39942a,a39943a,a39944a,a39948a,a39949a,a39953a,a39954a,a39955a,a39959a,a39960a,a39964a,a39965a,a39966a,a39970a,a39971a,a39975a,a39976a,a39977a,a39981a,a39982a,a39986a,a39987a,a39988a,a39992a,a39993a,a39997a,a39998a,a39999a,a40003a,a40004a,a40008a,a40009a,a40010a,a40014a,a40015a,a40019a,a40020a,a40021a,a40025a,a40026a,a40030a,a40031a,a40032a,a40036a,a40037a,a40041a,a40042a,a40043a,a40047a,a40048a,a40052a,a40053a,a40054a,a40058a,a40059a,a40063a,a40064a,a40065a,a40069a,a40070a,a40074a,a40075a,a40076a,a40080a,a40081a,a40085a,a40086a,a40087a,a40091a,a40092a,a40096a,a40097a,a40098a,a40102a,a40103a,a40107a,a40108a,a40109a,a40113a,a40114a,a40118a,a40119a,a40120a,a40124a,a40125a,a40129a,a40130a,a40131a,a40135a,a40136a,a40140a,a40141a,a40142a,a40146a,a40147a,a40151a,a40152a,a40153a,a40157a,a40158a,a40162a,a40163a,a40164a,a40168a,a40169a,a40173a,a40174a,a40175a,a40179a,a40180a,a40184a,a40185a,a40186a,a40190a,a40191a,a40195a,a40196a,a40197a,a40201a,a40202a,a40206a,a40207a,a40208a,a40212a,a40213a,a40217a,a40218a,a40219a,a40223a,a40224a,a40228a,a40229a,a40230a,a40234a,a40235a,a40239a,a40240a,a40241a,a40245a,a40246a,a40250a,a40251a,a40252a,a40256a,a40257a,a40261a,a40262a,a40263a,a40267a,a40268a,a40272a,a40273a,a40274a,a40278a,a40279a,a40283a,a40284a,a40285a,a40289a,a40290a,a40294a,a40295a,a40296a,a40300a,a40301a,a40305a,a40306a,a40307a,a40311a,a40312a,a40316a,a40317a,a40318a,a40322a,a40323a,a40327a,a40328a,a40329a,a40333a,a40334a,a40338a,a40339a,a40340a,a40344a,a40345a,a40349a,a40350a,a40351a,a40355a,a40356a,a40360a,a40361a,a40362a,a40366a,a40367a,a40371a,a40372a,a40373a,a40377a,a40378a,a40382a,a40383a,a40384a,a40388a,a40389a,a40393a,a40394a,a40395a,a40399a,a40400a,a40404a,a40405a,a40406a,a40410a,a40411a,a40415a,a40416a,a40417a,a40421a,a40422a,a40426a,a40427a,a40428a,a40432a,a40433a,a40437a,a40438a,a40439a,a40443a,a40444a,a40448a,a40449a,a40450a,a40454a,a40455a,a40459a,a40460a,a40461a,a40465a,a40466a,a40470a,a40471a,a40472a,a40476a,a40477a,a40481a,a40482a,a40483a,a40487a,a40488a,a40492a,a40493a,a40494a,a40498a,a40499a,a40503a,a40504a,a40505a,a40509a,a40510a,a40514a,a40515a,a40516a,a40520a,a40521a,a40525a,a40526a,a40527a,a40531a,a40532a,a40536a,a40537a,a40538a,a40542a,a40543a,a40547a,a40548a,a40549a,a40553a,a40554a,a40558a,a40559a,a40560a,a40564a,a40565a,a40569a,a40570a,a40571a,a40575a,a40576a,a40580a,a40581a,a40582a,a40586a,a40587a,a40591a,a40592a,a40593a,a40597a,a40598a,a40602a,a40603a,a40604a,a40608a,a40609a,a40613a,a40614a,a40615a,a40619a,a40620a,a40624a,a40625a,a40626a,a40630a,a40631a,a40635a,a40636a,a40637a,a40641a,a40642a,a40646a,a40647a,a40648a,a40652a,a40653a,a40657a,a40658a,a40659a,a40663a,a40664a,a40668a,a40669a,a40670a,a40674a,a40675a,a40679a,a40680a,a40681a,a40685a,a40686a,a40690a,a40691a,a40692a,a40696a,a40697a,a40701a,a40702a,a40703a,a40707a,a40708a,a40712a,a40713a,a40714a,a40718a,a40719a,a40723a,a40724a,a40725a,a40729a,a40730a,a40734a,a40735a,a40736a,a40740a,a40741a,a40745a,a40746a,a40747a,a40751a,a40752a,a40756a,a40757a,a40758a,a40762a,a40763a,a40767a,a40768a,a40769a,a40773a,a40774a,a40778a,a40779a,a40780a,a40784a,a40785a,a40789a,a40790a,a40791a,a40795a,a40796a,a40800a,a40801a,a40802a,a40806a,a40807a,a40811a,a40812a,a40813a,a40817a,a40818a,a40822a,a40823a,a40824a,a40828a,a40829a,a40833a,a40834a,a40835a,a40839a,a40840a,a40844a,a40845a,a40846a,a40850a,a40851a,a40855a,a40856a,a40857a,a40861a,a40862a,a40866a,a40867a,a40868a,a40872a,a40873a,a40877a,a40878a,a40879a,a40883a,a40884a,a40888a,a40889a,a40890a,a40894a,a40895a,a40899a,a40900a,a40901a,a40905a,a40906a,a40910a,a40911a,a40912a,a40916a,a40917a,a40921a,a40922a,a40923a,a40927a,a40928a,a40932a,a40933a,a40934a,a40938a,a40939a,a40943a,a40944a,a40945a,a40949a,a40950a,a40954a,a40955a,a40956a,a40960a,a40961a,a40965a,a40966a,a40967a,a40971a,a40972a,a40976a,a40977a,a40978a,a40982a,a40983a,a40987a,a40988a,a40989a,a40993a,a40994a,a40998a,a40999a,a41000a,a41004a,a41005a,a41009a,a41010a,a41011a,a41015a,a41016a,a41020a,a41021a,a41022a,a41026a,a41027a,a41031a,a41032a,a41033a,a41037a,a41038a,a41042a,a41043a,a41044a,a41048a,a41049a,a41053a,a41054a,a41055a,a41059a,a41060a,a41064a,a41065a,a41066a,a41070a,a41071a,a41075a,a41076a,a41077a,a41081a,a41082a,a41086a,a41087a,a41088a,a41092a,a41093a,a41097a,a41098a,a41099a,a41103a,a41104a,a41108a,a41109a,a41110a,a41114a,a41115a,a41119a,a41120a,a41121a,a41125a,a41126a,a41130a,a41131a,a41132a,a41136a,a41137a,a41141a,a41142a,a41143a,a41147a,a41148a,a41152a,a41153a,a41154a,a41158a,a41159a,a41163a,a41164a,a41165a,a41169a,a41170a,a41174a,a41175a,a41176a,a41180a,a41181a,a41185a,a41186a,a41187a,a41191a,a41192a,a41196a,a41197a,a41198a,a41202a,a41203a,a41207a,a41208a,a41209a,a41213a,a41214a,a41218a,a41219a,a41220a,a41224a,a41225a,a41229a,a41230a,a41231a,a41235a,a41236a,a41240a,a41241a,a41242a,a41246a,a41247a,a41251a,a41252a,a41253a,a41257a,a41258a,a41262a,a41263a,a41264a,a41268a,a41269a,a41273a,a41274a,a41275a,a41279a,a41280a,a41284a,a41285a,a41286a,a41290a,a41291a,a41295a,a41296a,a41297a,a41301a,a41302a,a41306a,a41307a,a41308a,a41312a,a41313a,a41317a,a41318a,a41319a,a41323a,a41324a,a41328a,a41329a,a41330a,a41334a,a41335a,a41339a,a41340a,a41341a,a41345a,a41346a,a41350a,a41351a,a41352a,a41356a,a41357a,a41361a,a41362a,a41363a,a41367a,a41368a,a41372a,a41373a,a41374a,a41378a,a41379a,a41383a,a41384a,a41385a,a41389a,a41390a,a41394a,a41395a,a41396a,a41400a,a41401a,a41405a,a41406a,a41407a,a41411a,a41412a,a41416a,a41417a,a41418a,a41422a,a41423a,a41427a,a41428a,a41429a,a41433a,a41434a,a41438a,a41439a,a41440a,a41444a,a41445a,a41449a,a41450a,a41451a,a41455a,a41456a,a41460a,a41461a,a41462a,a41466a,a41467a,a41471a,a41472a,a41473a,a41477a,a41478a,a41482a,a41483a,a41484a,a41488a,a41489a,a41493a,a41494a,a41495a,a41499a,a41500a,a41504a,a41505a,a41506a,a41510a,a41511a,a41515a,a41516a,a41517a,a41521a,a41522a,a41526a,a41527a,a41528a,a41532a,a41533a,a41537a,a41538a,a41539a,a41543a,a41544a,a41548a,a41549a,a41550a,a41554a,a41555a,a41559a,a41560a,a41561a,a41565a,a41566a,a41570a,a41571a,a41572a,a41576a,a41577a,a41581a,a41582a,a41583a,a41587a,a41588a,a41592a,a41593a,a41594a,a41598a,a41599a,a41603a,a41604a,a41605a,a41609a,a41610a,a41614a,a41615a,a41616a,a41620a,a41621a,a41625a,a41626a,a41627a,a41631a,a41632a,a41636a,a41637a,a41638a,a41642a,a41643a,a41647a,a41648a,a41649a,a41653a,a41654a,a41658a,a41659a,a41660a,a41664a,a41665a,a41669a,a41670a,a41671a,a41675a,a41676a,a41680a,a41681a,a41682a,a41686a,a41687a,a41691a,a41692a,a41693a,a41697a,a41698a,a41702a,a41703a,a41704a,a41708a,a41709a,a41713a,a41714a,a41715a,a41719a,a41720a,a41724a,a41725a,a41726a,a41730a,a41731a,a41735a,a41736a,a41737a,a41741a,a41742a,a41746a,a41747a,a41748a,a41752a,a41753a,a41757a,a41758a,a41759a,a41763a,a41764a,a41768a,a41769a,a41770a,a41774a,a41775a,a41779a,a41780a,a41781a,a41785a,a41786a,a41790a,a41791a,a41792a,a41796a,a41797a,a41801a,a41802a,a41803a,a41807a,a41808a,a41812a,a41813a,a41814a,a41818a,a41819a,a41823a,a41824a,a41825a,a41829a,a41830a,a41834a,a41835a,a41836a,a41840a,a41841a,a41845a,a41846a,a41847a,a41851a,a41852a,a41856a,a41857a,a41858a,a41862a,a41863a,a41867a,a41868a,a41869a,a41873a,a41874a,a41878a,a41879a,a41880a,a41884a,a41885a,a41889a,a41890a,a41891a,a41895a,a41896a,a41900a,a41901a,a41902a,a41906a,a41907a,a41911a,a41912a,a41913a,a41917a,a41918a,a41922a,a41923a,a41924a,a41928a,a41929a,a41933a,a41934a,a41935a,a41939a,a41940a,a41944a,a41945a,a41946a,a41950a,a41951a,a41955a,a41956a,a41957a,a41961a,a41962a,a41966a,a41967a,a41968a,a41972a,a41973a,a41977a,a41978a,a41979a,a41983a,a41984a,a41988a,a41989a,a41990a,a41994a,a41995a,a41999a,a42000a,a42001a,a42005a,a42006a,a42010a,a42011a,a42012a,a42016a,a42017a,a42021a,a42022a,a42023a,a42027a,a42028a,a42032a,a42033a,a42034a,a42038a,a42039a,a42043a,a42044a,a42045a,a42049a,a42050a,a42054a,a42055a,a42056a,a42060a,a42061a,a42065a,a42066a,a42067a,a42071a,a42072a,a42076a,a42077a,a42078a,a42082a,a42083a,a42087a,a42088a,a42089a,a42093a,a42094a,a42098a,a42099a,a42100a,a42104a,a42105a,a42109a,a42110a,a42111a,a42115a,a42116a,a42120a,a42121a,a42122a,a42126a,a42127a,a42131a,a42132a,a42133a,a42137a,a42138a,a42142a,a42143a,a42144a,a42148a,a42149a,a42153a,a42154a,a42155a,a42159a,a42160a,a42164a,a42165a,a42166a,a42170a,a42171a,a42175a,a42176a,a42177a,a42181a,a42182a,a42186a,a42187a,a42188a,a42192a,a42193a,a42197a,a42198a,a42199a,a42203a,a42204a,a42208a,a42209a,a42210a,a42214a,a42215a,a42219a,a42220a,a42221a,a42225a,a42226a,a42230a,a42231a,a42232a,a42236a,a42237a,a42241a,a42242a,a42243a,a42247a,a42248a,a42252a,a42253a,a42254a,a42258a,a42259a,a42263a,a42264a,a42265a,a42269a,a42270a,a42274a,a42275a,a42276a,a42280a,a42281a,a42285a,a42286a,a42287a,a42291a,a42292a,a42296a,a42297a,a42298a,a42302a,a42303a,a42307a,a42308a,a42309a,a42313a,a42314a,a42318a,a42319a,a42320a,a42324a,a42325a,a42329a,a42330a,a42331a,a42335a,a42336a,a42340a,a42341a,a42342a,a42346a,a42347a,a42351a,a42352a,a42353a,a42357a,a42358a,a42362a,a42363a,a42364a,a42368a,a42369a,a42373a,a42374a,a42375a,a42379a,a42380a,a42384a,a42385a,a42386a,a42390a,a42391a,a42395a,a42396a,a42397a,a42401a,a42402a,a42406a,a42407a,a42408a,a42412a,a42413a,a42417a,a42418a,a42419a,a42423a,a42424a,a42428a,a42429a,a42430a,a42434a,a42435a,a42439a,a42440a,a42441a,a42445a,a42446a,a42450a,a42451a,a42452a,a42456a,a42457a,a42461a,a42462a,a42463a,a42467a,a42468a,a42472a,a42473a,a42474a,a42478a,a42479a,a42483a,a42484a,a42485a,a42489a,a42490a,a42494a,a42495a,a42496a,a42500a,a42501a,a42505a,a42506a,a42507a,a42511a,a42512a,a42516a,a42517a,a42518a,a42522a,a42523a,a42527a,a42528a,a42529a,a42533a,a42534a,a42538a,a42539a,a42540a,a42544a,a42545a,a42549a,a42550a,a42551a,a42555a,a42556a,a42560a,a42561a,a42562a,a42566a,a42567a,a42571a,a42572a,a42573a,a42577a,a42578a,a42582a,a42583a,a42584a,a42588a,a42589a,a42593a,a42594a,a42595a,a42599a,a42600a,a42604a,a42605a,a42606a,a42610a,a42611a,a42615a,a42616a,a42617a,a42621a,a42622a,a42626a,a42627a,a42628a,a42632a,a42633a,a42637a,a42638a,a42639a,a42643a,a42644a,a42648a,a42649a,a42650a,a42654a,a42655a,a42659a,a42660a,a42661a,a42665a,a42666a,a42670a,a42671a,a42672a,a42676a,a42677a,a42681a,a42682a,a42683a,a42687a,a42688a,a42692a,a42693a,a42694a,a42698a,a42699a,a42703a,a42704a,a42705a,a42709a,a42710a,a42714a,a42715a,a42716a,a42720a,a42721a,a42725a,a42726a,a42727a,a42731a,a42732a,a42736a,a42737a,a42738a,a42742a,a42743a,a42747a,a42748a,a42749a,a42753a,a42754a,a42758a,a42759a,a42760a,a42764a,a42765a,a42769a,a42770a,a42771a,a42775a,a42776a,a42780a,a42781a,a42782a,a42786a,a42787a,a42791a,a42792a,a42793a,a42797a,a42798a,a42802a,a42803a,a42804a,a42808a,a42809a,a42813a,a42814a,a42815a,a42819a,a42820a,a42824a,a42825a,a42826a,a42830a,a42831a,a42835a,a42836a,a42837a,a42841a,a42842a,a42846a,a42847a,a42848a,a42852a,a42853a,a42857a,a42858a,a42859a,a42863a,a42864a,a42868a,a42869a,a42870a,a42874a,a42875a,a42879a,a42880a,a42881a,a42885a,a42886a,a42890a,a42891a,a42892a,a42896a,a42897a,a42901a,a42902a,a42903a,a42907a,a42908a,a42912a,a42913a,a42914a,a42918a,a42919a,a42923a,a42924a,a42925a,a42929a,a42930a,a42934a,a42935a,a42936a,a42940a,a42941a,a42945a,a42946a,a42947a,a42951a,a42952a,a42956a,a42957a,a42958a,a42962a,a42963a,a42967a,a42968a,a42969a,a42973a,a42974a,a42978a,a42979a,a42980a,a42984a,a42985a,a42989a,a42990a,a42991a,a42995a,a42996a,a43000a,a43001a,a43002a,a43006a,a43007a,a43011a,a43012a,a43013a,a43017a,a43018a,a43022a,a43023a,a43024a,a43028a,a43029a,a43033a,a43034a,a43035a,a43039a,a43040a,a43044a,a43045a,a43046a,a43050a,a43051a,a43055a,a43056a,a43057a,a43061a,a43062a,a43066a,a43067a,a43068a,a43072a,a43073a,a43077a,a43078a,a43079a,a43083a,a43084a,a43088a,a43089a,a43090a,a43094a,a43095a,a43099a,a43100a,a43101a,a43105a,a43106a,a43110a,a43111a,a43112a,a43116a,a43117a,a43121a,a43122a,a43123a,a43127a,a43128a,a43132a,a43133a,a43134a,a43138a,a43139a,a43143a,a43144a,a43145a,a43149a,a43150a,a43154a,a43155a,a43156a,a43160a,a43161a,a43165a,a43166a,a43167a,a43171a,a43172a,a43176a,a43177a,a43178a,a43182a,a43183a,a43187a,a43188a,a43189a,a43193a,a43194a,a43198a,a43199a,a43200a,a43204a,a43205a,a43209a,a43210a,a43211a,a43215a,a43216a,a43220a,a43221a,a43222a,a43226a,a43227a,a43231a,a43232a,a43233a,a43237a,a43238a,a43242a,a43243a,a43244a,a43248a,a43249a,a43253a,a43254a,a43255a,a43259a,a43260a,a43264a,a43265a,a43266a,a43270a,a43271a,a43275a,a43276a,a43277a,a43281a,a43282a,a43286a,a43287a,a43288a,a43292a,a43293a,a43297a,a43298a,a43299a,a43303a,a43304a,a43308a,a43309a,a43310a,a43314a,a43315a,a43319a,a43320a,a43321a,a43325a,a43326a,a43330a,a43331a,a43332a,a43336a,a43337a,a43341a,a43342a,a43343a,a43347a,a43348a,a43352a,a43353a,a43354a,a43358a,a43359a,a43363a,a43364a,a43365a,a43369a,a43370a,a43374a,a43375a,a43376a,a43380a,a43381a,a43385a,a43386a,a43387a,a43391a,a43392a,a43396a,a43397a,a43398a,a43402a,a43403a,a43407a,a43408a,a43409a,a43413a,a43414a,a43418a,a43419a,a43420a,a43424a,a43425a,a43429a,a43430a,a43431a,a43435a,a43436a,a43440a,a43441a,a43442a,a43446a,a43447a,a43451a,a43452a,a43453a,a43457a,a43458a,a43462a,a43463a,a43464a,a43468a,a43469a,a43473a,a43474a,a43475a,a43479a,a43480a,a43484a,a43485a,a43486a,a43490a,a43491a,a43495a,a43496a,a43497a,a43501a,a43502a,a43506a,a43507a,a43508a,a43512a,a43513a,a43517a,a43518a,a43519a,a43523a,a43524a,a43528a,a43529a,a43530a,a43534a,a43535a,a43539a,a43540a,a43541a,a43545a,a43546a,a43550a,a43551a,a43552a,a43556a,a43557a,a43561a,a43562a,a43563a,a43567a,a43568a,a43572a,a43573a,a43574a,a43578a,a43579a,a43583a,a43584a,a43585a,a43589a,a43590a,a43594a,a43595a,a43596a,a43600a,a43601a,a43605a,a43606a,a43607a,a43611a,a43612a,a43616a,a43617a,a43618a,a43622a,a43623a,a43627a,a43628a,a43629a,a43633a,a43634a,a43638a,a43639a,a43640a,a43644a,a43645a,a43649a,a43650a,a43651a,a43655a,a43656a,a43660a,a43661a,a43662a,a43666a,a43667a,a43671a,a43672a,a43673a,a43677a,a43678a,a43682a,a43683a,a43684a,a43688a,a43689a,a43693a,a43694a,a43695a,a43699a,a43700a,a43704a,a43705a,a43706a,a43710a,a43711a,a43715a,a43716a,a43717a,a43721a,a43722a,a43726a,a43727a,a43728a,a43732a,a43733a,a43737a,a43738a,a43739a,a43743a,a43744a,a43748a,a43749a,a43750a,a43754a,a43755a,a43759a,a43760a,a43761a,a43765a,a43766a,a43770a,a43771a,a43772a,a43776a,a43777a,a43781a,a43782a,a43783a,a43787a,a43788a,a43792a,a43793a,a43794a,a43798a,a43799a,a43803a,a43804a,a43805a,a43809a,a43810a,a43814a,a43815a,a43816a,a43820a,a43821a,a43825a,a43826a,a43827a,a43831a,a43832a,a43836a,a43837a,a43838a,a43842a,a43843a,a43847a,a43848a,a43849a,a43853a,a43854a,a43858a,a43859a,a43860a,a43864a,a43865a,a43869a,a43870a,a43871a,a43875a,a43876a,a43880a,a43881a,a43882a,a43886a,a43887a,a43891a,a43892a,a43893a,a43897a,a43898a,a43902a,a43903a,a43904a,a43908a,a43909a,a43913a,a43914a,a43915a,a43919a,a43920a,a43924a,a43925a,a43926a,a43930a,a43931a,a43935a,a43936a,a43937a,a43941a,a43942a,a43946a,a43947a,a43948a,a43952a,a43953a,a43957a,a43958a,a43959a,a43963a,a43964a,a43968a,a43969a,a43970a,a43974a,a43975a,a43979a,a43980a,a43981a,a43985a,a43986a,a43990a,a43991a,a43992a,a43996a,a43997a,a44001a,a44002a,a44003a,a44007a,a44008a,a44012a,a44013a,a44014a,a44018a,a44019a,a44023a,a44024a,a44025a,a44029a,a44030a,a44034a,a44035a,a44036a,a44040a,a44041a,a44045a,a44046a,a44047a,a44051a,a44052a,a44056a,a44057a,a44058a,a44062a,a44063a,a44067a,a44068a,a44069a,a44073a,a44074a,a44078a,a44079a,a44080a,a44084a,a44085a,a44089a,a44090a,a44091a,a44095a,a44096a,a44100a,a44101a,a44102a,a44106a,a44107a,a44111a,a44112a,a44113a,a44117a,a44118a,a44122a,a44123a,a44124a,a44128a,a44129a,a44133a,a44134a,a44135a,a44139a,a44140a,a44144a,a44145a,a44146a,a44150a,a44151a,a44155a,a44156a,a44157a,a44161a,a44162a,a44166a,a44167a,a44168a,a44172a,a44173a,a44177a,a44178a,a44179a,a44183a,a44184a,a44188a,a44189a,a44190a,a44194a,a44195a,a44199a,a44200a,a44201a,a44205a,a44206a,a44210a,a44211a,a44212a,a44216a,a44217a,a44221a,a44222a,a44223a,a44227a,a44228a,a44232a,a44233a,a44234a,a44238a,a44239a,a44243a,a44244a,a44245a,a44249a,a44250a,a44254a,a44255a,a44256a,a44260a,a44261a,a44265a,a44266a,a44267a,a44271a,a44272a,a44276a,a44277a,a44278a,a44282a,a44283a,a44287a,a44288a,a44289a,a44293a,a44294a,a44298a,a44299a,a44300a,a44304a,a44305a,a44309a,a44310a,a44311a,a44315a,a44316a,a44320a,a44321a,a44322a,a44326a,a44327a,a44331a,a44332a,a44333a,a44337a,a44338a,a44342a,a44343a,a44344a,a44348a,a44349a,a44353a,a44354a,a44355a,a44359a,a44360a,a44364a,a44365a,a44366a,a44370a,a44371a,a44375a,a44376a,a44377a,a44381a,a44382a,a44386a,a44387a,a44388a,a44392a,a44393a,a44397a,a44398a,a44399a,a44403a,a44404a,a44408a,a44409a,a44410a,a44414a,a44415a,a44419a,a44420a,a44421a,a44425a,a44426a,a44430a,a44431a,a44432a,a44436a,a44437a,a44441a,a44442a,a44443a,a44447a,a44448a,a44452a,a44453a,a44454a,a44458a,a44459a,a44463a,a44464a,a44465a,a44469a,a44470a,a44474a,a44475a,a44476a,a44480a,a44481a,a44485a,a44486a,a44487a,a44491a,a44492a,a44496a,a44497a,a44498a,a44502a,a44503a,a44507a,a44508a,a44509a,a44513a,a44514a,a44518a,a44519a,a44520a,a44524a,a44525a,a44529a,a44530a,a44531a,a44535a,a44536a,a44540a,a44541a,a44542a,a44546a,a44547a,a44551a,a44552a,a44553a,a44557a,a44558a,a44562a,a44563a,a44564a,a44568a,a44569a,a44573a,a44574a,a44575a,a44579a,a44580a,a44583a,a44586a,a44587a,a44588a,a44592a,a44593a,a44597a,a44598a,a44599a,a44603a,a44604a,a44607a,a44610a,a44611a,a44612a,a44616a,a44617a,a44621a,a44622a,a44623a,a44627a,a44628a,a44631a,a44634a,a44635a,a44636a,a44640a,a44641a,a44645a,a44646a,a44647a,a44651a,a44652a,a44655a,a44658a,a44659a,a44660a,a44664a,a44665a,a44669a,a44670a,a44671a,a44675a,a44676a,a44679a,a44682a,a44683a,a44684a,a44688a,a44689a,a44693a,a44694a,a44695a,a44699a,a44700a,a44703a,a44706a,a44707a,a44708a,a44712a,a44713a,a44717a,a44718a,a44719a,a44723a,a44724a,a44727a,a44730a,a44731a,a44732a,a44736a,a44737a,a44741a,a44742a,a44743a,a44747a,a44748a,a44751a,a44754a,a44755a,a44756a,a44760a,a44761a,a44765a,a44766a,a44767a,a44771a,a44772a,a44775a,a44778a,a44779a,a44780a,a44784a,a44785a,a44789a,a44790a,a44791a,a44795a,a44796a,a44799a,a44802a,a44803a,a44804a,a44808a,a44809a,a44813a,a44814a,a44815a,a44819a,a44820a,a44823a,a44826a,a44827a,a44828a,a44832a,a44833a,a44837a,a44838a,a44839a,a44843a,a44844a,a44847a,a44850a,a44851a,a44852a,a44856a,a44857a,a44861a,a44862a,a44863a,a44867a,a44868a,a44871a,a44874a,a44875a,a44876a,a44880a,a44881a,a44885a,a44886a,a44887a,a44891a,a44892a,a44895a,a44898a,a44899a,a44900a,a44904a,a44905a,a44909a,a44910a,a44911a,a44915a,a44916a,a44919a,a44922a,a44923a,a44924a,a44928a,a44929a,a44933a,a44934a,a44935a,a44939a,a44940a,a44943a,a44946a,a44947a,a44948a,a44952a,a44953a,a44957a,a44958a,a44959a,a44963a,a44964a,a44967a,a44970a,a44971a,a44972a,a44976a,a44977a,a44981a,a44982a,a44983a,a44987a,a44988a,a44991a,a44994a,a44995a,a44996a,a45000a,a45001a,a45005a,a45006a,a45007a,a45011a,a45012a,a45015a,a45018a,a45019a,a45020a,a45024a,a45025a,a45029a,a45030a,a45031a,a45035a,a45036a,a45039a,a45042a,a45043a,a45044a,a45048a,a45049a,a45053a,a45054a,a45055a,a45059a,a45060a,a45063a,a45066a,a45067a,a45068a,a45072a,a45073a,a45077a,a45078a,a45079a,a45083a,a45084a,a45087a,a45090a,a45091a,a45092a,a45096a,a45097a,a45101a,a45102a,a45103a,a45107a,a45108a,a45111a,a45114a,a45115a,a45116a,a45120a,a45121a,a45125a,a45126a,a45127a,a45131a,a45132a,a45135a,a45138a,a45139a,a45140a,a45144a,a45145a,a45149a,a45150a,a45151a,a45155a,a45156a,a45159a,a45162a,a45163a,a45164a,a45168a,a45169a,a45173a,a45174a,a45175a,a45179a,a45180a,a45183a,a45186a,a45187a,a45188a,a45192a,a45193a,a45197a,a45198a,a45199a,a45203a,a45204a,a45207a,a45210a,a45211a,a45212a,a45216a,a45217a,a45221a,a45222a,a45223a,a45227a,a45228a,a45231a,a45234a,a45235a,a45236a,a45240a,a45241a,a45245a,a45246a,a45247a,a45251a,a45252a,a45255a,a45258a,a45259a,a45260a,a45264a,a45265a,a45269a,a45270a,a45271a,a45275a,a45276a,a45279a,a45282a,a45283a,a45284a,a45288a,a45289a,a45293a,a45294a,a45295a,a45299a,a45300a,a45303a,a45306a,a45307a,a45308a,a45312a,a45313a,a45317a,a45318a,a45319a,a45323a,a45324a,a45327a,a45330a,a45331a,a45332a,a45336a,a45337a,a45341a,a45342a,a45343a,a45347a,a45348a,a45351a,a45354a,a45355a,a45356a,a45360a,a45361a,a45365a,a45366a,a45367a,a45371a,a45372a,a45375a,a45378a,a45379a,a45380a,a45384a,a45385a,a45389a,a45390a,a45391a,a45395a,a45396a,a45399a,a45402a,a45403a,a45404a,a45408a,a45409a,a45413a,a45414a,a45415a,a45419a,a45420a,a45423a,a45426a,a45427a,a45428a,a45432a,a45433a,a45437a,a45438a,a45439a,a45443a,a45444a,a45447a,a45450a,a45451a,a45452a,a45456a,a45457a,a45461a,a45462a,a45463a,a45467a,a45468a,a45471a,a45474a,a45475a,a45476a,a45480a,a45481a,a45485a,a45486a,a45487a,a45491a,a45492a,a45495a,a45498a,a45499a,a45500a,a45504a,a45505a,a45509a,a45510a,a45511a,a45515a,a45516a,a45519a,a45522a,a45523a,a45524a,a45528a,a45529a,a45533a,a45534a,a45535a,a45539a,a45540a,a45543a,a45546a,a45547a,a45548a,a45552a,a45553a,a45557a,a45558a,a45559a,a45563a,a45564a,a45567a,a45570a,a45571a,a45572a,a45576a,a45577a,a45581a,a45582a,a45583a,a45587a,a45588a,a45591a,a45594a,a45595a,a45596a,a45600a,a45601a,a45605a,a45606a,a45607a,a45611a,a45612a,a45615a,a45618a,a45619a,a45620a,a45624a,a45625a,a45629a,a45630a,a45631a,a45635a,a45636a,a45639a,a45642a,a45643a,a45644a,a45648a,a45649a,a45653a,a45654a,a45655a,a45659a,a45660a,a45663a,a45666a,a45667a,a45668a,a45672a,a45673a,a45677a,a45678a,a45679a,a45683a,a45684a,a45687a,a45690a,a45691a,a45692a,a45696a,a45697a,a45701a,a45702a,a45703a,a45707a,a45708a,a45711a,a45714a,a45715a,a45716a,a45720a,a45721a,a45725a,a45726a,a45727a,a45731a,a45732a,a45735a,a45738a,a45739a,a45740a,a45744a,a45745a,a45749a,a45750a,a45751a,a45755a,a45756a,a45759a,a45762a,a45763a,a45764a,a45768a,a45769a,a45773a,a45774a,a45775a,a45779a,a45780a,a45783a,a45786a,a45787a,a45788a,a45792a,a45793a,a45797a,a45798a,a45799a,a45803a,a45804a,a45807a,a45810a,a45811a,a45812a,a45816a,a45817a,a45821a,a45822a,a45823a,a45827a,a45828a,a45831a,a45834a,a45835a,a45836a,a45840a,a45841a,a45845a,a45846a,a45847a,a45851a,a45852a,a45855a,a45858a,a45859a,a45860a,a45864a,a45865a,a45869a,a45870a,a45871a,a45875a,a45876a,a45879a,a45882a,a45883a,a45884a,a45888a,a45889a,a45893a,a45894a,a45895a,a45899a,a45900a,a45903a,a45906a,a45907a,a45908a,a45912a,a45913a,a45917a,a45918a,a45919a,a45923a,a45924a,a45927a,a45930a,a45931a,a45932a,a45936a,a45937a,a45941a,a45942a,a45943a,a45947a,a45948a,a45951a,a45954a,a45955a,a45956a,a45960a,a45961a,a45965a,a45966a,a45967a,a45971a,a45972a,a45975a,a45978a,a45979a,a45980a,a45984a,a45985a,a45989a,a45990a,a45991a,a45995a,a45996a,a45999a,a46002a,a46003a,a46004a,a46008a,a46009a,a46013a,a46014a,a46015a,a46019a,a46020a,a46023a,a46026a,a46027a,a46028a,a46032a,a46033a,a46037a,a46038a,a46039a,a46043a,a46044a,a46047a,a46050a,a46051a,a46052a,a46056a,a46057a,a46061a,a46062a,a46063a,a46067a,a46068a,a46071a,a46074a,a46075a,a46076a,a46080a,a46081a,a46085a,a46086a,a46087a,a46091a,a46092a,a46095a,a46098a,a46099a,a46100a,a46104a,a46105a,a46109a,a46110a,a46111a,a46115a,a46116a,a46119a,a46122a,a46123a,a46124a,a46128a,a46129a,a46133a,a46134a,a46135a,a46139a,a46140a,a46143a,a46146a,a46147a,a46148a,a46152a,a46153a,a46157a,a46158a,a46159a,a46163a,a46164a,a46167a,a46170a,a46171a,a46172a,a46176a,a46177a,a46181a,a46182a,a46183a,a46187a,a46188a,a46191a,a46194a,a46195a,a46196a,a46200a,a46201a,a46205a,a46206a,a46207a,a46211a,a46212a,a46215a,a46218a,a46219a,a46220a,a46224a,a46225a,a46229a,a46230a,a46231a,a46235a,a46236a,a46239a,a46242a,a46243a,a46244a,a46248a,a46249a,a46253a,a46254a,a46255a,a46259a,a46260a,a46263a,a46266a,a46267a,a46268a,a46272a,a46273a,a46277a,a46278a,a46279a,a46283a,a46284a,a46287a,a46290a,a46291a,a46292a,a46296a,a46297a,a46301a,a46302a,a46303a,a46307a,a46308a,a46311a,a46314a,a46315a,a46316a,a46320a,a46321a,a46325a,a46326a,a46327a,a46331a,a46332a,a46335a,a46338a,a46339a,a46340a,a46344a,a46345a,a46349a,a46350a,a46351a,a46355a,a46356a,a46359a,a46362a,a46363a,a46364a,a46368a,a46369a,a46373a,a46374a,a46375a,a46379a,a46380a,a46383a,a46386a,a46387a,a46388a,a46392a,a46393a,a46397a,a46398a,a46399a,a46403a,a46404a,a46407a,a46410a,a46411a,a46412a,a46416a,a46417a,a46421a,a46422a,a46423a,a46427a,a46428a,a46431a,a46434a,a46435a,a46436a,a46440a,a46441a,a46445a,a46446a,a46447a,a46451a,a46452a,a46455a,a46458a,a46459a,a46460a,a46464a,a46465a,a46469a,a46470a,a46471a,a46475a,a46476a,a46479a,a46482a,a46483a,a46484a,a46488a,a46489a,a46493a,a46494a,a46495a,a46499a,a46500a,a46503a,a46506a,a46507a,a46508a,a46512a,a46513a,a46517a,a46518a,a46519a,a46523a,a46524a,a46527a,a46530a,a46531a,a46532a,a46536a,a46537a,a46541a,a46542a,a46543a,a46547a,a46548a,a46551a,a46554a,a46555a,a46556a,a46560a,a46561a,a46565a,a46566a,a46567a,a46571a,a46572a,a46575a,a46578a,a46579a,a46580a,a46584a,a46585a,a46589a,a46590a,a46591a,a46595a,a46596a,a46599a,a46602a,a46603a,a46604a,a46608a,a46609a,a46613a,a46614a,a46615a,a46619a,a46620a,a46623a,a46626a,a46627a,a46628a,a46632a,a46633a,a46637a,a46638a,a46639a,a46643a,a46644a,a46647a,a46650a,a46651a,a46652a,a46656a,a46657a,a46661a,a46662a,a46663a,a46667a,a46668a,a46671a,a46674a,a46675a,a46676a,a46680a,a46681a,a46685a,a46686a,a46687a,a46691a,a46692a,a46695a,a46698a,a46699a,a46700a,a46704a,a46705a,a46709a,a46710a,a46711a,a46715a,a46716a,a46719a,a46722a,a46723a,a46724a,a46728a,a46729a,a46733a,a46734a,a46735a,a46739a,a46740a,a46743a,a46746a,a46747a,a46748a,a46752a,a46753a,a46757a,a46758a,a46759a,a46763a,a46764a,a46767a,a46770a,a46771a,a46772a,a46776a,a46777a,a46781a,a46782a,a46783a,a46787a,a46788a,a46791a,a46794a,a46795a,a46796a,a46800a,a46801a,a46805a,a46806a,a46807a,a46811a,a46812a,a46815a,a46818a,a46819a,a46820a,a46824a,a46825a,a46829a,a46830a,a46831a,a46835a,a46836a,a46839a,a46842a,a46843a,a46844a,a46848a,a46849a,a46853a,a46854a,a46855a,a46859a,a46860a,a46863a,a46866a,a46867a,a46868a,a46872a,a46873a,a46877a,a46878a,a46879a,a46883a,a46884a,a46887a,a46890a,a46891a,a46892a,a46896a,a46897a,a46901a,a46902a,a46903a,a46907a,a46908a,a46911a,a46914a,a46915a,a46916a,a46920a,a46921a,a46925a,a46926a,a46927a,a46931a,a46932a,a46935a,a46938a,a46939a,a46940a,a46944a,a46945a,a46949a,a46950a,a46951a,a46955a,a46956a,a46959a,a46962a,a46963a,a46964a,a46968a,a46969a,a46973a,a46974a,a46975a,a46979a,a46980a,a46983a,a46986a,a46987a,a46988a,a46992a,a46993a,a46997a,a46998a,a46999a,a47003a,a47004a,a47007a,a47010a,a47011a,a47012a,a47016a,a47017a,a47021a,a47022a,a47023a,a47027a,a47028a,a47031a,a47034a,a47035a,a47036a,a47040a,a47041a,a47045a,a47046a,a47047a,a47051a,a47052a,a47055a,a47058a,a47059a,a47060a,a47064a,a47065a,a47069a,a47070a,a47071a,a47075a,a47076a,a47079a,a47082a,a47083a,a47084a,a47088a,a47089a,a47093a,a47094a,a47095a,a47099a,a47100a,a47103a,a47106a,a47107a,a47108a,a47112a,a47113a,a47117a,a47118a,a47119a,a47123a,a47124a,a47127a,a47130a,a47131a,a47132a,a47136a,a47137a,a47141a,a47142a,a47143a,a47147a,a47148a,a47151a,a47154a,a47155a,a47156a,a47160a,a47161a,a47165a,a47166a,a47167a,a47171a,a47172a,a47175a,a47178a,a47179a,a47180a,a47184a,a47185a,a47189a,a47190a,a47191a,a47195a,a47196a,a47199a,a47202a,a47203a,a47204a,a47208a,a47209a,a47213a,a47214a,a47215a,a47219a,a47220a,a47223a,a47226a,a47227a,a47228a,a47232a,a47233a,a47237a,a47238a,a47239a,a47243a,a47244a,a47247a,a47250a,a47251a,a47252a,a47256a,a47257a,a47261a,a47262a,a47263a,a47267a,a47268a,a47271a,a47274a,a47275a,a47276a,a47280a,a47281a,a47285a,a47286a,a47287a,a47291a,a47292a,a47295a,a47298a,a47299a,a47300a,a47304a,a47305a,a47309a,a47310a,a47311a,a47315a,a47316a,a47319a,a47322a,a47323a,a47324a,a47328a,a47329a,a47333a,a47334a,a47335a,a47339a,a47340a,a47343a,a47346a,a47347a,a47348a,a47352a,a47353a,a47357a,a47358a,a47359a,a47363a,a47364a,a47367a,a47370a,a47371a,a47372a,a47376a,a47377a,a47381a,a47382a,a47383a,a47387a,a47388a,a47391a,a47394a,a47395a,a47396a,a47400a,a47401a,a47405a,a47406a,a47407a,a47411a,a47412a,a47415a,a47418a,a47419a,a47420a,a47424a,a47425a,a47429a,a47430a,a47431a,a47435a,a47436a,a47439a,a47442a,a47443a,a47444a,a47448a,a47449a,a47453a,a47454a,a47455a,a47459a,a47460a,a47463a,a47466a,a47467a,a47468a,a47472a,a47473a,a47477a,a47478a,a47479a,a47483a,a47484a,a47487a,a47490a,a47491a,a47492a,a47496a,a47497a,a47501a,a47502a,a47503a,a47507a,a47508a,a47511a,a47514a,a47515a,a47516a,a47520a,a47521a,a47525a,a47526a,a47527a,a47531a,a47532a,a47535a,a47538a,a47539a,a47540a,a47544a,a47545a,a47549a,a47550a,a47551a,a47555a,a47556a,a47559a,a47562a,a47563a,a47564a,a47568a,a47569a,a47573a,a47574a,a47575a,a47579a,a47580a,a47583a,a47586a,a47587a,a47588a,a47592a,a47593a,a47597a,a47598a,a47599a,a47603a,a47604a,a47607a,a47610a,a47611a,a47612a,a47616a,a47617a,a47621a,a47622a,a47623a,a47627a,a47628a,a47631a,a47634a,a47635a,a47636a,a47640a,a47641a,a47645a,a47646a,a47647a,a47651a,a47652a,a47655a,a47658a,a47659a,a47660a,a47664a,a47665a,a47669a,a47670a,a47671a,a47675a,a47676a,a47679a,a47682a,a47683a,a47684a,a47688a,a47689a,a47693a,a47694a,a47695a,a47699a,a47700a,a47703a,a47706a,a47707a,a47708a,a47712a,a47713a,a47717a,a47718a,a47719a,a47723a,a47724a,a47727a,a47730a,a47731a,a47732a,a47736a,a47737a,a47741a,a47742a,a47743a,a47747a,a47748a,a47751a,a47754a,a47755a,a47756a,a47760a,a47761a,a47765a,a47766a,a47767a,a47771a,a47772a,a47775a,a47778a,a47779a,a47780a,a47784a,a47785a,a47789a,a47790a,a47791a,a47795a,a47796a,a47799a,a47802a,a47803a,a47804a,a47808a,a47809a,a47813a,a47814a,a47815a,a47819a,a47820a,a47823a,a47826a,a47827a,a47828a,a47832a,a47833a,a47837a,a47838a,a47839a,a47843a,a47844a,a47847a,a47850a,a47851a,a47852a,a47856a,a47857a,a47861a,a47862a,a47863a,a47867a,a47868a,a47871a,a47874a,a47875a,a47876a,a47880a,a47881a,a47885a,a47886a,a47887a,a47891a,a47892a,a47895a,a47898a,a47899a,a47900a,a47904a,a47905a,a47909a,a47910a,a47911a,a47915a,a47916a,a47919a,a47922a,a47923a,a47924a,a47928a,a47929a,a47933a,a47934a,a47935a,a47939a,a47940a,a47943a,a47946a,a47947a,a47948a,a47952a,a47953a,a47957a,a47958a,a47959a,a47963a,a47964a,a47967a,a47970a,a47971a,a47972a,a47976a,a47977a,a47981a,a47982a,a47983a,a47987a,a47988a,a47991a,a47994a,a47995a,a47996a,a48000a,a48001a,a48005a,a48006a,a48007a,a48011a,a48012a,a48015a,a48018a,a48019a,a48020a,a48024a,a48025a,a48029a,a48030a,a48031a,a48035a,a48036a,a48039a,a48042a,a48043a,a48044a,a48048a,a48049a,a48053a,a48054a,a48055a,a48059a,a48060a,a48063a,a48066a,a48067a,a48068a,a48072a,a48073a,a48077a,a48078a,a48079a,a48083a,a48084a,a48087a,a48090a,a48091a,a48092a,a48096a,a48097a,a48101a,a48102a,a48103a,a48107a,a48108a,a48111a,a48114a,a48115a,a48116a,a48120a,a48121a,a48125a,a48126a,a48127a,a48131a,a48132a,a48135a,a48138a,a48139a,a48140a,a48144a,a48145a,a48149a,a48150a,a48151a,a48155a,a48156a,a48159a,a48162a,a48163a,a48164a,a48168a,a48169a,a48173a,a48174a,a48175a,a48179a,a48180a,a48183a,a48186a,a48187a,a48188a,a48192a,a48193a,a48197a,a48198a,a48199a,a48203a,a48204a,a48207a,a48210a,a48211a,a48212a,a48216a,a48217a,a48221a,a48222a,a48223a,a48227a,a48228a,a48231a,a48234a,a48235a,a48236a,a48240a,a48241a,a48245a,a48246a,a48247a,a48251a,a48252a,a48255a,a48258a,a48259a,a48260a,a48264a,a48265a,a48269a,a48270a,a48271a,a48275a,a48276a,a48279a,a48282a,a48283a,a48284a,a48288a,a48289a,a48293a,a48294a,a48295a,a48299a,a48300a,a48303a,a48306a,a48307a,a48308a,a48312a,a48313a,a48317a,a48318a,a48319a,a48323a,a48324a,a48327a,a48330a,a48331a,a48332a,a48336a,a48337a,a48341a,a48342a,a48343a,a48347a,a48348a,a48351a,a48354a,a48355a,a48356a,a48360a,a48361a,a48365a,a48366a,a48367a,a48371a,a48372a,a48375a,a48378a,a48379a,a48380a,a48384a,a48385a,a48389a,a48390a,a48391a,a48395a,a48396a,a48399a,a48402a,a48403a,a48404a,a48408a,a48409a,a48413a,a48414a,a48415a,a48419a,a48420a,a48423a,a48426a,a48427a,a48428a,a48432a,a48433a,a48437a,a48438a,a48439a,a48443a,a48444a,a48447a,a48450a,a48451a,a48452a,a48456a,a48457a,a48461a,a48462a,a48463a,a48467a,a48468a,a48471a,a48474a,a48475a,a48476a,a48480a,a48481a,a48485a,a48486a,a48487a,a48491a,a48492a,a48495a,a48498a,a48499a,a48500a,a48504a,a48505a,a48509a,a48510a,a48511a,a48515a,a48516a,a48519a,a48522a,a48523a,a48524a,a48528a,a48529a,a48533a,a48534a,a48535a,a48539a,a48540a,a48543a,a48546a,a48547a,a48548a,a48552a,a48553a,a48557a,a48558a,a48559a,a48563a,a48564a,a48567a,a48570a,a48571a,a48572a,a48576a,a48577a,a48581a,a48582a,a48583a,a48587a,a48588a,a48591a,a48594a,a48595a,a48596a,a48600a,a48601a,a48605a,a48606a,a48607a,a48611a,a48612a,a48615a,a48618a,a48619a,a48620a,a48624a,a48625a,a48629a,a48630a,a48631a,a48635a,a48636a,a48639a,a48642a,a48643a,a48644a,a48648a,a48649a,a48653a,a48654a,a48655a,a48659a,a48660a,a48663a,a48666a,a48667a,a48668a,a48672a,a48673a,a48677a,a48678a,a48679a,a48683a,a48684a,a48687a,a48690a,a48691a,a48692a,a48696a,a48697a,a48701a,a48702a,a48703a,a48707a,a48708a,a48711a,a48714a,a48715a,a48716a,a48720a,a48721a,a48725a,a48726a,a48727a,a48731a,a48732a,a48735a,a48738a,a48739a,a48740a,a48744a,a48745a,a48749a,a48750a,a48751a,a48755a,a48756a,a48759a,a48762a,a48763a,a48764a,a48768a,a48769a,a48773a,a48774a,a48775a,a48779a,a48780a,a48783a,a48786a,a48787a,a48788a,a48792a,a48793a,a48797a,a48798a,a48799a,a48803a,a48804a,a48807a,a48810a,a48811a,a48812a,a48816a,a48817a,a48821a,a48822a,a48823a,a48827a,a48828a,a48831a,a48834a,a48835a,a48836a,a48840a,a48841a,a48845a,a48846a,a48847a,a48851a,a48852a,a48855a,a48858a,a48859a,a48860a,a48864a,a48865a,a48869a,a48870a,a48871a,a48875a,a48876a,a48879a,a48882a,a48883a,a48884a,a48888a,a48889a,a48893a,a48894a,a48895a,a48899a,a48900a,a48903a,a48906a,a48907a,a48908a,a48912a,a48913a,a48917a,a48918a,a48919a,a48923a,a48924a,a48927a,a48930a,a48931a,a48932a,a48936a,a48937a,a48941a,a48942a,a48943a,a48947a,a48948a,a48951a,a48954a,a48955a,a48956a,a48960a,a48961a,a48965a,a48966a,a48967a,a48971a,a48972a,a48975a,a48978a,a48979a,a48980a,a48984a,a48985a,a48989a,a48990a,a48991a,a48995a,a48996a,a48999a,a49002a,a49003a,a49004a,a49008a,a49009a,a49013a,a49014a,a49015a,a49019a,a49020a,a49023a,a49026a,a49027a,a49028a,a49032a,a49033a,a49037a,a49038a,a49039a,a49043a,a49044a,a49047a,a49050a,a49051a,a49052a,a49056a,a49057a,a49061a,a49062a,a49063a,a49067a,a49068a,a49071a,a49074a,a49075a,a49076a,a49080a,a49081a,a49085a,a49086a,a49087a,a49091a,a49092a,a49095a,a49098a,a49099a,a49100a,a49104a,a49105a,a49109a,a49110a,a49111a,a49115a,a49116a,a49119a,a49122a,a49123a,a49124a,a49128a,a49129a,a49133a,a49134a,a49135a,a49139a,a49140a,a49143a,a49146a,a49147a,a49148a,a49152a,a49153a,a49157a,a49158a,a49159a,a49163a,a49164a,a49167a,a49170a,a49171a,a49172a,a49176a,a49177a,a49181a,a49182a,a49183a,a49187a,a49188a,a49191a,a49194a,a49195a,a49196a,a49200a,a49201a,a49205a,a49206a,a49207a,a49211a,a49212a,a49215a,a49218a,a49219a,a49220a,a49224a,a49225a,a49229a,a49230a,a49231a,a49235a,a49236a,a49239a,a49242a,a49243a,a49244a,a49248a,a49249a,a49253a,a49254a,a49255a,a49259a,a49260a,a49263a,a49266a,a49267a,a49268a,a49272a,a49273a,a49277a,a49278a,a49279a,a49283a,a49284a,a49287a,a49290a,a49291a,a49292a,a49296a,a49297a,a49301a,a49302a,a49303a,a49307a,a49308a,a49311a,a49314a,a49315a,a49316a,a49320a,a49321a,a49325a,a49326a,a49327a,a49331a,a49332a,a49335a,a49338a,a49339a,a49340a,a49344a,a49345a,a49349a,a49350a,a49351a,a49355a,a49356a,a49359a,a49362a,a49363a,a49364a,a49368a,a49369a,a49373a,a49374a,a49375a,a49379a,a49380a,a49383a,a49386a,a49387a,a49388a,a49392a,a49393a,a49397a,a49398a,a49399a,a49403a,a49404a,a49407a,a49410a,a49411a,a49412a,a49416a,a49417a,a49421a,a49422a,a49423a,a49427a,a49428a,a49431a,a49434a,a49435a,a49436a,a49440a,a49441a,a49445a,a49446a,a49447a,a49451a,a49452a,a49455a,a49458a,a49459a,a49460a,a49464a,a49465a,a49469a,a49470a,a49471a,a49475a,a49476a,a49479a,a49482a,a49483a,a49484a,a49488a,a49489a,a49493a,a49494a,a49495a,a49499a,a49500a,a49503a,a49506a,a49507a,a49508a,a49512a,a49513a,a49517a,a49518a,a49519a,a49523a,a49524a,a49527a,a49530a,a49531a,a49532a,a49536a,a49537a,a49541a,a49542a,a49543a,a49547a,a49548a,a49551a,a49554a,a49555a,a49556a,a49560a,a49561a,a49565a,a49566a,a49567a,a49571a,a49572a,a49575a,a49578a,a49579a,a49580a,a49584a,a49585a,a49589a,a49590a,a49591a,a49595a,a49596a,a49599a,a49602a,a49603a,a49604a,a49608a,a49609a,a49613a,a49614a,a49615a,a49619a,a49620a,a49623a,a49626a,a49627a,a49628a,a49632a,a49633a,a49637a,a49638a,a49639a,a49643a,a49644a,a49647a,a49650a,a49651a,a49652a,a49656a,a49657a,a49661a,a49662a,a49663a,a49667a,a49668a,a49671a,a49674a,a49675a,a49676a,a49680a,a49681a,a49685a,a49686a,a49687a,a49691a,a49692a,a49695a,a49698a,a49699a,a49700a,a49704a,a49705a,a49709a,a49710a,a49711a,a49715a,a49716a,a49719a,a49722a,a49723a,a49724a,a49728a,a49729a,a49733a,a49734a,a49735a,a49739a,a49740a,a49743a,a49746a,a49747a,a49748a,a49752a,a49753a,a49757a,a49758a,a49759a,a49763a,a49764a,a49767a,a49770a,a49771a,a49772a,a49776a,a49777a,a49781a,a49782a,a49783a,a49787a,a49788a,a49791a,a49794a,a49795a,a49796a,a49800a,a49801a,a49805a,a49806a,a49807a,a49811a,a49812a,a49815a,a49818a,a49819a,a49820a,a49824a,a49825a,a49829a,a49830a,a49831a,a49835a,a49836a,a49839a,a49842a,a49843a,a49844a,a49848a,a49849a,a49853a,a49854a,a49855a,a49859a,a49860a,a49863a,a49866a,a49867a,a49868a,a49872a,a49873a,a49877a,a49878a,a49879a,a49883a,a49884a,a49887a,a49890a,a49891a,a49892a,a49896a,a49897a,a49901a,a49902a,a49903a,a49907a,a49908a,a49911a,a49914a,a49915a,a49916a,a49920a,a49921a,a49925a,a49926a,a49927a,a49931a,a49932a,a49935a,a49938a,a49939a,a49940a,a49944a,a49945a,a49949a,a49950a,a49951a,a49955a,a49956a,a49959a,a49962a,a49963a,a49964a,a49968a,a49969a,a49973a,a49974a,a49975a,a49979a,a49980a,a49983a,a49986a,a49987a,a49988a,a49992a,a49993a,a49997a,a49998a,a49999a,a50003a,a50004a,a50007a,a50010a,a50011a,a50012a,a50016a,a50017a,a50021a,a50022a,a50023a,a50027a,a50028a,a50031a,a50034a,a50035a,a50036a,a50040a,a50041a,a50045a,a50046a,a50047a,a50051a,a50052a,a50055a,a50058a,a50059a,a50060a,a50064a,a50065a,a50069a,a50070a,a50071a,a50075a,a50076a,a50079a,a50082a,a50083a,a50084a,a50088a,a50089a,a50093a,a50094a,a50095a,a50099a,a50100a,a50103a,a50106a,a50107a,a50108a,a50112a,a50113a,a50117a,a50118a,a50119a,a50123a,a50124a,a50127a,a50130a,a50131a,a50132a,a50136a,a50137a,a50141a,a50142a,a50143a,a50147a,a50148a,a50151a,a50154a,a50155a,a50156a,a50160a,a50161a,a50165a,a50166a,a50167a,a50171a,a50172a,a50175a,a50178a,a50179a,a50180a,a50184a,a50185a,a50189a,a50190a,a50191a,a50195a,a50196a,a50199a,a50202a,a50203a,a50204a,a50208a,a50209a,a50213a,a50214a,a50215a,a50219a,a50220a,a50223a,a50226a,a50227a,a50228a,a50232a,a50233a,a50237a,a50238a,a50239a,a50243a,a50244a,a50247a,a50250a,a50251a,a50252a,a50256a,a50257a,a50261a,a50262a,a50263a,a50267a,a50268a,a50271a,a50274a,a50275a,a50276a,a50280a,a50281a,a50285a,a50286a,a50287a,a50291a,a50292a,a50295a,a50298a,a50299a,a50300a,a50304a,a50305a,a50309a,a50310a,a50311a,a50315a,a50316a,a50319a,a50322a,a50323a,a50324a,a50328a,a50329a,a50333a,a50334a,a50335a,a50339a,a50340a,a50343a,a50346a,a50347a,a50348a,a50352a,a50353a,a50357a,a50358a,a50359a,a50363a,a50364a,a50367a,a50370a,a50371a,a50372a,a50376a,a50377a,a50381a,a50382a,a50383a,a50387a,a50388a,a50391a,a50394a,a50395a,a50396a,a50400a,a50401a,a50405a,a50406a,a50407a,a50411a,a50412a,a50415a,a50418a,a50419a,a50420a,a50424a,a50425a,a50429a,a50430a,a50431a,a50435a,a50436a,a50439a,a50442a,a50443a,a50444a,a50448a,a50449a,a50453a,a50454a,a50455a,a50459a,a50460a,a50463a,a50466a,a50467a,a50468a,a50472a,a50473a,a50477a,a50478a,a50479a,a50483a,a50484a,a50487a,a50490a,a50491a,a50492a,a50496a,a50497a,a50501a,a50502a,a50503a,a50507a,a50508a,a50511a,a50514a,a50515a,a50516a,a50520a,a50521a,a50525a,a50526a,a50527a,a50531a,a50532a,a50535a,a50538a,a50539a,a50540a,a50544a,a50545a,a50549a,a50550a,a50551a,a50555a,a50556a,a50559a,a50562a,a50563a,a50564a,a50568a,a50569a,a50573a,a50574a,a50575a,a50579a,a50580a,a50583a,a50586a,a50587a,a50588a,a50592a,a50593a,a50597a,a50598a,a50599a,a50603a,a50604a,a50607a,a50610a,a50611a,a50612a,a50616a,a50617a,a50621a,a50622a,a50623a,a50627a,a50628a,a50631a,a50634a,a50635a,a50636a,a50640a,a50641a,a50645a,a50646a,a50647a,a50651a,a50652a,a50655a,a50658a,a50659a,a50660a,a50664a,a50665a,a50669a,a50670a,a50671a,a50675a,a50676a,a50679a,a50682a,a50683a,a50684a,a50688a,a50689a,a50693a,a50694a,a50695a,a50699a,a50700a,a50703a,a50706a,a50707a,a50708a,a50712a,a50713a,a50717a,a50718a,a50719a,a50723a,a50724a,a50727a,a50730a,a50731a,a50732a,a50736a,a50737a,a50741a,a50742a,a50743a,a50747a,a50748a,a50751a,a50754a,a50755a,a50756a,a50760a,a50761a,a50765a,a50766a,a50767a,a50771a,a50772a,a50775a,a50778a,a50779a,a50780a,a50784a,a50785a,a50789a,a50790a,a50791a,a50795a,a50796a,a50799a,a50802a,a50803a,a50804a,a50808a,a50809a,a50813a,a50814a,a50815a,a50819a,a50820a,a50823a,a50826a,a50827a,a50828a,a50832a,a50833a,a50837a,a50838a,a50839a,a50843a,a50844a,a50847a,a50850a,a50851a,a50852a,a50856a,a50857a,a50861a,a50862a,a50863a,a50867a,a50868a,a50871a,a50874a,a50875a,a50876a,a50880a,a50881a,a50885a,a50886a,a50887a,a50891a,a50892a,a50895a,a50898a,a50899a,a50900a,a50904a,a50905a,a50909a,a50910a,a50911a,a50915a,a50916a,a50919a,a50922a,a50923a,a50924a,a50928a,a50929a,a50933a,a50934a,a50935a,a50939a,a50940a,a50943a,a50946a,a50947a,a50948a,a50952a,a50953a,a50957a,a50958a,a50959a,a50963a,a50964a,a50967a,a50970a,a50971a,a50972a,a50976a,a50977a,a50981a,a50982a,a50983a,a50987a,a50988a,a50991a,a50994a,a50995a,a50996a,a51000a,a51001a,a51005a,a51006a,a51007a,a51011a,a51012a,a51015a,a51018a,a51019a,a51020a,a51024a,a51025a,a51029a,a51030a,a51031a,a51035a,a51036a,a51039a,a51042a,a51043a,a51044a,a51048a,a51049a,a51053a,a51054a,a51055a,a51059a,a51060a,a51063a,a51066a,a51067a,a51068a,a51072a,a51073a,a51077a,a51078a,a51079a,a51083a,a51084a,a51087a,a51090a,a51091a,a51092a,a51096a,a51097a,a51101a,a51102a,a51103a,a51107a,a51108a,a51111a,a51114a,a51115a,a51116a,a51120a,a51121a,a51125a,a51126a,a51127a,a51131a,a51132a,a51135a,a51138a,a51139a,a51140a,a51144a,a51145a,a51149a,a51150a,a51151a,a51155a,a51156a,a51159a,a51162a,a51163a,a51164a,a51168a,a51169a,a51173a,a51174a,a51175a,a51179a,a51180a,a51183a,a51186a,a51187a,a51188a,a51192a,a51193a,a51197a,a51198a,a51199a,a51203a,a51204a,a51207a,a51210a,a51211a,a51212a,a51216a,a51217a,a51221a,a51222a,a51223a,a51227a,a51228a,a51231a,a51234a,a51235a,a51236a,a51240a,a51241a,a51245a,a51246a,a51247a,a51251a,a51252a,a51255a,a51258a,a51259a,a51260a,a51264a,a51265a,a51269a,a51270a,a51271a,a51275a,a51276a,a51279a,a51282a,a51283a,a51284a,a51288a,a51289a,a51293a,a51294a,a51295a,a51299a,a51300a,a51303a,a51306a,a51307a,a51308a,a51312a,a51313a,a51317a,a51318a,a51319a,a51323a,a51324a,a51327a,a51330a,a51331a,a51332a,a51336a,a51337a,a51341a,a51342a,a51343a,a51347a,a51348a,a51351a,a51354a,a51355a,a51356a,a51360a,a51361a,a51365a,a51366a,a51367a,a51371a,a51372a,a51375a,a51378a,a51379a,a51380a,a51384a,a51385a,a51389a,a51390a,a51391a,a51395a,a51396a,a51399a,a51402a,a51403a,a51404a,a51408a,a51409a,a51413a,a51414a,a51415a,a51419a,a51420a,a51423a,a51426a,a51427a,a51428a,a51432a,a51433a,a51437a,a51438a,a51439a,a51443a,a51444a,a51447a,a51450a,a51451a,a51452a,a51456a,a51457a,a51461a,a51462a,a51463a,a51467a,a51468a,a51471a,a51474a,a51475a,a51476a,a51480a,a51481a,a51485a,a51486a,a51487a,a51491a,a51492a,a51495a,a51498a,a51499a,a51500a,a51504a,a51505a,a51509a,a51510a,a51511a,a51515a,a51516a,a51519a,a51522a,a51523a,a51524a,a51528a,a51529a,a51533a,a51534a,a51535a,a51539a,a51540a,a51543a,a51546a,a51547a,a51548a,a51552a,a51553a,a51557a,a51558a,a51559a,a51563a,a51564a,a51567a,a51570a,a51571a,a51572a,a51576a,a51577a,a51581a,a51582a,a51583a,a51587a,a51588a,a51591a,a51594a,a51595a,a51596a,a51600a,a51601a,a51605a,a51606a,a51607a,a51611a,a51612a,a51615a,a51618a,a51619a,a51620a,a51624a,a51625a,a51629a,a51630a,a51631a,a51635a,a51636a,a51639a,a51642a,a51643a,a51644a,a51648a,a51649a,a51653a,a51654a,a51655a,a51659a,a51660a,a51663a,a51666a,a51667a,a51668a,a51672a,a51673a,a51677a,a51678a,a51679a,a51683a,a51684a,a51687a,a51690a,a51691a,a51692a,a51696a,a51697a,a51701a,a51702a,a51703a,a51707a,a51708a,a51711a,a51714a,a51715a,a51716a,a51720a,a51721a,a51725a,a51726a,a51727a,a51731a,a51732a,a51735a,a51738a,a51739a,a51740a,a51744a,a51745a,a51749a,a51750a,a51751a,a51755a,a51756a,a51759a,a51762a,a51763a,a51764a,a51768a,a51769a,a51773a,a51774a,a51775a,a51779a,a51780a,a51783a,a51786a,a51787a,a51788a,a51792a,a51793a,a51797a,a51798a,a51799a,a51803a,a51804a,a51807a,a51810a,a51811a,a51812a,a51816a,a51817a,a51821a,a51822a,a51823a,a51827a,a51828a,a51831a,a51834a,a51835a,a51836a,a51840a,a51841a,a51845a,a51846a,a51847a,a51851a,a51852a,a51855a,a51858a,a51859a,a51860a,a51864a,a51865a,a51869a,a51870a,a51871a,a51875a,a51876a,a51879a,a51882a,a51883a,a51884a,a51888a,a51889a,a51893a,a51894a,a51895a,a51899a,a51900a,a51903a,a51906a,a51907a,a51908a,a51912a,a51913a,a51917a,a51918a,a51919a,a51923a,a51924a,a51927a,a51930a,a51931a,a51932a,a51936a,a51937a,a51941a,a51942a,a51943a,a51947a,a51948a,a51951a,a51954a,a51955a,a51956a,a51960a,a51961a,a51965a,a51966a,a51967a,a51971a,a51972a,a51975a,a51978a,a51979a,a51980a,a51984a,a51985a,a51989a,a51990a,a51991a,a51995a,a51996a,a51999a,a52002a,a52003a,a52004a,a52008a,a52009a,a52013a,a52014a,a52015a,a52019a,a52020a,a52023a,a52026a,a52027a,a52028a,a52032a,a52033a,a52037a,a52038a,a52039a,a52043a,a52044a,a52047a,a52050a,a52051a,a52052a,a52056a,a52057a,a52061a,a52062a,a52063a,a52067a,a52068a,a52071a,a52074a,a52075a,a52076a,a52080a,a52081a,a52085a,a52086a,a52087a,a52091a,a52092a,a52095a,a52098a,a52099a,a52100a,a52104a,a52105a,a52109a,a52110a,a52111a,a52115a,a52116a,a52119a,a52122a,a52123a,a52124a,a52128a,a52129a,a52133a,a52134a,a52135a,a52139a,a52140a,a52143a,a52146a,a52147a,a52148a,a52152a,a52153a,a52157a,a52158a,a52159a,a52163a,a52164a,a52167a,a52170a,a52171a,a52172a,a52176a,a52177a,a52181a,a52182a,a52183a,a52187a,a52188a,a52191a,a52194a,a52195a,a52196a,a52200a,a52201a,a52205a,a52206a,a52207a,a52211a,a52212a,a52215a,a52218a,a52219a,a52220a,a52224a,a52225a,a52229a,a52230a,a52231a,a52235a,a52236a,a52239a,a52242a,a52243a,a52244a,a52248a,a52249a,a52253a,a52254a,a52255a,a52259a,a52260a,a52263a,a52266a,a52267a,a52268a,a52272a,a52273a,a52277a,a52278a,a52279a,a52283a,a52284a,a52287a,a52290a,a52291a,a52292a,a52296a,a52297a,a52301a,a52302a,a52303a,a52307a,a52308a,a52311a,a52314a,a52315a,a52316a,a52320a,a52321a,a52325a,a52326a,a52327a,a52331a,a52332a,a52335a,a52338a,a52339a,a52340a,a52344a,a52345a,a52349a,a52350a,a52351a,a52355a,a52356a,a52359a,a52362a,a52363a,a52364a,a52368a,a52369a,a52373a,a52374a,a52375a,a52379a,a52380a,a52383a,a52386a,a52387a,a52388a,a52392a,a52393a,a52397a,a52398a,a52399a,a52403a,a52404a,a52407a,a52410a,a52411a,a52412a,a52416a,a52417a,a52421a,a52422a,a52423a,a52427a,a52428a,a52431a,a52434a,a52435a,a52436a,a52440a,a52441a,a52445a,a52446a,a52447a,a52451a,a52452a,a52455a,a52458a,a52459a,a52460a,a52464a,a52465a,a52469a,a52470a,a52471a,a52475a,a52476a,a52479a,a52482a,a52483a,a52484a,a52488a,a52489a,a52493a,a52494a,a52495a,a52499a,a52500a,a52503a,a52506a,a52507a,a52508a,a52512a,a52513a,a52517a,a52518a,a52519a,a52523a,a52524a,a52527a,a52530a,a52531a,a52532a,a52536a,a52537a,a52541a,a52542a,a52543a,a52547a,a52548a,a52551a,a52554a,a52555a,a52556a,a52560a,a52561a,a52565a,a52566a,a52567a,a52571a,a52572a,a52575a,a52578a,a52579a,a52580a,a52584a,a52585a,a52589a,a52590a,a52591a,a52595a,a52596a,a52599a,a52602a,a52603a,a52604a,a52608a,a52609a,a52613a,a52614a,a52615a,a52619a,a52620a,a52623a,a52626a,a52627a,a52628a,a52632a,a52633a,a52637a,a52638a,a52639a,a52643a,a52644a,a52647a,a52650a,a52651a,a52652a,a52656a,a52657a,a52661a,a52662a,a52663a,a52667a,a52668a,a52671a,a52674a,a52675a,a52676a,a52680a,a52681a,a52685a,a52686a,a52687a,a52691a,a52692a,a52695a,a52698a,a52699a,a52700a,a52704a,a52705a,a52709a,a52710a,a52711a,a52715a,a52716a,a52719a,a52722a,a52723a,a52724a,a52728a,a52729a,a52733a,a52734a,a52735a,a52739a,a52740a,a52743a,a52746a,a52747a,a52748a,a52752a,a52753a,a52757a,a52758a,a52759a,a52763a,a52764a,a52767a,a52770a,a52771a,a52772a,a52776a,a52777a,a52781a,a52782a,a52783a,a52787a,a52788a,a52791a,a52794a,a52795a,a52796a,a52800a,a52801a,a52805a,a52806a,a52807a,a52811a,a52812a,a52815a,a52818a,a52819a,a52820a,a52824a,a52825a,a52829a,a52830a,a52831a,a52835a,a52836a,a52839a,a52842a,a52843a,a52844a,a52848a,a52849a,a52853a,a52854a,a52855a,a52859a,a52860a,a52863a,a52866a,a52867a,a52868a,a52872a,a52873a,a52877a,a52878a,a52879a,a52883a,a52884a,a52887a,a52890a,a52891a,a52892a,a52896a,a52897a,a52901a,a52902a,a52903a,a52907a,a52908a,a52911a,a52914a,a52915a,a52916a,a52920a,a52921a,a52925a,a52926a,a52927a,a52931a,a52932a,a52935a,a52938a,a52939a,a52940a,a52944a,a52945a,a52949a,a52950a,a52951a,a52955a,a52956a,a52959a,a52962a,a52963a,a52964a,a52968a,a52969a,a52973a,a52974a,a52975a,a52979a,a52980a,a52983a,a52986a,a52987a,a52988a,a52992a,a52993a,a52997a,a52998a,a52999a,a53003a,a53004a,a53007a,a53010a,a53011a,a53012a,a53016a,a53017a,a53021a,a53022a,a53023a,a53027a,a53028a,a53031a,a53034a,a53035a,a53036a,a53040a,a53041a,a53045a,a53046a,a53047a,a53051a,a53052a,a53055a,a53058a,a53059a,a53060a,a53064a,a53065a,a53069a,a53070a,a53071a,a53075a,a53076a,a53079a,a53082a,a53083a,a53084a,a53088a,a53089a,a53093a,a53094a,a53095a,a53099a,a53100a,a53103a,a53106a,a53107a,a53108a,a53112a,a53113a,a53117a,a53118a,a53119a,a53123a,a53124a,a53127a,a53130a,a53131a,a53132a,a53136a,a53137a,a53141a,a53142a,a53143a,a53147a,a53148a,a53151a,a53154a,a53155a,a53156a,a53160a,a53161a,a53165a,a53166a,a53167a,a53171a,a53172a,a53175a,a53178a,a53179a,a53180a,a53184a,a53185a,a53189a,a53190a,a53191a,a53195a,a53196a,a53199a,a53202a,a53203a,a53204a,a53208a,a53209a,a53213a,a53214a,a53215a,a53219a,a53220a,a53223a,a53226a,a53227a,a53228a,a53232a,a53233a,a53237a,a53238a,a53239a,a53243a,a53244a,a53247a,a53250a,a53251a,a53252a,a53256a,a53257a,a53261a,a53262a,a53263a,a53267a,a53268a,a53271a,a53274a,a53275a,a53276a,a53280a,a53281a,a53285a,a53286a,a53287a,a53291a,a53292a,a53295a,a53298a,a53299a,a53300a,a53304a,a53305a,a53309a,a53310a,a53311a,a53315a,a53316a,a53319a,a53322a,a53323a,a53324a,a53328a,a53329a,a53333a,a53334a,a53335a,a53339a,a53340a,a53343a,a53346a,a53347a,a53348a,a53352a,a53353a,a53357a,a53358a,a53359a,a53363a,a53364a,a53367a,a53370a,a53371a,a53372a,a53376a,a53377a,a53381a,a53382a,a53383a,a53387a,a53388a,a53391a,a53394a,a53395a,a53396a,a53400a,a53401a,a53405a,a53406a,a53407a,a53411a,a53412a,a53415a,a53418a,a53419a,a53420a,a53424a,a53425a,a53429a,a53430a,a53431a,a53435a,a53436a,a53439a,a53442a,a53443a,a53444a,a53448a,a53449a,a53453a,a53454a,a53455a,a53459a,a53460a,a53463a,a53466a,a53467a,a53468a,a53472a,a53473a,a53477a,a53478a,a53479a,a53483a,a53484a,a53487a,a53490a,a53491a,a53492a,a53496a,a53497a,a53501a,a53502a,a53503a,a53507a,a53508a,a53511a,a53514a,a53515a,a53516a,a53520a,a53521a,a53525a,a53526a,a53527a,a53531a,a53532a,a53535a,a53538a,a53539a,a53540a,a53544a,a53545a,a53549a,a53550a,a53551a,a53555a,a53556a,a53559a,a53562a,a53563a,a53564a,a53568a,a53569a,a53573a,a53574a,a53575a,a53579a,a53580a,a53583a,a53586a,a53587a,a53588a,a53592a,a53593a,a53597a,a53598a,a53599a,a53603a,a53604a,a53607a,a53610a,a53611a,a53612a,a53616a,a53617a,a53621a,a53622a,a53623a,a53627a,a53628a,a53631a,a53634a,a53635a,a53636a,a53640a,a53641a,a53645a,a53646a,a53647a,a53651a,a53652a,a53655a,a53658a,a53659a,a53660a,a53664a,a53665a,a53669a,a53670a,a53671a,a53675a,a53676a,a53679a,a53682a,a53683a,a53684a,a53688a,a53689a,a53693a,a53694a,a53695a,a53699a,a53700a,a53703a,a53706a,a53707a,a53708a,a53712a,a53713a,a53717a,a53718a,a53719a,a53723a,a53724a,a53727a,a53730a,a53731a,a53732a,a53736a,a53737a,a53741a,a53742a,a53743a,a53747a,a53748a,a53751a,a53754a,a53755a,a53756a,a53760a,a53761a,a53765a,a53766a,a53767a,a53771a,a53772a,a53775a,a53778a,a53779a,a53780a,a53784a,a53785a,a53789a,a53790a,a53791a,a53795a,a53796a,a53799a,a53802a,a53803a,a53804a,a53808a,a53809a,a53813a,a53814a,a53815a,a53819a,a53820a,a53823a,a53826a,a53827a,a53828a,a53832a,a53833a,a53837a,a53838a,a53839a,a53843a,a53844a,a53847a,a53850a,a53851a,a53852a,a53856a,a53857a,a53861a,a53862a,a53863a,a53867a,a53868a,a53871a,a53874a,a53875a,a53876a,a53880a,a53881a,a53885a,a53886a,a53887a,a53891a,a53892a,a53895a,a53898a,a53899a,a53900a,a53904a,a53905a,a53909a,a53910a,a53911a,a53915a,a53916a,a53919a,a53922a,a53923a,a53924a,a53928a,a53929a,a53933a,a53934a,a53935a,a53939a,a53940a,a53943a,a53946a,a53947a,a53948a,a53952a,a53953a,a53957a,a53958a,a53959a,a53963a,a53964a,a53967a,a53970a,a53971a,a53972a,a53976a,a53977a,a53981a,a53982a,a53983a,a53987a,a53988a,a53991a,a53994a,a53995a,a53996a,a54000a,a54001a,a54005a,a54006a,a54007a,a54011a,a54012a,a54015a,a54018a,a54019a,a54020a,a54024a,a54025a,a54029a,a54030a,a54031a,a54035a,a54036a,a54039a,a54042a,a54043a,a54044a,a54048a,a54049a,a54053a,a54054a,a54055a,a54059a,a54060a,a54063a,a54066a,a54067a,a54068a,a54072a,a54073a,a54077a,a54078a,a54079a,a54083a,a54084a,a54087a,a54090a,a54091a,a54092a,a54096a,a54097a,a54101a,a54102a,a54103a,a54107a,a54108a,a54111a,a54114a,a54115a,a54116a,a54120a,a54121a,a54125a,a54126a,a54127a,a54131a,a54132a,a54135a,a54138a,a54139a,a54140a,a54144a,a54145a,a54149a,a54150a,a54151a,a54155a,a54156a,a54159a,a54162a,a54163a,a54164a,a54168a,a54169a,a54173a,a54174a,a54175a,a54179a,a54180a,a54183a,a54186a,a54187a,a54188a,a54192a,a54193a,a54197a,a54198a,a54199a,a54203a,a54204a,a54207a,a54210a,a54211a,a54212a,a54216a,a54217a,a54221a,a54222a,a54223a,a54227a,a54228a,a54231a,a54234a,a54235a,a54236a,a54240a,a54241a,a54245a,a54246a,a54247a,a54251a,a54252a,a54255a,a54258a,a54259a,a54260a,a54264a,a54265a,a54269a,a54270a,a54271a,a54275a,a54276a,a54279a,a54282a,a54283a,a54284a,a54288a,a54289a,a54293a,a54294a,a54295a,a54299a,a54300a,a54303a,a54306a,a54307a,a54308a,a54312a,a54313a,a54317a,a54318a,a54319a,a54323a,a54324a,a54327a,a54330a,a54331a,a54332a,a54336a,a54337a,a54341a,a54342a,a54343a,a54347a,a54348a,a54351a,a54354a,a54355a,a54356a,a54360a,a54361a,a54365a,a54366a,a54367a,a54371a,a54372a,a54375a,a54378a,a54379a,a54380a,a54384a,a54385a,a54389a,a54390a,a54391a,a54395a,a54396a,a54399a,a54402a,a54403a,a54404a,a54408a,a54409a,a54413a,a54414a,a54415a,a54419a,a54420a,a54423a,a54426a,a54427a,a54428a,a54432a,a54433a,a54437a,a54438a,a54439a,a54443a,a54444a,a54447a,a54450a,a54451a,a54452a,a54456a,a54457a,a54461a,a54462a,a54463a,a54467a,a54468a,a54471a,a54474a,a54475a,a54476a,a54480a,a54481a,a54485a,a54486a,a54487a,a54491a,a54492a,a54495a,a54498a,a54499a,a54500a,a54504a,a54505a,a54509a,a54510a,a54511a,a54515a,a54516a,a54519a,a54522a,a54523a,a54524a,a54528a,a54529a,a54533a,a54534a,a54535a,a54539a,a54540a,a54543a,a54546a,a54547a,a54548a,a54552a,a54553a,a54557a,a54558a,a54559a,a54563a,a54564a,a54567a,a54570a,a54571a,a54572a,a54576a,a54577a,a54581a,a54582a,a54583a,a54587a,a54588a,a54591a,a54594a,a54595a,a54596a,a54600a,a54601a,a54605a,a54606a,a54607a,a54611a,a54612a,a54615a,a54618a,a54619a,a54620a,a54624a,a54625a,a54629a,a54630a,a54631a,a54635a,a54636a,a54639a,a54642a,a54643a,a54644a,a54648a,a54649a,a54653a,a54654a,a54655a,a54659a,a54660a,a54663a,a54666a,a54667a,a54668a,a54672a,a54673a,a54677a,a54678a,a54679a,a54683a,a54684a,a54687a,a54690a,a54691a,a54692a,a54696a,a54697a,a54701a,a54702a,a54703a,a54707a,a54708a,a54711a,a54714a,a54715a,a54716a,a54720a,a54721a,a54725a,a54726a,a54727a,a54731a,a54732a,a54735a,a54738a,a54739a,a54740a,a54744a,a54745a,a54749a,a54750a,a54751a,a54755a,a54756a,a54759a,a54762a,a54763a,a54764a,a54768a,a54769a,a54773a,a54774a,a54775a,a54779a,a54780a,a54783a,a54786a,a54787a,a54788a,a54792a,a54793a,a54797a,a54798a,a54799a,a54803a,a54804a,a54807a,a54810a,a54811a,a54812a,a54816a,a54817a,a54821a,a54822a,a54823a,a54827a,a54828a,a54831a,a54834a,a54835a,a54836a,a54840a,a54841a,a54845a,a54846a,a54847a,a54851a,a54852a,a54855a,a54858a,a54859a,a54860a,a54864a,a54865a,a54869a,a54870a,a54871a,a54875a,a54876a,a54879a,a54882a,a54883a,a54884a,a54888a,a54889a,a54893a,a54894a,a54895a,a54899a,a54900a,a54903a,a54906a,a54907a,a54908a,a54912a,a54913a,a54917a,a54918a,a54919a,a54923a,a54924a,a54927a,a54930a,a54931a,a54932a,a54936a,a54937a,a54941a,a54942a,a54943a,a54947a,a54948a,a54951a,a54954a,a54955a,a54956a,a54960a,a54961a,a54965a,a54966a,a54967a,a54971a,a54972a,a54975a,a54978a,a54979a,a54980a,a54984a,a54985a,a54989a,a54990a,a54991a,a54995a,a54996a,a54999a,a55002a,a55003a,a55004a,a55008a,a55009a,a55013a,a55014a,a55015a,a55019a,a55020a,a55023a,a55026a,a55027a,a55028a,a55032a,a55033a,a55037a,a55038a,a55039a,a55043a,a55044a,a55047a,a55050a,a55051a,a55052a,a55056a,a55057a,a55061a,a55062a,a55063a,a55067a,a55068a,a55071a,a55074a,a55075a,a55076a,a55080a,a55081a,a55085a,a55086a,a55087a,a55091a,a55092a,a55095a,a55098a,a55099a,a55100a,a55104a,a55105a,a55109a,a55110a,a55111a,a55115a,a55116a,a55119a,a55122a,a55123a,a55124a,a55128a,a55129a,a55133a,a55134a,a55135a,a55139a,a55140a,a55143a,a55146a,a55147a,a55148a,a55152a,a55153a,a55157a,a55158a,a55159a,a55163a,a55164a,a55167a,a55170a,a55171a,a55172a,a55176a,a55177a,a55181a,a55182a,a55183a,a55187a,a55188a,a55191a,a55194a,a55195a,a55196a,a55200a,a55201a,a55205a,a55206a,a55207a,a55211a,a55212a,a55215a,a55218a,a55219a,a55220a,a55224a,a55225a,a55229a,a55230a,a55231a,a55235a,a55236a,a55239a,a55242a,a55243a,a55244a,a55248a,a55249a,a55253a,a55254a,a55255a,a55259a,a55260a,a55263a,a55266a,a55267a,a55268a,a55272a,a55273a,a55277a,a55278a,a55279a,a55283a,a55284a,a55287a,a55290a,a55291a,a55292a,a55296a,a55297a,a55301a,a55302a,a55303a,a55307a,a55308a,a55311a,a55314a,a55315a,a55316a,a55320a,a55321a,a55325a,a55326a,a55327a,a55331a,a55332a,a55335a,a55338a,a55339a,a55340a,a55344a,a55345a,a55349a,a55350a,a55351a,a55355a,a55356a,a55359a,a55362a,a55363a,a55364a,a55368a,a55369a,a55373a,a55374a,a55375a,a55379a,a55380a,a55383a,a55386a,a55387a,a55388a,a55392a,a55393a,a55397a,a55398a,a55399a,a55403a,a55404a,a55407a,a55410a,a55411a,a55412a,a55416a,a55417a,a55421a,a55422a,a55423a,a55427a,a55428a,a55431a,a55434a,a55435a,a55436a,a55440a,a55441a,a55445a,a55446a,a55447a,a55451a,a55452a,a55455a,a55458a,a55459a,a55460a,a55464a,a55465a,a55469a,a55470a,a55471a,a55475a,a55476a,a55479a,a55482a,a55483a,a55484a,a55488a,a55489a,a55493a,a55494a,a55495a,a55499a,a55500a,a55503a,a55506a,a55507a,a55508a,a55512a,a55513a,a55517a,a55518a,a55519a,a55523a,a55524a,a55527a,a55530a,a55531a,a55532a,a55536a,a55537a,a55541a,a55542a,a55543a,a55547a,a55548a,a55551a,a55554a,a55555a,a55556a,a55560a,a55561a,a55565a,a55566a,a55567a,a55571a,a55572a,a55575a,a55578a,a55579a,a55580a,a55584a,a55585a,a55589a,a55590a,a55591a,a55595a,a55596a,a55599a,a55602a,a55603a,a55604a,a55608a,a55609a,a55613a,a55614a,a55615a,a55619a,a55620a,a55623a,a55626a,a55627a,a55628a,a55632a,a55633a,a55637a,a55638a,a55639a,a55643a,a55644a,a55647a,a55650a,a55651a,a55652a,a55656a,a55657a,a55661a,a55662a,a55663a,a55667a,a55668a,a55671a,a55674a,a55675a,a55676a,a55680a,a55681a,a55685a,a55686a,a55687a,a55691a,a55692a,a55695a,a55698a,a55699a,a55700a,a55704a,a55705a,a55709a,a55710a,a55711a,a55715a,a55716a,a55719a,a55722a,a55723a,a55724a,a55728a,a55729a,a55733a,a55734a,a55735a,a55739a,a55740a,a55743a,a55746a,a55747a,a55748a,a55752a,a55753a,a55757a,a55758a,a55759a,a55763a,a55764a,a55767a,a55770a,a55771a,a55772a,a55776a,a55777a,a55781a,a55782a,a55783a,a55787a,a55788a,a55791a,a55794a,a55795a,a55796a,a55800a,a55801a,a55805a,a55806a,a55807a,a55811a,a55812a,a55815a,a55818a,a55819a,a55820a,a55824a,a55825a,a55829a,a55830a,a55831a,a55835a,a55836a,a55839a,a55842a,a55843a,a55844a,a55848a,a55849a,a55853a,a55854a,a55855a,a55859a,a55860a,a55863a,a55866a,a55867a,a55868a,a55872a,a55873a,a55877a,a55878a,a55879a,a55883a,a55884a,a55887a,a55890a,a55891a,a55892a,a55896a,a55897a,a55901a,a55902a,a55903a,a55907a,a55908a,a55911a,a55914a,a55915a,a55916a,a55920a,a55921a,a55925a,a55926a,a55927a,a55931a,a55932a,a55935a,a55938a,a55939a,a55940a,a55944a,a55945a,a55949a,a55950a,a55951a,a55955a,a55956a,a55959a,a55962a,a55963a,a55964a,a55968a,a55969a,a55973a,a55974a,a55975a,a55979a,a55980a,a55983a,a55986a,a55987a,a55988a,a55992a,a55993a,a55997a,a55998a,a55999a,a56003a,a56004a,a56007a,a56010a,a56011a,a56012a,a56016a,a56017a,a56021a,a56022a,a56023a,a56027a,a56028a,a56031a,a56034a,a56035a,a56036a,a56040a,a56041a,a56045a,a56046a,a56047a,a56051a,a56052a,a56055a,a56058a,a56059a,a56060a,a56064a,a56065a,a56069a,a56070a,a56071a,a56075a,a56076a,a56079a,a56082a,a56083a,a56084a,a56088a,a56089a,a56093a,a56094a,a56095a,a56099a,a56100a,a56103a,a56106a,a56107a,a56108a,a56112a,a56113a,a56117a,a56118a,a56119a,a56123a,a56124a,a56127a,a56130a,a56131a,a56132a,a56136a,a56137a,a56141a,a56142a,a56143a,a56147a,a56148a,a56151a,a56154a,a56155a,a56156a,a56160a,a56161a,a56165a,a56166a,a56167a,a56171a,a56172a,a56175a,a56178a,a56179a,a56180a,a56184a,a56185a,a56189a,a56190a,a56191a,a56195a,a56196a,a56199a,a56202a,a56203a,a56204a,a56208a,a56209a,a56213a,a56214a,a56215a,a56219a,a56220a,a56223a,a56226a,a56227a,a56228a,a56232a,a56233a,a56237a,a56238a,a56239a,a56243a,a56244a,a56247a,a56250a,a56251a,a56252a,a56256a,a56257a,a56261a,a56262a,a56263a,a56267a,a56268a,a56271a,a56274a,a56275a,a56276a,a56280a,a56281a,a56285a,a56286a,a56287a,a56291a,a56292a,a56295a,a56298a,a56299a,a56300a,a56304a,a56305a,a56309a,a56310a,a56311a,a56315a,a56316a,a56319a,a56322a,a56323a,a56324a,a56328a,a56329a,a56333a,a56334a,a56335a,a56339a,a56340a,a56343a,a56346a,a56347a,a56348a,a56352a,a56353a,a56357a,a56358a,a56359a,a56363a,a56364a,a56367a,a56370a,a56371a,a56372a,a56376a,a56377a,a56381a,a56382a,a56383a,a56387a,a56388a,a56391a,a56394a,a56395a,a56396a,a56400a,a56401a,a56405a,a56406a,a56407a,a56411a,a56412a,a56415a,a56418a,a56419a,a56420a,a56424a,a56425a,a56429a,a56430a,a56431a,a56435a,a56436a,a56439a,a56442a,a56443a,a56444a,a56448a,a56449a,a56453a,a56454a,a56455a,a56459a,a56460a,a56463a,a56466a,a56467a,a56468a,a56472a,a56473a,a56477a,a56478a,a56479a,a56483a,a56484a,a56487a,a56490a,a56491a,a56492a,a56496a,a56497a,a56501a,a56502a,a56503a,a56507a,a56508a,a56511a,a56514a,a56515a,a56516a,a56520a,a56521a,a56525a,a56526a,a56527a,a56531a,a56532a,a56535a,a56538a,a56539a,a56540a,a56544a,a56545a,a56549a,a56550a,a56551a,a56555a,a56556a,a56559a,a56562a,a56563a,a56564a,a56568a,a56569a,a56573a,a56574a,a56575a,a56579a,a56580a,a56583a,a56586a,a56587a,a56588a,a56592a,a56593a,a56597a,a56598a,a56599a,a56603a,a56604a,a56607a,a56610a,a56611a,a56612a,a56616a,a56617a,a56621a,a56622a,a56623a,a56627a,a56628a,a56631a,a56634a,a56635a,a56636a,a56640a,a56641a,a56645a,a56646a,a56647a,a56651a,a56652a,a56655a,a56658a,a56659a,a56660a,a56664a,a56665a,a56669a,a56670a,a56671a,a56675a,a56676a,a56679a,a56682a,a56683a,a56684a,a56688a,a56689a,a56693a,a56694a,a56695a,a56699a,a56700a,a56703a,a56706a,a56707a,a56708a,a56712a,a56713a,a56717a,a56718a,a56719a,a56723a,a56724a,a56727a,a56730a,a56731a,a56732a,a56736a,a56737a,a56741a,a56742a,a56743a,a56747a,a56748a,a56751a,a56754a,a56755a,a56756a,a56760a,a56761a,a56765a,a56766a,a56767a,a56771a,a56772a,a56775a,a56778a,a56779a,a56780a,a56784a,a56785a,a56789a,a56790a,a56791a,a56795a,a56796a,a56799a,a56802a,a56803a,a56804a,a56808a,a56809a,a56813a,a56814a,a56815a,a56819a,a56820a,a56823a,a56826a,a56827a,a56828a,a56832a,a56833a,a56837a,a56838a,a56839a,a56843a,a56844a,a56847a,a56850a,a56851a,a56852a,a56856a,a56857a,a56861a,a56862a,a56863a,a56867a,a56868a,a56871a,a56874a,a56875a,a56876a,a56880a,a56881a,a56885a,a56886a,a56887a,a56891a,a56892a,a56895a,a56898a,a56899a,a56900a,a56904a,a56905a,a56909a,a56910a,a56911a,a56915a,a56916a,a56919a,a56922a,a56923a,a56924a,a56928a,a56929a,a56933a,a56934a,a56935a,a56939a,a56940a,a56943a,a56946a,a56947a,a56948a,a56952a,a56953a,a56957a,a56958a,a56959a,a56963a,a56964a,a56967a,a56970a,a56971a,a56972a,a56976a,a56977a,a56981a,a56982a,a56983a,a56987a,a56988a,a56991a,a56994a,a56995a,a56996a,a57000a,a57001a,a57005a,a57006a,a57007a,a57011a,a57012a,a57015a,a57018a,a57019a,a57020a,a57024a,a57025a,a57029a,a57030a,a57031a,a57035a,a57036a,a57039a,a57042a,a57043a,a57044a,a57048a,a57049a,a57053a,a57054a,a57055a,a57059a,a57060a,a57063a,a57066a,a57067a,a57068a,a57072a,a57073a,a57077a,a57078a,a57079a,a57083a,a57084a,a57087a,a57090a,a57091a,a57092a,a57096a,a57097a,a57101a,a57102a,a57103a,a57107a,a57108a,a57111a,a57114a,a57115a,a57116a,a57120a,a57121a,a57125a,a57126a,a57127a,a57131a,a57132a,a57135a,a57138a,a57139a,a57140a,a57144a,a57145a,a57149a,a57150a,a57151a,a57155a,a57156a,a57159a,a57162a,a57163a,a57164a,a57168a,a57169a,a57173a,a57174a,a57175a,a57179a,a57180a,a57183a,a57186a,a57187a,a57188a,a57192a,a57193a,a57197a,a57198a,a57199a,a57203a,a57204a,a57207a,a57210a,a57211a,a57212a,a57216a,a57217a,a57221a,a57222a,a57223a,a57227a,a57228a,a57231a,a57234a,a57235a,a57236a,a57240a,a57241a,a57245a,a57246a,a57247a,a57251a,a57252a,a57255a,a57258a,a57259a,a57260a,a57264a,a57265a,a57269a,a57270a,a57271a,a57275a,a57276a,a57279a,a57282a,a57283a,a57284a,a57288a,a57289a,a57293a,a57294a,a57295a,a57299a,a57300a,a57303a,a57306a,a57307a,a57308a,a57312a,a57313a,a57317a,a57318a,a57319a,a57323a,a57324a,a57327a,a57330a,a57331a,a57332a,a57336a,a57337a,a57341a,a57342a,a57343a,a57347a,a57348a,a57351a,a57354a,a57355a,a57356a,a57360a,a57361a,a57365a,a57366a,a57367a,a57371a,a57372a,a57375a,a57378a,a57379a,a57380a,a57384a,a57385a,a57389a,a57390a,a57391a,a57395a,a57396a,a57399a,a57402a,a57403a,a57404a,a57408a,a57409a,a57413a,a57414a,a57415a,a57419a,a57420a,a57423a,a57426a,a57427a,a57428a,a57432a,a57433a,a57437a,a57438a,a57439a,a57443a,a57444a,a57447a,a57450a,a57451a,a57452a,a57456a,a57457a,a57461a,a57462a,a57463a,a57467a,a57468a,a57471a,a57474a,a57475a,a57476a,a57480a,a57481a,a57485a,a57486a,a57487a,a57491a,a57492a,a57495a,a57498a,a57499a,a57500a,a57504a,a57505a,a57509a,a57510a,a57511a,a57515a,a57516a,a57519a,a57522a,a57523a,a57524a,a57528a,a57529a,a57533a,a57534a,a57535a,a57539a,a57540a,a57543a,a57546a,a57547a,a57548a,a57552a,a57553a,a57557a,a57558a,a57559a,a57563a,a57564a,a57567a,a57570a,a57571a,a57572a,a57576a,a57577a,a57581a,a57582a,a57583a,a57587a,a57588a,a57591a,a57594a,a57595a,a57596a,a57600a,a57601a,a57605a,a57606a,a57607a,a57611a,a57612a,a57615a,a57618a,a57619a,a57620a,a57624a,a57625a,a57629a,a57630a,a57631a,a57635a,a57636a,a57639a,a57642a,a57643a,a57644a,a57648a,a57649a,a57653a,a57654a,a57655a,a57659a,a57660a,a57663a,a57666a,a57667a,a57668a,a57672a,a57673a,a57677a,a57678a,a57679a,a57683a,a57684a,a57687a,a57690a,a57691a,a57692a,a57696a,a57697a,a57701a,a57702a,a57703a,a57707a,a57708a,a57711a,a57714a,a57715a,a57716a,a57720a,a57721a,a57725a,a57726a,a57727a,a57731a,a57732a,a57735a,a57738a,a57739a,a57740a,a57744a,a57745a,a57749a,a57750a,a57751a,a57755a,a57756a,a57759a,a57762a,a57763a,a57764a,a57768a,a57769a,a57773a,a57774a,a57775a,a57779a,a57780a,a57783a,a57786a,a57787a,a57788a,a57792a,a57793a,a57797a,a57798a,a57799a,a57803a,a57804a,a57807a,a57810a,a57811a,a57812a,a57816a,a57817a,a57821a,a57822a,a57823a,a57827a,a57828a,a57831a,a57834a,a57835a,a57836a,a57840a,a57841a,a57845a,a57846a,a57847a,a57851a,a57852a,a57855a,a57858a,a57859a,a57860a,a57864a,a57865a,a57869a,a57870a,a57871a,a57875a,a57876a,a57879a,a57882a,a57883a,a57884a,a57888a,a57889a,a57893a,a57894a,a57895a,a57899a,a57900a,a57903a,a57906a,a57907a,a57908a,a57912a,a57913a,a57917a,a57918a,a57919a,a57923a,a57924a,a57927a,a57930a,a57931a,a57932a,a57936a,a57937a,a57941a,a57942a,a57943a,a57947a,a57948a,a57951a,a57954a,a57955a,a57956a,a57960a,a57961a,a57965a,a57966a,a57967a,a57971a,a57972a,a57975a,a57978a,a57979a,a57980a,a57984a,a57985a,a57989a,a57990a,a57991a,a57995a,a57996a,a57999a,a58002a,a58003a,a58004a,a58008a,a58009a,a58013a,a58014a,a58015a,a58019a,a58020a,a58023a,a58026a,a58027a,a58028a,a58032a,a58033a,a58037a,a58038a,a58039a,a58043a,a58044a,a58047a,a58050a,a58051a,a58052a,a58056a,a58057a,a58061a,a58062a,a58063a,a58067a,a58068a,a58071a,a58074a,a58075a,a58076a,a58080a,a58081a,a58085a,a58086a,a58087a,a58091a,a58092a,a58095a,a58098a,a58099a,a58100a,a58104a,a58105a,a58109a,a58110a,a58111a,a58115a,a58116a,a58119a,a58122a,a58123a,a58124a,a58128a,a58129a,a58133a,a58134a,a58135a,a58139a,a58140a,a58143a,a58146a,a58147a,a58148a,a58152a,a58153a,a58157a,a58158a,a58159a,a58163a,a58164a,a58167a,a58170a,a58171a,a58172a,a58176a,a58177a,a58181a,a58182a,a58183a,a58187a,a58188a,a58191a,a58194a,a58195a,a58196a,a58200a,a58201a,a58205a,a58206a,a58207a,a58211a,a58212a,a58215a,a58218a,a58219a,a58220a,a58224a,a58225a,a58229a,a58230a,a58231a,a58235a,a58236a,a58239a,a58242a,a58243a,a58244a,a58248a,a58249a,a58253a,a58254a,a58255a,a58259a,a58260a,a58263a,a58266a,a58267a,a58268a,a58272a,a58273a,a58277a,a58278a,a58279a,a58283a,a58284a,a58287a,a58290a,a58291a,a58292a,a58296a,a58297a,a58301a,a58302a,a58303a,a58307a,a58308a,a58311a,a58314a,a58315a,a58316a,a58320a,a58321a,a58325a,a58326a,a58327a,a58331a,a58332a,a58335a,a58338a,a58339a,a58340a,a58344a,a58345a,a58349a,a58350a,a58351a,a58355a,a58356a,a58359a,a58362a,a58363a,a58364a,a58368a,a58369a,a58373a,a58374a,a58375a,a58379a,a58380a,a58383a,a58386a,a58387a,a58388a,a58392a,a58393a,a58397a,a58398a,a58399a,a58403a,a58404a,a58407a,a58410a,a58411a,a58412a,a58416a,a58417a,a58421a,a58422a,a58423a,a58427a,a58428a,a58431a,a58434a,a58435a,a58436a,a58440a,a58441a,a58445a,a58446a,a58447a,a58451a,a58452a,a58455a,a58458a,a58459a,a58460a,a58464a,a58465a,a58469a,a58470a,a58471a,a58475a,a58476a,a58479a,a58482a,a58483a,a58484a,a58488a,a58489a,a58493a,a58494a,a58495a,a58499a,a58500a,a58503a,a58506a,a58507a,a58508a,a58512a,a58513a,a58517a,a58518a,a58519a,a58523a,a58524a,a58527a,a58530a,a58531a,a58532a,a58536a,a58537a,a58541a,a58542a,a58543a,a58547a,a58548a,a58551a,a58554a,a58555a,a58556a,a58560a,a58561a,a58565a,a58566a,a58567a,a58571a,a58572a,a58575a,a58578a,a58579a,a58580a,a58584a,a58585a,a58589a,a58590a,a58591a,a58595a,a58596a,a58599a,a58602a,a58603a,a58604a,a58608a,a58609a,a58613a,a58614a,a58615a,a58619a,a58620a,a58623a,a58626a,a58627a,a58628a,a58632a,a58633a,a58637a,a58638a,a58639a,a58643a,a58644a,a58647a,a58650a,a58651a,a58652a,a58656a,a58657a,a58661a,a58662a,a58663a,a58667a,a58668a,a58671a,a58674a,a58675a,a58676a,a58680a,a58681a,a58685a,a58686a,a58687a,a58691a,a58692a,a58695a,a58698a,a58699a,a58700a,a58704a,a58705a,a58709a,a58710a,a58711a,a58715a,a58716a,a58719a,a58722a,a58723a,a58724a,a58728a,a58729a,a58733a,a58734a,a58735a,a58739a,a58740a,a58743a,a58746a,a58747a,a58748a,a58752a,a58753a,a58757a,a58758a,a58759a,a58763a,a58764a,a58767a,a58770a,a58771a,a58772a,a58776a,a58777a,a58781a,a58782a,a58783a,a58787a,a58788a,a58791a,a58794a,a58795a,a58796a,a58800a,a58801a,a58805a,a58806a,a58807a,a58811a,a58812a,a58815a,a58818a,a58819a,a58820a,a58824a,a58825a,a58829a,a58830a,a58831a,a58835a,a58836a,a58839a,a58842a,a58843a,a58844a,a58848a,a58849a,a58853a,a58854a,a58855a,a58859a,a58860a,a58863a,a58866a,a58867a,a58868a,a58872a,a58873a,a58877a,a58878a,a58879a,a58883a,a58884a,a58887a,a58890a,a58891a,a58892a,a58896a,a58897a,a58901a,a58902a,a58903a,a58907a,a58908a,a58911a,a58914a,a58915a,a58916a,a58920a,a58921a,a58925a,a58926a,a58927a,a58931a,a58932a,a58935a,a58938a,a58939a,a58940a,a58944a,a58945a,a58949a,a58950a,a58951a,a58955a,a58956a,a58959a,a58962a,a58963a,a58964a,a58968a,a58969a,a58973a,a58974a,a58975a,a58979a,a58980a,a58983a,a58986a,a58987a,a58988a,a58992a,a58993a,a58997a,a58998a,a58999a,a59003a,a59004a,a59007a,a59010a,a59011a,a59012a,a59016a,a59017a,a59021a,a59022a,a59023a,a59027a,a59028a,a59031a,a59034a,a59035a,a59036a,a59040a,a59041a,a59045a,a59046a,a59047a,a59051a,a59052a,a59055a,a59058a,a59059a,a59060a,a59064a,a59065a,a59069a,a59070a,a59071a,a59075a,a59076a,a59079a,a59082a,a59083a,a59084a,a59088a,a59089a,a59093a,a59094a,a59095a,a59099a,a59100a,a59103a,a59106a,a59107a,a59108a,a59112a,a59113a,a59117a,a59118a,a59119a,a59123a,a59124a,a59127a,a59130a,a59131a,a59132a,a59136a,a59137a,a59141a,a59142a,a59143a,a59147a,a59148a,a59151a,a59154a,a59155a,a59156a,a59160a,a59161a,a59165a,a59166a,a59167a,a59171a,a59172a,a59175a,a59178a,a59179a,a59180a,a59184a,a59185a,a59189a,a59190a,a59191a,a59195a,a59196a,a59199a,a59202a,a59203a,a59204a,a59208a,a59209a,a59213a,a59214a,a59215a,a59219a,a59220a,a59223a,a59226a,a59227a,a59228a,a59232a,a59233a,a59237a,a59238a,a59239a,a59243a,a59244a,a59247a,a59250a,a59251a,a59252a,a59256a,a59257a,a59261a,a59262a,a59263a,a59267a,a59268a,a59271a,a59274a,a59275a,a59276a,a59280a,a59281a,a59285a,a59286a,a59287a,a59291a,a59292a,a59295a,a59298a,a59299a,a59300a,a59304a,a59305a,a59309a,a59310a,a59311a,a59315a,a59316a,a59319a,a59322a,a59323a,a59324a,a59328a,a59329a,a59333a,a59334a,a59335a,a59339a,a59340a,a59343a,a59346a,a59347a,a59348a,a59352a,a59353a,a59357a,a59358a,a59359a,a59363a,a59364a,a59367a,a59370a,a59371a,a59372a,a59376a,a59377a,a59381a,a59382a,a59383a,a59387a,a59388a,a59391a,a59394a,a59395a,a59396a,a59400a,a59401a,a59405a,a59406a,a59407a,a59411a,a59412a,a59415a,a59418a,a59419a,a59420a,a59424a,a59425a,a59429a,a59430a,a59431a,a59435a,a59436a,a59439a,a59442a,a59443a,a59444a,a59448a,a59449a,a59453a,a59454a,a59455a,a59459a,a59460a,a59463a,a59466a,a59467a,a59468a,a59472a,a59473a,a59477a,a59478a,a59479a,a59483a,a59484a,a59487a,a59490a,a59491a,a59492a,a59496a,a59497a,a59501a,a59502a,a59503a,a59507a,a59508a,a59511a,a59514a,a59515a,a59516a,a59520a,a59521a,a59525a,a59526a,a59527a,a59531a,a59532a,a59535a,a59538a,a59539a,a59540a,a59544a,a59545a,a59549a,a59550a,a59551a,a59555a,a59556a,a59559a,a59562a,a59563a,a59564a,a59568a,a59569a,a59573a,a59574a,a59575a,a59579a,a59580a,a59583a,a59586a,a59587a,a59588a,a59592a,a59593a,a59597a,a59598a,a59599a,a59603a,a59604a,a59607a,a59610a,a59611a,a59612a,a59616a,a59617a,a59621a,a59622a,a59623a,a59627a,a59628a,a59631a,a59634a,a59635a,a59636a,a59640a,a59641a,a59645a,a59646a,a59647a,a59651a,a59652a,a59655a,a59658a,a59659a,a59660a,a59664a,a59665a,a59669a,a59670a,a59671a,a59675a,a59676a,a59679a,a59682a,a59683a,a59684a,a59688a,a59689a,a59693a,a59694a,a59695a,a59699a,a59700a,a59703a,a59706a,a59707a,a59708a,a59712a,a59713a,a59717a,a59718a,a59719a,a59723a,a59724a,a59727a,a59730a,a59731a,a59732a,a59736a,a59737a,a59741a,a59742a,a59743a,a59747a,a59748a,a59751a,a59754a,a59755a,a59756a,a59760a,a59761a,a59765a,a59766a,a59767a,a59771a,a59772a,a59775a,a59778a,a59779a,a59780a,a59784a,a59785a,a59789a,a59790a,a59791a,a59795a,a59796a,a59799a,a59802a,a59803a,a59804a,a59808a,a59809a,a59813a,a59814a,a59815a,a59819a,a59820a,a59823a,a59826a,a59827a,a59828a,a59832a,a59833a,a59837a,a59838a,a59839a,a59843a,a59844a,a59847a,a59850a,a59851a,a59852a,a59856a,a59857a,a59861a,a59862a,a59863a,a59867a,a59868a,a59871a,a59874a,a59875a,a59876a,a59880a,a59881a,a59885a,a59886a,a59887a,a59891a,a59892a,a59895a,a59898a,a59899a,a59900a,a59904a,a59905a,a59909a,a59910a,a59911a,a59915a,a59916a,a59919a,a59922a,a59923a,a59924a,a59928a,a59929a,a59933a,a59934a,a59935a,a59939a,a59940a,a59943a,a59946a,a59947a,a59948a,a59952a,a59953a,a59957a,a59958a,a59959a,a59963a,a59964a,a59967a,a59970a,a59971a,a59972a,a59976a,a59977a,a59981a,a59982a,a59983a,a59987a,a59988a,a59991a,a59994a,a59995a,a59996a,a60000a,a60001a,a60005a,a60006a,a60007a,a60011a,a60012a,a60015a,a60018a,a60019a,a60020a,a60024a,a60025a,a60029a,a60030a,a60031a,a60035a,a60036a,a60039a,a60042a,a60043a,a60044a,a60048a,a60049a,a60053a,a60054a,a60055a,a60059a,a60060a,a60063a,a60066a,a60067a,a60068a,a60072a,a60073a,a60077a,a60078a,a60079a,a60083a,a60084a,a60087a,a60090a,a60091a,a60092a,a60096a,a60097a,a60101a,a60102a,a60103a,a60107a,a60108a,a60111a,a60114a,a60115a,a60116a,a60120a,a60121a,a60125a,a60126a,a60127a,a60131a,a60132a,a60135a,a60138a,a60139a,a60140a,a60144a,a60145a,a60149a,a60150a,a60151a,a60155a,a60156a,a60159a,a60162a,a60163a,a60164a,a60168a,a60169a,a60173a,a60174a,a60175a,a60179a,a60180a,a60183a,a60186a,a60187a,a60188a,a60192a,a60193a,a60197a,a60198a,a60199a,a60203a,a60204a,a60207a,a60210a,a60211a,a60212a,a60216a,a60217a,a60221a,a60222a,a60223a,a60227a,a60228a,a60231a,a60234a,a60235a,a60236a,a60240a,a60241a,a60245a,a60246a,a60247a,a60251a,a60252a,a60255a,a60258a,a60259a,a60260a,a60264a,a60265a,a60269a,a60270a,a60271a,a60275a,a60276a,a60279a,a60282a,a60283a,a60284a,a60288a,a60289a,a60293a,a60294a,a60295a,a60299a,a60300a,a60303a,a60306a,a60307a,a60308a,a60312a,a60313a,a60317a,a60318a,a60319a,a60323a,a60324a,a60327a,a60330a,a60331a,a60332a,a60336a,a60337a,a60341a,a60342a,a60343a,a60347a,a60348a,a60351a,a60354a,a60355a,a60356a,a60360a,a60361a,a60365a,a60366a,a60367a,a60371a,a60372a,a60375a,a60378a,a60379a,a60380a,a60384a,a60385a,a60389a,a60390a,a60391a,a60395a,a60396a,a60399a,a60402a,a60403a,a60404a,a60408a,a60409a,a60413a,a60414a,a60415a,a60419a,a60420a,a60423a,a60426a,a60427a,a60428a,a60432a,a60433a,a60437a,a60438a,a60439a,a60443a,a60444a,a60447a,a60450a,a60451a,a60452a,a60456a,a60457a,a60461a,a60462a,a60463a,a60467a,a60468a,a60471a,a60474a,a60475a,a60476a,a60480a,a60481a,a60485a,a60486a,a60487a,a60491a,a60492a,a60495a,a60498a,a60499a,a60500a,a60504a,a60505a,a60509a,a60510a,a60511a,a60515a,a60516a,a60519a,a60522a,a60523a,a60524a,a60528a,a60529a,a60533a,a60534a,a60535a,a60539a,a60540a,a60543a,a60546a,a60547a,a60548a,a60552a,a60553a,a60557a,a60558a,a60559a,a60563a,a60564a,a60567a,a60570a,a60571a,a60572a,a60576a,a60577a,a60581a,a60582a,a60583a,a60587a,a60588a,a60591a,a60594a,a60595a,a60596a,a60600a,a60601a,a60605a,a60606a,a60607a,a60611a,a60612a,a60615a,a60618a,a60619a,a60620a,a60624a,a60625a,a60629a,a60630a,a60631a,a60635a,a60636a,a60639a,a60642a,a60643a,a60644a,a60648a,a60649a,a60653a,a60654a,a60655a,a60659a,a60660a,a60663a,a60666a,a60667a,a60668a,a60672a,a60673a,a60677a,a60678a,a60679a,a60683a,a60684a,a60687a,a60690a,a60691a,a60692a,a60696a,a60697a,a60701a,a60702a,a60703a,a60707a,a60708a,a60711a,a60714a,a60715a,a60716a,a60720a,a60721a,a60725a,a60726a,a60727a,a60731a,a60732a,a60735a,a60738a,a60739a,a60740a,a60744a,a60745a,a60749a,a60750a,a60751a,a60755a,a60756a,a60759a,a60762a,a60763a,a60764a,a60768a,a60769a,a60773a,a60774a,a60775a,a60779a,a60780a,a60783a,a60786a,a60787a,a60788a,a60792a,a60793a,a60797a,a60798a,a60799a,a60803a,a60804a,a60807a,a60810a,a60811a,a60812a,a60816a,a60817a,a60821a,a60822a,a60823a,a60827a,a60828a,a60831a,a60834a,a60835a,a60836a,a60840a,a60841a,a60845a,a60846a,a60847a,a60851a,a60852a,a60855a,a60858a,a60859a,a60860a,a60864a,a60865a,a60869a,a60870a,a60871a,a60875a,a60876a,a60879a,a60882a,a60883a,a60884a,a60888a,a60889a,a60893a,a60894a,a60895a,a60899a,a60900a,a60903a,a60906a,a60907a,a60908a,a60912a,a60913a,a60917a,a60918a,a60919a,a60923a,a60924a,a60927a,a60930a,a60931a,a60932a,a60936a,a60937a,a60941a,a60942a,a60943a,a60947a,a60948a,a60951a,a60954a,a60955a,a60956a,a60960a,a60961a,a60965a,a60966a,a60967a,a60971a,a60972a,a60975a,a60978a,a60979a,a60980a,a60984a,a60985a,a60989a,a60990a,a60991a,a60995a,a60996a,a60999a,a61002a,a61003a,a61004a,a61008a,a61009a,a61013a,a61014a,a61015a,a61019a,a61020a,a61023a,a61026a,a61027a,a61028a,a61032a,a61033a,a61037a,a61038a,a61039a,a61043a,a61044a,a61047a,a61050a,a61051a,a61052a,a61056a,a61057a,a61061a,a61062a,a61063a,a61067a,a61068a,a61071a,a61074a,a61075a,a61076a,a61080a,a61081a,a61085a,a61086a,a61087a,a61091a,a61092a,a61095a,a61098a,a61099a,a61100a,a61104a,a61105a,a61109a,a61110a,a61111a,a61115a,a61116a,a61119a,a61122a,a61123a,a61124a,a61128a,a61129a,a61133a,a61134a,a61135a,a61139a,a61140a,a61143a,a61146a,a61147a,a61148a,a61152a,a61153a,a61157a,a61158a,a61159a,a61163a,a61164a,a61167a,a61170a,a61171a,a61172a,a61176a,a61177a,a61181a,a61182a,a61183a,a61187a,a61188a,a61191a,a61194a,a61195a,a61196a,a61200a,a61201a,a61205a,a61206a,a61207a,a61211a,a61212a,a61215a,a61218a,a61219a,a61220a,a61224a,a61225a,a61229a,a61230a,a61231a,a61235a,a61236a,a61239a,a61242a,a61243a,a61244a,a61248a,a61249a,a61253a,a61254a,a61255a,a61259a,a61260a,a61263a,a61266a,a61267a,a61268a,a61272a,a61273a,a61277a,a61278a,a61279a,a61283a,a61284a,a61287a,a61290a,a61291a,a61292a,a61296a,a61297a,a61301a,a61302a,a61303a,a61307a,a61308a,a61311a,a61314a,a61315a,a61316a,a61320a,a61321a,a61325a,a61326a,a61327a,a61331a,a61332a,a61335a,a61338a,a61339a,a61340a,a61344a,a61345a,a61349a,a61350a,a61351a,a61355a,a61356a,a61359a,a61362a,a61363a,a61364a,a61368a,a61369a,a61373a,a61374a,a61375a,a61379a,a61380a,a61383a,a61386a,a61387a,a61388a,a61392a,a61393a,a61397a,a61398a,a61399a,a61403a,a61404a,a61407a,a61410a,a61411a,a61412a,a61416a,a61417a,a61421a,a61422a,a61423a,a61427a,a61428a,a61431a,a61434a,a61435a,a61436a,a61440a,a61441a,a61445a,a61446a,a61447a,a61451a,a61452a,a61455a,a61458a,a61459a,a61460a,a61464a,a61465a,a61469a,a61470a,a61471a,a61475a,a61476a,a61479a,a61482a,a61483a,a61484a,a61488a,a61489a,a61493a,a61494a,a61495a,a61499a,a61500a,a61503a,a61506a,a61507a,a61508a,a61512a,a61513a,a61517a,a61518a,a61519a,a61523a,a61524a,a61527a,a61530a,a61531a,a61532a,a61536a,a61537a,a61541a,a61542a,a61543a,a61547a,a61548a,a61551a,a61554a,a61555a,a61556a,a61560a,a61561a,a61565a,a61566a,a61567a,a61571a,a61572a,a61575a,a61578a,a61579a,a61580a,a61584a,a61585a,a61589a,a61590a,a61591a,a61595a,a61596a,a61599a,a61602a,a61603a,a61604a,a61608a,a61609a,a61613a,a61614a,a61615a,a61619a,a61620a,a61623a,a61626a,a61627a,a61628a,a61632a,a61633a,a61637a,a61638a,a61639a,a61643a,a61644a,a61647a,a61650a,a61651a,a61652a,a61656a,a61657a,a61661a,a61662a,a61663a,a61667a,a61668a,a61671a,a61674a,a61675a,a61676a,a61680a,a61681a,a61685a,a61686a,a61687a,a61691a,a61692a,a61695a,a61698a,a61699a,a61700a,a61704a,a61705a,a61709a,a61710a,a61711a,a61715a,a61716a,a61719a,a61722a,a61723a,a61724a,a61728a,a61729a,a61733a,a61734a,a61735a,a61739a,a61740a,a61743a,a61746a,a61747a,a61748a,a61752a,a61753a,a61757a,a61758a,a61759a,a61763a,a61764a,a61767a,a61770a,a61771a,a61772a,a61776a,a61777a,a61781a,a61782a,a61783a,a61787a,a61788a,a61791a,a61794a,a61795a,a61796a,a61800a,a61801a,a61805a,a61806a,a61807a,a61811a,a61812a,a61815a,a61818a,a61819a,a61820a,a61824a,a61825a,a61829a,a61830a,a61831a,a61835a,a61836a,a61839a,a61842a,a61843a,a61844a,a61848a,a61849a,a61853a,a61854a,a61855a,a61859a,a61860a,a61863a,a61866a,a61867a,a61868a,a61872a,a61873a,a61877a,a61878a,a61879a,a61883a,a61884a,a61887a,a61890a,a61891a,a61892a,a61896a,a61897a,a61901a,a61902a,a61903a,a61907a,a61908a,a61911a,a61914a,a61915a,a61916a,a61920a,a61921a,a61925a,a61926a,a61927a,a61931a,a61932a,a61935a,a61938a,a61939a,a61940a,a61944a,a61945a,a61949a,a61950a,a61951a,a61955a,a61956a,a61959a,a61962a,a61963a,a61964a,a61968a,a61969a,a61973a,a61974a,a61975a,a61979a,a61980a,a61983a,a61986a,a61987a,a61988a,a61992a,a61993a,a61997a,a61998a,a61999a,a62003a,a62004a,a62007a,a62010a,a62011a,a62012a,a62016a,a62017a,a62021a,a62022a,a62023a,a62027a,a62028a,a62031a,a62034a,a62035a,a62036a,a62040a,a62041a,a62045a,a62046a,a62047a,a62051a,a62052a,a62055a,a62058a,a62059a,a62060a,a62064a,a62065a,a62069a,a62070a,a62071a,a62075a,a62076a,a62079a,a62082a,a62083a,a62084a,a62088a,a62089a,a62093a,a62094a,a62095a,a62099a,a62100a,a62103a,a62106a,a62107a,a62108a,a62112a,a62113a,a62117a,a62118a,a62119a,a62123a,a62124a,a62127a,a62130a,a62131a,a62132a,a62136a,a62137a,a62141a,a62142a,a62143a,a62147a,a62148a,a62151a,a62154a,a62155a,a62156a,a62160a,a62161a,a62165a,a62166a,a62167a,a62171a,a62172a,a62175a,a62178a,a62179a,a62180a,a62184a,a62185a,a62189a,a62190a,a62191a,a62195a,a62196a,a62199a,a62202a,a62203a,a62204a,a62208a,a62209a,a62213a,a62214a,a62215a,a62219a,a62220a,a62223a,a62226a,a62227a,a62228a,a62232a,a62233a,a62237a,a62238a,a62239a,a62243a,a62244a,a62247a,a62250a,a62251a,a62252a,a62256a,a62257a,a62261a,a62262a,a62263a,a62267a,a62268a,a62271a,a62274a,a62275a,a62276a,a62280a,a62281a,a62285a,a62286a,a62287a,a62291a,a62292a,a62295a,a62298a,a62299a,a62300a,a62304a,a62305a,a62309a,a62310a,a62311a,a62315a,a62316a,a62319a,a62322a,a62323a,a62324a,a62328a,a62329a,a62333a,a62334a,a62335a,a62339a,a62340a,a62343a,a62346a,a62347a,a62348a,a62352a,a62353a,a62357a,a62358a,a62359a,a62363a,a62364a,a62367a,a62370a,a62371a,a62372a,a62376a,a62377a,a62381a,a62382a,a62383a,a62387a,a62388a,a62391a,a62394a,a62395a,a62396a,a62400a,a62401a,a62405a,a62406a,a62407a,a62411a,a62412a,a62415a,a62418a,a62419a,a62420a,a62424a,a62425a,a62429a,a62430a,a62431a,a62435a,a62436a,a62439a,a62442a,a62443a,a62444a,a62448a,a62449a,a62453a,a62454a,a62455a,a62459a,a62460a,a62463a,a62466a,a62467a,a62468a,a62472a,a62473a,a62477a,a62478a,a62479a,a62483a,a62484a,a62487a,a62490a,a62491a,a62492a,a62496a,a62497a,a62501a,a62502a,a62503a,a62507a,a62508a,a62511a,a62514a,a62515a,a62516a,a62520a,a62521a,a62525a,a62526a,a62527a,a62531a,a62532a,a62535a,a62538a,a62539a,a62540a,a62544a,a62545a,a62549a,a62550a,a62551a,a62555a,a62556a,a62559a,a62562a,a62563a,a62564a,a62568a,a62569a,a62573a,a62574a,a62575a,a62579a,a62580a,a62583a,a62586a,a62587a,a62588a,a62592a,a62593a,a62597a,a62598a,a62599a,a62603a,a62604a,a62607a,a62610a,a62611a,a62612a,a62616a,a62617a,a62621a,a62622a,a62623a,a62627a,a62628a,a62631a,a62634a,a62635a,a62636a,a62640a,a62641a,a62645a,a62646a,a62647a,a62651a,a62652a,a62655a,a62658a,a62659a,a62660a,a62664a,a62665a,a62669a,a62670a,a62671a,a62675a,a62676a,a62679a,a62682a,a62683a,a62684a,a62688a,a62689a,a62693a,a62694a,a62695a,a62699a,a62700a,a62703a,a62706a,a62707a,a62708a,a62712a,a62713a,a62717a,a62718a,a62719a,a62723a,a62724a,a62727a,a62730a,a62731a,a62732a,a62736a,a62737a,a62741a,a62742a,a62743a,a62747a,a62748a,a62751a,a62754a,a62755a,a62756a,a62760a,a62761a,a62765a,a62766a,a62767a,a62771a,a62772a,a62775a,a62778a,a62779a,a62780a,a62784a,a62785a,a62789a,a62790a,a62791a,a62795a,a62796a,a62799a,a62802a,a62803a,a62804a,a62808a,a62809a,a62813a,a62814a,a62815a,a62819a,a62820a,a62823a,a62826a,a62827a,a62828a,a62832a,a62833a,a62837a,a62838a,a62839a,a62843a,a62844a,a62847a,a62850a,a62851a,a62852a,a62856a,a62857a,a62861a,a62862a,a62863a,a62867a,a62868a,a62871a,a62874a,a62875a,a62876a,a62880a,a62881a,a62885a,a62886a,a62887a,a62891a,a62892a,a62895a,a62898a,a62899a,a62900a,a62904a,a62905a,a62909a,a62910a,a62911a,a62915a,a62916a,a62919a,a62922a,a62923a,a62924a,a62928a,a62929a,a62933a,a62934a,a62935a,a62939a,a62940a,a62943a,a62946a,a62947a,a62948a,a62952a,a62953a,a62957a,a62958a,a62959a,a62963a,a62964a,a62967a,a62970a,a62971a,a62972a,a62976a,a62977a,a62981a,a62982a,a62983a,a62987a,a62988a,a62991a,a62994a,a62995a,a62996a,a63000a,a63001a,a63005a,a63006a,a63007a,a63011a,a63012a,a63015a,a63018a,a63019a,a63020a,a63024a,a63025a,a63029a,a63030a,a63031a,a63035a,a63036a,a63039a,a63042a,a63043a,a63044a,a63048a,a63049a,a63053a,a63054a,a63055a,a63059a,a63060a,a63063a,a63066a,a63067a,a63068a,a63072a,a63073a,a63077a,a63078a,a63079a,a63083a,a63084a,a63087a,a63090a,a63091a,a63092a,a63096a,a63097a,a63101a,a63102a,a63103a,a63107a,a63108a,a63111a,a63114a,a63115a,a63116a,a63120a,a63121a,a63125a,a63126a,a63127a,a63131a,a63132a,a63135a,a63138a,a63139a,a63140a,a63144a,a63145a,a63149a,a63150a,a63151a,a63155a,a63156a,a63159a,a63162a,a63163a,a63164a,a63168a,a63169a,a63173a,a63174a,a63175a,a63179a,a63180a,a63183a,a63186a,a63187a,a63188a,a63192a,a63193a,a63197a,a63198a,a63199a,a63203a,a63204a,a63207a,a63210a,a63211a,a63212a,a63216a,a63217a,a63221a,a63222a,a63223a,a63227a,a63228a,a63231a,a63234a,a63235a,a63236a,a63240a,a63241a,a63245a,a63246a,a63247a,a63251a,a63252a,a63255a,a63258a,a63259a,a63260a,a63264a,a63265a,a63269a,a63270a,a63271a,a63275a,a63276a,a63279a,a63282a,a63283a,a63284a,a63288a,a63289a,a63293a,a63294a,a63295a,a63299a,a63300a,a63303a,a63306a,a63307a,a63308a,a63312a,a63313a,a63317a,a63318a,a63319a,a63323a,a63324a,a63327a,a63330a,a63331a,a63332a,a63336a,a63337a,a63341a,a63342a,a63343a,a63347a,a63348a,a63351a,a63354a,a63355a,a63356a,a63360a,a63361a,a63365a,a63366a,a63367a,a63371a,a63372a,a63375a,a63378a,a63379a,a63380a,a63384a,a63385a,a63389a,a63390a,a63391a,a63395a,a63396a,a63399a,a63402a,a63403a,a63404a,a63408a,a63409a,a63413a,a63414a,a63415a,a63419a,a63420a,a63423a,a63426a,a63427a,a63428a,a63432a,a63433a,a63437a,a63438a,a63439a,a63443a,a63444a,a63447a,a63450a,a63451a,a63452a,a63456a,a63457a,a63461a,a63462a,a63463a,a63467a,a63468a,a63471a,a63474a,a63475a,a63476a,a63480a,a63481a,a63485a,a63486a,a63487a,a63491a,a63492a,a63495a,a63498a,a63499a,a63500a,a63504a,a63505a,a63509a,a63510a,a63511a,a63515a,a63516a,a63519a,a63522a,a63523a,a63524a,a63528a,a63529a,a63533a,a63534a,a63535a,a63539a,a63540a,a63543a,a63546a,a63547a,a63548a,a63552a,a63553a,a63557a,a63558a,a63559a,a63563a,a63564a,a63567a,a63570a,a63571a,a63572a,a63576a,a63577a,a63581a,a63582a,a63583a,a63587a,a63588a,a63591a,a63594a,a63595a,a63596a,a63600a,a63601a,a63605a,a63606a,a63607a,a63611a,a63612a,a63615a,a63618a,a63619a,a63620a,a63624a,a63625a,a63629a,a63630a,a63631a,a63635a,a63636a,a63639a,a63642a,a63643a,a63644a,a63648a,a63649a,a63653a,a63654a,a63655a,a63659a,a63660a,a63663a,a63666a,a63667a,a63668a,a63672a,a63673a,a63677a,a63678a,a63679a,a63683a,a63684a,a63687a,a63690a,a63691a,a63692a,a63696a,a63697a,a63701a,a63702a,a63703a,a63707a,a63708a,a63711a,a63714a,a63715a,a63716a,a63720a,a63721a,a63725a,a63726a,a63727a,a63731a,a63732a,a63735a,a63738a,a63739a,a63740a,a63744a,a63745a,a63749a,a63750a,a63751a,a63755a,a63756a,a63759a,a63762a,a63763a,a63764a,a63768a,a63769a,a63773a,a63774a,a63775a,a63779a,a63780a,a63783a,a63786a,a63787a,a63788a,a63792a,a63793a,a63797a,a63798a,a63799a,a63803a,a63804a,a63807a,a63810a,a63811a,a63812a,a63816a,a63817a,a63821a,a63822a,a63823a,a63827a,a63828a,a63831a,a63834a,a63835a,a63836a,a63840a,a63841a,a63845a,a63846a,a63847a,a63851a,a63852a,a63855a,a63858a,a63859a,a63860a,a63864a,a63865a,a63869a,a63870a,a63871a,a63875a,a63876a,a63879a,a63882a,a63883a,a63884a,a63888a,a63889a,a63893a,a63894a,a63895a,a63899a,a63900a,a63903a,a63906a,a63907a,a63908a,a63912a,a63913a,a63917a,a63918a,a63919a,a63923a,a63924a,a63927a,a63930a,a63931a,a63932a,a63936a,a63937a,a63941a,a63942a,a63943a,a63947a,a63948a,a63951a,a63954a,a63955a,a63956a,a63960a,a63961a,a63965a,a63966a,a63967a,a63971a,a63972a,a63975a,a63978a,a63979a,a63980a,a63984a,a63985a,a63989a,a63990a,a63991a,a63995a,a63996a,a63999a,a64002a,a64003a,a64004a,a64008a,a64009a,a64013a,a64014a,a64015a,a64019a,a64020a,a64023a,a64026a,a64027a,a64028a,a64032a,a64033a,a64037a,a64038a,a64039a,a64043a,a64044a,a64047a,a64050a,a64051a,a64052a,a64056a,a64057a,a64061a,a64062a,a64063a,a64067a,a64068a,a64071a,a64074a,a64075a,a64076a,a64080a,a64081a,a64085a,a64086a,a64087a,a64091a,a64092a,a64095a,a64098a,a64099a,a64100a,a64104a,a64105a,a64109a,a64110a,a64111a,a64115a,a64116a,a64119a,a64122a,a64123a,a64124a,a64128a,a64129a,a64133a,a64134a,a64135a,a64139a,a64140a,a64143a,a64146a,a64147a,a64148a,a64152a,a64153a,a64157a,a64158a,a64159a,a64163a,a64164a,a64167a,a64170a,a64171a,a64172a,a64176a,a64177a,a64181a,a64182a,a64183a,a64187a,a64188a,a64191a,a64194a,a64195a,a64196a,a64200a,a64201a,a64205a,a64206a,a64207a,a64211a,a64212a,a64215a,a64218a,a64219a,a64220a,a64224a,a64225a,a64229a,a64230a,a64231a,a64235a,a64236a,a64239a,a64242a,a64243a,a64244a,a64248a,a64249a,a64253a,a64254a,a64255a,a64259a,a64260a,a64263a,a64266a,a64267a,a64268a,a64272a,a64273a,a64277a,a64278a,a64279a,a64283a,a64284a,a64287a,a64290a,a64291a,a64292a,a64296a,a64297a,a64301a,a64302a,a64303a,a64307a,a64308a,a64311a,a64314a,a64315a,a64316a,a64320a,a64321a,a64325a,a64326a,a64327a,a64331a,a64332a,a64335a,a64338a,a64339a,a64340a,a64344a,a64345a,a64349a,a64350a,a64351a,a64355a,a64356a,a64359a,a64362a,a64363a,a64364a,a64368a,a64369a,a64373a,a64374a,a64375a,a64379a,a64380a,a64383a,a64386a,a64387a,a64388a,a64392a,a64393a,a64397a,a64398a,a64399a,a64403a,a64404a,a64407a,a64410a,a64411a,a64412a,a64416a,a64417a,a64421a,a64422a,a64423a,a64427a,a64428a,a64431a,a64434a,a64435a,a64436a,a64440a,a64441a,a64445a,a64446a,a64447a,a64451a,a64452a,a64455a,a64458a,a64459a,a64460a,a64464a,a64465a,a64469a,a64470a,a64471a,a64475a,a64476a,a64479a,a64482a,a64483a,a64484a,a64488a,a64489a,a64493a,a64494a,a64495a,a64499a,a64500a,a64503a,a64506a,a64507a,a64508a,a64512a,a64513a,a64517a,a64518a,a64519a,a64523a,a64524a,a64527a,a64530a,a64531a,a64532a,a64536a,a64537a,a64541a,a64542a,a64543a,a64547a,a64548a,a64551a,a64554a,a64555a,a64556a,a64560a,a64561a,a64565a,a64566a,a64567a,a64571a,a64572a,a64575a,a64578a,a64579a,a64580a,a64584a,a64585a,a64589a,a64590a,a64591a,a64595a,a64596a,a64599a,a64602a,a64603a,a64604a,a64608a,a64609a,a64613a,a64614a,a64615a,a64619a,a64620a,a64623a,a64626a,a64627a,a64628a,a64632a,a64633a,a64637a,a64638a,a64639a,a64643a,a64644a,a64647a,a64650a,a64651a,a64652a,a64656a,a64657a,a64661a,a64662a,a64663a,a64667a,a64668a,a64671a,a64674a,a64675a,a64676a,a64680a,a64681a,a64685a,a64686a,a64687a,a64691a,a64692a,a64695a,a64698a,a64699a,a64700a,a64704a,a64705a,a64709a,a64710a,a64711a,a64715a,a64716a,a64719a,a64722a,a64723a,a64724a,a64728a,a64729a,a64733a,a64734a,a64735a,a64739a,a64740a,a64743a,a64746a,a64747a,a64748a,a64752a,a64753a,a64757a,a64758a,a64759a,a64763a,a64764a,a64767a,a64770a,a64771a,a64772a,a64776a,a64777a,a64781a,a64782a,a64783a,a64787a,a64788a,a64791a,a64794a,a64795a,a64796a,a64800a,a64801a,a64805a,a64806a,a64807a,a64811a,a64812a,a64815a,a64818a,a64819a,a64820a,a64824a,a64825a,a64829a,a64830a,a64831a,a64835a,a64836a,a64839a,a64842a,a64843a,a64844a,a64848a,a64849a,a64853a,a64854a,a64855a,a64859a,a64860a,a64863a,a64866a,a64867a,a64868a,a64872a,a64873a,a64877a,a64878a,a64879a,a64883a,a64884a,a64887a,a64890a,a64891a,a64892a,a64896a,a64897a,a64901a,a64902a,a64903a,a64907a,a64908a,a64911a,a64914a,a64915a,a64916a,a64920a,a64921a,a64925a,a64926a,a64927a,a64931a,a64932a,a64935a,a64938a,a64939a,a64940a,a64944a,a64945a,a64949a,a64950a,a64951a,a64955a,a64956a,a64959a,a64962a,a64963a,a64964a,a64968a,a64969a,a64973a,a64974a,a64975a,a64979a,a64980a,a64983a,a64986a,a64987a,a64988a,a64992a,a64993a,a64997a,a64998a,a64999a,a65003a,a65004a,a65007a,a65010a,a65011a,a65012a,a65016a,a65017a,a65021a,a65022a,a65023a,a65027a,a65028a,a65031a,a65034a,a65035a,a65036a,a65040a,a65041a,a65045a,a65046a,a65047a,a65051a,a65052a,a65055a,a65058a,a65059a,a65060a,a65064a,a65065a,a65069a,a65070a,a65071a,a65075a,a65076a,a65079a,a65082a,a65083a,a65084a,a65088a,a65089a,a65093a,a65094a,a65095a,a65099a,a65100a,a65103a,a65106a,a65107a,a65108a,a65112a,a65113a,a65116a,a65119a,a65120a,a65121a,a65125a,a65126a,a65129a,a65132a,a65133a,a65134a,a65138a,a65139a,a65142a,a65145a,a65146a,a65147a,a65151a,a65152a,a65155a,a65158a,a65159a,a65160a,a65164a,a65165a,a65168a,a65171a,a65172a,a65173a,a65177a,a65178a,a65181a,a65184a,a65185a,a65186a,a65190a,a65191a,a65194a,a65197a,a65198a,a65199a,a65203a,a65204a,a65207a,a65210a,a65211a,a65212a,a65216a,a65217a,a65220a,a65223a,a65224a,a65225a,a65229a,a65230a,a65233a,a65236a,a65237a,a65238a,a65242a,a65243a,a65246a,a65249a,a65250a,a65251a,a65255a,a65256a,a65259a,a65262a,a65263a,a65264a,a65268a,a65269a,a65272a,a65275a,a65276a,a65277a,a65281a,a65282a,a65285a,a65288a,a65289a,a65290a,a65294a,a65295a,a65298a,a65301a,a65302a,a65303a,a65307a,a65308a,a65311a,a65314a,a65315a,a65316a,a65320a,a65321a,a65324a,a65327a,a65328a,a65329a,a65333a,a65334a,a65337a,a65340a,a65341a,a65342a,a65346a,a65347a,a65350a,a65353a,a65354a,a65355a,a65359a,a65360a,a65363a,a65366a,a65367a,a65368a,a65372a,a65373a,a65376a,a65379a,a65380a,a65381a,a65385a,a65386a,a65389a,a65392a,a65393a,a65394a,a65398a,a65399a,a65402a,a65405a,a65406a,a65407a,a65411a,a65412a,a65415a,a65418a,a65419a,a65420a,a65424a,a65425a,a65428a,a65431a,a65432a,a65433a,a65437a,a65438a,a65441a,a65444a,a65445a,a65446a,a65450a,a65451a,a65454a,a65457a,a65458a,a65459a,a65463a,a65464a,a65467a,a65470a,a65471a,a65472a,a65476a,a65477a,a65480a,a65483a,a65484a,a65485a,a65489a,a65490a,a65493a,a65496a,a65497a,a65498a,a65502a,a65503a,a65506a,a65509a,a65510a,a65511a,a65515a,a65516a,a65519a,a65522a,a65523a,a65524a,a65528a,a65529a,a65532a,a65535a,a65536a,a65537a,a65541a,a65542a,a65545a,a65548a,a65549a,a65550a,a65554a,a65555a,a65558a,a65561a,a65562a,a65563a,a65567a,a65568a,a65571a,a65574a,a65575a,a65576a,a65580a,a65581a,a65584a,a65587a,a65588a,a65589a,a65593a,a65594a,a65597a,a65600a,a65601a,a65602a,a65606a,a65607a,a65610a,a65613a,a65614a,a65615a,a65619a,a65620a,a65623a,a65626a,a65627a,a65628a,a65632a,a65633a,a65636a,a65639a,a65640a,a65641a,a65645a,a65646a,a65649a,a65652a,a65653a,a65654a,a65658a,a65659a,a65662a,a65665a,a65666a,a65667a,a65671a,a65672a,a65675a,a65678a,a65679a,a65680a,a65684a,a65685a,a65688a,a65691a,a65692a,a65693a,a65697a,a65698a,a65701a,a65704a,a65705a,a65706a,a65710a,a65711a,a65714a,a65717a,a65718a,a65719a,a65723a,a65724a,a65727a,a65730a,a65731a,a65732a,a65736a,a65737a,a65740a,a65743a,a65744a,a65745a,a65749a,a65750a,a65753a,a65756a,a65757a,a65758a,a65762a,a65763a,a65766a,a65769a,a65770a,a65771a,a65775a,a65776a,a65779a,a65782a,a65783a,a65784a,a65788a,a65789a,a65792a,a65795a,a65796a,a65797a,a65801a,a65802a,a65805a,a65808a,a65809a,a65810a,a65814a,a65815a,a65818a,a65821a,a65822a,a65823a,a65827a,a65828a,a65831a,a65834a,a65835a,a65836a,a65840a,a65841a,a65844a,a65847a,a65848a,a65849a,a65853a,a65854a,a65857a,a65860a,a65861a,a65862a,a65866a,a65867a,a65870a,a65873a,a65874a,a65875a,a65879a,a65880a,a65883a,a65886a,a65887a,a65888a,a65892a,a65893a,a65896a,a65899a,a65900a,a65901a,a65905a,a65906a,a65909a,a65912a,a65913a,a65914a,a65918a,a65919a,a65922a,a65925a,a65926a,a65927a,a65931a,a65932a,a65935a,a65938a,a65939a,a65940a,a65944a,a65945a,a65948a,a65951a,a65952a,a65953a,a65957a,a65958a,a65961a,a65964a,a65965a,a65966a,a65970a,a65971a,a65974a,a65977a,a65978a,a65979a,a65983a,a65984a,a65987a,a65990a,a65991a,a65992a,a65996a,a65997a,a66000a,a66003a,a66004a,a66005a,a66009a,a66010a,a66013a,a66016a,a66017a,a66018a,a66022a,a66023a,a66026a,a66029a,a66030a,a66031a,a66035a,a66036a,a66039a,a66042a,a66043a,a66044a,a66048a,a66049a,a66052a,a66055a,a66056a,a66057a,a66061a,a66062a,a66065a,a66068a,a66069a,a66070a,a66074a,a66075a,a66078a,a66081a,a66082a,a66083a,a66087a,a66088a,a66091a,a66094a,a66095a,a66096a,a66100a,a66101a,a66104a,a66107a,a66108a,a66109a,a66113a,a66114a,a66117a,a66120a,a66121a,a66122a,a66126a,a66127a,a66130a,a66133a,a66134a,a66135a,a66139a,a66140a,a66143a,a66146a,a66147a,a66148a,a66152a,a66153a,a66156a,a66159a,a66160a,a66161a,a66165a,a66166a,a66169a,a66172a,a66173a,a66174a,a66178a,a66179a,a66182a,a66185a,a66186a,a66187a,a66191a,a66192a,a66195a,a66198a,a66199a,a66200a,a66204a,a66205a,a66208a,a66211a,a66212a,a66213a,a66217a,a66218a,a66221a,a66224a,a66225a,a66226a,a66230a,a66231a,a66234a,a66237a,a66238a,a66239a,a66243a,a66244a,a66247a,a66250a,a66251a,a66252a,a66256a,a66257a,a66260a,a66263a,a66264a,a66265a,a66269a,a66270a,a66273a,a66276a,a66277a,a66278a,a66282a,a66283a,a66286a,a66289a,a66290a,a66291a,a66295a,a66296a,a66299a,a66302a,a66303a,a66304a,a66308a,a66309a,a66312a,a66315a,a66316a,a66317a,a66321a,a66322a,a66325a,a66328a,a66329a,a66330a,a66334a,a66335a,a66338a,a66341a,a66342a,a66343a,a66347a,a66348a,a66351a,a66354a,a66355a,a66356a,a66360a,a66361a,a66364a,a66367a,a66368a,a66369a,a66373a,a66374a,a66377a,a66380a,a66381a,a66382a,a66386a,a66387a,a66390a,a66393a,a66394a,a66395a,a66399a,a66400a,a66403a,a66406a,a66407a,a66408a,a66412a,a66413a,a66416a,a66419a,a66420a,a66421a,a66425a,a66426a,a66429a,a66432a,a66433a,a66434a,a66438a,a66439a,a66442a,a66445a,a66446a,a66447a,a66451a,a66452a,a66455a,a66458a,a66459a,a66460a,a66464a,a66465a,a66468a,a66471a,a66472a,a66473a,a66477a,a66478a,a66481a,a66484a,a66485a,a66486a,a66490a,a66491a,a66494a,a66497a,a66498a,a66499a,a66503a,a66504a,a66507a,a66510a,a66511a,a66512a,a66516a,a66517a,a66520a,a66523a,a66524a,a66525a,a66529a,a66530a,a66533a,a66536a,a66537a,a66538a,a66542a,a66543a,a66546a,a66549a,a66550a,a66551a,a66555a,a66556a,a66559a,a66562a,a66563a,a66564a,a66568a,a66569a,a66572a,a66575a,a66576a,a66577a,a66581a,a66582a,a66585a,a66588a,a66589a,a66590a,a66594a,a66595a,a66598a,a66601a,a66602a,a66603a,a66607a,a66608a,a66611a,a66614a,a66615a,a66616a,a66620a,a66621a,a66624a,a66627a,a66628a,a66629a,a66633a,a66634a,a66637a,a66640a,a66641a,a66642a,a66646a,a66647a,a66650a,a66653a,a66654a,a66655a,a66659a,a66660a,a66663a,a66666a,a66667a,a66668a,a66672a,a66673a,a66676a,a66679a,a66680a,a66681a,a66685a,a66686a,a66689a,a66692a,a66693a,a66694a,a66698a,a66699a,a66702a,a66705a,a66706a,a66707a,a66711a,a66712a,a66715a,a66718a,a66719a,a66720a,a66724a,a66725a,a66728a,a66731a,a66732a,a66733a,a66737a,a66738a,a66741a,a66744a,a66745a,a66746a,a66750a,a66751a,a66754a,a66757a,a66758a,a66759a,a66763a,a66764a,a66767a,a66770a,a66771a,a66772a,a66776a,a66777a,a66780a,a66783a,a66784a,a66785a,a66789a,a66790a,a66793a,a66796a,a66797a,a66798a,a66802a,a66803a,a66806a,a66809a,a66810a,a66811a,a66815a,a66816a,a66819a,a66822a,a66823a,a66824a,a66828a,a66829a,a66832a,a66835a,a66836a,a66837a,a66841a,a66842a,a66845a,a66848a,a66849a,a66850a,a66854a,a66855a,a66858a,a66861a,a66862a,a66863a,a66867a,a66868a,a66871a,a66874a,a66875a,a66876a,a66880a,a66881a,a66884a,a66887a,a66888a,a66889a,a66893a,a66894a,a66897a,a66900a,a66901a,a66902a,a66906a,a66907a,a66910a,a66913a,a66914a,a66915a,a66919a,a66920a,a66923a,a66926a,a66927a,a66928a,a66932a,a66933a,a66936a,a66939a,a66940a,a66941a,a66945a,a66946a,a66949a,a66952a,a66953a,a66954a,a66958a,a66959a,a66962a,a66965a,a66966a,a66967a,a66971a,a66972a,a66975a,a66978a,a66979a,a66980a,a66984a,a66985a,a66988a,a66991a,a66992a,a66993a,a66997a,a66998a,a67001a,a67004a,a67005a,a67006a,a67010a,a67011a,a67014a,a67017a,a67018a,a67019a,a67023a,a67024a,a67027a,a67030a,a67031a,a67032a,a67036a,a67037a,a67040a,a67043a,a67044a,a67045a,a67049a,a67050a,a67053a,a67056a,a67057a,a67058a,a67062a,a67063a,a67066a,a67069a,a67070a,a67071a,a67075a,a67076a,a67079a,a67082a,a67083a,a67084a,a67088a,a67089a,a67092a,a67095a,a67096a,a67097a,a67101a,a67102a,a67105a,a67108a,a67109a,a67110a,a67114a,a67115a,a67118a,a67121a,a67122a,a67123a,a67127a,a67128a,a67131a,a67134a,a67135a,a67136a,a67140a,a67141a,a67144a,a67147a,a67148a,a67149a,a67153a,a67154a,a67157a,a67160a,a67161a,a67162a,a67166a,a67167a,a67170a,a67173a,a67174a,a67175a,a67179a,a67180a,a67183a,a67186a,a67187a,a67188a,a67192a,a67193a,a67196a,a67199a,a67200a,a67201a,a67205a,a67206a,a67209a,a67212a,a67213a,a67214a,a67218a,a67219a,a67222a,a67225a,a67226a,a67227a,a67231a,a67232a,a67235a,a67238a,a67239a,a67240a,a67244a,a67245a,a67248a,a67251a,a67252a,a67253a,a67257a,a67258a,a67261a,a67264a,a67265a,a67266a,a67270a,a67271a,a67274a,a67277a,a67278a,a67279a,a67283a,a67284a,a67287a,a67290a,a67291a,a67292a,a67296a,a67297a,a67300a,a67303a,a67304a,a67305a,a67309a,a67310a,a67313a,a67316a,a67317a,a67318a,a67322a,a67323a,a67326a,a67329a,a67330a,a67331a,a67335a,a67336a,a67339a,a67342a,a67343a,a67344a,a67348a,a67349a,a67352a,a67355a,a67356a,a67357a,a67361a,a67362a,a67365a,a67368a,a67369a,a67370a,a67374a,a67375a,a67378a,a67381a,a67382a,a67383a,a67387a,a67388a,a67391a,a67394a,a67395a,a67396a,a67400a,a67401a,a67404a,a67407a,a67408a,a67409a,a67413a,a67414a,a67417a,a67420a,a67421a,a67422a,a67426a,a67427a,a67430a,a67433a,a67434a,a67435a,a67439a,a67440a,a67443a,a67446a,a67447a,a67448a,a67452a,a67453a,a67456a,a67459a,a67460a,a67461a,a67465a,a67466a,a67469a,a67472a,a67473a,a67474a,a67478a,a67479a,a67482a,a67485a,a67486a,a67487a,a67491a,a67492a,a67495a,a67498a,a67499a,a67500a,a67504a,a67505a,a67508a,a67511a,a67512a,a67513a,a67517a,a67518a,a67521a,a67524a,a67525a,a67526a,a67530a,a67531a,a67534a,a67537a,a67538a,a67539a,a67543a,a67544a,a67547a,a67550a,a67551a,a67552a,a67556a,a67557a,a67560a,a67563a,a67564a,a67565a,a67569a,a67570a,a67573a,a67576a,a67577a,a67578a,a67582a,a67583a,a67586a,a67589a,a67590a,a67591a,a67595a,a67596a,a67599a,a67602a,a67603a,a67604a,a67608a,a67609a,a67612a,a67615a,a67616a,a67617a,a67621a,a67622a,a67625a,a67628a,a67629a,a67630a,a67634a,a67635a,a67638a,a67641a,a67642a,a67643a,a67647a,a67648a,a67651a,a67654a,a67655a,a67656a,a67660a,a67661a,a67664a,a67667a,a67668a,a67669a,a67673a,a67674a,a67677a,a67680a,a67681a,a67682a,a67686a,a67687a,a67690a,a67693a,a67694a,a67695a,a67699a,a67700a,a67703a,a67706a,a67707a,a67708a,a67712a,a67713a,a67716a,a67719a,a67720a,a67721a,a67725a,a67726a,a67729a,a67732a,a67733a,a67734a,a67738a,a67739a,a67742a,a67745a,a67746a,a67747a,a67751a,a67752a,a67755a,a67758a,a67759a,a67760a,a67764a,a67765a,a67768a,a67771a,a67772a,a67773a,a67777a,a67778a,a67781a,a67784a,a67785a,a67786a,a67790a,a67791a,a67794a,a67797a,a67798a,a67799a,a67803a,a67804a,a67807a,a67810a,a67811a,a67812a,a67816a,a67817a,a67820a,a67823a,a67824a,a67825a,a67829a,a67830a,a67833a,a67836a,a67837a,a67838a,a67842a,a67843a,a67846a,a67849a,a67850a,a67851a,a67855a,a67856a,a67859a,a67862a,a67863a,a67864a,a67868a,a67869a,a67872a,a67875a,a67876a,a67877a,a67881a,a67882a,a67885a,a67888a,a67889a,a67890a,a67894a,a67895a,a67898a,a67901a,a67902a,a67903a,a67907a,a67908a,a67911a,a67914a,a67915a,a67916a,a67920a,a67921a,a67924a,a67927a,a67928a,a67929a,a67933a,a67934a,a67937a,a67940a,a67941a,a67942a,a67946a,a67947a,a67950a,a67953a,a67954a,a67955a,a67959a,a67960a,a67963a,a67966a,a67967a,a67968a,a67972a,a67973a,a67976a,a67979a,a67980a,a67981a,a67985a,a67986a,a67989a,a67992a,a67993a,a67994a,a67998a,a67999a,a68002a,a68005a,a68006a,a68007a,a68011a,a68012a,a68015a,a68018a,a68019a,a68020a,a68024a,a68025a,a68028a,a68031a,a68032a,a68033a,a68037a,a68038a,a68041a,a68044a,a68045a,a68046a,a68050a,a68051a,a68054a,a68057a,a68058a,a68059a,a68063a,a68064a,a68067a,a68070a,a68071a,a68072a,a68076a,a68077a,a68080a,a68083a,a68084a,a68085a,a68089a,a68090a,a68093a,a68096a,a68097a,a68098a,a68102a,a68103a,a68106a,a68109a,a68110a,a68111a,a68115a,a68116a,a68119a,a68122a,a68123a,a68124a,a68128a,a68129a,a68132a,a68135a,a68136a,a68137a,a68141a,a68142a,a68145a,a68148a,a68149a,a68150a,a68154a,a68155a,a68158a,a68161a,a68162a,a68163a,a68167a,a68168a,a68171a,a68174a,a68175a,a68176a,a68180a,a68181a,a68184a,a68187a,a68188a,a68189a,a68193a,a68194a,a68197a,a68200a,a68201a,a68202a,a68206a,a68207a,a68210a,a68213a,a68214a,a68215a,a68219a,a68220a,a68223a,a68226a,a68227a,a68228a,a68232a,a68233a,a68236a,a68239a,a68240a,a68241a,a68245a,a68246a,a68249a,a68252a,a68253a,a68254a,a68258a,a68259a,a68262a,a68265a,a68266a,a68267a,a68271a,a68272a,a68275a,a68278a,a68279a,a68280a,a68284a,a68285a,a68288a,a68291a,a68292a,a68293a,a68297a,a68298a,a68301a,a68304a,a68305a,a68306a,a68310a,a68311a,a68314a,a68317a,a68318a,a68319a,a68323a,a68324a,a68327a,a68330a,a68331a,a68332a,a68336a,a68337a,a68340a,a68343a,a68344a,a68345a,a68349a,a68350a,a68353a,a68356a,a68357a,a68358a,a68362a,a68363a,a68366a,a68369a,a68370a,a68371a,a68375a,a68376a,a68379a,a68382a,a68383a,a68384a,a68388a,a68389a,a68392a,a68395a,a68396a,a68397a,a68401a,a68402a,a68405a,a68408a,a68409a,a68410a,a68414a,a68415a,a68418a,a68421a,a68422a,a68423a,a68427a,a68428a,a68431a,a68434a,a68435a,a68436a,a68440a,a68441a,a68444a,a68447a,a68448a,a68449a,a68453a,a68454a,a68457a,a68460a,a68461a,a68462a,a68466a,a68467a,a68470a,a68473a,a68474a,a68475a,a68479a,a68480a,a68483a,a68486a,a68487a,a68488a,a68492a,a68493a,a68496a,a68499a,a68500a,a68501a,a68505a,a68506a,a68509a,a68512a,a68513a,a68514a,a68518a,a68519a,a68522a,a68525a,a68526a,a68527a,a68531a,a68532a,a68535a,a68538a,a68539a,a68540a,a68544a,a68545a,a68548a,a68551a,a68552a,a68553a,a68557a,a68558a,a68561a,a68564a,a68565a,a68566a,a68570a,a68571a,a68574a,a68577a,a68578a,a68579a,a68583a,a68584a,a68587a,a68590a,a68591a,a68592a,a68596a,a68597a,a68600a,a68603a,a68604a,a68605a,a68609a,a68610a,a68613a,a68616a,a68617a,a68618a,a68622a,a68623a,a68626a,a68629a,a68630a,a68631a,a68635a,a68636a,a68639a,a68642a,a68643a,a68644a,a68648a,a68649a,a68652a,a68655a,a68656a,a68657a,a68661a,a68662a,a68665a,a68668a,a68669a,a68670a,a68674a,a68675a,a68678a,a68681a,a68682a,a68683a,a68687a,a68688a,a68691a,a68694a,a68695a,a68696a,a68700a,a68701a,a68704a,a68707a,a68708a,a68709a,a68713a,a68714a,a68717a,a68720a,a68721a,a68722a,a68726a,a68727a,a68730a,a68733a,a68734a,a68735a,a68739a,a68740a,a68743a,a68746a,a68747a,a68748a,a68752a,a68753a,a68756a,a68759a,a68760a,a68761a,a68765a,a68766a,a68769a,a68772a,a68773a,a68774a,a68778a,a68779a,a68782a,a68785a,a68786a,a68787a,a68791a,a68792a,a68795a,a68798a,a68799a,a68800a,a68804a,a68805a,a68808a,a68811a,a68812a,a68813a,a68817a,a68818a,a68821a,a68824a,a68825a,a68826a,a68830a,a68831a,a68834a,a68837a,a68838a,a68839a,a68843a,a68844a,a68847a,a68850a,a68851a,a68852a,a68856a,a68857a,a68860a,a68863a,a68864a,a68865a,a68869a,a68870a,a68873a,a68876a,a68877a,a68878a,a68882a,a68883a,a68886a,a68889a,a68890a,a68891a,a68895a,a68896a,a68899a,a68902a,a68903a,a68904a,a68908a,a68909a,a68912a,a68915a,a68916a,a68917a,a68921a,a68922a,a68925a,a68928a,a68929a,a68930a,a68934a,a68935a,a68938a,a68941a,a68942a,a68943a,a68947a,a68948a,a68951a,a68954a,a68955a,a68956a,a68960a,a68961a,a68964a,a68967a,a68968a,a68969a,a68973a,a68974a,a68977a,a68980a,a68981a,a68982a,a68986a,a68987a,a68990a,a68993a,a68994a,a68995a,a68999a,a69000a,a69003a,a69006a,a69007a,a69008a,a69012a,a69013a,a69016a,a69019a,a69020a,a69021a,a69025a,a69026a,a69029a,a69032a,a69033a,a69034a,a69038a,a69039a,a69042a,a69045a,a69046a,a69047a,a69051a,a69052a,a69055a,a69058a,a69059a,a69060a,a69064a,a69065a,a69068a,a69071a,a69072a,a69073a,a69077a,a69078a,a69081a,a69084a,a69085a,a69086a,a69090a,a69091a,a69094a,a69097a,a69098a,a69099a,a69103a,a69104a,a69107a,a69110a,a69111a,a69112a,a69116a,a69117a,a69120a,a69123a,a69124a,a69125a,a69129a,a69130a,a69133a,a69136a,a69137a,a69138a,a69142a,a69143a,a69146a,a69149a,a69150a,a69151a,a69155a,a69156a,a69159a,a69162a,a69163a,a69164a,a69168a,a69169a,a69172a,a69175a,a69176a,a69177a,a69181a,a69182a,a69185a,a69188a,a69189a,a69190a,a69194a,a69195a,a69198a,a69201a,a69202a,a69203a,a69207a,a69208a,a69211a,a69214a,a69215a,a69216a,a69220a,a69221a,a69224a,a69227a,a69228a,a69229a,a69233a,a69234a,a69237a,a69240a,a69241a,a69242a,a69246a,a69247a,a69250a,a69253a,a69254a,a69255a,a69259a,a69260a,a69263a,a69266a,a69267a,a69268a,a69272a,a69273a,a69276a,a69279a,a69280a,a69281a,a69285a,a69286a,a69289a,a69292a,a69293a,a69294a,a69298a,a69299a,a69302a,a69305a,a69306a,a69307a,a69311a,a69312a,a69315a,a69318a,a69319a,a69320a,a69324a,a69325a,a69328a,a69331a,a69332a,a69333a,a69337a,a69338a,a69341a,a69344a,a69345a,a69346a,a69350a,a69351a,a69354a,a69357a,a69358a,a69359a,a69363a,a69364a,a69367a,a69370a,a69371a,a69372a,a69376a,a69377a,a69380a,a69383a,a69384a,a69385a,a69389a,a69390a,a69393a,a69396a,a69397a,a69398a,a69402a,a69403a,a69406a,a69409a,a69410a,a69411a,a69415a,a69416a,a69419a,a69422a,a69423a,a69424a,a69428a,a69429a,a69432a,a69435a,a69436a,a69437a,a69441a,a69442a,a69445a,a69448a,a69449a,a69450a,a69454a,a69455a,a69458a,a69461a,a69462a,a69463a,a69467a,a69468a,a69471a,a69474a,a69475a,a69476a,a69480a,a69481a,a69484a,a69487a,a69488a,a69489a,a69493a,a69494a,a69497a,a69500a,a69501a,a69502a,a69506a,a69507a,a69510a,a69513a,a69514a,a69515a,a69519a,a69520a,a69523a,a69526a,a69527a,a69528a,a69532a,a69533a,a69536a,a69539a,a69540a,a69541a,a69545a,a69546a,a69549a,a69552a,a69553a,a69554a,a69558a,a69559a,a69562a,a69565a,a69566a,a69567a,a69571a,a69572a,a69575a,a69578a,a69579a,a69580a,a69584a,a69585a,a69588a,a69591a,a69592a,a69593a,a69597a,a69598a,a69601a,a69604a,a69605a,a69606a,a69610a,a69611a,a69614a,a69617a,a69618a,a69619a,a69623a,a69624a,a69627a,a69630a,a69631a,a69632a,a69636a,a69637a,a69640a,a69643a,a69644a,a69645a,a69649a,a69650a,a69653a,a69656a,a69657a,a69658a,a69662a,a69663a,a69666a,a69669a,a69670a,a69671a,a69675a,a69676a,a69679a,a69682a,a69683a,a69684a,a69688a,a69689a,a69692a,a69695a,a69696a,a69697a,a69701a,a69702a,a69705a,a69708a,a69709a,a69710a,a69714a,a69715a,a69718a,a69721a,a69722a,a69723a,a69727a,a69728a,a69731a,a69734a,a69735a,a69736a,a69740a,a69741a,a69744a,a69747a,a69748a,a69749a,a69753a,a69754a,a69757a,a69760a,a69761a,a69762a,a69766a,a69767a,a69770a,a69773a,a69774a,a69775a,a69779a,a69780a,a69783a,a69786a,a69787a,a69788a,a69792a,a69793a,a69796a,a69799a,a69800a,a69801a,a69805a,a69806a,a69809a,a69812a,a69813a,a69814a,a69818a,a69819a,a69822a,a69825a,a69826a,a69827a,a69831a,a69832a,a69835a,a69838a,a69839a,a69840a,a69844a,a69845a,a69848a,a69851a,a69852a,a69853a,a69857a,a69858a,a69861a,a69864a,a69865a,a69866a,a69870a,a69871a,a69874a,a69877a,a69878a,a69879a,a69883a,a69884a,a69887a,a69890a,a69891a,a69892a,a69896a,a69897a,a69900a,a69903a,a69904a,a69905a,a69909a,a69910a,a69913a,a69916a,a69917a,a69918a,a69922a,a69923a,a69926a,a69929a,a69930a,a69931a,a69935a,a69936a,a69939a,a69942a,a69943a,a69944a,a69948a,a69949a,a69952a,a69955a,a69956a,a69957a,a69961a,a69962a,a69965a,a69968a,a69969a,a69970a,a69974a,a69975a,a69978a,a69981a,a69982a,a69983a,a69987a,a69988a,a69991a,a69994a,a69995a,a69996a,a70000a,a70001a,a70004a,a70007a,a70008a,a70009a,a70013a,a70014a,a70017a,a70020a,a70021a,a70022a,a70026a,a70027a,a70030a,a70033a,a70034a,a70035a,a70039a,a70040a,a70043a,a70046a,a70047a,a70048a,a70052a,a70053a,a70056a,a70059a,a70060a,a70061a,a70065a,a70066a,a70069a,a70072a,a70073a,a70074a,a70078a,a70079a,a70082a,a70085a,a70086a,a70087a,a70091a,a70092a,a70095a,a70098a,a70099a,a70100a,a70104a,a70105a,a70108a,a70111a,a70112a,a70113a,a70117a,a70118a,a70121a,a70124a,a70125a,a70126a,a70130a,a70131a,a70134a,a70137a,a70138a,a70139a,a70143a,a70144a,a70147a,a70150a,a70151a,a70152a,a70156a,a70157a,a70160a,a70163a,a70164a,a70165a,a70169a,a70170a,a70173a,a70176a,a70177a,a70178a,a70182a,a70183a,a70186a,a70189a,a70190a,a70191a,a70195a,a70196a,a70199a,a70202a,a70203a,a70204a,a70208a,a70209a,a70212a,a70215a,a70216a,a70217a,a70221a,a70222a,a70225a,a70228a,a70229a,a70230a,a70234a,a70235a,a70238a,a70241a,a70242a,a70243a,a70247a,a70248a,a70251a,a70254a,a70255a,a70256a,a70260a,a70261a,a70264a,a70267a,a70268a,a70269a,a70273a,a70274a,a70277a,a70280a,a70281a,a70282a,a70286a,a70287a,a70290a,a70293a,a70294a,a70295a,a70299a,a70300a,a70303a,a70306a,a70307a,a70308a,a70312a,a70313a,a70316a,a70319a,a70320a,a70321a,a70325a,a70326a,a70329a,a70332a,a70333a,a70334a,a70338a,a70339a,a70342a,a70345a,a70346a,a70347a,a70351a,a70352a,a70355a,a70358a,a70359a,a70360a,a70364a,a70365a,a70368a,a70371a,a70372a,a70373a,a70377a,a70378a,a70381a,a70384a,a70385a,a70386a,a70390a,a70391a,a70394a,a70397a,a70398a,a70399a,a70403a,a70404a,a70407a,a70410a,a70411a,a70412a,a70416a,a70417a,a70420a,a70423a,a70424a,a70425a,a70429a,a70430a,a70433a,a70436a,a70437a,a70438a,a70442a,a70443a,a70446a,a70449a,a70450a,a70451a,a70455a,a70456a,a70459a,a70462a,a70463a,a70464a,a70468a,a70469a,a70472a,a70475a,a70476a,a70477a,a70481a,a70482a,a70485a,a70488a,a70489a,a70490a,a70494a,a70495a,a70498a,a70501a,a70502a,a70503a,a70507a,a70508a,a70511a,a70514a,a70515a,a70516a,a70520a,a70521a,a70524a,a70527a,a70528a,a70529a,a70533a,a70534a,a70537a,a70540a,a70541a,a70542a,a70546a,a70547a,a70550a,a70553a,a70554a,a70555a,a70559a,a70560a,a70563a,a70566a,a70567a,a70568a,a70572a,a70573a,a70576a,a70579a,a70580a,a70581a,a70585a,a70586a,a70589a,a70592a,a70593a,a70594a,a70598a,a70599a,a70602a,a70605a,a70606a,a70607a,a70611a,a70612a,a70615a,a70618a,a70619a,a70620a,a70624a,a70625a,a70628a,a70631a,a70632a,a70633a,a70637a,a70638a,a70641a,a70644a,a70645a,a70646a,a70650a,a70651a,a70654a,a70657a,a70658a,a70659a,a70663a,a70664a,a70667a,a70670a,a70671a,a70672a,a70676a,a70677a,a70680a,a70683a,a70684a,a70685a,a70689a,a70690a,a70693a,a70696a,a70697a,a70698a,a70702a,a70703a,a70706a,a70709a,a70710a,a70711a,a70715a,a70716a,a70719a,a70722a,a70723a,a70724a,a70728a,a70729a,a70732a,a70735a,a70736a,a70737a,a70741a,a70742a,a70745a,a70748a,a70749a,a70750a,a70754a,a70755a,a70758a,a70761a,a70762a,a70763a,a70767a,a70768a,a70771a,a70774a,a70775a,a70776a,a70780a,a70781a,a70784a,a70787a,a70788a,a70789a,a70793a,a70794a,a70797a,a70800a,a70801a,a70802a,a70806a,a70807a,a70810a,a70813a,a70814a,a70815a,a70819a,a70820a,a70823a,a70826a,a70827a,a70828a,a70832a,a70833a,a70836a,a70839a,a70840a,a70841a,a70845a,a70846a,a70849a,a70852a,a70853a,a70854a,a70858a,a70859a,a70862a,a70865a,a70866a,a70867a,a70871a,a70872a,a70875a,a70878a,a70879a,a70880a,a70884a,a70885a,a70888a,a70891a,a70892a,a70893a,a70897a,a70898a,a70901a,a70904a,a70905a,a70906a,a70910a,a70911a,a70914a,a70917a,a70918a,a70919a,a70923a,a70924a,a70927a,a70930a,a70931a,a70932a,a70936a,a70937a,a70940a,a70943a,a70944a,a70945a,a70949a,a70950a,a70953a,a70956a,a70957a,a70958a,a70962a,a70963a,a70966a,a70969a,a70970a,a70971a,a70975a,a70976a,a70979a,a70982a,a70983a,a70984a,a70988a,a70989a,a70992a,a70995a,a70996a,a70997a,a71001a,a71002a,a71005a,a71008a,a71009a,a71010a,a71014a,a71015a,a71018a,a71021a,a71022a,a71023a,a71027a,a71028a,a71031a,a71034a,a71035a,a71036a,a71040a,a71041a,a71044a,a71047a,a71048a,a71049a,a71053a,a71054a,a71057a,a71060a,a71061a,a71062a,a71066a,a71067a,a71070a,a71073a,a71074a,a71075a,a71079a,a71080a,a71083a,a71086a,a71087a,a71088a,a71092a,a71093a,a71096a,a71099a,a71100a,a71101a,a71105a,a71106a,a71109a,a71112a,a71113a,a71114a,a71118a,a71119a,a71122a,a71125a,a71126a,a71127a,a71131a,a71132a,a71135a,a71138a,a71139a,a71140a,a71144a,a71145a,a71148a,a71151a,a71152a,a71153a,a71157a,a71158a,a71161a,a71164a,a71165a,a71166a,a71170a,a71171a,a71174a,a71177a,a71178a,a71179a,a71183a,a71184a,a71187a,a71190a,a71191a,a71192a,a71196a,a71197a,a71200a,a71203a,a71204a,a71205a,a71209a,a71210a,a71213a,a71216a,a71217a,a71218a,a71222a,a71223a,a71226a,a71229a,a71230a,a71231a,a71235a,a71236a,a71239a,a71242a,a71243a,a71244a,a71248a,a71249a,a71252a,a71255a,a71256a,a71257a,a71261a,a71262a,a71265a,a71268a,a71269a,a71270a,a71274a,a71275a,a71278a,a71281a,a71282a,a71283a,a71287a,a71288a,a71291a,a71294a,a71295a,a71296a,a71300a,a71301a,a71304a,a71307a,a71308a,a71309a,a71313a,a71314a,a71317a,a71320a,a71321a,a71322a,a71326a,a71327a,a71330a,a71333a,a71334a,a71335a,a71339a,a71340a,a71343a,a71346a,a71347a,a71348a,a71352a,a71353a,a71356a,a71359a,a71360a,a71361a,a71365a,a71366a,a71369a,a71372a,a71373a,a71374a,a71378a,a71379a,a71382a,a71385a,a71386a,a71387a,a71391a,a71392a,a71395a,a71398a,a71399a,a71400a,a71404a,a71405a,a71408a,a71411a,a71412a,a71413a,a71417a,a71418a,a71421a,a71424a,a71425a,a71426a,a71430a,a71431a,a71434a,a71437a,a71438a,a71439a,a71443a,a71444a,a71447a,a71450a,a71451a,a71452a,a71456a,a71457a,a71460a,a71463a,a71464a,a71465a,a71469a,a71470a,a71473a,a71476a,a71477a,a71478a,a71482a,a71483a,a71486a,a71489a,a71490a,a71491a,a71495a,a71496a,a71499a,a71502a,a71503a,a71504a,a71508a,a71509a,a71512a,a71515a,a71516a,a71517a,a71521a,a71522a,a71525a,a71528a,a71529a,a71530a,a71534a,a71535a,a71538a,a71541a,a71542a,a71543a,a71547a,a71548a,a71551a,a71554a,a71555a,a71556a,a71560a,a71561a,a71564a,a71567a,a71568a,a71569a,a71573a,a71574a,a71577a,a71580a,a71581a,a71582a,a71586a,a71587a,a71590a,a71593a,a71594a,a71595a,a71599a,a71600a,a71603a,a71606a,a71607a,a71608a,a71612a,a71613a,a71616a,a71619a,a71620a,a71621a,a71625a,a71626a,a71629a,a71632a,a71633a,a71634a,a71638a,a71639a,a71642a,a71645a,a71646a,a71647a,a71651a,a71652a,a71655a,a71658a,a71659a,a71660a,a71664a,a71665a,a71668a,a71671a,a71672a,a71673a,a71677a,a71678a,a71681a,a71684a,a71685a,a71686a,a71690a,a71691a,a71694a,a71697a,a71698a,a71699a,a71703a,a71704a,a71707a,a71710a,a71711a,a71712a,a71716a,a71717a,a71720a,a71723a,a71724a,a71725a,a71729a,a71730a,a71733a,a71736a,a71737a,a71738a,a71742a,a71743a,a71746a,a71749a,a71750a,a71751a,a71755a,a71756a,a71759a,a71762a,a71763a,a71764a,a71768a,a71769a,a71772a,a71775a,a71776a,a71777a,a71781a,a71782a,a71785a,a71788a,a71789a,a71790a,a71794a,a71795a,a71798a,a71801a,a71802a,a71803a,a71807a,a71808a,a71811a,a71814a,a71815a,a71816a,a71820a,a71821a,a71824a,a71827a,a71828a,a71829a,a71833a,a71834a,a71837a,a71840a,a71841a,a71842a,a71846a,a71847a,a71850a,a71853a,a71854a,a71855a,a71859a,a71860a,a71863a,a71866a,a71867a,a71868a,a71872a,a71873a,a71876a,a71879a,a71880a,a71881a,a71885a,a71886a,a71889a,a71892a,a71893a,a71894a,a71898a,a71899a,a71902a,a71905a,a71906a,a71907a,a71911a,a71912a,a71915a,a71918a,a71919a,a71920a,a71924a,a71925a,a71928a,a71931a,a71932a,a71933a,a71937a,a71938a,a71941a,a71944a,a71945a,a71946a,a71950a,a71951a,a71954a,a71957a,a71958a,a71959a,a71963a,a71964a,a71967a,a71970a,a71971a,a71972a,a71976a,a71977a,a71980a,a71983a,a71984a,a71985a,a71989a,a71990a,a71993a,a71996a,a71997a,a71998a,a72002a,a72003a,a72006a,a72009a,a72010a,a72011a,a72015a,a72016a,a72019a,a72022a,a72023a,a72024a,a72028a,a72029a,a72032a,a72035a,a72036a,a72037a,a72041a,a72042a,a72045a,a72048a,a72049a,a72050a,a72054a,a72055a,a72058a,a72061a,a72062a,a72063a,a72067a,a72068a,a72071a,a72074a,a72075a,a72076a,a72080a,a72081a,a72084a,a72087a,a72088a,a72089a,a72093a,a72094a,a72097a,a72100a,a72101a,a72102a,a72106a,a72107a,a72110a,a72113a,a72114a,a72115a,a72119a,a72120a,a72123a,a72126a,a72127a,a72128a,a72132a,a72133a,a72136a,a72139a,a72140a,a72141a,a72145a,a72146a,a72149a,a72152a,a72153a,a72154a,a72158a,a72159a,a72162a,a72165a,a72166a,a72167a,a72171a,a72172a,a72175a,a72178a,a72179a,a72180a,a72184a,a72185a,a72188a,a72191a,a72192a,a72193a,a72197a,a72198a,a72201a,a72204a,a72205a,a72206a,a72210a,a72211a,a72214a,a72217a,a72218a,a72219a,a72223a,a72224a,a72227a,a72230a,a72231a,a72232a,a72236a,a72237a,a72240a,a72243a,a72244a,a72245a,a72249a,a72250a,a72253a,a72256a,a72257a,a72258a,a72262a,a72263a,a72266a,a72269a,a72270a,a72271a,a72275a,a72276a,a72279a,a72282a,a72283a,a72284a,a72288a,a72289a,a72292a,a72295a,a72296a,a72297a,a72301a,a72302a,a72305a,a72308a,a72309a,a72310a,a72314a,a72315a,a72318a,a72321a,a72322a,a72323a,a72327a,a72328a,a72331a,a72334a,a72335a,a72336a,a72340a,a72341a,a72344a,a72347a,a72348a,a72349a,a72353a,a72354a,a72357a,a72360a,a72361a,a72362a,a72366a,a72367a,a72370a,a72373a,a72374a,a72375a,a72379a,a72380a,a72383a,a72386a,a72387a,a72388a,a72392a,a72393a,a72396a,a72399a,a72400a,a72401a,a72405a,a72406a,a72409a,a72412a,a72413a,a72414a,a72418a,a72419a,a72422a,a72425a,a72426a,a72427a,a72431a,a72432a,a72435a,a72438a,a72439a,a72440a,a72444a,a72445a,a72448a,a72451a,a72452a,a72453a,a72457a,a72458a,a72461a,a72464a,a72465a,a72466a,a72470a,a72471a,a72474a,a72477a,a72478a,a72479a,a72483a,a72484a,a72487a,a72490a,a72491a,a72492a,a72496a,a72497a,a72500a,a72503a,a72504a,a72505a,a72509a,a72510a,a72513a,a72516a,a72517a,a72518a,a72522a,a72523a,a72526a,a72529a,a72530a,a72531a,a72535a,a72536a,a72539a,a72542a,a72543a,a72544a,a72548a,a72549a,a72552a,a72555a,a72556a,a72557a,a72561a,a72562a,a72565a,a72568a,a72569a,a72570a,a72574a,a72575a,a72578a,a72581a,a72582a,a72583a,a72587a,a72588a,a72591a,a72594a,a72595a,a72596a,a72600a,a72601a,a72604a,a72607a,a72608a,a72609a,a72613a,a72614a,a72617a,a72620a,a72621a,a72622a,a72626a,a72627a,a72630a,a72633a,a72634a,a72635a,a72639a,a72640a,a72643a,a72646a,a72647a,a72648a,a72652a,a72653a,a72656a,a72659a,a72660a,a72661a,a72665a,a72666a,a72669a,a72672a,a72673a,a72674a,a72678a,a72679a,a72682a,a72685a,a72686a,a72687a,a72691a,a72692a,a72695a,a72698a,a72699a,a72700a,a72704a,a72705a,a72708a,a72711a,a72712a,a72713a,a72717a,a72718a,a72721a,a72724a,a72725a,a72726a,a72730a,a72731a,a72734a,a72737a,a72738a,a72739a,a72743a,a72744a,a72747a,a72750a,a72751a,a72752a,a72756a,a72757a,a72760a,a72763a,a72764a,a72765a,a72769a,a72770a,a72773a,a72776a,a72777a,a72778a,a72782a,a72783a,a72786a,a72789a,a72790a,a72791a,a72795a,a72796a,a72799a,a72802a,a72803a,a72804a,a72808a,a72809a,a72812a,a72815a,a72816a,a72817a,a72821a,a72822a,a72825a,a72828a,a72829a,a72830a,a72834a,a72835a,a72838a,a72841a,a72842a,a72843a,a72847a,a72848a,a72851a,a72854a,a72855a,a72856a,a72860a,a72861a,a72864a,a72867a,a72868a,a72869a,a72873a,a72874a,a72877a,a72880a,a72881a,a72882a,a72886a,a72887a,a72890a,a72893a,a72894a,a72895a,a72899a,a72900a,a72903a,a72906a,a72907a,a72908a,a72912a,a72913a,a72916a,a72919a,a72920a,a72921a,a72925a,a72926a,a72929a,a72932a,a72933a,a72934a,a72938a,a72939a,a72942a,a72945a,a72946a,a72947a,a72951a,a72952a,a72955a,a72958a,a72959a,a72960a,a72964a,a72965a,a72968a,a72971a,a72972a,a72973a,a72977a,a72978a,a72981a,a72984a,a72985a,a72986a,a72990a,a72991a,a72994a,a72997a,a72998a,a72999a,a73003a,a73004a,a73007a,a73010a,a73011a,a73012a,a73016a,a73017a,a73020a,a73023a,a73024a,a73025a,a73029a,a73030a,a73033a,a73036a,a73037a,a73038a,a73042a,a73043a,a73046a,a73049a,a73050a,a73051a,a73055a,a73056a,a73059a,a73062a,a73063a,a73064a,a73068a,a73069a,a73072a,a73075a,a73076a,a73077a,a73081a,a73082a,a73085a,a73088a,a73089a,a73090a,a73094a,a73095a,a73098a,a73101a,a73102a,a73103a,a73107a,a73108a,a73111a,a73114a,a73115a,a73116a,a73120a,a73121a,a73124a,a73127a,a73128a,a73129a,a73133a,a73134a,a73137a,a73140a,a73141a,a73142a,a73146a,a73147a,a73150a,a73153a,a73154a,a73155a,a73159a,a73160a,a73163a,a73166a,a73167a,a73168a,a73172a,a73173a,a73176a,a73179a,a73180a,a73181a,a73185a,a73186a,a73189a,a73192a,a73193a,a73194a,a73198a,a73199a,a73202a,a73205a,a73206a,a73207a,a73211a,a73212a,a73215a,a73218a,a73219a,a73220a,a73224a,a73225a,a73228a,a73231a,a73232a,a73233a,a73237a,a73238a,a73241a,a73244a,a73245a,a73246a,a73250a,a73251a,a73254a,a73257a,a73258a,a73259a,a73263a,a73264a,a73267a,a73270a,a73271a,a73272a,a73276a,a73277a,a73280a,a73283a,a73284a,a73285a,a73289a,a73290a,a73293a,a73296a,a73297a,a73298a,a73302a,a73303a,a73306a,a73309a,a73310a,a73311a,a73315a,a73316a,a73319a,a73322a,a73323a,a73324a,a73328a,a73329a,a73332a,a73335a,a73336a,a73337a,a73341a,a73342a,a73345a,a73348a,a73349a,a73350a,a73354a,a73355a,a73358a,a73361a,a73362a,a73363a,a73367a,a73368a,a73371a,a73374a,a73375a,a73376a,a73380a,a73381a,a73384a,a73387a,a73388a,a73389a,a73393a,a73394a,a73397a,a73400a,a73401a,a73402a,a73406a,a73407a,a73410a,a73413a,a73414a,a73415a,a73419a,a73420a,a73423a,a73426a,a73427a,a73428a,a73432a,a73433a,a73436a,a73439a,a73440a,a73441a,a73445a,a73446a,a73449a,a73452a,a73453a,a73454a,a73458a,a73459a,a73462a,a73465a,a73466a,a73467a,a73471a,a73472a,a73475a,a73478a,a73479a,a73480a,a73484a,a73485a,a73488a,a73491a,a73492a,a73493a,a73497a,a73498a,a73501a,a73504a,a73505a,a73506a,a73510a,a73511a,a73514a,a73517a,a73518a,a73519a,a73523a,a73524a,a73527a,a73530a,a73531a,a73532a,a73536a,a73537a,a73540a,a73543a,a73544a,a73545a,a73549a,a73550a,a73553a,a73556a,a73557a,a73558a,a73562a,a73563a,a73566a,a73569a,a73570a,a73571a,a73575a,a73576a,a73579a,a73582a,a73583a,a73584a,a73588a,a73589a,a73592a,a73595a,a73596a,a73597a,a73601a,a73602a,a73605a,a73608a,a73609a,a73610a,a73614a,a73615a,a73618a,a73621a,a73622a,a73623a,a73627a,a73628a,a73631a,a73634a,a73635a,a73636a,a73640a,a73641a,a73644a,a73647a,a73648a,a73649a,a73653a,a73654a,a73657a,a73660a,a73661a,a73662a,a73666a,a73667a,a73670a,a73673a,a73674a,a73675a,a73679a,a73680a,a73683a,a73686a,a73687a,a73688a,a73692a,a73693a,a73696a,a73699a,a73700a,a73701a,a73705a,a73706a,a73709a,a73712a,a73713a,a73714a,a73718a,a73719a,a73722a,a73725a,a73726a,a73727a,a73731a,a73732a,a73735a,a73738a,a73739a,a73740a,a73744a,a73745a,a73748a,a73751a,a73752a,a73753a,a73757a,a73758a,a73761a,a73764a,a73765a,a73766a,a73770a,a73771a,a73774a,a73777a,a73778a,a73779a,a73783a,a73784a,a73787a,a73790a,a73791a,a73792a,a73796a,a73797a,a73800a,a73803a,a73804a,a73805a,a73809a,a73810a,a73813a,a73816a,a73817a,a73818a,a73822a,a73823a,a73826a,a73829a,a73830a,a73831a,a73835a,a73836a,a73839a,a73842a,a73843a,a73844a,a73848a,a73849a,a73852a,a73855a,a73856a,a73857a,a73861a,a73862a,a73865a,a73868a,a73869a,a73870a,a73874a,a73875a,a73878a,a73881a,a73882a,a73883a,a73887a,a73888a,a73891a,a73894a,a73895a,a73896a,a73900a,a73901a,a73904a,a73907a,a73908a,a73909a,a73913a,a73914a,a73917a,a73920a,a73921a,a73922a,a73926a,a73927a,a73930a,a73933a,a73934a,a73935a,a73939a,a73940a,a73943a,a73946a,a73947a,a73948a,a73952a,a73953a,a73956a,a73959a,a73960a,a73961a,a73965a,a73966a,a73969a,a73972a,a73973a,a73974a,a73978a,a73979a,a73982a,a73985a,a73986a,a73987a,a73991a,a73992a,a73995a,a73998a,a73999a,a74000a,a74004a,a74005a,a74008a,a74011a,a74012a,a74013a,a74017a,a74018a,a74021a,a74024a,a74025a,a74026a,a74030a,a74031a,a74034a,a74037a,a74038a,a74039a,a74043a,a74044a,a74047a,a74050a,a74051a,a74052a,a74056a,a74057a,a74060a,a74063a,a74064a,a74065a,a74069a,a74070a,a74073a,a74076a,a74077a,a74078a,a74082a,a74083a,a74086a,a74089a,a74090a,a74091a,a74095a,a74096a,a74099a,a74102a,a74103a,a74104a,a74108a,a74109a,a74112a,a74115a,a74116a,a74117a,a74121a,a74122a,a74125a,a74128a,a74129a,a74130a,a74134a,a74135a,a74138a,a74141a,a74142a,a74143a,a74147a,a74148a,a74151a,a74154a,a74155a,a74156a,a74160a,a74161a,a74164a,a74167a,a74168a,a74169a,a74173a,a74174a,a74177a,a74180a,a74181a,a74182a,a74186a,a74187a,a74190a,a74193a,a74194a,a74195a,a74199a,a74200a,a74203a,a74206a,a74207a,a74208a,a74212a,a74213a,a74216a,a74219a,a74220a,a74221a,a74225a,a74226a,a74229a,a74232a,a74233a,a74234a,a74238a,a74239a,a74242a,a74245a,a74246a,a74247a,a74251a,a74252a,a74255a,a74258a,a74259a,a74260a,a74264a,a74265a,a74268a,a74271a,a74272a,a74273a,a74277a,a74278a,a74281a,a74284a,a74285a,a74286a,a74290a,a74291a,a74294a,a74297a,a74298a,a74299a,a74303a,a74304a,a74307a,a74310a,a74311a,a74312a,a74316a,a74317a,a74320a,a74323a,a74324a,a74325a,a74329a,a74330a,a74333a,a74336a,a74337a,a74338a,a74342a,a74343a,a74346a,a74349a,a74350a,a74351a,a74355a,a74356a,a74359a,a74362a,a74363a,a74364a,a74368a,a74369a,a74372a,a74375a,a74376a,a74377a,a74381a,a74382a,a74385a,a74388a,a74389a,a74390a,a74394a,a74395a,a74398a,a74401a,a74402a,a74403a,a74407a,a74408a,a74411a,a74414a,a74415a,a74416a,a74420a,a74421a,a74424a,a74427a,a74428a,a74429a,a74433a,a74434a,a74437a,a74440a,a74441a,a74442a,a74446a,a74447a,a74450a,a74453a,a74454a,a74455a,a74459a,a74460a,a74463a,a74466a,a74467a,a74468a,a74472a,a74473a,a74476a,a74479a,a74480a,a74481a,a74485a,a74486a,a74489a,a74492a,a74493a,a74494a,a74498a,a74499a,a74502a,a74505a,a74506a,a74507a,a74511a,a74512a,a74515a,a74518a,a74519a,a74520a,a74524a,a74525a,a74528a,a74531a,a74532a,a74533a,a74537a,a74538a,a74541a,a74544a,a74545a,a74546a,a74550a,a74551a,a74554a,a74557a,a74558a,a74559a,a74563a,a74564a,a74567a,a74570a,a74571a,a74572a,a74576a,a74577a,a74580a,a74583a,a74584a,a74585a,a74589a,a74590a,a74593a,a74596a,a74597a,a74598a,a74602a,a74603a,a74606a,a74609a,a74610a,a74611a,a74615a,a74616a,a74619a,a74622a,a74623a,a74624a,a74628a,a74629a,a74632a,a74635a,a74636a,a74637a,a74641a,a74642a,a74645a,a74648a,a74649a,a74650a,a74654a,a74655a,a74658a,a74661a,a74662a,a74663a,a74667a,a74668a,a74671a,a74674a,a74675a,a74676a,a74680a,a74681a,a74684a,a74687a,a74688a,a74689a,a74693a,a74694a,a74697a,a74700a,a74701a,a74702a,a74706a,a74707a,a74710a,a74713a,a74714a,a74715a,a74719a,a74720a,a74723a,a74726a,a74727a,a74728a,a74732a,a74733a,a74736a,a74739a,a74740a,a74741a,a74745a,a74746a,a74749a,a74752a,a74753a,a74754a,a74758a,a74759a,a74762a,a74765a,a74766a,a74767a,a74771a,a74772a,a74775a,a74778a,a74779a,a74780a,a74784a,a74785a,a74788a,a74791a,a74792a,a74793a,a74797a,a74798a,a74801a,a74804a,a74805a,a74806a,a74810a,a74811a,a74814a,a74817a,a74818a,a74819a,a74823a,a74824a,a74827a,a74830a,a74831a,a74832a,a74836a,a74837a,a74840a,a74843a,a74844a,a74845a,a74849a,a74850a,a74853a,a74856a,a74857a,a74858a,a74862a,a74863a,a74866a,a74869a,a74870a,a74871a,a74875a,a74876a,a74879a,a74882a,a74883a,a74884a,a74888a,a74889a,a74892a,a74895a,a74896a,a74897a,a74901a,a74902a,a74905a,a74908a,a74909a,a74910a,a74914a,a74915a,a74918a,a74921a,a74922a,a74923a,a74927a,a74928a,a74931a,a74934a,a74935a,a74936a,a74940a,a74941a,a74944a,a74947a,a74948a,a74949a,a74953a,a74954a,a74957a,a74960a,a74961a,a74962a,a74966a,a74967a,a74970a,a74973a,a74974a,a74975a,a74979a,a74980a,a74983a,a74986a,a74987a,a74988a,a74992a,a74993a,a74996a,a74999a,a75000a,a75001a,a75005a,a75006a,a75009a,a75012a,a75013a,a75014a,a75018a,a75019a,a75022a,a75025a,a75026a,a75027a,a75031a,a75032a,a75035a,a75038a,a75039a,a75040a,a75044a,a75045a,a75048a,a75051a,a75052a,a75053a,a75057a,a75058a,a75061a,a75064a,a75065a,a75066a,a75070a,a75071a,a75074a,a75077a,a75078a,a75079a,a75083a,a75084a,a75087a,a75090a,a75091a,a75092a,a75096a,a75097a,a75100a,a75103a,a75104a,a75105a,a75109a,a75110a,a75113a,a75116a,a75117a,a75118a,a75122a,a75123a,a75126a,a75129a,a75130a,a75131a,a75135a,a75136a,a75139a,a75142a,a75143a,a75144a,a75148a,a75149a,a75152a,a75155a,a75156a,a75157a,a75161a,a75162a,a75165a,a75168a,a75169a,a75170a,a75174a,a75175a,a75178a,a75181a,a75182a,a75183a,a75187a,a75188a,a75191a,a75194a,a75195a,a75196a,a75200a,a75201a,a75204a,a75207a,a75208a,a75209a,a75213a,a75214a,a75217a,a75220a,a75221a,a75222a,a75226a,a75227a,a75230a,a75233a,a75234a,a75235a,a75239a,a75240a,a75243a,a75246a,a75247a,a75248a,a75252a,a75253a,a75256a,a75259a,a75260a,a75261a,a75265a,a75266a,a75269a,a75272a,a75273a,a75274a,a75278a,a75279a,a75282a,a75285a,a75286a,a75287a,a75291a,a75292a,a75295a,a75298a,a75299a,a75300a,a75304a,a75305a,a75308a,a75311a,a75312a,a75313a,a75317a,a75318a,a75321a,a75324a,a75325a,a75326a,a75330a,a75331a,a75334a,a75337a,a75338a,a75339a,a75343a,a75344a,a75347a,a75350a,a75351a,a75352a,a75356a,a75357a,a75360a,a75363a,a75364a,a75365a,a75369a,a75370a,a75373a,a75376a,a75377a,a75378a,a75382a,a75383a,a75386a,a75389a,a75390a,a75391a,a75395a,a75396a,a75399a,a75402a,a75403a,a75404a,a75408a,a75409a,a75412a,a75415a,a75416a,a75417a,a75421a,a75422a,a75425a,a75428a,a75429a,a75430a,a75434a,a75435a,a75438a,a75441a,a75442a,a75443a,a75447a,a75448a,a75451a,a75454a,a75455a,a75456a,a75460a,a75461a,a75464a,a75467a,a75468a,a75469a,a75473a,a75474a,a75477a,a75480a,a75481a,a75482a,a75486a,a75487a,a75490a,a75493a,a75494a,a75495a,a75499a,a75500a,a75503a,a75506a,a75507a,a75508a,a75512a,a75513a,a75516a,a75519a,a75520a,a75521a,a75525a,a75526a,a75529a,a75532a,a75533a,a75534a,a75538a,a75539a,a75542a,a75545a,a75546a,a75547a,a75551a,a75552a,a75555a,a75558a,a75559a,a75560a,a75564a,a75565a,a75568a,a75571a,a75572a,a75573a,a75577a,a75578a,a75581a,a75584a,a75585a,a75586a,a75590a,a75591a,a75594a,a75597a,a75598a,a75599a,a75603a,a75604a,a75607a,a75610a,a75611a,a75612a,a75616a,a75617a,a75620a,a75623a,a75624a,a75625a,a75629a,a75630a,a75633a,a75636a,a75637a,a75638a,a75642a,a75643a,a75646a,a75649a,a75650a,a75651a,a75655a,a75656a,a75659a,a75662a,a75663a,a75664a,a75668a,a75669a,a75672a,a75675a,a75676a,a75677a,a75681a,a75682a,a75685a,a75688a,a75689a,a75690a,a75694a,a75695a,a75698a,a75701a,a75702a,a75703a,a75707a,a75708a,a75711a,a75714a,a75715a,a75716a,a75720a,a75721a,a75724a,a75727a,a75728a,a75729a,a75733a,a75734a,a75737a,a75740a,a75741a,a75742a,a75746a,a75747a,a75750a,a75753a,a75754a,a75755a,a75759a,a75760a,a75763a,a75766a,a75767a,a75768a,a75772a,a75773a,a75776a,a75779a,a75780a,a75781a,a75785a,a75786a,a75789a,a75792a,a75793a,a75794a,a75798a,a75799a,a75802a,a75805a,a75806a,a75807a,a75811a,a75812a,a75815a,a75818a,a75819a,a75820a,a75824a,a75825a,a75828a,a75831a,a75832a,a75833a,a75837a,a75838a,a75841a,a75844a,a75845a,a75846a,a75850a,a75851a,a75854a,a75857a,a75858a,a75859a,a75863a,a75864a,a75867a,a75870a,a75871a,a75872a,a75876a,a75877a,a75880a,a75883a,a75884a,a75885a,a75889a,a75890a,a75893a,a75896a,a75897a,a75898a,a75902a,a75903a,a75906a,a75909a,a75910a,a75911a,a75915a,a75916a,a75919a,a75922a,a75923a,a75924a,a75928a,a75929a,a75932a,a75935a,a75936a,a75937a,a75941a,a75942a,a75945a,a75948a,a75949a,a75950a,a75954a,a75955a,a75958a,a75961a,a75962a,a75963a,a75967a,a75968a,a75971a,a75974a,a75975a,a75976a,a75980a,a75981a,a75984a,a75987a,a75988a,a75989a,a75993a,a75994a,a75997a,a76000a,a76001a,a76002a,a76006a,a76007a,a76010a,a76013a,a76014a,a76015a,a76019a,a76020a,a76023a,a76026a,a76027a,a76028a,a76032a,a76033a,a76036a,a76039a,a76040a,a76041a,a76045a,a76046a,a76049a,a76052a,a76053a,a76054a,a76058a,a76059a,a76062a,a76065a,a76066a,a76067a,a76071a,a76072a,a76075a,a76078a,a76079a,a76080a,a76084a,a76085a,a76088a,a76091a,a76092a,a76093a,a76097a,a76098a,a76101a,a76104a,a76105a,a76106a,a76110a,a76111a,a76114a,a76117a,a76118a,a76119a,a76123a,a76124a,a76127a,a76130a,a76131a,a76132a,a76136a,a76137a,a76140a,a76143a,a76144a,a76145a,a76149a,a76150a,a76153a,a76156a,a76157a,a76158a,a76162a,a76163a,a76166a,a76169a,a76170a,a76171a,a76175a,a76176a,a76179a,a76182a,a76183a,a76184a,a76188a,a76189a,a76192a,a76195a,a76196a,a76197a,a76201a,a76202a,a76205a,a76208a,a76209a,a76210a,a76214a,a76215a,a76218a,a76221a,a76222a,a76223a,a76227a,a76228a,a76231a,a76234a,a76235a,a76236a,a76240a,a76241a,a76244a,a76247a,a76248a,a76249a,a76253a,a76254a,a76257a,a76260a,a76261a,a76262a,a76266a,a76267a,a76270a,a76273a,a76274a,a76275a,a76279a,a76280a,a76283a,a76286a,a76287a,a76288a,a76292a,a76293a,a76296a,a76299a,a76300a,a76301a,a76305a,a76306a,a76309a,a76312a,a76313a,a76314a,a76318a,a76319a,a76322a,a76325a,a76326a,a76327a,a76331a,a76332a,a76335a,a76338a,a76339a,a76340a,a76344a,a76345a,a76348a,a76351a,a76352a,a76353a,a76357a,a76358a,a76361a,a76364a,a76365a,a76366a,a76370a,a76371a,a76374a,a76377a,a76378a,a76379a,a76383a,a76384a,a76387a,a76390a,a76391a,a76392a,a76396a,a76397a,a76400a,a76403a,a76404a,a76405a,a76409a,a76410a,a76413a,a76416a,a76417a,a76418a,a76422a,a76423a,a76426a,a76429a,a76430a,a76431a,a76435a,a76436a,a76439a,a76442a,a76443a,a76444a,a76448a,a76449a,a76452a,a76455a,a76456a,a76457a,a76461a,a76462a,a76465a,a76468a,a76469a,a76470a,a76474a,a76475a,a76478a,a76481a,a76482a,a76483a,a76487a,a76488a,a76491a,a76494a,a76495a,a76496a,a76500a,a76501a,a76504a,a76507a,a76508a,a76509a,a76513a,a76514a,a76517a,a76520a,a76521a,a76522a,a76526a,a76527a,a76530a,a76533a,a76534a,a76535a,a76539a,a76540a,a76543a,a76546a,a76547a,a76548a,a76552a,a76553a,a76556a,a76559a,a76560a,a76561a,a76565a,a76566a,a76569a,a76572a,a76573a,a76574a,a76578a,a76579a,a76582a,a76585a,a76586a,a76587a,a76591a,a76592a,a76595a,a76598a,a76599a,a76600a,a76604a,a76605a,a76608a,a76611a,a76612a,a76613a,a76617a,a76618a,a76621a,a76624a,a76625a,a76626a,a76630a,a76631a,a76634a,a76637a,a76638a,a76639a,a76643a,a76644a,a76647a,a76650a,a76651a,a76652a,a76656a,a76657a,a76660a,a76663a,a76664a,a76665a,a76669a,a76670a,a76673a,a76676a,a76677a,a76678a,a76682a,a76683a,a76686a,a76689a,a76690a,a76691a,a76695a,a76696a,a76699a,a76702a,a76703a,a76704a,a76708a,a76709a,a76712a,a76715a,a76716a,a76717a,a76721a,a76722a,a76725a,a76728a,a76729a,a76730a,a76734a,a76735a,a76738a,a76741a,a76742a,a76743a,a76747a,a76748a,a76751a,a76754a,a76755a,a76756a,a76760a,a76761a,a76764a,a76767a,a76768a,a76769a,a76773a,a76774a,a76777a,a76780a,a76781a,a76782a,a76786a,a76787a,a76790a,a76793a,a76794a,a76795a,a76799a,a76800a,a76803a,a76806a,a76807a,a76808a,a76812a,a76813a,a76816a,a76819a,a76820a,a76821a,a76825a,a76826a,a76829a,a76832a,a76833a,a76834a,a76838a,a76839a,a76842a,a76845a,a76846a,a76847a,a76851a,a76852a,a76855a,a76858a,a76859a,a76860a,a76864a,a76865a,a76868a,a76871a,a76872a,a76873a,a76877a,a76878a,a76881a,a76884a,a76885a,a76886a,a76890a,a76891a,a76894a,a76897a,a76898a,a76899a,a76903a,a76904a,a76907a,a76910a,a76911a,a76912a,a76916a,a76917a,a76920a,a76923a,a76924a,a76925a,a76929a,a76930a,a76933a,a76936a,a76937a,a76938a,a76942a,a76943a,a76946a,a76949a,a76950a,a76951a,a76955a,a76956a,a76959a,a76962a,a76963a,a76964a,a76968a,a76969a,a76972a,a76975a,a76976a,a76977a,a76981a,a76982a,a76985a,a76988a,a76989a,a76990a,a76994a,a76995a,a76998a,a77001a,a77002a,a77003a,a77007a,a77008a,a77011a,a77014a,a77015a,a77016a,a77020a,a77021a,a77024a,a77027a,a77028a,a77029a,a77033a,a77034a,a77037a,a77040a,a77041a,a77042a,a77046a,a77047a,a77050a,a77053a,a77054a,a77055a,a77059a,a77060a,a77063a,a77066a,a77067a,a77068a,a77072a,a77073a,a77076a,a77079a,a77080a,a77081a,a77085a,a77086a,a77089a,a77092a,a77093a,a77094a,a77098a,a77099a,a77102a,a77105a,a77106a,a77107a,a77111a,a77112a,a77115a,a77118a,a77119a,a77120a,a77124a,a77125a,a77128a,a77131a,a77132a,a77133a,a77137a,a77138a,a77141a,a77144a,a77145a,a77146a,a77150a,a77151a,a77154a,a77157a,a77158a,a77159a,a77163a,a77164a,a77167a,a77170a,a77171a,a77172a,a77176a,a77177a,a77180a,a77183a,a77184a,a77185a,a77189a,a77190a,a77193a,a77196a,a77197a,a77198a,a77202a,a77203a,a77206a,a77209a,a77210a,a77211a,a77215a,a77216a,a77219a,a77222a,a77223a,a77224a,a77228a,a77229a,a77232a,a77235a,a77236a,a77237a,a77241a,a77242a,a77245a,a77248a,a77249a,a77250a,a77254a,a77255a,a77258a,a77261a,a77262a,a77263a,a77267a,a77268a,a77271a,a77274a,a77275a,a77276a,a77280a,a77281a,a77284a,a77287a,a77288a,a77289a,a77293a,a77294a,a77297a,a77300a,a77301a,a77302a,a77306a,a77307a,a77310a,a77313a,a77314a,a77315a,a77319a,a77320a,a77323a,a77326a,a77327a,a77328a,a77332a,a77333a,a77336a,a77339a,a77340a,a77341a,a77345a,a77346a,a77349a,a77352a,a77353a,a77354a,a77358a,a77359a,a77362a,a77365a,a77366a,a77367a,a77371a,a77372a,a77375a,a77378a,a77379a,a77380a,a77384a,a77385a,a77388a,a77391a,a77392a,a77393a,a77397a,a77398a,a77401a,a77404a,a77405a,a77406a,a77410a,a77411a,a77414a,a77417a,a77418a,a77419a,a77423a,a77424a,a77427a,a77430a,a77431a,a77432a,a77436a,a77437a,a77440a,a77443a,a77444a,a77445a,a77449a,a77450a,a77453a,a77456a,a77457a,a77458a,a77462a,a77463a,a77466a,a77469a,a77470a,a77471a,a77475a,a77476a,a77479a,a77482a,a77483a,a77484a,a77488a,a77489a,a77492a,a77495a,a77496a,a77497a,a77501a,a77502a,a77505a,a77508a,a77509a,a77510a,a77514a,a77515a,a77518a,a77521a,a77522a,a77523a,a77527a,a77528a,a77531a,a77534a,a77535a,a77536a,a77540a,a77541a,a77544a,a77547a,a77548a,a77549a,a77553a,a77554a,a77557a,a77560a,a77561a,a77562a,a77566a,a77567a,a77570a,a77573a,a77574a,a77575a,a77579a,a77580a,a77583a,a77586a,a77587a,a77588a,a77592a,a77593a,a77596a,a77599a,a77600a,a77601a,a77605a,a77606a,a77609a,a77612a,a77613a,a77614a,a77618a,a77619a,a77622a,a77625a,a77626a,a77627a,a77631a,a77632a,a77635a,a77638a,a77639a,a77640a,a77644a,a77645a,a77648a,a77651a,a77652a,a77653a,a77657a,a77658a,a77661a,a77664a,a77665a,a77666a,a77670a,a77671a,a77674a,a77677a,a77678a,a77679a,a77683a,a77684a,a77687a,a77690a,a77691a,a77692a,a77696a,a77697a,a77700a,a77703a,a77704a,a77705a,a77709a,a77710a,a77713a,a77716a,a77717a,a77718a,a77722a,a77723a,a77726a,a77729a,a77730a,a77731a,a77735a,a77736a,a77739a,a77742a,a77743a,a77744a,a77748a,a77749a,a77752a,a77755a,a77756a,a77757a,a77761a,a77762a,a77765a,a77768a,a77769a,a77770a,a77774a,a77775a,a77778a,a77781a,a77782a,a77783a,a77787a,a77788a,a77791a,a77794a,a77795a,a77796a,a77800a,a77801a,a77804a,a77807a,a77808a,a77809a,a77813a,a77814a,a77817a,a77820a,a77821a,a77822a,a77826a,a77827a,a77830a,a77833a,a77834a,a77835a,a77839a,a77840a,a77843a,a77846a,a77847a,a77848a,a77852a,a77853a,a77856a,a77859a,a77860a,a77861a,a77865a,a77866a,a77869a,a77872a,a77873a,a77874a,a77878a,a77879a,a77882a,a77885a,a77886a,a77887a,a77891a,a77892a,a77895a,a77898a,a77899a,a77900a,a77904a,a77905a,a77908a,a77911a,a77912a,a77913a,a77917a,a77918a,a77921a,a77924a,a77925a,a77926a,a77930a,a77931a,a77934a,a77937a,a77938a,a77939a,a77943a,a77944a,a77947a,a77950a,a77951a,a77952a,a77956a,a77957a,a77960a,a77963a,a77964a,a77965a,a77969a,a77970a,a77973a,a77976a,a77977a,a77978a,a77982a,a77983a,a77986a,a77989a,a77990a,a77991a,a77995a,a77996a,a77999a,a78002a,a78003a,a78004a,a78008a,a78009a,a78012a,a78015a,a78016a,a78017a,a78021a,a78022a,a78025a,a78028a,a78029a,a78030a,a78034a,a78035a,a78038a,a78041a,a78042a,a78043a,a78047a,a78048a,a78051a,a78054a,a78055a,a78056a,a78060a,a78061a,a78064a,a78067a,a78068a,a78069a,a78073a,a78074a,a78077a,a78080a,a78081a,a78082a,a78086a,a78087a,a78090a,a78093a,a78094a,a78095a,a78099a,a78100a,a78103a,a78106a,a78107a,a78108a,a78112a,a78113a,a78116a,a78119a,a78120a,a78121a,a78125a,a78126a,a78129a,a78132a,a78133a,a78134a,a78138a,a78139a,a78142a,a78145a,a78146a,a78147a,a78151a,a78152a,a78155a,a78158a,a78159a,a78160a,a78164a,a78165a,a78168a,a78171a,a78172a,a78173a,a78177a,a78178a,a78181a,a78184a,a78185a,a78186a,a78190a,a78191a,a78194a,a78197a,a78198a,a78199a,a78203a,a78204a,a78207a,a78210a,a78211a,a78212a,a78216a,a78217a,a78220a,a78223a,a78224a,a78225a,a78229a,a78230a,a78233a,a78236a,a78237a,a78238a,a78242a,a78243a,a78246a,a78249a,a78250a,a78251a,a78255a,a78256a,a78259a,a78262a,a78263a,a78264a,a78268a,a78269a,a78272a,a78275a,a78276a,a78277a,a78281a,a78282a,a78285a,a78288a,a78289a,a78290a,a78294a,a78295a,a78298a,a78301a,a78302a,a78303a,a78307a,a78308a,a78311a,a78314a,a78315a,a78316a,a78320a,a78321a,a78324a,a78327a,a78328a,a78329a,a78333a,a78334a,a78337a,a78340a,a78341a,a78342a,a78346a,a78347a,a78350a,a78353a,a78354a,a78355a,a78359a,a78360a,a78363a,a78366a,a78367a,a78368a,a78372a,a78373a,a78376a,a78379a,a78380a,a78381a,a78385a,a78386a,a78389a,a78392a,a78393a,a78394a,a78398a,a78399a,a78402a,a78405a,a78406a,a78407a,a78411a,a78412a,a78415a,a78418a,a78419a,a78420a,a78424a,a78425a,a78428a,a78431a,a78432a,a78433a,a78437a,a78438a,a78441a,a78444a,a78445a,a78446a,a78450a,a78451a,a78454a,a78457a,a78458a,a78459a,a78463a,a78464a,a78467a,a78470a,a78471a,a78472a,a78476a,a78477a,a78480a,a78483a,a78484a,a78485a,a78489a,a78490a,a78493a,a78496a,a78497a,a78498a,a78502a,a78503a,a78506a,a78509a,a78510a,a78511a,a78515a,a78516a,a78519a,a78522a,a78523a,a78524a,a78528a,a78529a,a78532a,a78535a,a78536a,a78537a,a78541a,a78542a,a78545a,a78548a,a78549a,a78550a,a78554a,a78555a,a78558a,a78561a,a78562a,a78563a,a78567a,a78568a,a78571a,a78574a,a78575a,a78576a,a78580a,a78581a,a78584a,a78587a,a78588a,a78589a,a78593a,a78594a,a78597a,a78600a,a78601a,a78602a,a78606a,a78607a,a78610a,a78613a,a78614a,a78615a,a78619a,a78620a,a78623a,a78626a,a78627a,a78628a,a78632a,a78633a,a78636a,a78639a,a78640a,a78641a,a78645a,a78646a,a78649a,a78652a,a78653a,a78654a,a78658a,a78659a,a78662a,a78665a,a78666a,a78667a,a78671a,a78672a,a78675a,a78678a,a78679a,a78680a,a78684a,a78685a,a78688a,a78691a,a78692a,a78693a,a78697a,a78698a,a78701a,a78704a,a78705a,a78706a,a78710a,a78711a,a78714a,a78717a,a78718a,a78719a,a78723a,a78724a,a78727a,a78730a,a78731a,a78732a,a78736a,a78737a,a78740a,a78743a,a78744a,a78745a,a78749a,a78750a,a78753a,a78756a,a78757a,a78758a,a78762a,a78763a,a78766a,a78769a,a78770a,a78771a,a78775a,a78776a,a78779a,a78782a,a78783a,a78784a,a78788a,a78789a,a78792a,a78795a,a78796a,a78797a,a78801a,a78802a,a78805a,a78808a,a78809a,a78810a,a78814a,a78815a,a78818a,a78821a,a78822a,a78823a,a78827a,a78828a,a78831a,a78834a,a78835a,a78836a,a78840a,a78841a,a78844a,a78847a,a78848a,a78849a,a78853a,a78854a,a78857a,a78860a,a78861a,a78862a,a78866a,a78867a,a78870a,a78873a,a78874a,a78875a,a78879a,a78880a,a78883a,a78886a,a78887a,a78888a,a78892a,a78893a,a78896a,a78899a,a78900a,a78901a,a78905a,a78906a,a78909a,a78912a,a78913a,a78914a,a78918a,a78919a,a78922a,a78925a,a78926a,a78927a,a78931a,a78932a,a78935a,a78938a,a78939a,a78940a,a78944a,a78945a,a78948a,a78951a,a78952a,a78953a,a78957a,a78958a,a78961a,a78964a,a78965a,a78966a,a78970a,a78971a,a78974a,a78977a,a78978a,a78979a,a78983a,a78984a,a78987a,a78990a,a78991a,a78992a,a78996a,a78997a,a79000a,a79003a,a79004a,a79005a,a79009a,a79010a,a79013a,a79016a,a79017a,a79018a,a79022a,a79023a,a79026a,a79029a,a79030a,a79031a,a79035a,a79036a,a79039a,a79042a,a79043a,a79044a,a79048a,a79049a,a79052a,a79055a,a79056a,a79057a,a79061a,a79062a,a79065a,a79068a,a79069a,a79070a,a79074a,a79075a,a79078a,a79081a,a79082a,a79083a,a79087a,a79088a,a79091a,a79094a,a79095a,a79096a,a79100a,a79101a,a79104a,a79107a,a79108a,a79109a,a79113a,a79114a,a79117a,a79120a,a79121a,a79122a,a79126a,a79127a,a79130a,a79133a,a79134a,a79135a,a79139a,a79140a,a79143a,a79146a,a79147a,a79148a,a79152a,a79153a,a79156a,a79159a,a79160a,a79161a,a79165a,a79166a,a79169a,a79172a,a79173a,a79174a,a79178a,a79179a,a79182a,a79185a,a79186a,a79187a,a79191a,a79192a,a79195a,a79198a,a79199a,a79200a,a79204a,a79205a,a79208a,a79211a,a79212a,a79213a,a79217a,a79218a,a79221a,a79224a,a79225a,a79226a,a79230a,a79231a,a79234a,a79237a,a79238a,a79239a,a79243a,a79244a,a79247a,a79250a,a79251a,a79252a,a79256a,a79257a,a79260a,a79263a,a79264a,a79265a,a79269a,a79270a,a79273a,a79276a,a79277a,a79278a,a79282a,a79283a,a79286a,a79289a,a79290a,a79291a,a79295a,a79296a,a79299a,a79302a,a79303a,a79304a,a79308a,a79309a,a79312a,a79315a,a79316a,a79317a,a79321a,a79322a,a79325a,a79328a,a79329a,a79330a,a79334a,a79335a,a79338a,a79341a,a79342a,a79343a,a79347a,a79348a,a79351a,a79354a,a79355a,a79356a,a79360a,a79361a,a79364a,a79367a,a79368a,a79369a,a79373a,a79374a,a79377a,a79380a,a79381a,a79382a,a79386a,a79387a,a79390a,a79393a,a79394a,a79395a,a79399a,a79400a,a79403a,a79406a,a79407a,a79408a,a79412a,a79413a,a79416a,a79419a,a79420a,a79421a,a79425a,a79426a,a79429a,a79432a,a79433a,a79434a,a79438a,a79439a,a79442a,a79445a,a79446a,a79447a,a79451a,a79452a,a79455a,a79458a,a79459a,a79460a,a79464a,a79465a,a79468a,a79471a,a79472a,a79473a,a79477a,a79478a,a79481a,a79484a,a79485a,a79486a,a79490a,a79491a,a79494a,a79497a,a79498a,a79499a,a79503a,a79504a,a79507a,a79510a,a79511a,a79512a,a79516a,a79517a,a79520a,a79523a,a79524a,a79525a,a79529a,a79530a,a79533a,a79536a,a79537a,a79538a,a79542a,a79543a,a79546a,a79549a,a79550a,a79551a,a79555a,a79556a,a79559a,a79562a,a79563a,a79564a,a79568a,a79569a,a79572a,a79575a,a79576a,a79577a,a79581a,a79582a,a79585a,a79588a,a79589a,a79590a,a79594a,a79595a,a79598a,a79601a,a79602a,a79603a,a79607a,a79608a,a79611a,a79614a,a79615a,a79616a,a79620a,a79621a,a79624a,a79627a,a79628a,a79629a,a79633a,a79634a,a79637a,a79640a,a79641a,a79642a,a79646a,a79647a,a79650a,a79653a,a79654a,a79655a,a79659a,a79660a,a79663a,a79666a,a79667a,a79668a,a79672a,a79673a,a79676a,a79679a,a79680a,a79681a,a79685a,a79686a,a79689a,a79692a,a79693a,a79694a,a79698a,a79699a,a79702a,a79705a,a79706a,a79707a,a79711a,a79712a,a79715a,a79718a,a79719a,a79720a,a79724a,a79725a,a79728a,a79731a,a79732a,a79733a,a79737a,a79738a,a79741a,a79744a,a79745a,a79746a,a79750a,a79751a,a79754a,a79757a,a79758a,a79759a,a79763a,a79764a,a79767a,a79770a,a79771a,a79772a,a79776a,a79777a,a79780a,a79783a,a79784a,a79785a,a79789a,a79790a,a79793a,a79796a,a79797a,a79798a,a79802a,a79803a,a79806a,a79809a,a79810a,a79811a,a79815a,a79816a,a79819a,a79822a,a79823a,a79824a,a79828a,a79829a,a79832a,a79835a,a79836a,a79837a,a79841a,a79842a,a79845a,a79848a,a79849a,a79850a,a79854a,a79855a,a79858a,a79861a,a79862a,a79863a,a79867a,a79868a,a79871a,a79874a,a79875a,a79876a,a79880a,a79881a,a79884a,a79887a,a79888a,a79889a,a79893a,a79894a,a79897a,a79900a,a79901a,a79902a,a79906a,a79907a,a79910a,a79913a,a79914a,a79915a,a79919a,a79920a,a79923a,a79926a,a79927a,a79928a,a79932a,a79933a,a79936a,a79939a,a79940a,a79941a,a79945a,a79946a,a79949a,a79952a,a79953a,a79954a,a79958a,a79959a,a79962a,a79965a,a79966a,a79967a,a79971a,a79972a,a79975a,a79978a,a79979a,a79980a,a79984a,a79985a,a79988a,a79991a,a79992a,a79993a,a79997a,a79998a,a80001a,a80004a,a80005a,a80006a,a80010a,a80011a,a80014a,a80017a,a80018a,a80019a,a80023a,a80024a,a80027a,a80030a,a80031a,a80032a,a80036a,a80037a,a80040a,a80043a,a80044a,a80045a,a80049a,a80050a,a80053a,a80056a,a80057a,a80058a,a80062a,a80063a,a80066a,a80069a,a80070a,a80071a,a80075a,a80076a,a80079a,a80082a,a80083a,a80084a,a80088a,a80089a,a80092a,a80095a,a80096a,a80097a,a80101a,a80102a,a80105a,a80108a,a80109a,a80110a,a80114a,a80115a,a80118a,a80121a,a80122a,a80123a,a80127a,a80128a,a80131a,a80134a,a80135a,a80136a,a80140a,a80141a,a80144a,a80147a,a80148a,a80149a,a80153a,a80154a,a80157a,a80160a,a80161a,a80162a,a80166a,a80167a,a80170a,a80173a,a80174a,a80175a,a80179a,a80180a,a80183a,a80186a,a80187a,a80188a,a80192a,a80193a,a80196a,a80199a,a80200a,a80201a,a80205a,a80206a,a80209a,a80212a,a80213a,a80214a,a80218a,a80219a,a80222a,a80225a,a80226a,a80227a,a80231a,a80232a,a80235a,a80238a,a80239a,a80240a,a80244a,a80245a,a80248a,a80251a,a80252a,a80253a,a80257a,a80258a,a80261a,a80264a,a80265a,a80266a,a80270a,a80271a,a80274a,a80277a,a80278a,a80279a,a80283a,a80284a,a80287a,a80290a,a80291a,a80292a,a80296a,a80297a,a80300a,a80303a,a80304a,a80305a,a80309a,a80310a,a80313a,a80316a,a80317a,a80318a,a80322a,a80323a,a80326a,a80329a,a80330a,a80331a,a80335a,a80336a,a80339a,a80342a,a80343a,a80344a,a80348a,a80349a,a80352a,a80355a,a80356a,a80357a,a80361a,a80362a,a80365a,a80368a,a80369a,a80370a,a80374a,a80375a,a80378a,a80381a,a80382a,a80383a,a80387a,a80388a,a80391a,a80394a,a80395a,a80396a,a80400a,a80401a,a80404a,a80407a,a80408a,a80409a,a80413a,a80414a,a80417a,a80420a,a80421a,a80422a,a80426a,a80427a,a80430a,a80433a,a80434a,a80435a,a80439a,a80440a,a80443a,a80446a,a80447a,a80448a,a80452a,a80453a,a80456a,a80459a,a80460a,a80461a,a80465a,a80466a,a80469a,a80472a,a80473a,a80474a,a80478a,a80479a,a80482a,a80485a,a80486a,a80487a,a80491a,a80492a,a80495a,a80498a,a80499a,a80500a,a80504a,a80505a,a80508a,a80511a,a80512a,a80513a,a80517a,a80518a,a80521a,a80524a,a80525a,a80526a,a80530a,a80531a,a80534a,a80537a,a80538a,a80539a,a80543a,a80544a,a80547a,a80550a,a80551a,a80552a,a80556a,a80557a,a80560a,a80563a,a80564a,a80565a,a80569a,a80570a,a80573a,a80576a,a80577a,a80578a,a80582a,a80583a,a80586a,a80589a,a80590a,a80591a,a80595a,a80596a,a80599a,a80602a,a80603a,a80604a,a80608a,a80609a,a80612a,a80615a,a80616a,a80617a,a80621a,a80622a,a80625a,a80628a,a80629a,a80630a,a80634a,a80635a,a80638a,a80641a,a80642a,a80643a,a80647a,a80648a,a80651a,a80654a,a80655a,a80656a,a80660a,a80661a,a80664a,a80667a,a80668a,a80669a,a80673a,a80674a,a80677a,a80680a,a80681a,a80682a,a80686a,a80687a,a80690a,a80693a,a80694a,a80695a,a80699a,a80700a,a80703a,a80706a,a80707a,a80708a,a80712a,a80713a,a80716a,a80719a,a80720a,a80721a,a80725a,a80726a,a80729a,a80732a,a80733a,a80734a,a80738a,a80739a,a80742a,a80745a,a80746a,a80747a,a80751a,a80752a,a80755a,a80758a,a80759a,a80760a,a80764a,a80765a,a80768a,a80771a,a80772a,a80773a,a80777a,a80778a,a80781a,a80784a,a80785a,a80786a,a80790a,a80791a,a80794a,a80797a,a80798a,a80799a,a80803a,a80804a,a80807a,a80810a,a80811a,a80812a,a80816a,a80817a,a80820a,a80823a,a80824a,a80825a,a80829a,a80830a,a80833a,a80836a,a80837a,a80838a,a80842a,a80843a,a80846a,a80849a,a80850a,a80851a,a80855a,a80856a,a80859a,a80862a,a80863a,a80864a,a80868a,a80869a,a80872a,a80875a,a80876a,a80877a,a80881a,a80882a,a80885a,a80888a,a80889a,a80890a,a80894a,a80895a,a80898a,a80901a,a80902a,a80903a,a80907a,a80908a,a80911a,a80914a,a80915a,a80916a,a80920a,a80921a,a80924a,a80927a,a80928a,a80929a,a80933a,a80934a,a80937a,a80940a,a80941a,a80942a,a80946a,a80947a,a80950a,a80953a,a80954a,a80955a,a80959a,a80960a,a80963a,a80966a,a80967a,a80968a,a80972a,a80973a,a80976a,a80979a,a80980a,a80981a,a80985a,a80986a,a80989a,a80992a,a80993a,a80994a,a80998a,a80999a,a81002a,a81005a,a81006a,a81007a,a81011a,a81012a,a81015a,a81018a,a81019a,a81020a,a81024a,a81025a,a81028a,a81031a,a81032a,a81033a,a81037a,a81038a,a81041a,a81044a,a81045a,a81046a,a81050a,a81051a,a81054a,a81057a,a81058a,a81059a,a81063a,a81064a,a81067a,a81070a,a81071a,a81072a,a81076a,a81077a,a81080a,a81083a,a81084a,a81085a,a81089a,a81090a,a81093a,a81096a,a81097a,a81098a,a81102a,a81103a,a81106a,a81109a,a81110a,a81111a,a81115a,a81116a,a81119a,a81122a,a81123a,a81124a,a81128a,a81129a,a81132a,a81135a,a81136a,a81137a,a81141a,a81142a,a81145a,a81148a,a81149a,a81150a,a81154a,a81155a,a81158a,a81161a,a81162a,a81163a,a81167a,a81168a,a81171a,a81174a,a81175a,a81176a,a81180a,a81181a,a81184a,a81187a,a81188a,a81189a,a81193a,a81194a,a81197a,a81200a,a81201a,a81202a,a81206a,a81207a,a81210a,a81213a,a81214a,a81215a,a81219a,a81220a,a81223a,a81226a,a81227a,a81228a,a81232a,a81233a,a81236a,a81239a,a81240a,a81241a,a81245a,a81246a,a81249a,a81252a,a81253a,a81254a,a81258a,a81259a,a81262a,a81265a,a81266a,a81267a,a81271a,a81272a,a81275a,a81278a,a81279a,a81280a,a81284a,a81285a,a81288a,a81291a,a81292a,a81293a,a81297a,a81298a,a81301a,a81304a,a81305a,a81306a,a81310a,a81311a,a81314a,a81317a,a81318a,a81319a,a81323a,a81324a,a81327a,a81330a,a81331a,a81332a,a81336a,a81337a,a81340a,a81343a,a81344a,a81345a,a81349a,a81350a,a81353a,a81356a,a81357a,a81358a,a81362a,a81363a,a81366a,a81369a,a81370a,a81371a,a81375a,a81376a,a81379a,a81382a,a81383a,a81384a,a81388a,a81389a,a81392a,a81395a,a81396a,a81397a,a81401a,a81402a,a81405a,a81408a,a81409a,a81410a,a81414a,a81415a,a81418a,a81421a,a81422a,a81423a,a81427a,a81428a,a81431a,a81434a,a81435a,a81436a,a81440a,a81441a,a81444a,a81447a,a81448a,a81449a,a81453a,a81454a,a81457a,a81460a,a81461a,a81462a,a81466a,a81467a,a81470a,a81473a,a81474a,a81475a,a81479a,a81480a,a81483a,a81486a,a81487a,a81488a,a81492a,a81493a,a81496a,a81499a,a81500a,a81501a,a81505a,a81506a,a81509a,a81512a,a81513a,a81514a,a81518a,a81519a,a81522a,a81525a,a81526a,a81527a,a81531a,a81532a,a81535a,a81538a,a81539a,a81540a,a81544a,a81545a,a81548a,a81551a,a81552a,a81553a,a81557a,a81558a,a81561a,a81564a,a81565a,a81566a,a81570a,a81571a,a81574a,a81577a,a81578a,a81579a,a81583a,a81584a,a81587a,a81590a,a81591a,a81592a,a81596a,a81597a,a81600a,a81603a,a81604a,a81605a,a81609a,a81610a,a81613a,a81616a,a81617a,a81618a,a81622a,a81623a,a81626a,a81629a,a81630a,a81631a,a81635a,a81636a,a81639a,a81642a,a81643a,a81644a,a81648a,a81649a,a81652a,a81655a,a81656a,a81657a,a81661a,a81662a,a81665a,a81668a,a81669a,a81670a,a81674a,a81675a,a81678a,a81681a,a81682a,a81683a,a81687a,a81688a,a81691a,a81694a,a81695a,a81696a,a81700a,a81701a,a81704a,a81707a,a81708a,a81709a,a81713a,a81714a,a81717a,a81720a,a81721a,a81722a,a81726a,a81727a,a81730a,a81733a,a81734a,a81735a,a81739a,a81740a,a81743a,a81746a,a81747a,a81748a,a81752a,a81753a,a81756a,a81759a,a81760a,a81761a,a81765a,a81766a,a81769a,a81772a,a81773a,a81774a,a81778a,a81779a,a81782a,a81785a,a81786a,a81787a,a81791a,a81792a,a81795a,a81798a,a81799a,a81800a,a81804a,a81805a,a81808a,a81811a,a81812a,a81813a,a81817a,a81818a,a81821a,a81824a,a81825a,a81826a,a81830a,a81831a,a81834a,a81837a,a81838a,a81839a,a81843a,a81844a,a81847a,a81850a,a81851a,a81852a,a81856a,a81857a,a81860a,a81863a,a81864a,a81865a,a81869a,a81870a,a81873a,a81876a,a81877a,a81878a,a81882a,a81883a,a81886a,a81889a,a81890a,a81891a,a81895a,a81896a,a81899a,a81902a,a81903a,a81904a,a81908a,a81909a,a81912a,a81915a,a81916a,a81917a,a81921a,a81922a,a81925a,a81928a,a81929a,a81930a,a81934a,a81935a,a81938a,a81941a,a81942a,a81943a,a81947a,a81948a,a81951a,a81954a,a81955a,a81956a,a81960a,a81961a,a81964a,a81967a,a81968a,a81969a,a81973a,a81974a,a81977a,a81980a,a81981a,a81982a,a81986a,a81987a,a81990a,a81993a,a81994a,a81995a,a81999a,a82000a,a82003a,a82006a,a82007a,a82008a,a82012a,a82013a,a82016a,a82019a,a82020a,a82021a,a82025a,a82026a,a82029a,a82032a,a82033a,a82034a,a82038a,a82039a,a82042a,a82045a,a82046a,a82047a,a82051a,a82052a,a82055a,a82058a,a82059a,a82060a,a82064a,a82065a,a82068a,a82071a,a82072a,a82073a,a82077a,a82078a,a82081a,a82084a,a82085a,a82086a,a82090a,a82091a,a82094a,a82097a,a82098a,a82099a,a82103a,a82104a,a82107a,a82110a,a82111a,a82112a,a82116a,a82117a,a82120a,a82123a,a82124a,a82125a,a82129a,a82130a,a82133a,a82136a,a82137a,a82138a,a82142a,a82143a,a82146a,a82149a,a82150a,a82151a,a82155a,a82156a,a82159a,a82162a,a82163a,a82164a,a82168a,a82169a,a82172a,a82175a,a82176a,a82177a,a82181a,a82182a,a82185a,a82188a,a82189a,a82190a,a82194a,a82195a,a82198a,a82201a,a82202a,a82203a,a82207a,a82208a,a82211a,a82214a,a82215a,a82216a,a82220a,a82221a,a82224a,a82227a,a82228a,a82229a,a82233a,a82234a,a82237a,a82240a,a82241a,a82242a,a82246a,a82247a,a82250a,a82253a,a82254a,a82255a,a82259a,a82260a,a82263a,a82266a,a82267a,a82268a,a82272a,a82273a,a82276a,a82279a,a82280a,a82281a,a82285a,a82286a,a82289a,a82292a,a82293a,a82294a,a82298a,a82299a,a82302a,a82305a,a82306a,a82307a,a82311a,a82312a,a82315a,a82318a,a82319a,a82320a,a82324a,a82325a,a82328a,a82331a,a82332a,a82333a,a82337a,a82338a,a82341a,a82344a,a82345a,a82346a,a82350a,a82351a,a82354a,a82357a,a82358a,a82359a,a82363a,a82364a,a82367a,a82370a,a82371a,a82372a,a82376a,a82377a,a82380a,a82383a,a82384a,a82385a,a82389a,a82390a,a82393a,a82396a,a82397a,a82398a,a82402a,a82403a,a82406a,a82409a,a82410a,a82411a,a82415a,a82416a,a82419a,a82422a,a82423a,a82424a,a82428a,a82429a,a82432a,a82435a,a82436a,a82437a,a82441a,a82442a,a82445a,a82448a,a82449a,a82450a,a82454a,a82455a,a82458a,a82461a,a82462a,a82463a,a82467a,a82468a,a82471a,a82474a,a82475a,a82476a,a82480a,a82481a,a82484a,a82487a,a82488a,a82489a,a82493a,a82494a,a82497a,a82500a,a82501a,a82502a,a82506a,a82507a,a82510a,a82513a,a82514a,a82515a,a82519a,a82520a,a82523a,a82526a,a82527a,a82528a,a82532a,a82533a,a82536a,a82539a,a82540a,a82541a,a82545a,a82546a,a82549a,a82552a,a82553a,a82554a,a82558a,a82559a,a82562a,a82565a,a82566a,a82567a,a82571a,a82572a,a82575a,a82578a,a82579a,a82580a,a82584a,a82585a,a82588a,a82591a,a82592a,a82593a,a82597a,a82598a,a82601a,a82604a,a82605a,a82606a,a82610a,a82611a,a82614a,a82617a,a82618a,a82619a,a82623a,a82624a,a82627a,a82630a,a82631a,a82632a,a82636a,a82637a,a82640a,a82643a,a82644a,a82645a,a82649a,a82650a,a82653a,a82656a,a82657a,a82658a,a82662a,a82663a,a82666a,a82669a,a82670a,a82671a,a82675a,a82676a,a82679a,a82682a,a82683a,a82684a,a82688a,a82689a,a82692a,a82695a,a82696a,a82697a,a82701a,a82702a,a82705a,a82708a,a82709a,a82710a,a82714a,a82715a,a82718a,a82721a,a82722a,a82723a,a82727a,a82728a,a82731a,a82734a,a82735a,a82736a,a82740a,a82741a,a82744a,a82747a,a82748a,a82749a,a82753a,a82754a,a82757a,a82760a,a82761a,a82762a,a82766a,a82767a,a82770a,a82773a,a82774a,a82775a,a82779a,a82780a,a82783a,a82786a,a82787a,a82788a,a82792a,a82793a,a82796a,a82799a,a82800a,a82801a,a82805a,a82806a,a82809a,a82812a,a82813a,a82814a,a82818a,a82819a,a82822a,a82825a,a82826a,a82827a,a82831a,a82832a,a82835a,a82838a,a82839a,a82840a,a82844a,a82845a,a82848a,a82851a,a82852a,a82853a,a82857a,a82858a,a82861a,a82864a,a82865a,a82866a,a82870a,a82871a,a82874a,a82877a,a82878a,a82879a,a82883a,a82884a,a82887a,a82890a,a82891a,a82892a,a82896a,a82897a,a82900a,a82903a,a82904a,a82905a,a82909a,a82910a,a82913a,a82916a,a82917a,a82918a,a82922a,a82923a,a82926a,a82929a,a82930a,a82931a,a82935a,a82936a,a82939a,a82942a,a82943a,a82944a,a82948a,a82949a,a82952a,a82955a,a82956a,a82957a,a82961a,a82962a,a82965a,a82968a,a82969a,a82970a,a82974a,a82975a,a82978a,a82981a,a82982a,a82983a,a82987a,a82988a,a82991a,a82994a,a82995a,a82996a,a83000a,a83001a,a83004a,a83007a,a83008a,a83009a,a83013a,a83014a,a83017a,a83020a,a83021a,a83022a,a83026a,a83027a,a83030a,a83033a,a83034a,a83035a,a83039a,a83040a,a83043a,a83046a,a83047a,a83048a,a83052a,a83053a,a83056a,a83059a,a83060a,a83061a,a83065a,a83066a,a83069a,a83072a,a83073a,a83074a,a83078a,a83079a,a83082a,a83085a,a83086a,a83087a,a83091a,a83092a,a83095a,a83098a,a83099a,a83100a,a83104a,a83105a,a83108a,a83111a,a83112a,a83113a,a83117a,a83118a,a83121a,a83124a,a83125a,a83126a,a83130a,a83131a,a83134a,a83137a,a83138a,a83139a,a83143a,a83144a,a83147a,a83150a,a83151a,a83152a,a83156a,a83157a,a83160a,a83163a,a83164a,a83165a,a83169a,a83170a,a83173a,a83176a,a83177a,a83178a,a83182a,a83183a,a83186a,a83189a,a83190a,a83191a,a83195a,a83196a,a83199a,a83202a,a83203a,a83204a,a83208a,a83209a,a83212a,a83215a,a83216a,a83217a,a83221a,a83222a,a83225a,a83228a,a83229a,a83230a,a83234a,a83235a,a83238a,a83241a,a83242a,a83243a,a83247a,a83248a,a83251a,a83254a,a83255a,a83256a,a83260a,a83261a,a83264a,a83267a,a83268a,a83269a,a83273a,a83274a,a83277a,a83280a,a83281a,a83282a,a83286a,a83287a,a83290a,a83293a,a83294a,a83295a,a83299a,a83300a,a83303a,a83306a,a83307a,a83308a,a83312a,a83313a,a83316a,a83319a,a83320a,a83321a,a83325a,a83326a,a83329a,a83332a,a83333a,a83334a,a83338a,a83339a,a83342a,a83345a,a83346a,a83347a,a83351a,a83352a,a83355a,a83358a,a83359a,a83360a,a83364a,a83365a,a83368a,a83371a,a83372a,a83373a,a83377a,a83378a,a83381a,a83384a,a83385a,a83386a,a83390a,a83391a,a83394a,a83397a,a83398a,a83399a,a83403a,a83404a,a83407a,a83410a,a83411a,a83412a,a83416a,a83417a,a83420a,a83423a,a83424a,a83425a,a83429a,a83430a,a83433a,a83436a,a83437a,a83438a,a83442a,a83443a,a83446a,a83449a,a83450a,a83451a,a83455a,a83456a,a83459a,a83462a,a83463a,a83464a,a83468a,a83469a,a83472a,a83475a,a83476a,a83477a,a83481a,a83482a,a83485a,a83488a,a83489a,a83490a,a83494a,a83495a,a83498a,a83501a,a83502a,a83503a,a83507a,a83508a,a83511a,a83514a,a83515a,a83516a,a83520a,a83521a,a83524a,a83527a,a83528a,a83529a,a83533a,a83534a,a83537a,a83540a,a83541a,a83542a,a83546a,a83547a,a83550a,a83553a,a83554a,a83555a,a83559a,a83560a,a83563a,a83566a,a83567a,a83568a,a83572a,a83573a,a83576a,a83579a,a83580a,a83581a,a83585a,a83586a,a83589a,a83592a,a83593a,a83594a,a83598a,a83599a,a83602a,a83605a,a83606a,a83607a,a83611a,a83612a,a83615a,a83618a,a83619a,a83620a,a83624a,a83625a,a83628a,a83631a,a83632a,a83633a,a83637a,a83638a,a83641a,a83644a,a83645a,a83646a,a83650a,a83651a,a83654a,a83657a,a83658a,a83659a,a83663a,a83664a,a83667a,a83670a,a83671a,a83672a,a83676a,a83677a,a83680a,a83683a,a83684a,a83685a,a83689a,a83690a,a83693a,a83696a,a83697a,a83698a,a83702a,a83703a,a83706a,a83709a,a83710a,a83711a,a83715a,a83716a,a83719a,a83722a,a83723a,a83724a,a83728a,a83729a,a83732a,a83735a,a83736a,a83737a,a83741a,a83742a,a83745a,a83748a,a83749a,a83750a,a83754a,a83755a,a83758a,a83761a,a83762a,a83763a,a83767a,a83768a,a83771a,a83774a,a83775a,a83776a,a83780a,a83781a,a83784a,a83787a,a83788a,a83789a,a83793a,a83794a,a83797a,a83800a,a83801a,a83802a,a83806a,a83807a,a83810a,a83813a,a83814a,a83815a,a83819a,a83820a,a83823a,a83826a,a83827a,a83828a,a83832a,a83833a,a83836a,a83839a,a83840a,a83841a,a83845a,a83846a,a83849a,a83852a,a83853a,a83854a,a83858a,a83859a,a83862a,a83865a,a83866a,a83867a,a83871a,a83872a,a83875a,a83878a,a83879a,a83880a,a83884a,a83885a,a83888a,a83891a,a83892a,a83893a,a83897a,a83898a,a83901a,a83904a,a83905a,a83906a,a83910a,a83911a,a83914a,a83917a,a83918a,a83919a,a83923a,a83924a,a83927a,a83930a,a83931a,a83932a,a83936a,a83937a,a83940a,a83943a,a83944a,a83945a,a83949a,a83950a,a83953a,a83956a,a83957a,a83958a,a83962a,a83963a,a83966a,a83969a,a83970a,a83971a,a83975a,a83976a,a83979a,a83982a,a83983a,a83984a,a83988a,a83989a,a83992a,a83995a,a83996a,a83997a,a84001a,a84002a,a84005a,a84008a,a84009a,a84010a,a84014a,a84015a,a84018a,a84021a,a84022a,a84023a,a84027a,a84028a,a84031a,a84034a,a84035a,a84036a,a84040a,a84041a,a84044a,a84047a,a84048a,a84049a,a84053a,a84054a,a84057a,a84060a,a84061a,a84062a,a84066a,a84067a,a84070a,a84073a,a84074a,a84075a,a84079a,a84080a,a84083a,a84086a,a84087a,a84088a,a84092a,a84093a,a84096a,a84099a,a84100a,a84101a,a84105a,a84106a,a84109a,a84112a,a84113a,a84114a,a84118a,a84119a,a84122a,a84125a,a84126a,a84127a,a84131a,a84132a,a84135a,a84138a,a84139a,a84140a,a84144a,a84145a,a84148a,a84151a,a84152a,a84153a,a84157a,a84158a,a84161a,a84164a,a84165a,a84166a,a84170a,a84171a,a84174a,a84177a,a84178a,a84179a,a84183a,a84184a,a84187a,a84190a,a84191a,a84192a,a84196a,a84197a,a84200a,a84203a,a84204a,a84205a,a84209a,a84210a,a84213a,a84216a,a84217a,a84218a,a84222a,a84223a,a84226a,a84229a,a84230a,a84231a,a84235a,a84236a,a84239a,a84242a,a84243a,a84244a,a84248a,a84249a,a84252a,a84255a,a84256a,a84257a,a84261a,a84262a,a84265a,a84268a,a84269a,a84270a,a84274a,a84275a,a84278a,a84281a,a84282a,a84283a,a84287a,a84288a,a84291a,a84294a,a84295a,a84296a,a84300a,a84301a,a84304a,a84307a,a84308a,a84309a,a84313a,a84314a,a84317a,a84320a,a84321a,a84322a,a84326a,a84327a,a84330a,a84333a,a84334a,a84335a,a84339a,a84340a,a84343a,a84346a,a84347a,a84348a,a84352a,a84353a,a84356a,a84359a,a84360a,a84361a,a84365a,a84366a,a84369a,a84372a,a84373a,a84374a,a84378a,a84379a,a84382a,a84385a,a84386a,a84387a,a84391a,a84392a,a84395a,a84398a,a84399a,a84400a,a84404a,a84405a,a84408a,a84411a,a84412a,a84413a,a84417a,a84418a,a84421a,a84424a,a84425a,a84426a,a84430a,a84431a,a84434a,a84437a,a84438a,a84439a,a84443a,a84444a,a84447a,a84450a,a84451a,a84452a,a84456a,a84457a,a84460a,a84463a,a84464a,a84465a,a84469a,a84470a,a84473a,a84476a,a84477a,a84478a,a84482a,a84483a,a84486a,a84489a,a84490a,a84491a,a84495a,a84496a,a84499a,a84502a,a84503a,a84504a,a84508a,a84509a,a84512a,a84515a,a84516a,a84517a,a84521a,a84522a,a84525a,a84528a,a84529a,a84530a,a84534a,a84535a,a84538a,a84541a,a84542a,a84543a,a84547a,a84548a,a84551a,a84554a,a84555a,a84556a,a84560a,a84561a,a84564a,a84567a,a84568a,a84569a,a84573a,a84574a,a84577a,a84580a,a84581a,a84582a,a84586a,a84587a,a84590a,a84593a,a84594a,a84595a,a84599a,a84600a,a84603a,a84606a,a84607a,a84608a,a84612a,a84613a,a84616a,a84619a,a84620a,a84621a,a84625a,a84626a,a84629a,a84632a,a84633a,a84634a,a84638a,a84639a,a84642a,a84645a,a84646a,a84647a,a84651a,a84652a,a84655a,a84658a,a84659a,a84660a,a84664a,a84665a,a84668a,a84671a,a84672a,a84673a,a84677a,a84678a,a84681a,a84684a,a84685a,a84686a,a84690a,a84691a,a84694a,a84697a,a84698a,a84699a,a84703a,a84704a,a84707a,a84710a,a84711a,a84712a,a84716a,a84717a,a84720a,a84723a,a84724a,a84725a,a84729a,a84730a,a84733a,a84736a,a84737a,a84738a,a84742a,a84743a,a84746a,a84749a,a84750a,a84751a,a84755a,a84756a,a84759a,a84762a,a84763a,a84764a,a84768a,a84769a,a84772a,a84775a,a84776a,a84777a,a84781a,a84782a,a84785a,a84788a,a84789a,a84790a,a84794a,a84795a,a84798a,a84801a,a84802a,a84803a,a84807a,a84808a,a84811a,a84814a,a84815a,a84816a,a84820a,a84821a,a84824a,a84827a,a84828a,a84829a,a84833a,a84834a,a84837a,a84840a,a84841a,a84842a,a84846a,a84847a,a84850a,a84853a,a84854a,a84855a,a84859a,a84860a,a84863a,a84866a,a84867a,a84868a,a84872a,a84873a,a84876a,a84879a,a84880a,a84881a,a84885a,a84886a,a84889a,a84892a,a84893a,a84894a,a84898a,a84899a,a84902a,a84905a,a84906a,a84907a,a84911a,a84912a,a84915a,a84918a,a84919a,a84920a,a84924a,a84925a,a84928a,a84931a,a84932a,a84933a,a84937a,a84938a,a84941a,a84944a,a84945a,a84946a,a84950a,a84951a,a84954a,a84957a,a84958a,a84959a,a84963a,a84964a,a84967a,a84970a,a84971a,a84972a,a84976a,a84977a,a84980a,a84983a,a84984a,a84985a,a84989a,a84990a,a84993a,a84996a,a84997a,a84998a,a85002a,a85003a,a85006a,a85009a,a85010a,a85011a,a85015a,a85016a,a85019a,a85022a,a85023a,a85024a,a85028a,a85029a,a85032a,a85035a,a85036a,a85037a,a85041a,a85042a,a85045a,a85048a,a85049a,a85050a,a85054a,a85055a,a85058a,a85061a,a85062a,a85063a,a85067a,a85068a,a85071a,a85074a,a85075a,a85076a,a85080a,a85081a,a85084a,a85087a,a85088a,a85089a,a85093a,a85094a,a85097a,a85100a,a85101a,a85102a,a85106a,a85107a,a85110a,a85113a,a85114a,a85115a,a85119a,a85120a,a85123a,a85126a,a85127a,a85128a,a85132a,a85133a,a85136a,a85139a,a85140a,a85141a,a85145a,a85146a,a85149a,a85152a,a85153a,a85154a,a85158a,a85159a,a85162a,a85165a,a85166a,a85167a,a85171a,a85172a,a85175a,a85178a,a85179a,a85180a,a85184a,a85185a,a85188a,a85191a,a85192a,a85193a,a85197a,a85198a,a85201a,a85204a,a85205a,a85206a,a85210a,a85211a,a85214a,a85217a,a85218a,a85219a,a85223a,a85224a,a85227a,a85230a,a85231a,a85232a,a85236a,a85237a,a85240a,a85243a,a85244a,a85245a,a85249a,a85250a,a85253a,a85256a,a85257a,a85258a,a85262a,a85263a,a85266a,a85269a,a85270a,a85271a,a85275a,a85276a,a85279a,a85282a,a85283a,a85284a,a85288a,a85289a,a85292a,a85295a,a85296a,a85297a,a85301a,a85302a,a85305a,a85308a,a85309a,a85310a,a85314a,a85315a,a85318a,a85321a,a85322a,a85323a,a85327a,a85328a,a85331a,a85334a,a85335a,a85336a,a85340a,a85341a,a85344a,a85347a,a85348a,a85349a,a85353a,a85354a,a85357a,a85360a,a85361a,a85362a,a85366a,a85367a,a85370a,a85373a,a85374a,a85375a,a85379a,a85380a,a85383a,a85386a,a85387a,a85388a,a85392a,a85393a,a85396a,a85399a,a85400a,a85401a,a85405a,a85406a,a85409a,a85412a,a85413a,a85414a,a85418a,a85419a,a85422a,a85425a,a85426a,a85427a,a85431a,a85432a,a85435a,a85438a,a85439a,a85440a,a85444a,a85445a,a85448a,a85451a,a85452a,a85453a,a85457a,a85458a,a85461a,a85464a,a85465a,a85466a,a85470a,a85471a,a85474a,a85477a,a85478a,a85479a,a85483a,a85484a,a85487a,a85490a,a85491a,a85492a,a85496a,a85497a,a85500a,a85503a,a85504a,a85505a,a85509a,a85510a,a85513a,a85516a,a85517a,a85518a,a85522a,a85523a,a85526a,a85529a,a85530a,a85531a,a85535a,a85536a,a85539a,a85542a,a85543a,a85544a,a85548a,a85549a,a85552a,a85555a,a85556a,a85557a,a85561a,a85562a,a85565a,a85568a,a85569a,a85570a,a85574a,a85575a,a85578a,a85581a,a85582a,a85583a,a85587a,a85588a,a85591a,a85594a,a85595a,a85596a,a85600a,a85601a,a85604a,a85607a,a85608a,a85609a,a85613a,a85614a,a85617a,a85620a,a85621a,a85622a,a85626a,a85627a,a85630a,a85633a,a85634a,a85635a,a85639a,a85640a,a85643a,a85646a,a85647a,a85648a,a85652a,a85653a,a85656a,a85659a,a85660a,a85661a,a85665a,a85666a,a85669a,a85672a,a85673a,a85674a,a85678a,a85679a,a85682a,a85685a,a85686a,a85687a,a85691a,a85692a,a85695a,a85698a,a85699a,a85700a,a85704a,a85705a,a85708a,a85711a,a85712a,a85713a,a85717a,a85718a,a85721a,a85724a,a85725a,a85726a,a85730a,a85731a,a85734a,a85737a,a85738a,a85739a,a85743a,a85744a,a85747a,a85750a,a85751a,a85752a,a85756a,a85757a,a85760a,a85763a,a85764a,a85765a,a85769a,a85770a,a85773a,a85776a,a85777a,a85778a,a85782a,a85783a,a85786a,a85789a,a85790a,a85791a,a85795a,a85796a,a85799a,a85802a,a85803a,a85804a,a85808a,a85809a,a85812a,a85815a,a85816a,a85817a,a85821a,a85822a,a85825a,a85828a,a85829a,a85830a,a85834a,a85835a,a85838a,a85841a,a85842a,a85843a,a85847a,a85848a,a85851a,a85854a,a85855a,a85856a,a85860a,a85861a,a85864a,a85867a,a85868a,a85869a,a85873a,a85874a,a85877a,a85880a,a85881a,a85882a,a85886a,a85887a,a85890a,a85893a,a85894a,a85895a,a85899a,a85900a,a85903a,a85906a,a85907a,a85908a,a85912a,a85913a,a85916a,a85919a,a85920a,a85921a,a85925a,a85926a,a85929a,a85932a,a85933a,a85934a,a85938a,a85939a,a85942a,a85945a,a85946a,a85947a,a85951a,a85952a,a85955a,a85958a,a85959a,a85960a,a85964a,a85965a,a85968a,a85971a,a85972a,a85973a,a85977a,a85978a,a85981a,a85984a,a85985a,a85986a,a85990a,a85991a,a85994a,a85997a,a85998a,a85999a,a86003a,a86004a,a86007a,a86010a,a86011a,a86012a,a86016a,a86017a,a86020a,a86023a,a86024a,a86025a,a86029a,a86030a,a86033a,a86036a,a86037a,a86038a,a86042a,a86043a,a86046a,a86049a,a86050a,a86051a,a86055a,a86056a,a86059a,a86062a,a86063a,a86064a,a86068a,a86069a,a86072a,a86075a,a86076a,a86077a,a86081a,a86082a,a86085a,a86088a,a86089a,a86090a,a86094a,a86095a,a86098a,a86101a,a86102a,a86103a,a86107a,a86108a,a86111a,a86114a,a86115a,a86116a,a86120a,a86121a,a86124a,a86127a,a86128a,a86129a,a86133a,a86134a,a86137a,a86140a,a86141a,a86142a,a86146a,a86147a,a86150a,a86153a,a86154a,a86155a,a86159a,a86160a,a86163a,a86166a,a86167a,a86168a,a86172a,a86173a,a86176a,a86179a,a86180a,a86181a,a86185a,a86186a,a86189a,a86192a,a86193a,a86194a,a86198a,a86199a,a86202a,a86205a,a86206a,a86207a,a86211a,a86212a,a86215a,a86218a,a86219a,a86220a,a86224a,a86225a,a86228a,a86231a,a86232a,a86233a,a86237a,a86238a,a86241a,a86244a,a86245a,a86246a,a86250a,a86251a,a86254a,a86257a,a86258a,a86259a,a86263a,a86264a,a86267a,a86270a,a86271a,a86272a,a86276a,a86277a,a86280a,a86283a,a86284a,a86285a,a86289a,a86290a,a86293a,a86296a,a86297a,a86298a,a86302a,a86303a,a86306a,a86309a,a86310a,a86311a,a86315a,a86316a,a86319a,a86322a,a86323a,a86324a,a86328a,a86329a,a86332a,a86335a,a86336a,a86337a,a86341a,a86342a,a86345a,a86348a,a86349a,a86350a,a86354a,a86355a,a86358a,a86361a,a86362a,a86363a,a86367a,a86368a,a86371a,a86374a,a86375a,a86376a,a86380a,a86381a,a86384a,a86387a,a86388a,a86389a,a86393a,a86394a,a86397a,a86400a,a86401a,a86402a,a86406a,a86407a,a86410a,a86413a,a86414a,a86415a,a86419a,a86420a,a86423a,a86426a,a86427a,a86428a,a86432a,a86433a,a86436a,a86439a,a86440a,a86441a,a86445a,a86446a,a86449a,a86452a,a86453a,a86454a,a86458a,a86459a,a86462a,a86465a,a86466a,a86467a,a86471a,a86472a,a86475a,a86478a,a86479a,a86480a,a86484a,a86485a,a86488a,a86491a,a86492a,a86493a,a86497a,a86498a,a86501a,a86504a,a86505a,a86506a,a86510a,a86511a,a86514a,a86517a,a86518a,a86519a,a86523a,a86524a,a86527a,a86530a,a86531a,a86532a,a86536a,a86537a,a86540a,a86543a,a86544a,a86545a,a86549a,a86550a,a86553a,a86556a,a86557a,a86558a,a86562a,a86563a,a86566a,a86569a,a86570a,a86571a,a86575a,a86576a,a86579a,a86582a,a86583a,a86584a,a86588a,a86589a,a86592a,a86595a,a86596a,a86597a,a86601a,a86602a,a86605a,a86608a,a86609a,a86610a,a86614a,a86615a,a86618a,a86621a,a86622a,a86623a,a86627a,a86628a,a86631a,a86634a,a86635a,a86636a,a86640a,a86641a,a86644a,a86647a,a86648a,a86649a,a86653a,a86654a,a86657a,a86660a,a86661a,a86662a,a86666a,a86667a,a86670a,a86673a,a86674a,a86675a,a86679a,a86680a,a86683a,a86686a,a86687a,a86688a,a86692a,a86693a,a86696a,a86699a,a86700a,a86701a,a86705a,a86706a,a86709a,a86712a,a86713a,a86714a,a86718a,a86719a,a86722a,a86725a,a86726a,a86727a,a86731a,a86732a,a86735a,a86738a,a86739a,a86740a,a86744a,a86745a,a86748a,a86751a,a86752a,a86753a,a86757a,a86758a,a86761a,a86764a,a86765a,a86766a,a86770a,a86771a,a86774a,a86777a,a86778a,a86779a,a86783a,a86784a,a86787a,a86790a,a86791a,a86792a,a86796a,a86797a,a86800a,a86803a,a86804a,a86805a,a86809a,a86810a,a86813a,a86816a,a86817a,a86818a,a86822a,a86823a,a86826a,a86829a,a86830a,a86831a,a86835a,a86836a,a86839a,a86842a,a86843a,a86844a,a86848a,a86849a,a86852a,a86855a,a86856a,a86857a,a86861a,a86862a,a86865a,a86868a,a86869a,a86870a,a86874a,a86875a,a86878a,a86881a,a86882a,a86883a,a86887a,a86888a,a86891a,a86894a,a86895a,a86896a,a86900a,a86901a,a86904a,a86907a,a86908a,a86909a,a86913a,a86914a,a86917a,a86920a,a86921a,a86922a,a86926a,a86927a,a86930a,a86933a,a86934a,a86935a,a86939a,a86940a,a86943a,a86946a,a86947a,a86948a,a86952a,a86953a,a86956a,a86959a,a86960a,a86961a,a86965a,a86966a,a86969a,a86972a,a86973a,a86974a,a86978a,a86979a,a86982a,a86985a,a86986a,a86987a,a86991a,a86992a,a86995a,a86998a,a86999a,a87000a,a87004a,a87005a,a87008a,a87011a,a87012a,a87013a,a87017a,a87018a,a87021a,a87024a,a87025a,a87026a,a87030a,a87031a,a87034a,a87037a,a87038a,a87039a,a87043a,a87044a,a87047a,a87050a,a87051a,a87052a,a87056a,a87057a,a87060a,a87063a,a87064a,a87065a,a87069a,a87070a,a87073a,a87076a,a87077a,a87078a,a87082a,a87083a,a87086a,a87089a,a87090a,a87091a,a87095a,a87096a,a87099a,a87102a,a87103a,a87104a,a87108a,a87109a,a87112a,a87115a,a87116a,a87117a,a87121a,a87122a,a87125a,a87128a,a87129a,a87130a,a87134a,a87135a,a87138a,a87141a,a87142a,a87143a,a87147a,a87148a,a87151a,a87154a,a87155a,a87156a,a87160a,a87161a,a87164a,a87167a,a87168a,a87169a,a87173a,a87174a,a87177a,a87180a,a87181a,a87182a,a87186a,a87187a,a87190a,a87193a,a87194a,a87195a,a87199a,a87200a,a87203a,a87206a,a87207a,a87208a,a87212a,a87213a,a87216a,a87219a,a87220a,a87221a,a87225a,a87226a,a87229a,a87232a,a87233a,a87234a,a87238a,a87239a,a87242a,a87245a,a87246a,a87247a,a87251a,a87252a,a87255a,a87258a,a87259a,a87260a,a87264a,a87265a,a87268a,a87271a,a87272a,a87273a,a87277a,a87278a,a87281a,a87284a,a87285a,a87286a,a87290a,a87291a,a87294a,a87297a,a87298a,a87299a,a87303a,a87304a,a87307a,a87310a,a87311a,a87312a,a87316a,a87317a,a87320a,a87323a,a87324a,a87325a,a87329a,a87330a,a87333a,a87336a,a87337a,a87338a,a87342a,a87343a,a87346a,a87349a,a87350a,a87351a,a87355a,a87356a,a87359a,a87362a,a87363a,a87364a,a87368a,a87369a,a87372a,a87375a,a87376a,a87377a,a87381a,a87382a,a87385a,a87388a,a87389a,a87390a,a87394a,a87395a,a87398a,a87401a,a87402a,a87403a,a87407a,a87408a,a87411a,a87414a,a87415a,a87416a,a87420a,a87421a,a87424a,a87427a,a87428a,a87429a,a87433a,a87434a,a87437a,a87440a,a87441a,a87442a,a87446a,a87447a,a87450a,a87453a,a87454a,a87455a,a87459a,a87460a,a87463a,a87466a,a87467a,a87468a,a87472a,a87473a,a87476a,a87479a,a87480a,a87481a,a87485a,a87486a,a87489a,a87492a,a87493a,a87494a,a87498a,a87499a,a87502a,a87505a,a87506a,a87507a,a87511a,a87512a,a87515a,a87518a,a87519a,a87520a,a87524a,a87525a,a87528a,a87531a,a87532a,a87533a,a87537a,a87538a,a87541a,a87544a,a87545a,a87546a,a87550a,a87551a,a87554a,a87557a,a87558a,a87559a,a87563a,a87564a,a87567a,a87570a,a87571a,a87572a,a87576a,a87577a,a87580a,a87583a,a87584a,a87585a,a87589a,a87590a,a87593a,a87596a,a87597a,a87598a,a87602a,a87603a,a87606a,a87609a,a87610a,a87611a,a87615a,a87616a,a87619a,a87622a,a87623a,a87624a,a87628a,a87629a,a87632a,a87635a,a87636a,a87637a,a87641a,a87642a,a87645a,a87648a,a87649a,a87650a,a87654a,a87655a,a87658a,a87661a,a87662a,a87663a,a87667a,a87668a,a87671a,a87674a,a87675a,a87676a,a87680a,a87681a,a87684a,a87687a,a87688a,a87689a,a87693a,a87694a,a87697a,a87700a,a87701a,a87702a,a87706a,a87707a,a87710a,a87713a,a87714a,a87715a,a87719a,a87720a,a87723a,a87726a,a87727a,a87728a,a87732a,a87733a,a87736a,a87739a,a87740a,a87741a,a87745a,a87746a,a87749a,a87752a,a87753a,a87754a,a87758a,a87759a,a87762a,a87765a,a87766a,a87767a,a87771a,a87772a,a87775a,a87778a,a87779a,a87780a,a87784a,a87785a,a87788a,a87791a,a87792a,a87793a,a87797a,a87798a,a87801a,a87804a,a87805a,a87806a,a87810a,a87811a,a87814a,a87817a,a87818a,a87819a,a87823a,a87824a,a87827a,a87830a,a87831a,a87832a,a87836a,a87837a,a87840a,a87843a,a87844a,a87845a,a87849a,a87850a,a87853a,a87856a,a87857a,a87858a,a87862a,a87863a,a87866a,a87869a,a87870a,a87871a,a87875a,a87876a,a87879a,a87882a,a87883a,a87884a,a87888a,a87889a,a87892a,a87895a,a87896a,a87897a,a87901a,a87902a,a87905a,a87908a,a87909a,a87910a,a87914a,a87915a,a87918a,a87921a,a87922a,a87923a,a87927a,a87928a,a87931a,a87934a,a87935a,a87936a,a87940a,a87941a,a87944a,a87947a,a87948a,a87949a,a87953a,a87954a,a87957a,a87960a,a87961a,a87962a,a87966a,a87967a,a87970a,a87973a,a87974a,a87975a,a87979a,a87980a,a87983a,a87986a,a87987a,a87988a,a87992a,a87993a,a87996a,a87999a,a88000a,a88001a,a88005a,a88006a,a88009a,a88012a,a88013a,a88014a,a88018a,a88019a,a88022a,a88025a,a88026a,a88027a,a88031a,a88032a,a88035a,a88038a,a88039a,a88040a,a88044a,a88045a,a88048a,a88051a,a88052a,a88053a,a88057a,a88058a,a88061a,a88064a,a88065a,a88066a,a88070a,a88071a,a88074a,a88077a,a88078a,a88079a,a88083a,a88084a,a88087a,a88090a,a88091a,a88092a,a88096a,a88097a,a88100a,a88103a,a88104a,a88105a,a88109a,a88110a,a88113a,a88116a,a88117a,a88118a,a88122a,a88123a,a88126a,a88129a,a88130a,a88131a,a88135a,a88136a,a88139a,a88142a,a88143a,a88144a,a88148a,a88149a,a88152a,a88155a,a88156a,a88157a,a88161a,a88162a,a88165a,a88168a,a88169a,a88170a,a88174a,a88175a,a88178a,a88181a,a88182a,a88183a,a88187a,a88188a,a88191a,a88194a,a88195a,a88196a,a88200a,a88201a,a88204a,a88207a,a88208a,a88209a,a88213a,a88214a,a88217a,a88220a,a88221a,a88222a,a88226a,a88227a,a88230a,a88233a,a88234a,a88235a,a88239a,a88240a,a88243a,a88246a,a88247a,a88248a,a88252a,a88253a,a88256a,a88259a,a88260a,a88261a,a88265a,a88266a,a88269a,a88272a,a88273a,a88274a,a88278a,a88279a,a88282a,a88285a,a88286a,a88287a,a88291a,a88292a,a88295a,a88298a,a88299a,a88300a,a88304a,a88305a,a88308a,a88311a,a88312a,a88313a,a88317a,a88318a,a88321a,a88324a,a88325a,a88326a,a88330a,a88331a,a88334a,a88337a,a88338a,a88339a,a88343a,a88344a,a88347a,a88350a,a88351a,a88352a,a88356a,a88357a,a88360a,a88363a,a88364a,a88365a,a88369a,a88370a,a88373a,a88376a,a88377a,a88378a,a88382a,a88383a,a88386a,a88389a,a88390a,a88391a,a88395a,a88396a,a88399a,a88402a,a88403a,a88404a,a88408a,a88409a,a88412a,a88415a,a88416a,a88417a,a88421a,a88422a,a88425a,a88428a,a88429a,a88430a,a88434a,a88435a,a88438a,a88441a,a88442a,a88443a,a88447a,a88448a,a88451a,a88454a,a88455a,a88456a,a88460a,a88461a,a88464a,a88467a,a88468a,a88469a,a88473a,a88474a,a88477a,a88480a,a88481a,a88482a,a88486a,a88487a,a88490a,a88493a,a88494a,a88495a,a88499a,a88500a,a88503a,a88506a,a88507a,a88508a,a88512a,a88513a,a88516a,a88519a,a88520a,a88521a,a88525a,a88526a,a88529a,a88532a,a88533a,a88534a,a88538a,a88539a,a88542a,a88545a,a88546a,a88547a,a88551a,a88552a,a88555a,a88558a,a88559a,a88560a,a88564a,a88565a,a88568a,a88571a,a88572a,a88573a,a88577a,a88578a,a88581a,a88584a,a88585a,a88586a,a88590a,a88591a,a88594a,a88597a,a88598a,a88599a,a88603a,a88604a,a88607a,a88610a,a88611a,a88612a,a88616a,a88617a,a88620a,a88623a,a88624a,a88625a,a88629a,a88630a,a88633a,a88636a,a88637a,a88638a,a88642a,a88643a,a88646a,a88649a,a88650a,a88651a,a88655a,a88656a,a88659a,a88662a,a88663a,a88664a,a88668a,a88669a,a88672a,a88675a,a88676a,a88677a,a88681a,a88682a,a88685a,a88688a,a88689a,a88690a,a88694a,a88695a,a88698a,a88701a,a88702a,a88703a,a88707a,a88708a,a88711a,a88714a,a88715a,a88716a,a88720a,a88721a,a88724a,a88727a,a88728a,a88729a,a88733a,a88734a,a88737a,a88740a,a88741a,a88742a,a88746a,a88747a,a88750a,a88753a,a88754a,a88755a,a88759a,a88760a,a88763a,a88766a,a88767a,a88768a,a88772a,a88773a,a88776a,a88779a,a88780a,a88781a,a88785a,a88786a,a88789a,a88792a,a88793a,a88794a,a88798a,a88799a,a88802a,a88805a,a88806a,a88807a,a88811a,a88812a,a88815a,a88818a,a88819a,a88820a,a88824a,a88825a,a88828a,a88831a,a88832a,a88833a,a88837a,a88838a,a88841a,a88844a,a88845a,a88846a,a88850a,a88851a,a88854a,a88857a,a88858a,a88859a,a88863a,a88864a,a88867a,a88870a,a88871a,a88872a,a88876a,a88877a,a88880a,a88883a,a88884a,a88885a,a88889a,a88890a,a88893a,a88896a,a88897a,a88898a,a88902a,a88903a,a88906a,a88909a,a88910a,a88911a,a88915a,a88916a,a88919a,a88922a,a88923a,a88924a,a88928a,a88929a,a88932a,a88935a,a88936a,a88937a,a88941a,a88942a,a88945a,a88948a,a88949a,a88950a,a88954a,a88955a,a88958a,a88961a,a88962a,a88963a,a88967a,a88968a,a88971a,a88974a,a88975a,a88976a,a88980a,a88981a,a88984a,a88987a,a88988a,a88989a,a88993a,a88994a,a88997a,a89000a,a89001a,a89002a,a89006a,a89007a,a89010a,a89013a,a89014a,a89015a,a89019a,a89020a,a89023a,a89026a,a89027a,a89028a,a89032a,a89033a,a89036a,a89039a,a89040a,a89041a,a89045a,a89046a,a89049a,a89052a,a89053a,a89054a,a89058a,a89059a,a89062a,a89065a,a89066a,a89067a,a89071a,a89072a,a89075a,a89078a,a89079a,a89080a,a89084a,a89085a,a89088a,a89091a,a89092a,a89093a,a89097a,a89098a,a89101a,a89104a,a89105a,a89106a,a89110a,a89111a,a89114a,a89117a,a89118a,a89119a,a89123a,a89124a,a89127a,a89130a,a89131a,a89132a,a89136a,a89137a,a89140a,a89143a,a89144a,a89145a,a89149a,a89150a,a89153a,a89156a,a89157a,a89158a,a89162a,a89163a,a89166a,a89169a,a89170a,a89171a,a89175a,a89176a,a89179a,a89182a,a89183a,a89184a,a89188a,a89189a,a89192a,a89195a,a89196a,a89197a,a89201a,a89202a,a89205a,a89208a,a89209a,a89210a,a89214a,a89215a,a89218a,a89221a,a89222a,a89223a,a89227a,a89228a,a89231a,a89234a,a89235a,a89236a,a89240a,a89241a,a89244a,a89247a,a89248a,a89249a,a89253a,a89254a,a89257a,a89260a,a89261a,a89262a,a89266a,a89267a,a89270a,a89273a,a89274a,a89275a,a89279a,a89280a,a89283a,a89286a,a89287a,a89288a,a89292a,a89293a,a89296a,a89299a,a89300a,a89301a,a89305a,a89306a,a89309a,a89312a,a89313a,a89314a,a89318a,a89319a,a89322a,a89325a,a89326a,a89327a,a89331a,a89332a,a89335a,a89338a,a89339a,a89340a,a89344a,a89345a,a89348a,a89351a,a89352a,a89353a,a89357a,a89358a,a89361a,a89364a,a89365a,a89366a,a89370a,a89371a,a89374a,a89377a,a89378a,a89379a,a89383a,a89384a,a89387a,a89390a,a89391a,a89392a,a89396a,a89397a,a89400a,a89403a,a89404a,a89405a,a89409a,a89410a,a89413a,a89416a,a89417a,a89418a,a89422a,a89423a,a89426a,a89429a,a89430a,a89431a,a89435a,a89436a,a89439a,a89442a,a89443a,a89444a,a89448a,a89449a,a89452a,a89455a,a89456a,a89457a,a89461a,a89462a,a89465a,a89468a,a89469a,a89470a,a89474a,a89475a,a89478a,a89481a,a89482a,a89483a,a89487a,a89488a,a89491a,a89494a,a89495a,a89496a,a89500a,a89501a,a89504a,a89507a,a89508a,a89509a,a89513a,a89514a,a89517a,a89520a,a89521a,a89522a,a89526a,a89527a,a89530a,a89533a,a89534a,a89535a,a89539a,a89540a,a89543a,a89546a,a89547a,a89548a,a89552a,a89553a,a89556a,a89559a,a89560a,a89561a,a89565a,a89566a,a89569a,a89572a,a89573a,a89574a,a89578a,a89579a,a89582a,a89585a,a89586a,a89587a,a89591a,a89592a,a89595a,a89598a,a89599a,a89600a,a89604a,a89605a,a89608a,a89611a,a89612a,a89613a,a89617a,a89618a,a89621a,a89624a,a89625a,a89626a,a89630a,a89631a,a89634a,a89637a,a89638a,a89639a,a89643a,a89644a,a89647a,a89650a,a89651a,a89652a,a89656a,a89657a,a89660a,a89663a,a89664a,a89665a,a89669a,a89670a,a89673a,a89676a,a89677a,a89678a,a89682a,a89683a,a89686a,a89689a,a89690a,a89691a,a89695a,a89696a,a89699a,a89702a,a89703a,a89704a,a89708a,a89709a,a89712a,a89715a,a89716a,a89717a,a89721a,a89722a,a89725a,a89728a,a89729a,a89730a,a89734a,a89735a,a89738a,a89741a,a89742a,a89743a,a89747a,a89748a,a89751a,a89754a,a89755a,a89756a,a89760a,a89761a,a89764a,a89767a,a89768a,a89769a,a89773a,a89774a,a89777a,a89780a,a89781a,a89782a,a89786a,a89787a,a89790a,a89793a,a89794a,a89795a,a89799a,a89800a,a89803a,a89806a,a89807a,a89808a,a89812a,a89813a,a89816a,a89819a,a89820a,a89821a,a89825a,a89826a,a89829a,a89832a,a89833a,a89834a,a89838a,a89839a,a89842a,a89845a,a89846a,a89847a,a89851a,a89852a,a89855a,a89858a,a89859a,a89860a,a89864a,a89865a,a89868a,a89871a,a89872a,a89873a,a89877a,a89878a,a89881a,a89884a,a89885a,a89886a,a89890a,a89891a,a89894a,a89897a,a89898a,a89899a,a89903a,a89904a,a89907a,a89910a,a89911a,a89912a,a89916a,a89917a,a89920a,a89923a,a89924a,a89925a,a89929a,a89930a,a89933a,a89936a,a89937a,a89938a,a89942a,a89943a,a89946a,a89949a,a89950a,a89951a,a89955a,a89956a,a89959a,a89962a,a89963a,a89964a,a89968a,a89969a,a89972a,a89975a,a89976a,a89977a,a89981a,a89982a,a89985a,a89988a,a89989a,a89990a,a89994a,a89995a,a89998a,a90001a,a90002a,a90003a,a90007a,a90008a,a90011a,a90014a,a90015a,a90016a,a90020a,a90021a,a90024a,a90027a,a90028a,a90029a,a90033a,a90034a,a90037a,a90040a,a90041a,a90042a,a90046a,a90047a,a90050a,a90053a,a90054a,a90055a,a90059a,a90060a,a90063a,a90066a,a90067a,a90068a,a90072a,a90073a,a90076a,a90079a,a90080a,a90081a,a90085a,a90086a,a90089a,a90092a,a90093a,a90094a,a90098a,a90099a,a90102a,a90105a,a90106a,a90107a,a90111a,a90112a,a90115a,a90118a,a90119a,a90120a,a90124a,a90125a,a90128a,a90131a,a90132a,a90133a,a90137a,a90138a,a90141a,a90144a,a90145a,a90146a,a90150a,a90151a,a90154a,a90157a,a90158a,a90159a,a90163a,a90164a,a90167a,a90170a,a90171a,a90172a,a90176a,a90177a,a90180a,a90183a,a90184a,a90185a,a90189a,a90190a,a90193a,a90196a,a90197a,a90198a,a90202a,a90203a,a90206a,a90209a,a90210a,a90211a,a90215a,a90216a,a90219a,a90222a,a90223a,a90224a,a90228a,a90229a,a90232a,a90235a,a90236a,a90237a,a90241a,a90242a,a90245a,a90248a,a90249a,a90250a,a90254a,a90255a,a90258a,a90261a,a90262a,a90263a,a90267a,a90268a,a90271a,a90274a,a90275a,a90276a,a90280a,a90281a,a90284a,a90287a,a90288a,a90289a,a90293a,a90294a,a90297a,a90300a,a90301a,a90302a,a90306a,a90307a,a90310a,a90313a,a90314a,a90315a,a90319a,a90320a,a90323a,a90326a,a90327a,a90328a,a90332a,a90333a,a90336a,a90339a,a90340a,a90341a,a90345a,a90346a,a90349a,a90352a,a90353a,a90354a,a90358a,a90359a,a90362a,a90365a,a90366a,a90367a,a90371a,a90372a,a90375a,a90378a,a90379a,a90380a,a90384a,a90385a,a90388a,a90391a,a90392a,a90393a,a90397a,a90398a,a90401a,a90404a,a90405a,a90406a,a90410a,a90411a,a90414a,a90417a,a90418a,a90419a,a90423a,a90424a,a90427a,a90430a,a90431a,a90432a,a90436a,a90437a,a90440a,a90443a,a90444a,a90445a,a90449a,a90450a,a90453a,a90456a,a90457a,a90458a,a90462a,a90463a,a90466a,a90469a,a90470a,a90471a,a90475a,a90476a,a90479a,a90482a,a90483a,a90484a,a90488a,a90489a,a90492a,a90495a,a90496a,a90497a,a90501a,a90502a,a90505a,a90508a,a90509a,a90510a,a90514a,a90515a,a90518a,a90521a,a90522a,a90523a,a90527a,a90528a,a90531a,a90534a,a90535a,a90536a,a90540a,a90541a,a90544a,a90547a,a90548a,a90549a,a90553a,a90554a,a90557a,a90560a,a90561a,a90562a,a90566a,a90567a,a90570a,a90573a,a90574a,a90575a,a90579a,a90580a,a90583a,a90586a,a90587a,a90588a,a90592a,a90593a,a90596a,a90599a,a90600a,a90601a,a90605a,a90606a,a90609a,a90612a,a90613a,a90614a,a90618a,a90619a,a90622a,a90625a,a90626a,a90627a,a90631a,a90632a,a90635a,a90638a,a90639a,a90640a,a90644a,a90645a,a90648a,a90651a,a90652a,a90653a,a90657a,a90658a,a90661a,a90664a,a90665a,a90666a,a90670a,a90671a,a90674a,a90677a,a90678a,a90679a,a90683a,a90684a,a90687a,a90690a,a90691a,a90692a,a90696a,a90697a,a90700a,a90703a,a90704a,a90705a,a90709a,a90710a,a90713a,a90716a,a90717a,a90718a,a90722a,a90723a,a90726a,a90729a,a90730a,a90731a,a90735a,a90736a,a90739a,a90742a,a90743a,a90744a,a90748a,a90749a,a90752a,a90755a,a90756a,a90757a,a90761a,a90762a,a90765a,a90768a,a90769a,a90770a,a90774a,a90775a,a90778a,a90781a,a90782a,a90783a,a90787a,a90788a,a90791a,a90794a,a90795a,a90796a,a90800a,a90801a,a90804a,a90807a,a90808a,a90809a,a90813a,a90814a,a90817a,a90820a,a90821a,a90822a,a90826a,a90827a,a90830a,a90833a,a90834a,a90835a,a90839a,a90840a,a90843a,a90846a,a90847a,a90848a,a90852a,a90853a,a90856a,a90859a,a90860a,a90861a,a90865a,a90866a,a90869a,a90872a,a90873a,a90874a,a90878a,a90879a,a90882a,a90885a,a90886a,a90887a,a90891a,a90892a,a90895a,a90898a,a90899a,a90900a,a90904a,a90905a,a90908a,a90911a,a90912a,a90913a,a90917a,a90918a,a90921a,a90924a,a90925a,a90926a,a90930a,a90931a,a90934a,a90937a,a90938a,a90939a,a90943a,a90944a,a90947a,a90950a,a90951a,a90952a,a90956a,a90957a,a90960a,a90963a,a90964a,a90965a,a90969a,a90970a,a90973a,a90976a,a90977a,a90978a,a90982a,a90983a,a90986a,a90989a,a90990a,a90991a,a90995a,a90996a,a90999a,a91002a,a91003a,a91004a,a91008a,a91009a,a91012a,a91015a,a91016a,a91017a,a91021a,a91022a,a91025a,a91028a,a91029a,a91030a,a91034a,a91035a,a91038a,a91041a,a91042a,a91043a,a91047a,a91048a,a91051a,a91054a,a91055a,a91056a,a91060a,a91061a,a91064a,a91067a,a91068a,a91069a,a91073a,a91074a,a91077a,a91080a,a91081a,a91082a,a91086a,a91087a,a91090a,a91093a,a91094a,a91095a,a91099a,a91100a,a91103a,a91106a,a91107a,a91108a,a91112a,a91113a,a91116a,a91119a,a91120a,a91121a,a91125a,a91126a,a91129a,a91132a,a91133a,a91134a,a91138a,a91139a,a91142a,a91145a,a91146a,a91147a,a91151a,a91152a,a91155a,a91158a,a91159a,a91160a,a91164a,a91165a,a91168a,a91171a,a91172a,a91173a,a91177a,a91178a,a91181a,a91184a,a91185a,a91186a,a91190a,a91191a,a91194a,a91197a,a91198a,a91199a,a91203a,a91204a,a91207a,a91210a,a91211a,a91212a,a91216a,a91217a,a91220a,a91223a,a91224a,a91225a,a91229a,a91230a,a91233a,a91236a,a91237a,a91238a,a91242a,a91243a,a91246a,a91249a,a91250a,a91251a,a91255a,a91256a,a91259a,a91262a,a91263a,a91264a,a91268a,a91269a,a91272a,a91275a,a91276a,a91277a,a91281a,a91282a,a91285a,a91288a,a91289a,a91290a,a91294a,a91295a,a91298a,a91301a,a91302a,a91303a,a91307a,a91308a,a91311a,a91314a,a91315a,a91316a,a91320a,a91321a,a91324a,a91327a,a91328a,a91329a,a91333a,a91334a,a91337a,a91340a,a91341a,a91342a,a91346a,a91347a,a91350a,a91353a,a91354a,a91355a,a91359a,a91360a,a91363a,a91366a,a91367a,a91368a,a91372a,a91373a,a91376a,a91379a,a91380a,a91381a,a91385a,a91386a,a91389a,a91392a,a91393a,a91394a,a91398a,a91399a,a91402a,a91405a,a91406a,a91407a,a91411a,a91412a,a91415a,a91418a,a91419a,a91420a,a91424a,a91425a,a91428a,a91431a,a91432a,a91433a,a91437a,a91438a,a91441a,a91444a,a91445a,a91446a,a91450a,a91451a,a91454a,a91457a,a91458a,a91459a,a91463a,a91464a,a91467a,a91470a,a91471a,a91472a,a91476a,a91477a,a91480a,a91483a,a91484a,a91485a,a91489a,a91490a,a91493a,a91496a,a91497a,a91498a,a91502a,a91503a,a91506a,a91509a,a91510a,a91511a,a91515a,a91516a,a91519a,a91522a,a91523a,a91524a,a91528a,a91529a,a91532a,a91535a,a91536a,a91537a,a91541a,a91542a,a91545a,a91548a,a91549a,a91550a,a91554a,a91555a,a91558a,a91561a,a91562a,a91563a,a91567a,a91568a,a91571a,a91574a,a91575a,a91576a,a91580a,a91581a,a91584a,a91587a,a91588a,a91589a,a91593a,a91594a,a91597a,a91600a,a91601a,a91602a,a91606a,a91607a,a91610a,a91613a,a91614a,a91615a,a91619a,a91620a,a91623a,a91626a,a91627a,a91628a,a91632a,a91633a,a91636a,a91639a,a91640a,a91641a,a91645a,a91646a,a91649a,a91652a,a91653a,a91654a,a91658a,a91659a,a91662a,a91665a,a91666a,a91667a,a91671a,a91672a,a91675a,a91678a,a91679a,a91680a,a91684a,a91685a,a91688a,a91691a,a91692a,a91693a,a91697a,a91698a,a91701a,a91704a,a91705a,a91706a,a91710a,a91711a,a91714a,a91717a,a91718a,a91719a,a91723a,a91724a,a91727a,a91730a,a91731a,a91732a,a91736a,a91737a,a91740a,a91743a,a91744a,a91745a,a91749a,a91750a,a91753a,a91756a,a91757a,a91758a,a91762a,a91763a,a91766a,a91769a,a91770a,a91771a,a91775a,a91776a,a91779a,a91782a,a91783a,a91784a,a91788a,a91789a,a91792a,a91795a,a91796a,a91797a,a91801a,a91802a,a91805a,a91808a,a91809a,a91810a,a91814a,a91815a,a91818a,a91821a,a91822a,a91823a,a91827a,a91828a,a91831a,a91834a,a91835a,a91836a,a91840a,a91841a,a91844a,a91847a,a91848a,a91849a,a91853a,a91854a,a91857a,a91860a,a91861a,a91862a,a91866a,a91867a,a91870a,a91873a,a91874a,a91875a,a91879a,a91880a,a91883a,a91886a,a91887a,a91888a,a91892a,a91893a,a91896a,a91899a,a91900a,a91901a,a91905a,a91906a,a91909a,a91912a,a91913a,a91914a,a91918a,a91919a,a91922a,a91925a,a91926a,a91927a,a91931a,a91932a,a91935a,a91938a,a91939a,a91940a,a91944a,a91945a,a91948a,a91951a,a91952a,a91953a,a91957a,a91958a,a91961a,a91964a,a91965a,a91966a,a91970a,a91971a,a91974a,a91977a,a91978a,a91979a,a91983a,a91984a,a91987a,a91990a,a91991a,a91992a,a91996a,a91997a,a92000a,a92003a,a92004a,a92005a,a92009a,a92010a,a92013a,a92016a,a92017a,a92018a,a92022a,a92023a,a92026a,a92029a,a92030a,a92031a,a92035a,a92036a,a92039a,a92042a,a92043a,a92044a,a92048a,a92049a,a92052a,a92055a,a92056a,a92057a,a92061a,a92062a,a92065a,a92068a,a92069a,a92070a,a92074a,a92075a,a92078a,a92081a,a92082a,a92083a,a92087a,a92088a,a92091a,a92094a,a92095a,a92096a,a92100a,a92101a,a92104a,a92107a,a92108a,a92109a,a92113a,a92114a,a92117a,a92120a,a92121a,a92122a,a92126a,a92127a,a92130a,a92133a,a92134a,a92135a,a92139a,a92140a,a92143a,a92146a,a92147a,a92148a,a92152a,a92153a,a92156a,a92159a,a92160a,a92161a,a92165a,a92166a,a92169a,a92172a,a92173a,a92174a,a92178a,a92179a,a92182a,a92185a,a92186a,a92187a,a92191a,a92192a,a92195a,a92198a,a92199a,a92200a,a92204a,a92205a,a92208a,a92211a,a92212a,a92213a,a92217a,a92218a,a92221a,a92224a,a92225a,a92226a,a92230a,a92231a,a92234a,a92237a,a92238a,a92239a,a92243a,a92244a,a92247a,a92250a,a92251a,a92252a,a92256a,a92257a,a92260a,a92263a,a92264a,a92265a,a92269a,a92270a,a92273a,a92276a,a92277a,a92278a,a92282a,a92283a,a92286a,a92289a,a92290a,a92291a,a92295a,a92296a,a92299a,a92302a,a92303a,a92304a,a92308a,a92309a,a92312a,a92315a,a92316a,a92317a,a92321a,a92322a,a92325a,a92328a,a92329a,a92330a,a92334a,a92335a,a92338a,a92341a,a92342a,a92343a,a92347a,a92348a,a92351a,a92354a,a92355a,a92356a,a92360a,a92361a,a92364a,a92367a,a92368a,a92369a,a92373a,a92374a,a92377a,a92380a,a92381a,a92382a,a92386a,a92387a,a92390a,a92393a,a92394a,a92395a,a92399a,a92400a,a92403a,a92406a,a92407a,a92408a,a92412a,a92413a,a92416a,a92419a,a92420a,a92421a,a92425a,a92426a,a92429a,a92432a,a92433a,a92434a,a92438a,a92439a,a92442a,a92445a,a92446a,a92447a,a92451a,a92452a,a92455a,a92458a,a92459a,a92460a,a92464a,a92465a,a92468a,a92471a,a92472a,a92473a,a92477a,a92478a,a92481a,a92484a,a92485a,a92486a,a92490a,a92491a,a92494a,a92497a,a92498a,a92499a,a92503a,a92504a,a92507a,a92510a,a92511a,a92512a,a92516a,a92517a,a92520a,a92523a,a92524a,a92525a,a92529a,a92530a,a92533a,a92536a,a92537a,a92538a,a92542a,a92543a,a92546a,a92549a,a92550a,a92551a,a92555a,a92556a,a92559a,a92562a,a92563a,a92564a,a92568a,a92569a,a92572a,a92575a,a92576a,a92577a,a92581a,a92582a,a92585a,a92588a,a92589a,a92590a,a92594a,a92595a,a92598a,a92601a,a92602a,a92603a,a92607a,a92608a,a92611a,a92614a,a92615a,a92616a,a92620a,a92621a,a92624a,a92627a,a92628a,a92629a,a92633a,a92634a,a92637a,a92640a,a92641a,a92642a,a92646a,a92647a,a92650a,a92653a,a92654a,a92655a,a92659a,a92660a,a92663a,a92666a,a92667a,a92668a,a92672a,a92673a,a92676a,a92679a,a92680a,a92681a,a92685a,a92686a,a92689a,a92692a,a92693a,a92694a,a92698a,a92699a,a92702a,a92705a,a92706a,a92707a,a92711a,a92712a,a92715a,a92718a,a92719a,a92720a,a92724a,a92725a,a92728a,a92731a,a92732a,a92733a,a92737a,a92738a,a92741a,a92744a,a92745a,a92746a,a92750a,a92751a,a92754a,a92757a,a92758a,a92759a,a92763a,a92764a,a92767a,a92770a,a92771a,a92772a,a92776a,a92777a,a92780a,a92783a,a92784a,a92785a,a92789a,a92790a,a92793a,a92796a,a92797a,a92798a,a92802a,a92803a,a92806a,a92809a,a92810a,a92811a,a92815a,a92816a,a92819a,a92822a,a92823a,a92824a,a92828a,a92829a,a92832a,a92835a,a92836a,a92837a,a92841a,a92842a,a92845a,a92848a,a92849a,a92850a,a92854a,a92855a,a92858a,a92861a,a92862a,a92863a,a92867a,a92868a,a92871a,a92874a,a92875a,a92876a,a92880a,a92881a,a92884a,a92887a,a92888a,a92889a,a92893a,a92894a,a92897a,a92900a,a92901a,a92902a,a92906a,a92907a,a92910a,a92913a,a92914a,a92915a,a92919a,a92920a,a92923a,a92926a,a92927a,a92928a,a92932a,a92933a,a92936a,a92939a,a92940a,a92941a,a92945a,a92946a,a92949a,a92952a,a92953a,a92954a,a92958a,a92959a,a92962a,a92965a,a92966a,a92967a,a92971a,a92972a,a92975a,a92978a,a92979a,a92980a,a92984a,a92985a,a92988a,a92991a,a92992a,a92993a,a92997a,a92998a,a93001a,a93004a,a93005a,a93006a,a93010a,a93011a,a93014a,a93017a,a93018a,a93019a,a93023a,a93024a,a93027a,a93030a,a93031a,a93032a,a93036a,a93037a,a93040a,a93043a,a93044a,a93045a,a93049a,a93050a,a93053a,a93056a,a93057a,a93058a,a93062a,a93063a,a93066a,a93069a,a93070a,a93071a,a93075a,a93076a,a93079a,a93082a,a93083a,a93084a,a93088a,a93089a,a93092a,a93095a,a93096a,a93097a,a93101a,a93102a,a93105a,a93108a,a93109a,a93110a,a93114a,a93115a,a93118a,a93121a,a93122a,a93123a,a93127a,a93128a,a93131a,a93134a,a93135a,a93136a,a93140a,a93141a,a93144a,a93147a,a93148a,a93149a,a93153a,a93154a,a93157a,a93160a,a93161a,a93162a,a93166a,a93167a,a93170a,a93173a,a93174a,a93175a,a93179a,a93180a,a93183a,a93186a,a93187a,a93188a,a93192a,a93193a,a93196a,a93199a,a93200a,a93201a,a93205a,a93206a,a93209a,a93212a,a93213a,a93214a,a93218a,a93219a,a93222a,a93225a,a93226a,a93227a,a93231a,a93232a,a93235a,a93238a,a93239a,a93240a,a93244a,a93245a,a93248a,a93251a,a93252a,a93253a,a93257a,a93258a,a93261a,a93264a,a93265a,a93266a,a93270a,a93271a,a93274a,a93277a,a93278a,a93279a,a93283a,a93284a,a93287a,a93290a,a93291a,a93292a,a93296a,a93297a,a93300a,a93303a,a93304a,a93305a,a93309a,a93310a,a93313a,a93316a,a93317a,a93318a,a93322a,a93323a,a93326a,a93329a,a93330a,a93331a,a93335a,a93336a,a93339a,a93342a,a93343a,a93344a,a93348a,a93349a,a93352a,a93355a,a93356a,a93357a,a93361a,a93362a,a93365a,a93368a,a93369a,a93370a,a93374a,a93375a,a93378a,a93381a,a93382a,a93383a,a93387a,a93388a,a93391a,a93394a,a93395a,a93396a,a93400a,a93401a,a93404a,a93407a,a93408a,a93409a,a93413a,a93414a,a93417a,a93420a,a93421a,a93422a,a93426a,a93427a,a93430a,a93433a,a93434a,a93435a,a93439a,a93440a,a93443a,a93446a,a93447a,a93448a,a93452a,a93453a,a93456a,a93459a,a93460a,a93461a,a93465a,a93466a,a93469a,a93472a,a93473a,a93474a,a93478a,a93479a,a93482a,a93485a,a93486a,a93487a,a93491a,a93492a,a93495a,a93498a,a93499a,a93500a,a93504a,a93505a,a93508a,a93511a,a93512a,a93513a,a93517a,a93518a,a93521a,a93524a,a93525a,a93526a,a93530a,a93531a,a93534a,a93537a,a93538a,a93539a,a93543a,a93544a,a93547a,a93550a,a93551a,a93552a,a93556a,a93557a,a93560a,a93563a,a93564a,a93565a,a93569a,a93570a,a93573a,a93576a,a93577a,a93578a,a93582a,a93583a,a93586a,a93589a,a93590a,a93591a,a93595a,a93596a,a93599a,a93602a,a93603a,a93604a,a93608a,a93609a,a93612a,a93615a,a93616a,a93617a,a93621a,a93622a,a93625a,a93628a,a93629a,a93630a,a93634a,a93635a,a93638a,a93641a,a93642a,a93643a,a93647a,a93648a,a93651a,a93654a,a93655a,a93656a,a93660a,a93661a,a93664a,a93667a,a93668a,a93669a,a93673a,a93674a,a93677a,a93680a,a93681a,a93682a,a93686a,a93687a,a93690a,a93693a,a93694a,a93695a,a93699a,a93700a,a93703a,a93706a,a93707a,a93708a,a93712a,a93713a,a93716a,a93719a,a93720a,a93721a,a93725a,a93726a,a93729a,a93732a,a93733a,a93734a,a93738a,a93739a,a93742a,a93745a,a93746a,a93747a,a93751a,a93752a,a93755a,a93758a,a93759a,a93760a,a93764a,a93765a,a93768a,a93771a,a93772a,a93773a,a93777a,a93778a,a93781a,a93784a,a93785a,a93786a,a93790a,a93791a,a93794a,a93797a,a93798a,a93799a,a93803a,a93804a,a93807a,a93810a,a93811a,a93812a,a93816a,a93817a,a93820a,a93823a,a93824a,a93825a,a93829a,a93830a,a93833a,a93836a,a93837a,a93838a,a93842a,a93843a,a93846a,a93849a,a93850a,a93851a,a93855a,a93856a,a93859a,a93862a,a93863a,a93864a,a93868a,a93869a,a93872a,a93875a,a93876a,a93877a,a93881a,a93882a,a93885a,a93888a,a93889a,a93890a,a93894a,a93895a,a93898a,a93901a,a93902a,a93903a,a93907a,a93908a,a93911a,a93914a,a93915a,a93916a,a93920a,a93921a,a93924a,a93927a,a93928a,a93929a,a93933a,a93934a,a93937a,a93940a,a93941a,a93942a,a93946a,a93947a,a93950a,a93953a,a93954a,a93955a,a93959a,a93960a,a93963a,a93966a,a93967a,a93968a,a93972a,a93973a,a93976a,a93979a,a93980a,a93981a,a93985a,a93986a,a93989a,a93992a,a93993a,a93994a,a93998a,a93999a,a94002a,a94005a,a94006a,a94007a,a94011a,a94012a,a94015a,a94018a,a94019a,a94020a,a94024a,a94025a,a94028a,a94031a,a94032a,a94033a,a94037a,a94038a,a94041a,a94044a,a94045a,a94046a,a94050a,a94051a,a94054a,a94057a,a94058a,a94059a,a94063a,a94064a,a94067a,a94070a,a94071a,a94072a,a94076a,a94077a,a94080a,a94083a,a94084a,a94085a,a94089a,a94090a,a94093a,a94096a,a94097a,a94098a,a94102a,a94103a,a94106a,a94109a,a94110a,a94111a,a94115a,a94116a,a94119a,a94122a,a94123a,a94124a,a94128a,a94129a,a94132a,a94135a,a94136a,a94137a,a94141a,a94142a,a94145a,a94148a,a94149a,a94150a,a94154a,a94155a,a94158a,a94161a,a94162a,a94163a,a94167a,a94168a,a94171a,a94174a,a94175a,a94176a,a94180a,a94181a,a94184a,a94187a,a94188a,a94189a,a94193a,a94194a,a94197a,a94200a,a94201a,a94202a,a94206a,a94207a,a94210a,a94213a,a94214a,a94215a,a94219a,a94220a,a94223a,a94226a,a94227a,a94228a,a94232a,a94233a,a94236a,a94239a,a94240a,a94241a,a94245a,a94246a,a94249a,a94252a,a94253a,a94254a,a94258a,a94259a,a94262a,a94265a,a94266a,a94267a,a94271a,a94272a,a94275a,a94278a,a94279a,a94280a,a94284a,a94285a,a94288a,a94291a,a94292a,a94293a,a94297a,a94298a,a94301a,a94304a,a94305a,a94306a,a94310a,a94311a,a94314a,a94317a,a94318a,a94319a,a94323a,a94324a,a94327a,a94330a,a94331a,a94332a,a94336a,a94337a,a94340a,a94343a,a94344a,a94345a,a94349a,a94350a,a94353a,a94356a,a94357a,a94358a,a94362a,a94363a,a94366a,a94369a,a94370a,a94371a,a94375a,a94376a,a94379a,a94382a,a94383a,a94384a,a94388a,a94389a,a94392a,a94395a,a94396a,a94397a,a94401a,a94402a,a94405a,a94408a,a94409a,a94410a,a94414a,a94415a,a94418a,a94421a,a94422a,a94423a,a94427a,a94428a,a94431a,a94434a,a94435a,a94436a,a94440a,a94441a,a94444a,a94447a,a94448a,a94449a,a94453a,a94454a,a94457a,a94460a,a94461a,a94462a,a94466a,a94467a,a94470a,a94473a,a94474a,a94475a,a94479a,a94480a,a94483a,a94486a,a94487a,a94488a,a94492a,a94493a,a94496a,a94499a,a94500a,a94501a,a94505a,a94506a,a94509a,a94512a,a94513a,a94514a,a94518a,a94519a,a94522a,a94525a,a94526a,a94527a,a94531a,a94532a,a94535a,a94538a,a94539a,a94540a,a94544a,a94545a,a94548a,a94551a,a94552a,a94553a,a94557a,a94558a,a94561a,a94564a,a94565a,a94566a,a94570a,a94571a,a94574a,a94577a,a94578a,a94579a,a94583a,a94584a,a94587a,a94590a,a94591a,a94592a,a94596a,a94597a,a94600a,a94603a,a94604a,a94605a,a94609a,a94610a,a94613a,a94616a,a94617a,a94618a,a94622a,a94623a,a94626a,a94629a,a94630a,a94631a,a94635a,a94636a,a94639a,a94642a,a94643a,a94644a,a94648a,a94649a,a94652a,a94655a,a94656a,a94657a,a94661a,a94662a,a94665a,a94668a,a94669a,a94670a,a94674a,a94675a,a94678a,a94681a,a94682a,a94683a,a94687a,a94688a,a94691a,a94694a,a94695a,a94696a,a94700a,a94701a,a94704a,a94707a,a94708a,a94709a,a94713a,a94714a,a94717a,a94720a,a94721a,a94722a,a94726a,a94727a,a94730a,a94733a,a94734a,a94735a,a94739a,a94740a,a94743a,a94746a,a94747a,a94748a,a94752a,a94753a,a94756a,a94759a,a94760a,a94761a,a94765a,a94766a,a94769a,a94772a,a94773a,a94774a,a94778a,a94779a,a94782a,a94785a,a94786a,a94787a,a94791a,a94792a,a94795a,a94798a,a94799a,a94800a,a94804a,a94805a,a94808a,a94811a,a94812a,a94813a,a94817a,a94818a,a94821a,a94824a,a94825a,a94826a,a94830a,a94831a,a94834a,a94837a,a94838a,a94839a,a94843a,a94844a,a94847a,a94850a,a94851a,a94852a,a94856a,a94857a,a94860a,a94863a,a94864a,a94865a,a94869a,a94870a,a94873a,a94876a,a94877a,a94878a,a94882a,a94883a,a94886a,a94889a,a94890a,a94891a,a94895a,a94896a,a94899a,a94902a,a94903a,a94904a,a94908a,a94909a,a94912a,a94915a,a94916a,a94917a,a94921a,a94922a,a94925a,a94928a,a94929a,a94930a,a94934a,a94935a,a94938a,a94941a,a94942a,a94943a,a94947a,a94948a,a94951a,a94954a,a94955a,a94956a,a94960a,a94961a,a94964a,a94967a,a94968a,a94969a,a94973a,a94974a,a94977a,a94980a,a94981a,a94982a,a94986a,a94987a,a94990a,a94993a,a94994a,a94995a,a94999a,a95000a,a95003a,a95006a,a95007a,a95008a,a95012a,a95013a,a95016a,a95019a,a95020a,a95021a,a95025a,a95026a,a95029a,a95032a,a95033a,a95034a,a95038a,a95039a,a95042a,a95045a,a95046a,a95047a,a95051a,a95052a,a95055a,a95058a,a95059a,a95060a,a95064a,a95065a,a95068a,a95071a,a95072a,a95073a,a95077a,a95078a,a95081a,a95084a,a95085a,a95086a,a95090a,a95091a,a95094a,a95097a,a95098a,a95099a,a95103a,a95104a,a95107a,a95110a,a95111a,a95112a,a95116a,a95117a,a95120a,a95123a,a95124a,a95125a,a95129a,a95130a,a95133a,a95136a,a95137a,a95138a,a95142a,a95143a,a95146a,a95149a,a95150a,a95151a,a95155a,a95156a,a95159a,a95162a,a95163a,a95164a,a95168a,a95169a,a95172a,a95175a,a95176a,a95177a,a95181a,a95182a,a95185a,a95188a,a95189a,a95190a,a95194a,a95195a,a95198a,a95201a,a95202a,a95203a,a95207a,a95208a,a95211a,a95214a,a95215a,a95216a,a95220a,a95221a,a95224a,a95227a,a95228a,a95229a,a95233a,a95234a,a95237a,a95240a,a95241a,a95242a,a95246a,a95247a,a95250a,a95253a,a95254a,a95255a,a95259a,a95260a,a95263a,a95266a,a95267a,a95268a,a95272a,a95273a,a95276a,a95279a,a95280a,a95281a,a95285a,a95286a,a95289a,a95292a,a95293a,a95294a,a95298a,a95299a,a95302a,a95305a,a95306a,a95307a,a95311a,a95312a,a95315a,a95318a,a95319a,a95320a,a95324a,a95325a,a95328a,a95331a,a95332a,a95333a,a95337a,a95338a,a95341a,a95344a,a95345a,a95346a,a95350a,a95351a,a95354a,a95357a,a95358a,a95359a,a95363a,a95364a,a95367a,a95370a,a95371a,a95372a,a95376a,a95377a,a95380a,a95383a,a95384a,a95385a,a95389a,a95390a,a95393a,a95396a,a95397a,a95398a,a95402a,a95403a,a95406a,a95409a,a95410a,a95411a,a95415a,a95416a,a95419a,a95422a,a95423a,a95424a,a95428a,a95429a,a95432a,a95435a,a95436a,a95437a,a95441a,a95442a,a95445a,a95448a,a95449a,a95450a,a95454a,a95455a,a95458a,a95461a,a95462a,a95463a,a95467a,a95468a,a95471a,a95474a,a95475a,a95476a,a95480a,a95481a,a95484a,a95487a,a95488a,a95489a,a95493a,a95494a,a95497a,a95500a,a95501a,a95502a,a95506a,a95507a,a95510a,a95513a,a95514a,a95515a,a95519a,a95520a,a95523a,a95526a,a95527a,a95528a,a95532a,a95533a,a95536a,a95539a,a95540a,a95541a,a95545a,a95546a,a95549a,a95552a,a95553a,a95554a,a95558a,a95559a,a95562a,a95565a,a95566a,a95567a,a95571a,a95572a,a95575a,a95578a,a95579a,a95580a,a95584a,a95585a,a95588a,a95591a,a95592a,a95593a,a95597a,a95598a,a95601a,a95604a,a95605a,a95606a,a95610a,a95611a,a95614a,a95617a,a95618a,a95619a,a95623a,a95624a,a95627a,a95630a,a95631a,a95632a,a95636a,a95637a,a95640a,a95643a,a95644a,a95645a,a95649a,a95650a,a95653a,a95656a,a95657a,a95658a,a95662a,a95663a,a95666a,a95669a,a95670a,a95671a,a95675a,a95676a,a95679a,a95682a,a95683a,a95684a,a95688a,a95689a,a95692a,a95695a,a95696a,a95697a,a95701a,a95702a,a95705a,a95708a,a95709a,a95710a,a95714a,a95715a,a95718a,a95721a,a95722a,a95723a,a95727a,a95728a,a95731a,a95734a,a95735a,a95736a,a95740a,a95741a,a95744a,a95747a,a95748a,a95749a,a95753a,a95754a,a95757a,a95760a,a95761a,a95762a,a95766a,a95767a,a95770a,a95773a,a95774a,a95775a,a95779a,a95780a,a95783a,a95786a,a95787a,a95788a,a95792a,a95793a,a95796a,a95799a,a95800a,a95801a,a95805a,a95806a,a95809a,a95812a,a95813a,a95814a,a95818a,a95819a,a95822a,a95825a,a95826a,a95827a,a95831a,a95832a,a95835a,a95838a,a95839a,a95840a,a95844a,a95845a,a95848a,a95851a,a95852a,a95853a,a95857a,a95858a,a95861a,a95864a,a95865a,a95866a,a95870a,a95871a,a95874a,a95877a,a95878a,a95879a,a95883a,a95884a,a95887a,a95890a,a95891a,a95892a,a95896a,a95897a,a95900a,a95903a,a95904a,a95905a,a95909a,a95910a,a95913a,a95916a,a95917a,a95918a,a95922a,a95923a,a95926a,a95929a,a95930a,a95931a,a95935a,a95936a,a95939a,a95942a,a95943a,a95944a,a95948a,a95949a,a95952a,a95955a,a95956a,a95957a,a95961a,a95962a,a95965a,a95968a,a95969a,a95970a,a95974a,a95975a,a95978a,a95981a,a95982a,a95983a,a95987a,a95988a,a95991a,a95994a,a95995a,a95996a,a96000a,a96001a,a96004a,a96007a,a96008a,a96009a,a96013a,a96014a,a96017a,a96020a,a96021a,a96022a,a96026a,a96027a,a96030a,a96033a,a96034a,a96035a,a96039a,a96040a,a96043a,a96046a,a96047a,a96048a,a96052a,a96053a,a96056a,a96059a,a96060a,a96061a,a96065a,a96066a,a96069a,a96072a,a96073a,a96074a,a96078a,a96079a,a96082a,a96085a,a96086a,a96087a,a96091a,a96092a,a96095a,a96098a,a96099a,a96100a,a96104a,a96105a,a96108a,a96111a,a96112a,a96113a,a96117a,a96118a,a96121a,a96124a,a96125a,a96126a,a96130a,a96131a,a96134a,a96137a,a96138a,a96139a,a96143a,a96144a,a96147a,a96150a,a96151a,a96152a,a96156a,a96157a,a96160a,a96163a,a96164a,a96165a,a96169a,a96170a,a96173a,a96176a,a96177a,a96178a,a96182a,a96183a,a96186a,a96189a,a96190a,a96191a,a96195a,a96196a,a96199a,a96202a,a96203a,a96204a,a96208a,a96209a,a96212a,a96215a,a96216a,a96217a,a96221a,a96222a,a96225a,a96228a,a96229a,a96230a,a96234a,a96235a,a96238a,a96241a,a96242a,a96243a,a96247a,a96248a,a96251a,a96254a,a96255a,a96256a,a96260a,a96261a,a96264a,a96267a,a96268a,a96269a,a96273a,a96274a,a96277a,a96280a,a96281a,a96282a,a96286a,a96287a,a96290a,a96293a,a96294a,a96295a,a96299a,a96300a,a96303a,a96306a,a96307a,a96308a,a96312a,a96313a,a96316a,a96319a,a96320a,a96321a,a96325a,a96326a,a96329a,a96332a,a96333a,a96334a,a96338a,a96339a,a96342a,a96345a,a96346a,a96347a,a96351a,a96352a,a96355a,a96358a,a96359a,a96360a,a96364a,a96365a,a96368a,a96371a,a96372a,a96373a,a96377a,a96378a,a96381a,a96384a,a96385a,a96386a,a96390a,a96391a,a96394a,a96397a,a96398a,a96399a,a96403a,a96404a,a96407a,a96410a,a96411a,a96412a,a96416a,a96417a,a96420a,a96423a,a96424a,a96425a,a96429a,a96430a,a96433a,a96436a,a96437a,a96438a,a96442a,a96443a,a96446a,a96449a,a96450a,a96451a,a96455a,a96456a,a96459a,a96462a,a96463a,a96464a,a96468a,a96469a,a96472a,a96475a,a96476a,a96477a,a96481a,a96482a,a96485a,a96488a,a96489a,a96490a,a96494a,a96495a,a96498a,a96501a,a96502a,a96503a,a96507a,a96508a,a96511a,a96514a,a96515a,a96516a,a96520a,a96521a,a96524a,a96527a,a96528a,a96529a,a96533a,a96534a,a96537a,a96540a,a96541a,a96542a,a96546a,a96547a,a96550a,a96553a,a96554a,a96555a,a96559a,a96560a,a96563a,a96566a,a96567a,a96568a,a96572a,a96573a,a96576a,a96579a,a96580a,a96581a,a96585a,a96586a,a96589a,a96592a,a96593a,a96594a,a96598a,a96599a,a96602a,a96605a,a96606a,a96607a,a96611a,a96612a,a96615a,a96618a,a96619a,a96620a,a96624a,a96625a,a96628a,a96631a,a96632a,a96633a,a96637a,a96638a,a96641a,a96644a,a96645a,a96646a,a96650a,a96651a,a96654a,a96657a,a96658a,a96659a,a96663a,a96664a,a96667a,a96670a,a96671a,a96672a,a96676a,a96677a,a96680a,a96683a,a96684a,a96685a,a96689a,a96690a,a96693a,a96696a,a96697a,a96698a,a96702a,a96703a,a96706a,a96709a,a96710a,a96711a,a96715a,a96716a,a96719a,a96722a,a96723a,a96724a,a96728a,a96729a,a96732a,a96735a,a96736a,a96737a,a96741a,a96742a,a96745a,a96748a,a96749a,a96750a,a96754a,a96755a,a96758a,a96761a,a96762a,a96763a,a96767a,a96768a,a96771a,a96774a,a96775a,a96776a,a96780a,a96781a,a96784a,a96787a,a96788a,a96789a,a96793a,a96794a,a96797a,a96800a,a96801a,a96802a,a96806a,a96807a,a96810a,a96813a,a96814a,a96815a,a96819a,a96820a,a96823a,a96826a,a96827a,a96828a,a96832a,a96833a,a96836a,a96839a,a96840a,a96841a,a96845a,a96846a,a96849a,a96852a,a96853a,a96854a,a96858a,a96859a,a96862a,a96865a,a96866a,a96867a,a96871a,a96872a,a96875a,a96878a,a96879a,a96880a,a96884a,a96885a,a96888a,a96891a,a96892a,a96893a,a96897a,a96898a,a96901a,a96904a,a96905a,a96906a,a96910a,a96911a,a96914a,a96917a,a96918a,a96919a,a96923a,a96924a,a96927a,a96930a,a96931a,a96932a,a96936a,a96937a,a96940a,a96943a,a96944a,a96945a,a96949a,a96950a,a96953a,a96956a,a96957a,a96958a,a96962a,a96963a,a96966a,a96969a,a96970a,a96971a,a96975a,a96976a,a96979a,a96982a,a96983a,a96984a,a96988a,a96989a,a96992a,a96995a,a96996a,a96997a,a97001a,a97002a,a97005a,a97008a,a97009a,a97010a,a97014a,a97015a,a97018a,a97021a,a97022a,a97023a,a97027a,a97028a,a97031a,a97034a,a97035a,a97036a,a97040a,a97041a,a97044a,a97047a,a97048a,a97049a,a97053a,a97054a,a97057a,a97060a,a97061a,a97062a,a97066a,a97067a,a97070a,a97073a,a97074a,a97075a,a97079a,a97080a,a97083a,a97086a,a97087a,a97088a,a97092a,a97093a,a97096a,a97099a,a97100a,a97101a,a97105a,a97106a,a97109a,a97112a,a97113a,a97114a,a97118a,a97119a,a97122a,a97125a,a97126a,a97127a,a97131a,a97132a,a97135a,a97138a,a97139a,a97140a,a97144a,a97145a,a97148a,a97151a,a97152a,a97153a,a97157a,a97158a,a97161a,a97164a,a97165a,a97166a,a97170a,a97171a,a97174a,a97177a,a97178a,a97179a,a97183a,a97184a,a97187a,a97190a,a97191a,a97192a,a97196a,a97197a,a97200a,a97203a,a97204a,a97205a,a97209a,a97210a,a97213a,a97216a,a97217a,a97218a,a97222a,a97223a,a97226a,a97229a,a97230a,a97231a,a97235a,a97236a,a97239a,a97242a,a97243a,a97244a,a97248a,a97249a,a97252a,a97255a,a97256a,a97257a,a97261a,a97262a,a97265a,a97268a,a97269a,a97270a,a97274a,a97275a,a97278a,a97281a,a97282a,a97283a,a97287a,a97288a,a97291a,a97294a,a97295a,a97296a,a97300a,a97301a,a97304a,a97307a,a97308a,a97309a,a97313a,a97314a,a97317a,a97320a,a97321a,a97322a,a97326a,a97327a,a97330a,a97333a,a97334a,a97335a,a97339a,a97340a,a97343a,a97346a,a97347a,a97348a,a97352a,a97353a,a97356a,a97359a,a97360a,a97361a,a97365a,a97366a,a97369a,a97372a,a97373a,a97374a,a97378a,a97379a,a97382a,a97385a,a97386a,a97387a,a97391a,a97392a,a97395a,a97398a,a97399a,a97400a,a97404a,a97405a,a97408a,a97411a,a97412a,a97413a,a97417a,a97418a,a97421a,a97424a,a97425a,a97426a,a97430a,a97431a,a97434a,a97437a,a97438a,a97439a,a97443a,a97444a,a97447a,a97450a,a97451a,a97452a,a97456a,a97457a,a97460a,a97463a,a97464a,a97465a,a97469a,a97470a,a97473a,a97476a,a97477a,a97478a,a97482a,a97483a,a97486a,a97489a,a97490a,a97491a,a97495a,a97496a,a97499a,a97502a,a97503a,a97504a,a97508a,a97509a,a97512a,a97515a,a97516a,a97517a,a97521a,a97522a,a97525a,a97528a,a97529a,a97530a,a97534a,a97535a,a97538a,a97541a,a97542a,a97543a,a97547a,a97548a,a97551a,a97554a,a97555a,a97556a,a97560a,a97561a,a97564a,a97567a,a97568a,a97569a,a97573a,a97574a,a97577a,a97580a,a97581a,a97582a,a97586a,a97587a,a97590a,a97593a,a97594a,a97595a,a97599a,a97600a,a97603a,a97606a,a97607a,a97608a,a97612a,a97613a,a97616a,a97619a,a97620a,a97621a,a97625a,a97626a,a97629a,a97632a,a97633a,a97634a,a97638a,a97639a,a97642a,a97645a,a97646a,a97647a,a97651a,a97652a,a97655a,a97658a,a97659a,a97660a,a97664a,a97665a,a97668a,a97671a,a97672a,a97673a,a97677a,a97678a,a97681a,a97684a,a97685a,a97686a,a97690a,a97691a,a97694a,a97697a,a97698a,a97699a,a97703a,a97704a,a97707a,a97710a,a97711a,a97712a,a97716a,a97717a,a97720a,a97723a,a97724a,a97725a,a97729a,a97730a,a97733a,a97736a,a97737a,a97738a,a97742a,a97743a,a97746a,a97749a,a97750a,a97751a,a97755a,a97756a,a97759a,a97762a,a97763a,a97764a,a97768a,a97769a,a97772a,a97775a,a97776a,a97777a,a97781a,a97782a,a97785a,a97788a,a97789a,a97790a,a97794a,a97795a,a97798a,a97801a,a97802a,a97803a,a97807a,a97808a,a97811a,a97814a,a97815a,a97816a,a97820a,a97821a,a97824a,a97827a,a97828a,a97829a,a97833a,a97834a,a97837a,a97840a,a97841a,a97842a,a97846a,a97847a,a97850a,a97853a,a97854a,a97855a,a97859a,a97860a,a97863a,a97866a,a97867a,a97868a,a97872a,a97873a,a97876a,a97879a,a97880a,a97881a,a97885a,a97886a,a97889a,a97892a,a97893a,a97894a,a97898a,a97899a,a97902a,a97905a,a97906a,a97907a,a97911a,a97912a,a97915a,a97918a,a97919a,a97920a,a97924a,a97925a,a97928a,a97931a,a97932a,a97933a,a97937a,a97938a,a97941a,a97944a,a97945a,a97946a,a97950a,a97951a,a97954a,a97957a,a97958a,a97959a,a97963a,a97964a,a97967a,a97970a,a97971a,a97972a,a97976a,a97977a,a97980a,a97983a,a97984a,a97985a,a97989a,a97990a,a97993a,a97996a,a97997a,a97998a,a98002a,a98003a,a98006a,a98009a,a98010a,a98011a,a98015a,a98016a,a98019a,a98022a,a98023a,a98024a,a98028a,a98029a,a98032a,a98035a,a98036a,a98037a,a98041a,a98042a,a98045a,a98048a,a98049a,a98050a,a98054a,a98055a,a98058a,a98061a,a98062a,a98063a,a98067a,a98068a,a98071a,a98074a,a98075a,a98076a,a98080a,a98081a,a98084a,a98087a,a98088a,a98089a,a98093a,a98094a,a98097a,a98100a,a98101a,a98102a,a98106a,a98107a,a98110a,a98113a,a98114a,a98115a,a98119a,a98120a,a98123a,a98126a,a98127a,a98128a,a98132a,a98133a,a98136a,a98139a,a98140a,a98141a,a98145a,a98146a,a98149a,a98152a,a98153a,a98154a,a98158a,a98159a,a98162a,a98165a,a98166a,a98167a,a98171a,a98172a,a98175a,a98178a,a98179a,a98180a,a98184a,a98185a,a98188a,a98191a,a98192a,a98193a,a98197a,a98198a,a98201a,a98204a,a98205a,a98206a,a98210a,a98211a,a98214a,a98217a,a98218a,a98219a,a98223a,a98224a,a98227a,a98230a,a98231a,a98232a,a98236a,a98237a,a98240a,a98243a,a98244a,a98245a,a98249a,a98250a,a98253a,a98256a,a98257a,a98258a,a98262a,a98263a,a98266a,a98269a,a98270a,a98271a,a98275a,a98276a,a98279a,a98282a,a98283a,a98284a,a98288a,a98289a,a98292a,a98295a,a98296a,a98297a,a98301a,a98302a,a98305a,a98308a,a98309a,a98310a,a98314a,a98315a,a98318a,a98321a,a98322a,a98323a,a98327a,a98328a,a98331a,a98334a,a98335a,a98336a,a98340a,a98341a,a98344a,a98347a,a98348a,a98349a,a98353a,a98354a,a98357a,a98360a,a98361a,a98362a,a98366a,a98367a,a98370a,a98373a,a98374a,a98375a,a98379a,a98380a,a98383a,a98386a,a98387a,a98388a,a98392a,a98393a,a98396a,a98399a,a98400a,a98401a,a98405a,a98406a,a98409a,a98412a,a98413a,a98414a,a98418a,a98419a,a98422a,a98425a,a98426a,a98427a,a98431a,a98432a,a98435a,a98438a,a98439a,a98440a,a98444a,a98445a,a98448a,a98451a,a98452a,a98453a,a98457a,a98458a,a98461a,a98464a,a98465a,a98466a,a98470a,a98471a,a98474a,a98477a,a98478a,a98479a,a98483a,a98484a,a98487a,a98490a,a98491a,a98492a,a98496a,a98497a,a98500a,a98503a,a98504a,a98505a,a98509a,a98510a,a98513a,a98516a,a98517a,a98518a,a98522a,a98523a,a98526a,a98529a,a98530a,a98531a,a98535a,a98536a,a98539a,a98542a,a98543a,a98544a,a98548a,a98549a,a98552a,a98555a,a98556a,a98557a,a98561a,a98562a,a98565a,a98568a,a98569a,a98570a,a98574a,a98575a,a98578a,a98581a,a98582a,a98583a,a98587a,a98588a,a98591a,a98594a,a98595a,a98596a,a98600a,a98601a,a98604a,a98607a,a98608a,a98609a,a98613a,a98614a,a98617a,a98620a,a98621a,a98622a,a98626a,a98627a,a98630a,a98633a,a98634a,a98635a,a98639a,a98640a,a98643a,a98646a,a98647a,a98648a,a98652a,a98653a,a98656a,a98659a,a98660a,a98661a,a98665a,a98666a,a98669a,a98672a,a98673a,a98674a,a98678a,a98679a,a98682a,a98685a,a98686a,a98687a,a98691a,a98692a,a98695a,a98698a,a98699a,a98700a,a98704a,a98705a,a98708a,a98711a,a98712a,a98713a,a98717a,a98718a,a98721a,a98724a,a98725a,a98726a,a98730a,a98731a,a98734a,a98737a,a98738a,a98739a,a98743a,a98744a,a98747a,a98750a,a98751a,a98752a,a98756a,a98757a,a98760a,a98763a,a98764a,a98765a,a98769a,a98770a,a98773a,a98776a,a98777a,a98778a,a98782a,a98783a,a98786a,a98789a,a98790a,a98791a,a98795a,a98796a,a98799a,a98802a,a98803a,a98804a,a98808a,a98809a,a98812a,a98815a,a98816a,a98817a,a98821a,a98822a,a98825a,a98828a,a98829a,a98830a,a98834a,a98835a,a98838a,a98841a,a98842a,a98843a,a98847a,a98848a,a98851a,a98854a,a98855a,a98856a,a98860a,a98861a,a98864a,a98867a,a98868a,a98869a,a98873a,a98874a,a98877a,a98880a,a98881a,a98882a,a98886a,a98887a,a98890a,a98893a,a98894a,a98895a,a98899a,a98900a,a98903a,a98906a,a98907a,a98908a,a98912a,a98913a,a98916a,a98919a,a98920a,a98921a,a98925a,a98926a,a98929a,a98932a,a98933a,a98934a,a98938a,a98939a,a98942a,a98945a,a98946a,a98947a,a98951a,a98952a,a98955a,a98958a,a98959a,a98960a,a98964a,a98965a,a98968a,a98971a,a98972a,a98973a,a98977a,a98978a,a98981a,a98984a,a98985a,a98986a,a98990a,a98991a,a98994a,a98997a,a98998a,a98999a,a99003a,a99004a,a99007a,a99010a,a99011a,a99012a,a99016a,a99017a,a99020a,a99023a,a99024a,a99025a,a99029a,a99030a,a99033a,a99036a,a99037a,a99038a,a99042a,a99043a,a99046a,a99049a,a99050a,a99051a,a99055a,a99056a,a99059a,a99062a,a99063a,a99064a,a99068a,a99069a,a99072a,a99075a,a99076a,a99077a,a99081a,a99082a,a99085a,a99088a,a99089a,a99090a,a99094a,a99095a,a99098a,a99101a,a99102a,a99103a,a99107a,a99108a,a99111a,a99114a,a99115a,a99116a,a99120a,a99121a,a99124a,a99127a,a99128a,a99129a,a99133a,a99134a,a99137a,a99140a,a99141a,a99142a,a99146a,a99147a,a99150a,a99153a,a99154a,a99155a,a99159a,a99160a,a99163a,a99166a,a99167a,a99168a,a99172a,a99173a,a99176a,a99179a,a99180a,a99181a,a99185a,a99186a,a99189a,a99192a,a99193a,a99194a,a99198a,a99199a,a99202a,a99205a,a99206a,a99207a,a99211a,a99212a,a99215a,a99218a,a99219a,a99220a,a99224a,a99225a,a99228a,a99231a,a99232a,a99233a,a99237a,a99238a,a99241a,a99244a,a99245a,a99246a,a99250a,a99251a,a99254a,a99257a,a99258a,a99259a,a99263a,a99264a,a99267a,a99270a,a99271a,a99272a,a99276a,a99277a,a99280a,a99283a,a99284a,a99285a,a99289a,a99290a,a99293a,a99296a,a99297a,a99298a,a99302a,a99303a,a99306a,a99309a,a99310a,a99311a,a99315a,a99316a,a99319a,a99322a,a99323a,a99324a,a99328a,a99329a,a99332a,a99335a,a99336a,a99337a,a99341a,a99342a,a99345a,a99348a,a99349a,a99350a,a99354a,a99355a,a99358a,a99361a,a99362a,a99363a,a99367a,a99368a,a99371a,a99374a,a99375a,a99376a,a99380a,a99381a,a99384a,a99387a,a99388a,a99389a,a99393a,a99394a,a99397a,a99400a,a99401a,a99402a,a99406a,a99407a,a99410a,a99413a,a99414a,a99415a,a99419a,a99420a,a99423a,a99426a,a99427a,a99428a,a99432a,a99433a,a99436a,a99439a,a99440a,a99441a,a99445a,a99446a,a99449a,a99452a,a99453a,a99454a,a99458a,a99459a,a99462a,a99465a,a99466a,a99467a,a99471a,a99472a,a99475a,a99478a,a99479a,a99480a,a99484a,a99485a,a99488a,a99491a,a99492a,a99493a,a99497a,a99498a,a99501a,a99504a,a99505a,a99506a,a99510a,a99511a,a99514a,a99517a,a99518a,a99519a,a99523a,a99524a,a99527a,a99530a,a99531a,a99532a,a99536a,a99537a,a99540a,a99543a,a99544a,a99545a,a99549a,a99550a,a99553a,a99556a,a99557a,a99558a,a99562a,a99563a,a99566a,a99569a,a99570a,a99571a,a99575a,a99576a,a99579a,a99582a,a99583a,a99584a,a99588a,a99589a,a99592a,a99595a,a99596a,a99597a,a99601a,a99602a,a99605a,a99608a,a99609a,a99610a,a99614a,a99615a,a99618a,a99621a,a99622a,a99623a,a99627a,a99628a,a99631a,a99634a,a99635a,a99636a,a99640a,a99641a,a99644a,a99647a,a99648a,a99649a,a99653a,a99654a,a99657a,a99660a,a99661a,a99662a,a99666a,a99667a,a99670a,a99673a,a99674a,a99675a,a99679a,a99680a,a99683a,a99686a,a99687a,a99688a,a99692a,a99693a,a99696a,a99699a,a99700a,a99701a,a99705a,a99706a,a99709a,a99712a,a99713a,a99714a,a99718a,a99719a,a99722a,a99725a,a99726a,a99727a,a99731a,a99732a,a99735a,a99738a,a99739a,a99740a,a99744a,a99745a,a99748a,a99751a,a99752a,a99753a,a99757a,a99758a,a99761a,a99764a,a99765a,a99766a,a99770a,a99771a,a99774a,a99777a,a99778a,a99779a,a99783a,a99784a,a99787a,a99790a,a99791a,a99792a,a99796a,a99797a,a99800a,a99803a,a99804a,a99805a,a99809a,a99810a,a99813a,a99816a,a99817a,a99818a,a99822a,a99823a,a99826a,a99829a,a99830a,a99831a,a99835a,a99836a,a99839a,a99842a,a99843a,a99844a,a99848a,a99849a,a99852a,a99855a,a99856a,a99857a,a99861a,a99862a,a99865a,a99868a,a99869a,a99870a,a99874a,a99875a,a99878a,a99881a,a99882a,a99883a,a99887a,a99888a,a99891a,a99894a,a99895a,a99896a,a99900a,a99901a,a99904a,a99907a,a99908a,a99909a,a99913a,a99914a,a99917a,a99920a,a99921a,a99922a,a99926a,a99927a,a99930a,a99933a,a99934a,a99935a,a99939a,a99940a,a99943a,a99946a,a99947a,a99948a,a99952a,a99953a,a99956a,a99959a,a99960a,a99961a,a99965a,a99966a,a99969a,a99972a,a99973a,a99974a,a99978a,a99979a,a99982a,a99985a,a99986a,a99987a,a99991a,a99992a,a99995a,a99998a,a99999a,a100000a,a100004a,a100005a,a100008a,a100011a,a100012a,a100013a,a100017a,a100018a,a100021a,a100024a,a100025a,a100026a,a100030a,a100031a,a100034a,a100037a,a100038a,a100039a,a100043a,a100044a,a100047a,a100050a,a100051a,a100052a,a100056a,a100057a,a100060a,a100063a,a100064a,a100065a,a100069a,a100070a,a100073a,a100076a,a100077a,a100078a,a100082a,a100083a,a100086a,a100089a,a100090a,a100091a,a100095a,a100096a,a100099a,a100102a,a100103a,a100104a,a100108a,a100109a,a100112a,a100115a,a100116a,a100117a,a100121a,a100122a,a100125a,a100128a,a100129a,a100130a,a100134a,a100135a,a100138a,a100141a,a100142a,a100143a,a100147a,a100148a,a100151a,a100154a,a100155a,a100156a,a100160a,a100161a,a100164a,a100167a,a100168a,a100169a,a100173a,a100174a,a100177a,a100180a,a100181a,a100182a,a100186a,a100187a,a100190a,a100193a,a100194a,a100195a,a100199a,a100200a,a100203a,a100206a,a100207a,a100208a,a100212a,a100213a,a100216a,a100219a,a100220a,a100221a,a100225a,a100226a,a100229a,a100232a,a100233a,a100234a,a100238a,a100239a,a100242a,a100245a,a100246a,a100247a,a100251a,a100252a,a100255a,a100258a,a100259a,a100260a,a100264a,a100265a,a100268a,a100271a,a100272a,a100273a,a100277a,a100278a,a100281a,a100284a,a100285a,a100286a,a100290a,a100291a,a100294a,a100297a,a100298a,a100299a,a100303a,a100304a,a100307a,a100310a,a100311a,a100312a,a100316a,a100317a,a100320a,a100323a,a100324a,a100325a,a100329a,a100330a,a100333a,a100336a,a100337a,a100338a,a100342a,a100343a,a100346a,a100349a,a100350a,a100351a,a100355a,a100356a,a100359a,a100362a,a100363a,a100364a,a100368a,a100369a,a100372a,a100375a,a100376a,a100377a,a100381a,a100382a,a100385a,a100388a,a100389a,a100390a,a100394a,a100395a,a100398a,a100401a,a100402a,a100403a,a100407a,a100408a,a100411a,a100414a,a100415a,a100416a,a100420a,a100421a,a100424a,a100427a,a100428a,a100429a,a100433a,a100434a,a100437a,a100440a,a100441a,a100442a,a100446a,a100447a,a100450a,a100453a,a100454a,a100455a,a100459a,a100460a,a100463a,a100466a,a100467a,a100468a,a100472a,a100473a,a100476a,a100479a,a100480a,a100481a,a100485a,a100486a,a100489a,a100492a,a100493a,a100494a,a100498a,a100499a,a100502a,a100505a,a100506a,a100507a,a100511a,a100512a,a100515a,a100518a,a100519a,a100520a,a100524a,a100525a,a100528a,a100531a,a100532a,a100533a,a100537a,a100538a,a100541a,a100544a,a100545a,a100546a,a100550a,a100551a,a100554a,a100557a,a100558a,a100559a,a100563a,a100564a,a100567a,a100570a,a100571a,a100572a,a100576a,a100577a,a100580a,a100583a,a100584a,a100585a,a100589a,a100590a,a100593a,a100596a,a100597a,a100598a,a100602a,a100603a,a100606a,a100609a,a100610a,a100611a,a100615a,a100616a,a100619a,a100622a,a100623a,a100624a,a100628a,a100629a,a100632a,a100635a,a100636a,a100637a,a100641a,a100642a,a100645a,a100648a,a100649a,a100650a,a100654a,a100655a,a100658a,a100661a,a100662a,a100663a,a100667a,a100668a,a100671a,a100674a,a100675a,a100676a,a100680a,a100681a,a100684a,a100687a,a100688a,a100689a,a100693a,a100694a,a100697a,a100700a,a100701a,a100702a,a100706a,a100707a,a100710a,a100713a,a100714a,a100715a,a100719a,a100720a,a100723a,a100726a,a100727a,a100728a,a100732a,a100733a,a100736a,a100739a,a100740a,a100741a,a100745a,a100746a,a100749a,a100752a,a100753a,a100754a,a100758a,a100759a,a100762a,a100765a,a100766a,a100767a,a100771a,a100772a,a100775a,a100778a,a100779a,a100780a,a100784a,a100785a,a100788a,a100791a,a100792a,a100793a,a100797a,a100798a,a100801a,a100804a,a100805a,a100806a,a100810a,a100811a,a100814a,a100817a,a100818a,a100819a,a100823a,a100824a,a100827a,a100830a,a100831a,a100832a,a100836a,a100837a,a100840a,a100843a,a100844a,a100845a,a100849a,a100850a,a100853a,a100856a,a100857a,a100858a,a100862a,a100863a,a100866a,a100869a,a100870a,a100871a,a100875a,a100876a,a100879a,a100882a,a100883a,a100884a,a100888a,a100889a,a100892a,a100895a,a100896a,a100897a,a100901a,a100902a,a100905a,a100908a,a100909a,a100910a,a100914a,a100915a,a100918a,a100921a,a100922a,a100923a,a100927a,a100928a,a100931a,a100934a,a100935a,a100936a,a100940a,a100941a,a100944a,a100947a,a100948a,a100949a,a100953a,a100954a,a100957a,a100960a,a100961a,a100962a,a100966a,a100967a,a100970a,a100973a,a100974a,a100975a,a100979a,a100980a,a100983a,a100986a,a100987a,a100988a,a100992a,a100993a,a100996a,a100999a,a101000a,a101001a,a101005a,a101006a,a101009a,a101012a,a101013a,a101014a,a101018a,a101019a,a101022a,a101025a,a101026a,a101027a,a101031a,a101032a,a101035a,a101038a,a101039a,a101040a,a101044a,a101045a,a101048a,a101051a,a101052a,a101053a,a101057a,a101058a,a101061a,a101064a,a101065a,a101066a,a101070a,a101071a,a101074a,a101077a,a101078a,a101079a,a101083a,a101084a,a101087a,a101090a,a101091a,a101092a,a101096a,a101097a,a101100a,a101103a,a101104a,a101105a,a101109a,a101110a,a101113a,a101116a,a101117a,a101118a,a101122a,a101123a,a101126a,a101129a,a101130a,a101131a,a101135a,a101136a,a101139a,a101142a,a101143a,a101144a,a101148a,a101149a,a101152a,a101155a,a101156a,a101157a,a101161a,a101162a,a101165a,a101168a,a101169a,a101170a,a101174a,a101175a,a101178a,a101181a,a101182a,a101183a,a101187a,a101188a,a101191a,a101194a,a101195a,a101196a,a101200a,a101201a,a101204a,a101207a,a101208a,a101209a,a101213a,a101214a,a101217a,a101220a,a101221a,a101222a,a101226a,a101227a,a101230a,a101233a,a101234a,a101235a,a101239a,a101240a,a101243a,a101246a,a101247a,a101248a,a101252a,a101253a,a101256a,a101259a,a101260a,a101261a,a101265a,a101266a,a101269a,a101272a,a101273a,a101274a,a101278a,a101279a,a101282a,a101285a,a101286a,a101287a,a101291a,a101292a,a101295a,a101298a,a101299a,a101300a,a101304a,a101305a,a101308a,a101311a,a101312a,a101313a,a101317a,a101318a,a101321a,a101324a,a101325a,a101326a,a101330a,a101331a,a101334a,a101337a,a101338a,a101339a,a101343a,a101344a,a101347a,a101350a,a101351a,a101352a,a101356a,a101357a,a101360a,a101363a,a101364a,a101365a,a101369a,a101370a,a101373a,a101376a,a101377a,a101378a,a101382a,a101383a,a101386a,a101389a,a101390a,a101391a,a101395a,a101396a,a101399a,a101402a,a101403a,a101404a,a101408a,a101409a,a101412a,a101415a,a101416a,a101417a,a101421a,a101422a,a101425a,a101428a,a101429a,a101430a,a101434a,a101435a,a101438a,a101441a,a101442a,a101443a,a101447a,a101448a,a101451a,a101454a,a101455a,a101456a,a101460a,a101461a,a101464a,a101467a,a101468a,a101469a,a101473a,a101474a,a101477a,a101480a,a101481a,a101482a,a101486a,a101487a,a101490a,a101493a,a101494a,a101495a,a101499a,a101500a,a101503a,a101506a,a101507a,a101508a,a101512a,a101513a,a101516a,a101519a,a101520a,a101521a,a101525a,a101526a,a101529a,a101532a,a101533a,a101534a,a101538a,a101539a,a101542a,a101545a,a101546a,a101547a,a101551a,a101552a,a101555a,a101558a,a101559a,a101560a,a101564a,a101565a,a101568a,a101571a,a101572a,a101573a,a101577a,a101578a,a101581a,a101584a,a101585a,a101586a,a101590a,a101591a,a101594a,a101597a,a101598a,a101599a,a101603a,a101604a,a101607a,a101610a,a101611a,a101612a,a101616a,a101617a,a101620a,a101623a,a101624a,a101625a,a101629a,a101630a,a101633a,a101636a,a101637a,a101638a,a101642a,a101643a,a101646a,a101649a,a101650a,a101651a,a101655a,a101656a,a101659a,a101662a,a101663a,a101664a,a101668a,a101669a,a101672a,a101675a,a101676a,a101677a,a101681a,a101682a,a101685a,a101688a,a101689a,a101690a,a101694a,a101695a,a101698a,a101701a,a101702a,a101703a,a101707a,a101708a,a101711a,a101714a,a101715a,a101716a,a101720a,a101721a,a101724a,a101727a,a101728a,a101729a,a101733a,a101734a,a101737a,a101740a,a101741a,a101742a,a101746a,a101747a,a101750a,a101753a,a101754a,a101755a,a101759a,a101760a,a101763a,a101766a,a101767a,a101768a,a101772a,a101773a,a101776a,a101779a,a101780a,a101781a,a101785a,a101786a,a101789a,a101792a,a101793a,a101794a,a101798a,a101799a,a101802a,a101805a,a101806a,a101807a,a101811a,a101812a,a101815a,a101818a,a101819a,a101820a,a101824a,a101825a,a101828a,a101831a,a101832a,a101833a,a101837a,a101838a,a101841a,a101844a,a101845a,a101846a,a101850a,a101851a,a101854a,a101857a,a101858a,a101859a,a101863a,a101864a,a101867a,a101870a,a101871a,a101872a,a101876a,a101877a,a101880a,a101883a,a101884a,a101885a,a101889a,a101890a,a101893a,a101896a,a101897a,a101898a,a101902a,a101903a,a101906a,a101909a,a101910a,a101911a,a101915a,a101916a,a101919a,a101922a,a101923a,a101924a,a101928a,a101929a,a101932a,a101935a,a101936a,a101937a,a101941a,a101942a,a101945a,a101948a,a101949a,a101950a,a101954a,a101955a,a101958a,a101961a,a101962a,a101963a,a101967a,a101968a,a101971a,a101974a,a101975a,a101976a,a101980a,a101981a,a101984a,a101987a,a101988a,a101989a,a101993a,a101994a,a101997a,a102000a,a102001a,a102002a,a102006a,a102007a,a102010a,a102013a,a102014a,a102015a,a102019a,a102020a,a102023a,a102026a,a102027a,a102028a,a102032a,a102033a,a102036a,a102039a,a102040a,a102041a,a102045a,a102046a,a102049a,a102052a,a102053a,a102054a,a102058a,a102059a,a102062a,a102065a,a102066a,a102067a,a102071a,a102072a,a102075a,a102078a,a102079a,a102080a,a102084a,a102085a,a102088a,a102091a,a102092a,a102093a,a102097a,a102098a,a102101a,a102104a,a102105a,a102106a,a102110a,a102111a,a102114a,a102117a,a102118a,a102119a,a102123a,a102124a,a102127a,a102130a,a102131a,a102132a,a102136a,a102137a,a102140a,a102143a,a102144a,a102145a,a102149a,a102150a,a102153a,a102156a,a102157a,a102158a,a102162a,a102163a,a102166a,a102169a,a102170a,a102171a,a102175a,a102176a,a102179a,a102182a,a102183a,a102184a,a102188a,a102189a,a102192a,a102195a,a102196a,a102197a,a102201a,a102202a,a102205a,a102208a,a102209a,a102210a,a102214a,a102215a,a102218a,a102221a,a102222a,a102223a,a102227a,a102228a,a102231a,a102234a,a102235a,a102236a,a102240a,a102241a,a102244a,a102247a,a102248a,a102249a,a102253a,a102254a,a102257a,a102260a,a102261a,a102262a,a102266a,a102267a,a102270a,a102273a,a102274a,a102275a,a102279a,a102280a,a102283a,a102286a,a102287a,a102288a,a102292a,a102293a,a102296a,a102299a,a102300a,a102301a,a102305a,a102306a,a102309a,a102312a,a102313a,a102314a,a102318a,a102319a,a102322a,a102325a,a102326a,a102327a,a102331a,a102332a,a102335a,a102338a,a102339a,a102340a,a102344a,a102345a,a102348a,a102351a,a102352a,a102353a,a102357a,a102358a,a102361a,a102364a,a102365a,a102366a,a102370a,a102371a,a102374a,a102377a,a102378a,a102379a,a102383a,a102384a,a102387a,a102390a,a102391a,a102392a,a102396a,a102397a,a102400a,a102403a,a102404a,a102405a,a102409a,a102410a,a102413a,a102416a,a102417a,a102418a,a102422a,a102423a,a102426a,a102429a,a102430a,a102431a,a102435a,a102436a,a102439a,a102442a,a102443a,a102444a,a102448a,a102449a,a102452a,a102455a,a102456a,a102457a,a102461a,a102462a,a102465a,a102468a,a102469a,a102470a,a102474a,a102475a,a102478a,a102481a,a102482a,a102483a,a102487a,a102488a,a102491a,a102494a,a102495a,a102496a,a102500a,a102501a,a102504a,a102507a,a102508a,a102509a,a102513a,a102514a,a102517a,a102520a,a102521a,a102522a,a102526a,a102527a,a102530a,a102533a,a102534a,a102535a,a102539a,a102540a,a102543a,a102546a,a102547a,a102548a,a102552a,a102553a,a102556a,a102559a,a102560a,a102561a,a102565a,a102566a,a102569a,a102572a,a102573a,a102574a,a102578a,a102579a,a102582a,a102585a,a102586a,a102587a,a102591a,a102592a,a102595a,a102598a,a102599a,a102600a,a102604a,a102605a,a102608a,a102611a,a102612a,a102613a,a102617a,a102618a,a102621a,a102624a,a102625a,a102626a,a102630a,a102631a,a102634a,a102637a,a102638a,a102639a,a102643a,a102644a,a102647a,a102650a,a102651a,a102652a,a102656a,a102657a,a102660a,a102663a,a102664a,a102665a,a102669a,a102670a,a102673a,a102676a,a102677a,a102678a,a102682a,a102683a,a102686a,a102689a,a102690a,a102691a,a102695a,a102696a,a102699a,a102702a,a102703a,a102704a,a102708a,a102709a,a102712a,a102715a,a102716a,a102717a,a102721a,a102722a,a102725a,a102728a,a102729a,a102730a,a102734a,a102735a,a102738a,a102741a,a102742a,a102743a,a102747a,a102748a,a102751a,a102754a,a102755a,a102756a,a102760a,a102761a,a102764a,a102767a,a102768a,a102769a,a102773a,a102774a,a102777a,a102780a,a102781a,a102782a,a102786a,a102787a,a102790a,a102793a,a102794a,a102795a,a102799a,a102800a,a102803a,a102806a,a102807a,a102808a,a102812a,a102813a,a102816a,a102819a,a102820a,a102821a,a102825a,a102826a,a102829a,a102832a,a102833a,a102834a,a102838a,a102839a,a102842a,a102845a,a102846a,a102847a,a102851a,a102852a,a102855a,a102858a,a102859a,a102860a,a102864a,a102865a,a102868a,a102871a,a102872a,a102873a,a102877a,a102878a,a102881a,a102884a,a102885a,a102886a,a102890a,a102891a,a102894a,a102897a,a102898a,a102899a,a102903a,a102904a,a102907a,a102910a,a102911a,a102912a,a102916a,a102917a,a102920a,a102923a,a102924a,a102925a,a102929a,a102930a,a102933a,a102936a,a102937a,a102938a,a102942a,a102943a,a102946a,a102949a,a102950a,a102951a,a102955a,a102956a,a102959a,a102962a,a102963a,a102964a,a102968a,a102969a,a102972a,a102975a,a102976a,a102977a,a102980a,a102983a,a102984a,a102987a,a102990a,a102991a,a102992a,a102996a,a102997a,a103000a,a103003a,a103004a,a103005a,a103008a,a103011a,a103012a,a103015a,a103018a,a103019a,a103020a,a103024a,a103025a,a103028a,a103031a,a103032a,a103033a,a103036a,a103039a,a103040a,a103043a,a103046a,a103047a,a103048a,a103052a,a103053a,a103056a,a103059a,a103060a,a103061a,a103064a,a103067a,a103068a,a103071a,a103074a,a103075a,a103076a,a103080a,a103081a,a103084a,a103087a,a103088a,a103089a,a103092a,a103095a,a103096a,a103099a,a103102a,a103103a,a103104a,a103108a,a103109a,a103112a,a103115a,a103116a,a103117a,a103120a,a103123a,a103124a,a103127a,a103130a,a103131a,a103132a,a103136a,a103137a,a103140a,a103143a,a103144a,a103145a,a103148a,a103151a,a103152a,a103155a,a103158a,a103159a,a103160a,a103164a,a103165a,a103168a,a103171a,a103172a,a103173a,a103176a,a103179a,a103180a,a103183a,a103186a,a103187a,a103188a,a103192a,a103193a,a103196a,a103199a,a103200a,a103201a,a103204a,a103207a,a103208a,a103211a,a103214a,a103215a,a103216a,a103220a,a103221a,a103224a,a103227a,a103228a,a103229a,a103232a,a103235a,a103236a,a103239a,a103242a,a103243a,a103244a,a103248a,a103249a,a103252a,a103255a,a103256a,a103257a,a103260a,a103263a,a103264a,a103267a,a103270a,a103271a,a103272a,a103276a,a103277a,a103280a,a103283a,a103284a,a103285a,a103288a,a103291a,a103292a,a103295a,a103298a,a103299a,a103300a,a103304a,a103305a,a103308a,a103311a,a103312a,a103313a,a103316a,a103319a,a103320a,a103323a,a103326a,a103327a,a103328a,a103332a,a103333a,a103336a,a103339a,a103340a,a103341a,a103344a,a103347a,a103348a,a103351a,a103354a,a103355a,a103356a,a103360a,a103361a,a103364a,a103367a,a103368a,a103369a,a103372a,a103375a,a103376a,a103379a,a103382a,a103383a,a103384a,a103388a,a103389a,a103392a,a103395a,a103396a,a103397a,a103400a,a103403a,a103404a,a103407a,a103410a,a103411a,a103412a,a103416a,a103417a,a103420a,a103423a,a103424a,a103425a,a103428a,a103431a,a103432a,a103435a,a103438a,a103439a,a103440a,a103444a,a103445a,a103448a,a103451a,a103452a,a103453a,a103456a,a103459a,a103460a,a103463a,a103466a,a103467a,a103468a,a103472a,a103473a,a103476a,a103479a,a103480a,a103481a,a103484a,a103487a,a103488a,a103491a,a103494a,a103495a,a103496a,a103500a,a103501a,a103504a,a103507a,a103508a,a103509a,a103512a,a103515a,a103516a,a103519a,a103522a,a103523a,a103524a,a103528a,a103529a,a103532a,a103535a,a103536a,a103537a,a103540a,a103543a,a103544a,a103547a,a103550a,a103551a,a103552a,a103556a,a103557a,a103560a,a103563a,a103564a,a103565a,a103568a,a103571a,a103572a,a103575a,a103578a,a103579a,a103580a,a103584a,a103585a,a103588a,a103591a,a103592a,a103593a,a103596a,a103599a,a103600a,a103603a,a103606a,a103607a,a103608a,a103612a,a103613a,a103616a,a103619a,a103620a,a103621a,a103624a,a103627a,a103628a,a103631a,a103634a,a103635a,a103636a,a103640a,a103641a,a103644a,a103647a,a103648a,a103649a,a103652a,a103655a,a103656a,a103659a,a103662a,a103663a,a103664a,a103668a,a103669a,a103672a,a103675a,a103676a,a103677a,a103680a,a103683a,a103684a,a103687a,a103690a,a103691a,a103692a,a103696a,a103697a,a103700a,a103703a,a103704a,a103705a,a103708a,a103711a,a103712a,a103715a,a103718a,a103719a,a103720a,a103724a,a103725a,a103728a,a103731a,a103732a,a103733a,a103736a,a103739a,a103740a,a103743a,a103746a,a103747a,a103748a,a103752a,a103753a,a103756a,a103759a,a103760a,a103761a,a103764a,a103767a,a103768a,a103771a,a103774a,a103775a,a103776a,a103780a,a103781a,a103784a,a103787a,a103788a,a103789a,a103792a,a103795a,a103796a,a103799a,a103802a,a103803a,a103804a,a103808a,a103809a,a103812a,a103815a,a103816a,a103817a,a103820a,a103823a,a103824a,a103827a,a103830a,a103831a,a103832a,a103836a,a103837a,a103840a,a103843a,a103844a,a103845a,a103848a,a103851a,a103852a,a103855a,a103858a,a103859a,a103860a,a103864a,a103865a,a103868a,a103871a,a103872a,a103873a,a103876a,a103879a,a103880a,a103883a,a103886a,a103887a,a103888a,a103892a,a103893a,a103896a,a103899a,a103900a,a103901a,a103904a,a103907a,a103908a,a103911a,a103914a,a103915a,a103916a,a103920a,a103921a,a103924a,a103927a,a103928a,a103929a,a103932a,a103935a,a103936a,a103939a,a103942a,a103943a,a103944a,a103948a,a103949a,a103952a,a103955a,a103956a,a103957a,a103960a,a103963a,a103964a,a103967a,a103970a,a103971a,a103972a,a103976a,a103977a,a103980a,a103983a,a103984a,a103985a,a103988a,a103991a,a103992a,a103995a,a103998a,a103999a,a104000a,a104004a,a104005a,a104008a,a104011a,a104012a,a104013a,a104016a,a104019a,a104020a,a104023a,a104026a,a104027a,a104028a,a104032a,a104033a,a104036a,a104039a,a104040a,a104041a,a104044a,a104047a,a104048a,a104051a,a104054a,a104055a,a104056a,a104060a,a104061a,a104064a,a104067a,a104068a,a104069a,a104072a,a104075a,a104076a,a104079a,a104082a,a104083a,a104084a,a104088a,a104089a,a104092a,a104095a,a104096a,a104097a,a104100a,a104103a,a104104a,a104107a,a104110a,a104111a,a104112a,a104116a,a104117a,a104120a,a104123a,a104124a,a104125a,a104128a,a104131a,a104132a,a104135a,a104138a,a104139a,a104140a,a104144a,a104145a,a104148a,a104151a,a104152a,a104153a,a104156a,a104159a,a104160a,a104163a,a104166a,a104167a,a104168a,a104172a,a104173a,a104176a,a104179a,a104180a,a104181a,a104184a,a104187a,a104188a,a104191a,a104194a,a104195a,a104196a,a104200a,a104201a,a104204a,a104207a,a104208a,a104209a,a104212a,a104215a,a104216a,a104219a,a104222a,a104223a,a104224a,a104228a,a104229a,a104232a,a104235a,a104236a,a104237a,a104240a,a104243a,a104244a,a104247a,a104250a,a104251a,a104252a,a104256a,a104257a,a104260a,a104263a,a104264a,a104265a,a104268a,a104271a,a104272a,a104275a,a104278a,a104279a,a104280a,a104284a,a104285a,a104288a,a104291a,a104292a,a104293a,a104296a,a104299a,a104300a,a104303a,a104306a,a104307a,a104308a,a104312a,a104313a,a104316a,a104319a,a104320a,a104321a,a104324a,a104327a,a104328a,a104331a,a104334a,a104335a,a104336a,a104340a,a104341a,a104344a,a104347a,a104348a,a104349a,a104352a,a104355a,a104356a,a104359a,a104362a,a104363a,a104364a,a104368a,a104369a,a104372a,a104375a,a104376a,a104377a,a104380a,a104383a,a104384a,a104387a,a104390a,a104391a,a104392a,a104396a,a104397a,a104400a,a104403a,a104404a,a104405a,a104408a,a104411a,a104412a,a104415a,a104418a,a104419a,a104420a,a104424a,a104425a,a104428a,a104431a,a104432a,a104433a,a104436a,a104439a,a104440a,a104443a,a104446a,a104447a,a104448a,a104452a,a104453a,a104456a,a104459a,a104460a,a104461a,a104464a,a104467a,a104468a,a104471a,a104474a,a104475a,a104476a,a104480a,a104481a,a104484a,a104487a,a104488a,a104489a,a104492a,a104495a,a104496a,a104499a,a104502a,a104503a,a104504a,a104508a,a104509a,a104512a,a104515a,a104516a,a104517a,a104520a,a104523a,a104524a,a104527a,a104530a,a104531a,a104532a,a104536a,a104537a,a104540a,a104543a,a104544a,a104545a,a104548a,a104551a,a104552a,a104555a,a104558a,a104559a,a104560a,a104564a,a104565a,a104568a,a104571a,a104572a,a104573a,a104576a,a104579a,a104580a,a104583a,a104586a,a104587a,a104588a,a104592a,a104593a,a104596a,a104599a,a104600a,a104601a,a104604a,a104607a,a104608a,a104611a,a104614a,a104615a,a104616a,a104620a,a104621a,a104624a,a104627a,a104628a,a104629a,a104632a,a104635a,a104636a,a104639a,a104642a,a104643a,a104644a,a104648a,a104649a,a104652a,a104655a,a104656a,a104657a,a104660a,a104663a,a104664a,a104667a,a104670a,a104671a,a104672a,a104676a,a104677a,a104680a,a104683a,a104684a,a104685a,a104688a,a104691a,a104692a,a104695a,a104698a,a104699a,a104700a,a104704a,a104705a,a104708a,a104711a,a104712a,a104713a,a104716a,a104719a,a104720a,a104723a,a104726a,a104727a,a104728a,a104732a,a104733a,a104736a,a104739a,a104740a,a104741a,a104744a,a104747a,a104748a,a104751a,a104754a,a104755a,a104756a,a104760a,a104761a,a104764a,a104767a,a104768a,a104769a,a104772a,a104775a,a104776a,a104779a,a104782a,a104783a,a104784a,a104788a,a104789a,a104792a,a104795a,a104796a,a104797a,a104800a,a104803a,a104804a,a104807a,a104810a,a104811a,a104812a,a104816a,a104817a,a104820a,a104823a,a104824a,a104825a,a104828a,a104831a,a104832a,a104835a,a104838a,a104839a,a104840a,a104844a,a104845a,a104848a,a104851a,a104852a,a104853a,a104856a,a104859a,a104860a,a104863a,a104866a,a104867a,a104868a,a104872a,a104873a,a104876a,a104879a,a104880a,a104881a,a104884a,a104887a,a104888a,a104891a,a104894a,a104895a,a104896a,a104900a,a104901a,a104904a,a104907a,a104908a,a104909a,a104912a,a104915a,a104916a,a104919a,a104922a,a104923a,a104924a,a104928a,a104929a,a104932a,a104935a,a104936a,a104937a,a104940a,a104943a,a104944a,a104947a,a104950a,a104951a,a104952a,a104956a,a104957a,a104960a,a104963a,a104964a,a104965a,a104968a,a104971a,a104972a,a104975a,a104978a,a104979a,a104980a,a104984a,a104985a,a104988a,a104991a,a104992a,a104993a,a104996a,a104999a,a105000a,a105003a,a105006a,a105007a,a105008a,a105012a,a105013a,a105016a,a105019a,a105020a,a105021a,a105024a,a105027a,a105028a,a105031a,a105034a,a105035a,a105036a,a105040a,a105041a,a105044a,a105047a,a105048a,a105049a,a105052a,a105055a,a105056a,a105059a,a105062a,a105063a,a105064a,a105068a,a105069a,a105072a,a105075a,a105076a,a105077a,a105080a,a105083a,a105084a,a105087a,a105090a,a105091a,a105092a,a105096a,a105097a,a105100a,a105103a,a105104a,a105105a,a105108a,a105111a,a105112a,a105115a,a105118a,a105119a,a105120a,a105124a,a105125a,a105128a,a105131a,a105132a,a105133a,a105136a,a105139a,a105140a,a105143a,a105146a,a105147a,a105148a,a105152a,a105153a,a105156a,a105159a,a105160a,a105161a,a105164a,a105167a,a105168a,a105171a,a105174a,a105175a,a105176a,a105180a,a105181a,a105184a,a105187a,a105188a,a105189a,a105192a,a105195a,a105196a,a105199a,a105202a,a105203a,a105204a,a105208a,a105209a,a105212a,a105215a,a105216a,a105217a,a105220a,a105223a,a105224a,a105227a,a105230a,a105231a,a105232a,a105236a,a105237a,a105240a,a105243a,a105244a,a105245a,a105248a,a105251a,a105252a,a105255a,a105258a,a105259a,a105260a,a105264a,a105265a,a105268a,a105271a,a105272a,a105273a,a105276a,a105279a,a105280a,a105283a,a105286a,a105287a,a105288a,a105292a,a105293a,a105296a,a105299a,a105300a,a105301a,a105304a,a105307a,a105308a,a105311a,a105314a,a105315a,a105316a,a105320a,a105321a,a105324a,a105327a,a105328a,a105329a,a105332a,a105335a,a105336a,a105339a,a105342a,a105343a,a105344a,a105348a,a105349a,a105352a,a105355a,a105356a,a105357a,a105360a,a105363a,a105364a,a105367a,a105370a,a105371a,a105372a,a105376a,a105377a,a105380a,a105383a,a105384a,a105385a,a105388a,a105391a,a105392a,a105395a,a105398a,a105399a,a105400a,a105404a,a105405a,a105408a,a105411a,a105412a,a105413a,a105416a,a105419a,a105420a,a105423a,a105426a,a105427a,a105428a,a105432a,a105433a,a105436a,a105439a,a105440a,a105441a,a105444a,a105447a,a105448a,a105451a,a105454a,a105455a,a105456a,a105460a,a105461a,a105464a,a105467a,a105468a,a105469a,a105472a,a105475a,a105476a,a105479a,a105482a,a105483a,a105484a,a105488a,a105489a,a105492a,a105495a,a105496a,a105497a,a105500a,a105503a,a105504a,a105507a,a105510a,a105511a,a105512a,a105516a,a105517a,a105520a,a105523a,a105524a,a105525a,a105528a,a105531a,a105532a,a105535a,a105538a,a105539a,a105540a,a105544a,a105545a,a105548a,a105551a,a105552a,a105553a,a105556a,a105559a,a105560a,a105563a,a105566a,a105567a,a105568a,a105572a,a105573a,a105576a,a105579a,a105580a,a105581a,a105584a,a105587a,a105588a,a105591a,a105594a,a105595a,a105596a,a105600a,a105601a,a105604a,a105607a,a105608a,a105609a,a105612a,a105615a,a105616a,a105619a,a105622a,a105623a,a105624a,a105628a,a105629a,a105632a,a105635a,a105636a,a105637a,a105640a,a105643a,a105644a,a105647a,a105650a,a105651a,a105652a,a105656a,a105657a,a105660a,a105663a,a105664a,a105665a,a105668a,a105671a,a105672a,a105675a,a105678a,a105679a,a105680a,a105684a,a105685a,a105688a,a105691a,a105692a,a105693a,a105696a,a105699a,a105700a,a105703a,a105706a,a105707a,a105708a,a105712a,a105713a,a105716a,a105719a,a105720a,a105721a,a105724a,a105727a,a105728a,a105731a,a105734a,a105735a,a105736a,a105740a,a105741a,a105744a,a105747a,a105748a,a105749a,a105752a,a105755a,a105756a,a105759a,a105762a,a105763a,a105764a,a105768a,a105769a,a105772a,a105775a,a105776a,a105777a,a105780a,a105783a,a105784a,a105787a,a105790a,a105791a,a105792a,a105796a,a105797a,a105800a,a105803a,a105804a,a105805a,a105808a,a105811a,a105812a,a105815a,a105818a,a105819a,a105820a,a105824a,a105825a,a105828a,a105831a,a105832a,a105833a,a105836a,a105839a,a105840a,a105843a,a105846a,a105847a,a105848a,a105852a,a105853a,a105856a,a105859a,a105860a,a105861a,a105864a,a105867a,a105868a,a105871a,a105874a,a105875a,a105876a,a105880a,a105881a,a105884a,a105887a,a105888a,a105889a,a105892a,a105895a,a105896a,a105899a,a105902a,a105903a,a105904a,a105908a,a105909a,a105912a,a105915a,a105916a,a105917a,a105920a,a105923a,a105924a,a105927a,a105930a,a105931a,a105932a,a105936a,a105937a,a105940a,a105943a,a105944a,a105945a,a105948a,a105951a,a105952a,a105955a,a105958a,a105959a,a105960a,a105964a,a105965a,a105968a,a105971a,a105972a,a105973a,a105976a,a105979a,a105980a,a105983a,a105986a,a105987a,a105988a,a105992a,a105993a,a105996a,a105999a,a106000a,a106001a,a106004a,a106007a,a106008a,a106011a,a106014a,a106015a,a106016a,a106020a,a106021a,a106024a,a106027a,a106028a,a106029a,a106032a,a106035a,a106036a,a106039a,a106042a,a106043a,a106044a,a106048a,a106049a,a106052a,a106055a,a106056a,a106057a,a106060a,a106063a,a106064a,a106067a,a106070a,a106071a,a106072a,a106076a,a106077a,a106080a,a106083a,a106084a,a106085a,a106088a,a106091a,a106092a,a106095a,a106098a,a106099a,a106100a,a106104a,a106105a,a106108a,a106111a,a106112a,a106113a,a106116a,a106119a,a106120a,a106123a,a106126a,a106127a,a106128a,a106132a,a106133a,a106136a,a106139a,a106140a,a106141a,a106144a,a106147a,a106148a,a106151a,a106154a,a106155a,a106156a,a106160a,a106161a,a106164a,a106167a,a106168a,a106169a,a106172a,a106175a,a106176a,a106179a,a106182a,a106183a,a106184a,a106188a,a106189a,a106192a,a106195a,a106196a,a106197a,a106200a,a106203a,a106204a,a106207a,a106210a,a106211a,a106212a,a106216a,a106217a,a106220a,a106223a,a106224a,a106225a,a106228a,a106231a,a106232a,a106235a,a106238a,a106239a,a106240a,a106244a,a106245a,a106248a,a106251a,a106252a,a106253a,a106256a,a106259a,a106260a,a106263a,a106266a,a106267a,a106268a,a106272a,a106273a,a106276a,a106279a,a106280a,a106281a,a106284a,a106287a,a106288a,a106291a,a106294a,a106295a,a106296a,a106300a,a106301a,a106304a,a106307a,a106308a,a106309a,a106312a,a106315a,a106316a,a106319a,a106322a,a106323a,a106324a,a106328a,a106329a,a106332a,a106335a,a106336a,a106337a,a106340a,a106343a,a106344a,a106347a,a106350a,a106351a,a106352a,a106356a,a106357a,a106360a,a106363a,a106364a,a106365a,a106368a,a106371a,a106372a,a106375a,a106378a,a106379a,a106380a,a106384a,a106385a,a106388a,a106391a,a106392a,a106393a,a106396a,a106399a,a106400a,a106403a,a106406a,a106407a,a106408a,a106412a,a106413a,a106416a,a106419a,a106420a,a106421a,a106424a,a106427a,a106428a,a106431a,a106434a,a106435a,a106436a,a106440a,a106441a,a106444a,a106447a,a106448a,a106449a,a106452a,a106455a,a106456a,a106459a,a106462a,a106463a,a106464a,a106468a,a106469a,a106472a,a106475a,a106476a,a106477a,a106480a,a106483a,a106484a,a106487a,a106490a,a106491a,a106492a,a106496a,a106497a,a106500a,a106503a,a106504a,a106505a,a106508a,a106511a,a106512a,a106515a,a106518a,a106519a,a106520a,a106524a,a106525a,a106528a,a106531a,a106532a,a106533a,a106536a,a106539a,a106540a,a106543a,a106546a,a106547a,a106548a,a106552a,a106553a,a106556a,a106559a,a106560a,a106561a,a106564a,a106567a,a106568a,a106571a,a106574a,a106575a,a106576a,a106580a,a106581a,a106584a,a106587a,a106588a,a106589a,a106592a,a106595a,a106596a,a106599a,a106602a,a106603a,a106604a,a106608a,a106609a,a106612a,a106615a,a106616a,a106617a,a106620a,a106623a,a106624a,a106627a,a106630a,a106631a,a106632a,a106636a,a106637a,a106640a,a106643a,a106644a,a106645a,a106648a,a106651a,a106652a,a106655a,a106658a,a106659a,a106660a,a106664a,a106665a,a106668a,a106671a,a106672a,a106673a,a106676a,a106679a,a106680a,a106683a,a106686a,a106687a,a106688a,a106692a,a106693a,a106696a,a106699a,a106700a,a106701a,a106704a,a106707a,a106708a,a106711a,a106714a,a106715a,a106716a,a106720a,a106721a,a106724a,a106727a,a106728a,a106729a,a106732a,a106735a,a106736a,a106739a,a106742a,a106743a,a106744a,a106748a,a106749a,a106752a,a106755a,a106756a,a106757a,a106760a,a106763a,a106764a,a106767a,a106770a,a106771a,a106772a,a106776a,a106777a,a106780a,a106783a,a106784a,a106785a,a106788a,a106791a,a106792a,a106795a,a106798a,a106799a,a106800a,a106804a,a106805a,a106808a,a106811a,a106812a,a106813a,a106816a,a106819a,a106820a,a106823a,a106826a,a106827a,a106828a,a106832a,a106833a,a106836a,a106839a,a106840a,a106841a,a106844a,a106847a,a106848a,a106851a,a106854a,a106855a,a106856a,a106860a,a106861a,a106864a,a106867a,a106868a,a106869a,a106872a,a106875a,a106876a,a106879a,a106882a,a106883a,a106884a,a106888a,a106889a,a106892a,a106895a,a106896a,a106897a,a106900a,a106903a,a106904a,a106907a,a106910a,a106911a,a106912a,a106916a,a106917a,a106920a,a106923a,a106924a,a106925a,a106928a,a106931a,a106932a,a106935a,a106938a,a106939a,a106940a,a106944a,a106945a,a106948a,a106951a,a106952a,a106953a,a106956a,a106959a,a106960a,a106963a,a106966a,a106967a,a106968a,a106972a,a106973a,a106976a,a106979a,a106980a,a106981a,a106984a,a106987a,a106988a,a106991a,a106994a,a106995a,a106996a,a107000a,a107001a,a107004a,a107007a,a107008a,a107009a,a107012a,a107015a,a107016a,a107019a,a107022a,a107023a,a107024a,a107028a,a107029a,a107032a,a107035a,a107036a,a107037a,a107040a,a107043a,a107044a,a107047a,a107050a,a107051a,a107052a,a107056a,a107057a,a107060a,a107063a,a107064a,a107065a,a107068a,a107071a,a107072a,a107075a,a107078a,a107079a,a107080a,a107084a,a107085a,a107088a,a107091a,a107092a,a107093a,a107096a,a107099a,a107100a,a107103a,a107106a,a107107a,a107108a,a107112a,a107113a,a107116a,a107119a,a107120a,a107121a,a107124a,a107127a,a107128a,a107131a,a107134a,a107135a,a107136a,a107140a,a107141a,a107144a,a107147a,a107148a,a107149a,a107152a,a107155a,a107156a,a107159a,a107162a,a107163a,a107164a,a107168a,a107169a,a107172a,a107175a,a107176a,a107177a,a107180a,a107183a,a107184a,a107187a,a107190a,a107191a,a107192a,a107196a,a107197a,a107200a,a107203a,a107204a,a107205a,a107208a,a107211a,a107212a,a107215a,a107218a,a107219a,a107220a,a107224a,a107225a,a107228a,a107231a,a107232a,a107233a,a107236a,a107239a,a107240a,a107243a,a107246a,a107247a,a107248a,a107252a,a107253a,a107256a,a107259a,a107260a,a107261a,a107264a,a107267a,a107268a,a107271a,a107274a,a107275a,a107276a,a107280a,a107281a,a107284a,a107287a,a107288a,a107289a,a107292a,a107295a,a107296a,a107299a,a107302a,a107303a,a107304a,a107308a,a107309a,a107312a,a107315a,a107316a,a107317a,a107320a,a107323a,a107324a,a107327a,a107330a,a107331a,a107332a,a107336a,a107337a,a107340a,a107343a,a107344a,a107345a,a107348a,a107351a,a107352a,a107355a,a107358a,a107359a,a107360a,a107364a,a107365a,a107368a,a107371a,a107372a,a107373a,a107376a,a107379a,a107380a,a107383a,a107386a,a107387a,a107388a,a107392a,a107393a,a107396a,a107399a,a107400a,a107401a,a107404a,a107407a,a107408a,a107411a,a107414a,a107415a,a107416a,a107420a,a107421a,a107424a,a107427a,a107428a,a107429a,a107432a,a107435a,a107436a,a107439a,a107442a,a107443a,a107444a,a107448a,a107449a,a107452a,a107455a,a107456a,a107457a,a107460a,a107463a,a107464a,a107467a,a107470a,a107471a,a107472a,a107476a,a107477a,a107480a,a107483a,a107484a,a107485a,a107488a,a107491a,a107492a,a107495a,a107498a,a107499a,a107500a,a107504a,a107505a,a107508a,a107511a,a107512a,a107513a,a107516a,a107519a,a107520a,a107523a,a107526a,a107527a,a107528a,a107532a,a107533a,a107536a,a107539a,a107540a,a107541a,a107544a,a107547a,a107548a,a107551a,a107554a,a107555a,a107556a,a107560a,a107561a,a107564a,a107567a,a107568a,a107569a,a107572a,a107575a,a107576a,a107579a,a107582a,a107583a,a107584a,a107588a,a107589a,a107592a,a107595a,a107596a,a107597a,a107600a,a107603a,a107604a,a107607a,a107610a,a107611a,a107612a,a107616a,a107617a,a107620a,a107623a,a107624a,a107625a,a107628a,a107631a,a107632a,a107635a,a107638a,a107639a,a107640a,a107644a,a107645a,a107648a,a107651a,a107652a,a107653a,a107656a,a107659a,a107660a,a107663a,a107666a,a107667a,a107668a,a107672a,a107673a,a107676a,a107679a,a107680a,a107681a,a107684a,a107687a,a107688a,a107691a,a107694a,a107695a,a107696a,a107700a,a107701a,a107704a,a107707a,a107708a,a107709a,a107712a,a107715a,a107716a,a107719a,a107722a,a107723a,a107724a,a107728a,a107729a,a107732a,a107735a,a107736a,a107737a,a107740a,a107743a,a107744a,a107747a,a107750a,a107751a,a107752a,a107756a,a107757a,a107760a,a107763a,a107764a,a107765a,a107768a,a107771a,a107772a,a107775a,a107778a,a107779a,a107780a,a107784a,a107785a,a107788a,a107791a,a107792a,a107793a,a107796a,a107799a,a107800a,a107803a,a107806a,a107807a,a107808a,a107812a,a107813a,a107816a,a107819a,a107820a,a107821a,a107824a,a107827a,a107828a,a107831a,a107834a,a107835a,a107836a,a107840a,a107841a,a107844a,a107847a,a107848a,a107849a,a107852a,a107855a,a107856a,a107859a,a107862a,a107863a,a107864a,a107868a,a107869a,a107872a,a107875a,a107876a,a107877a,a107880a,a107883a,a107884a,a107887a,a107890a,a107891a,a107892a,a107896a,a107897a,a107900a,a107903a,a107904a,a107905a,a107908a,a107911a,a107912a,a107915a,a107918a,a107919a,a107920a,a107924a,a107925a,a107928a,a107931a,a107932a,a107933a,a107936a,a107939a,a107940a,a107943a,a107946a,a107947a,a107948a,a107952a,a107953a,a107956a,a107959a,a107960a,a107961a,a107964a,a107967a,a107968a,a107971a,a107974a,a107975a,a107976a,a107980a,a107981a,a107984a,a107987a,a107988a,a107989a,a107992a,a107995a,a107996a,a107999a,a108002a,a108003a,a108004a,a108008a,a108009a,a108012a,a108015a,a108016a,a108017a,a108020a,a108023a,a108024a,a108027a,a108030a,a108031a,a108032a,a108036a,a108037a,a108040a,a108043a,a108044a,a108045a,a108048a,a108051a,a108052a,a108055a,a108058a,a108059a,a108060a,a108064a,a108065a,a108068a,a108071a,a108072a,a108073a,a108076a,a108079a,a108080a,a108083a,a108086a,a108087a,a108088a,a108092a,a108093a,a108096a,a108099a,a108100a,a108101a,a108104a,a108107a,a108108a,a108111a,a108114a,a108115a,a108116a,a108120a,a108121a,a108124a,a108127a,a108128a,a108129a,a108132a,a108135a,a108136a,a108139a,a108142a,a108143a,a108144a,a108148a,a108149a,a108152a,a108155a,a108156a,a108157a,a108160a,a108163a,a108164a,a108167a,a108170a,a108171a,a108172a,a108176a,a108177a,a108180a,a108183a,a108184a,a108185a,a108188a,a108191a,a108192a,a108195a,a108198a,a108199a,a108200a,a108204a,a108205a,a108208a,a108211a,a108212a,a108213a,a108216a,a108219a,a108220a,a108223a,a108226a,a108227a,a108228a,a108232a,a108233a,a108236a,a108239a,a108240a,a108241a,a108244a,a108247a,a108248a,a108251a,a108254a,a108255a,a108256a,a108260a,a108261a,a108264a,a108267a,a108268a,a108269a,a108272a,a108275a,a108276a,a108279a,a108282a,a108283a,a108284a,a108288a,a108289a,a108292a,a108295a,a108296a,a108297a,a108300a,a108303a,a108304a,a108307a,a108310a,a108311a,a108312a,a108316a,a108317a,a108320a,a108323a,a108324a,a108325a,a108328a,a108331a,a108332a,a108335a,a108338a,a108339a,a108340a,a108344a,a108345a,a108348a,a108351a,a108352a,a108353a,a108356a,a108359a,a108360a,a108363a,a108366a,a108367a,a108368a,a108372a,a108373a,a108376a,a108379a,a108380a,a108381a,a108384a,a108387a,a108388a,a108391a,a108394a,a108395a,a108396a,a108400a,a108401a,a108404a,a108407a,a108408a,a108409a,a108412a,a108415a,a108416a,a108419a,a108422a,a108423a,a108424a,a108428a,a108429a,a108432a,a108435a,a108436a,a108437a,a108440a,a108443a,a108444a,a108447a,a108450a,a108451a,a108452a,a108456a,a108457a,a108460a,a108463a,a108464a,a108465a,a108468a,a108471a,a108472a,a108475a,a108478a,a108479a,a108480a,a108484a,a108485a,a108488a,a108491a,a108492a,a108493a,a108496a,a108499a,a108500a,a108503a,a108506a,a108507a,a108508a,a108512a,a108513a,a108516a,a108519a,a108520a,a108521a,a108524a,a108527a,a108528a,a108531a,a108534a,a108535a,a108536a,a108540a,a108541a,a108544a,a108547a,a108548a,a108549a,a108552a,a108555a,a108556a,a108559a,a108562a,a108563a,a108564a,a108568a,a108569a,a108572a,a108575a,a108576a,a108577a,a108580a,a108583a,a108584a,a108587a,a108590a,a108591a,a108592a,a108596a,a108597a,a108600a,a108603a,a108604a,a108605a,a108608a,a108611a,a108612a,a108615a,a108618a,a108619a,a108620a,a108624a,a108625a,a108628a,a108631a,a108632a,a108633a,a108636a,a108639a,a108640a,a108643a,a108646a,a108647a,a108648a,a108652a,a108653a,a108656a,a108659a,a108660a,a108661a,a108664a,a108667a,a108668a,a108671a,a108674a,a108675a,a108676a,a108680a,a108681a,a108684a,a108687a,a108688a,a108689a,a108692a,a108695a,a108696a,a108699a,a108702a,a108703a,a108704a,a108708a,a108709a,a108712a,a108715a,a108716a,a108717a,a108720a,a108723a,a108724a,a108727a,a108730a,a108731a,a108732a,a108736a,a108737a,a108740a,a108743a,a108744a,a108745a,a108748a,a108751a,a108752a,a108755a,a108758a,a108759a,a108760a,a108764a,a108765a,a108768a,a108771a,a108772a,a108773a,a108776a,a108779a,a108780a,a108783a,a108786a,a108787a,a108788a,a108792a,a108793a,a108796a,a108799a,a108800a,a108801a,a108804a,a108807a,a108808a,a108811a,a108814a,a108815a,a108816a,a108820a,a108821a,a108824a,a108827a,a108828a,a108829a,a108832a,a108835a,a108836a,a108839a,a108842a,a108843a,a108844a,a108848a,a108849a,a108852a,a108855a,a108856a,a108857a,a108860a,a108863a,a108864a,a108867a,a108870a,a108871a,a108872a,a108876a,a108877a,a108880a,a108883a,a108884a,a108885a,a108888a,a108891a,a108892a,a108895a,a108898a,a108899a,a108900a,a108904a,a108905a,a108908a,a108911a,a108912a,a108913a,a108916a,a108919a,a108920a,a108923a,a108926a,a108927a,a108928a,a108932a,a108933a,a108936a,a108939a,a108940a,a108941a,a108944a,a108947a,a108948a,a108951a,a108954a,a108955a,a108956a,a108960a,a108961a,a108964a,a108967a,a108968a,a108969a,a108972a,a108975a,a108976a,a108979a,a108982a,a108983a,a108984a,a108988a,a108989a,a108992a,a108995a,a108996a,a108997a,a109000a,a109003a,a109004a,a109007a,a109010a,a109011a,a109012a,a109016a,a109017a,a109020a,a109023a,a109024a,a109025a,a109028a,a109031a,a109032a,a109035a,a109038a,a109039a,a109040a,a109044a,a109045a,a109048a,a109051a,a109052a,a109053a,a109056a,a109059a,a109060a,a109063a,a109066a,a109067a,a109068a,a109072a,a109073a,a109076a,a109079a,a109080a,a109081a,a109084a,a109087a,a109088a,a109091a,a109094a,a109095a,a109096a,a109100a,a109101a,a109104a,a109107a,a109108a,a109109a,a109112a,a109115a,a109116a,a109119a,a109122a,a109123a,a109124a,a109128a,a109129a,a109132a,a109135a,a109136a,a109137a,a109140a,a109143a,a109144a,a109147a,a109150a,a109151a,a109152a,a109156a,a109157a,a109160a,a109163a,a109164a,a109165a,a109168a,a109171a,a109172a,a109175a,a109178a,a109179a,a109180a,a109184a,a109185a,a109188a,a109191a,a109192a,a109193a,a109196a,a109199a,a109200a,a109203a,a109206a,a109207a,a109208a,a109212a,a109213a,a109216a,a109219a,a109220a,a109221a,a109224a,a109227a,a109228a,a109231a,a109234a,a109235a,a109236a,a109240a,a109241a,a109244a,a109247a,a109248a,a109249a,a109252a,a109255a,a109256a,a109259a,a109262a,a109263a,a109264a,a109268a,a109269a,a109272a,a109275a,a109276a,a109277a,a109280a,a109283a,a109284a,a109287a,a109290a,a109291a,a109292a,a109296a,a109297a,a109300a,a109303a,a109304a,a109305a,a109308a,a109311a,a109312a,a109315a,a109318a,a109319a,a109320a,a109324a,a109325a,a109328a,a109331a,a109332a,a109333a,a109336a,a109339a,a109340a,a109343a,a109346a,a109347a,a109348a,a109352a,a109353a,a109356a,a109359a,a109360a,a109361a,a109364a,a109367a,a109368a,a109371a,a109374a,a109375a,a109376a,a109380a,a109381a,a109384a,a109387a,a109388a,a109389a,a109392a,a109395a,a109396a,a109399a,a109402a,a109403a,a109404a,a109408a,a109409a,a109412a,a109415a,a109416a,a109417a,a109420a,a109423a,a109424a,a109427a,a109430a,a109431a,a109432a,a109436a,a109437a,a109440a,a109443a,a109444a,a109445a,a109448a,a109451a,a109452a,a109455a,a109458a,a109459a,a109460a,a109464a,a109465a,a109468a,a109471a,a109472a,a109473a,a109476a,a109479a,a109480a,a109483a,a109486a,a109487a,a109488a,a109492a,a109493a,a109496a,a109499a,a109500a,a109501a,a109504a,a109507a,a109508a,a109511a,a109514a,a109515a,a109516a,a109520a,a109521a,a109524a,a109527a,a109528a,a109529a,a109532a,a109535a,a109536a,a109539a,a109542a,a109543a,a109544a,a109548a,a109549a,a109552a,a109555a,a109556a,a109557a,a109560a,a109563a,a109564a,a109567a,a109570a,a109571a,a109572a,a109576a,a109577a,a109580a,a109583a,a109584a,a109585a,a109588a,a109591a,a109592a,a109595a,a109598a,a109599a,a109600a,a109604a,a109605a,a109608a,a109611a,a109612a,a109613a,a109616a,a109619a,a109620a,a109623a,a109626a,a109627a,a109628a,a109632a,a109633a,a109636a,a109639a,a109640a,a109641a,a109644a,a109647a,a109648a,a109651a,a109654a,a109655a,a109656a,a109660a,a109661a,a109664a,a109667a,a109668a,a109669a,a109672a,a109675a,a109676a,a109679a,a109682a,a109683a,a109684a,a109688a,a109689a,a109692a,a109695a,a109696a,a109697a,a109700a,a109703a,a109704a,a109707a,a109710a,a109711a,a109712a,a109716a,a109717a,a109720a,a109723a,a109724a,a109725a,a109728a,a109731a,a109732a,a109735a,a109738a,a109739a,a109740a,a109744a,a109745a,a109748a,a109751a,a109752a,a109753a,a109756a,a109759a,a109760a,a109763a,a109766a,a109767a,a109768a,a109772a,a109773a,a109776a,a109779a,a109780a,a109781a,a109784a,a109787a,a109788a,a109791a,a109794a,a109795a,a109796a,a109800a,a109801a,a109804a,a109807a,a109808a,a109809a,a109812a,a109815a,a109816a,a109819a,a109822a,a109823a,a109824a,a109828a,a109829a,a109832a,a109835a,a109836a,a109837a,a109840a,a109843a,a109844a,a109847a,a109850a,a109851a,a109852a,a109856a,a109857a,a109860a,a109863a,a109864a,a109865a,a109868a,a109871a,a109872a,a109875a,a109878a,a109879a,a109880a,a109884a,a109885a,a109888a,a109891a,a109892a,a109893a,a109896a,a109899a,a109900a,a109903a,a109906a,a109907a,a109908a,a109912a,a109913a,a109916a,a109919a,a109920a,a109921a,a109924a,a109927a,a109928a,a109931a,a109934a,a109935a,a109936a,a109940a,a109941a,a109944a,a109947a,a109948a,a109949a,a109952a,a109955a,a109956a,a109959a,a109962a,a109963a,a109964a,a109968a,a109969a,a109972a,a109975a,a109976a,a109977a,a109980a,a109983a,a109984a,a109987a,a109990a,a109991a,a109992a,a109996a,a109997a,a110000a,a110003a,a110004a,a110005a,a110008a,a110011a,a110012a,a110015a,a110018a,a110019a,a110020a,a110024a,a110025a,a110028a,a110031a,a110032a,a110033a,a110036a,a110039a,a110040a,a110043a,a110046a,a110047a,a110048a,a110052a,a110053a,a110056a,a110059a,a110060a,a110061a,a110064a,a110067a,a110068a,a110071a,a110074a,a110075a,a110076a,a110080a,a110081a,a110084a,a110087a,a110088a,a110089a,a110092a,a110095a,a110096a,a110099a,a110102a,a110103a,a110104a,a110108a,a110109a,a110112a,a110115a,a110116a,a110117a,a110120a,a110123a,a110124a,a110127a,a110130a,a110131a,a110132a,a110136a,a110137a,a110140a,a110143a,a110144a,a110145a,a110148a,a110151a,a110152a,a110155a,a110158a,a110159a,a110160a,a110164a,a110165a,a110168a,a110171a,a110172a,a110173a,a110176a,a110179a,a110180a,a110183a,a110186a,a110187a,a110188a,a110192a,a110193a,a110196a,a110199a,a110200a,a110201a,a110204a,a110207a,a110208a,a110211a,a110214a,a110215a,a110216a,a110220a,a110221a,a110224a,a110227a,a110228a,a110229a,a110232a,a110235a,a110236a,a110239a,a110242a,a110243a,a110244a,a110248a,a110249a,a110252a,a110255a,a110256a,a110257a,a110260a,a110263a,a110264a,a110267a,a110270a,a110271a,a110272a,a110276a,a110277a,a110280a,a110283a,a110284a,a110285a,a110288a,a110291a,a110292a,a110295a,a110298a,a110299a,a110300a,a110304a,a110305a,a110308a,a110311a,a110312a,a110313a,a110316a,a110319a,a110320a,a110323a,a110326a,a110327a,a110328a,a110332a,a110333a,a110336a,a110339a,a110340a,a110341a,a110344a,a110347a,a110348a,a110351a,a110354a,a110355a,a110356a,a110360a,a110361a,a110364a,a110367a,a110368a,a110369a,a110372a,a110375a,a110376a,a110379a,a110382a,a110383a,a110384a,a110388a,a110389a,a110392a,a110395a,a110396a,a110397a,a110400a,a110403a,a110404a,a110407a,a110410a,a110411a,a110412a,a110416a,a110417a,a110420a,a110423a,a110424a,a110425a,a110428a,a110431a,a110432a,a110435a,a110438a,a110439a,a110440a,a110444a,a110445a,a110448a,a110451a,a110452a,a110453a,a110456a,a110459a,a110460a,a110463a,a110466a,a110467a,a110468a,a110472a,a110473a,a110476a,a110479a,a110480a,a110481a,a110484a,a110487a,a110488a,a110491a,a110494a,a110495a,a110496a,a110500a,a110501a,a110504a,a110507a,a110508a,a110509a,a110512a,a110515a,a110516a,a110519a,a110522a,a110523a,a110524a,a110528a,a110529a,a110532a,a110535a,a110536a,a110537a,a110540a,a110543a,a110544a,a110547a,a110550a,a110551a,a110552a,a110556a,a110557a,a110560a,a110563a,a110564a,a110565a,a110568a,a110571a,a110572a,a110575a,a110578a,a110579a,a110580a,a110584a,a110585a,a110588a,a110591a,a110592a,a110593a,a110596a,a110599a,a110600a,a110603a,a110606a,a110607a,a110608a,a110612a,a110613a,a110616a,a110619a,a110620a,a110621a,a110624a,a110627a,a110628a,a110631a,a110634a,a110635a,a110636a,a110640a,a110641a,a110644a,a110647a,a110648a,a110649a,a110652a,a110655a,a110656a,a110659a,a110662a,a110663a,a110664a,a110668a,a110669a,a110672a,a110675a,a110676a,a110677a,a110680a,a110683a,a110684a,a110687a,a110690a,a110691a,a110692a,a110696a,a110697a,a110700a,a110703a,a110704a,a110705a,a110708a,a110711a,a110712a,a110715a,a110718a,a110719a,a110720a,a110724a,a110725a,a110728a,a110731a,a110732a,a110733a,a110736a,a110739a,a110740a,a110743a,a110746a,a110747a,a110748a,a110752a,a110753a,a110756a,a110759a,a110760a,a110761a,a110764a,a110767a,a110768a,a110771a,a110774a,a110775a,a110776a,a110780a,a110781a,a110784a,a110787a,a110788a,a110789a,a110792a,a110795a,a110796a,a110799a,a110802a,a110803a,a110804a,a110808a,a110809a,a110812a,a110815a,a110816a,a110817a,a110820a,a110823a,a110824a,a110827a,a110830a,a110831a,a110832a,a110836a,a110837a,a110840a,a110843a,a110844a,a110845a,a110848a,a110851a,a110852a,a110855a,a110858a,a110859a,a110860a,a110864a,a110865a,a110868a,a110871a,a110872a,a110873a,a110876a,a110879a,a110880a,a110883a,a110886a,a110887a,a110888a,a110892a,a110893a,a110896a,a110899a,a110900a,a110901a,a110904a,a110907a,a110908a,a110911a,a110914a,a110915a,a110916a,a110920a,a110921a,a110924a,a110927a,a110928a,a110929a,a110932a,a110935a,a110936a,a110939a,a110942a,a110943a,a110944a,a110948a,a110949a,a110952a,a110955a,a110956a,a110957a,a110960a,a110963a,a110964a,a110967a,a110970a,a110971a,a110972a,a110976a,a110977a,a110980a,a110983a,a110984a,a110985a,a110988a,a110991a,a110992a,a110995a,a110998a,a110999a,a111000a,a111004a,a111005a,a111008a,a111011a,a111012a,a111013a,a111016a,a111019a,a111020a,a111023a,a111026a,a111027a,a111028a,a111032a,a111033a,a111036a,a111039a,a111040a,a111041a,a111044a,a111047a,a111048a,a111051a,a111054a,a111055a,a111056a,a111060a,a111061a,a111064a,a111067a,a111068a,a111069a,a111072a,a111075a,a111076a,a111079a,a111082a,a111083a,a111084a,a111088a,a111089a,a111092a,a111095a,a111096a,a111097a,a111100a,a111103a,a111104a,a111107a,a111110a,a111111a,a111112a,a111116a,a111117a,a111120a,a111123a,a111124a,a111125a,a111128a,a111131a,a111132a,a111135a,a111138a,a111139a,a111140a,a111144a,a111145a,a111148a,a111151a,a111152a,a111153a,a111156a,a111159a,a111160a,a111163a,a111166a,a111167a,a111168a,a111172a,a111173a,a111176a,a111179a,a111180a,a111181a,a111184a,a111187a,a111188a,a111191a,a111194a,a111195a,a111196a,a111200a,a111201a,a111204a,a111207a,a111208a,a111209a,a111212a,a111215a,a111216a,a111219a,a111222a,a111223a,a111224a,a111228a,a111229a,a111232a,a111235a,a111236a,a111237a,a111240a,a111243a,a111244a,a111247a,a111250a,a111251a,a111252a,a111256a,a111257a,a111260a,a111263a,a111264a,a111265a,a111268a,a111271a,a111272a,a111275a,a111278a,a111279a,a111280a,a111284a,a111285a,a111288a,a111291a,a111292a,a111293a,a111296a,a111299a,a111300a,a111303a,a111306a,a111307a,a111308a,a111312a,a111313a,a111316a,a111319a,a111320a,a111321a,a111324a,a111327a,a111328a,a111331a,a111334a,a111335a,a111336a,a111340a,a111341a,a111344a,a111347a,a111348a,a111349a,a111352a,a111355a,a111356a,a111359a,a111362a,a111363a,a111364a,a111368a,a111369a,a111372a,a111375a,a111376a,a111377a,a111380a,a111383a,a111384a,a111387a,a111390a,a111391a,a111392a,a111396a,a111397a,a111400a,a111403a,a111404a,a111405a,a111408a,a111411a,a111412a,a111415a,a111418a,a111419a,a111420a,a111424a,a111425a,a111428a,a111431a,a111432a,a111433a,a111436a,a111439a,a111440a,a111443a,a111446a,a111447a,a111448a,a111452a,a111453a,a111456a,a111459a,a111460a,a111461a,a111464a,a111467a,a111468a,a111471a,a111474a,a111475a,a111476a,a111480a,a111481a,a111484a,a111487a,a111488a,a111489a,a111492a,a111495a,a111496a,a111499a,a111502a,a111503a,a111504a,a111508a,a111509a,a111512a,a111515a,a111516a,a111517a,a111520a,a111523a,a111524a,a111527a,a111530a,a111531a,a111532a,a111536a,a111537a,a111540a,a111543a,a111544a,a111545a,a111548a,a111551a,a111552a,a111555a,a111558a,a111559a,a111560a,a111564a,a111565a,a111568a,a111571a,a111572a,a111573a,a111576a,a111579a,a111580a,a111583a,a111586a,a111587a,a111588a,a111592a,a111593a,a111596a,a111599a,a111600a,a111601a,a111604a,a111607a,a111608a,a111611a,a111614a,a111615a,a111616a,a111620a,a111621a,a111624a,a111627a,a111628a,a111629a,a111632a,a111635a,a111636a,a111639a,a111642a,a111643a,a111644a,a111648a,a111649a,a111652a,a111655a,a111656a,a111657a,a111660a,a111663a,a111664a,a111667a,a111670a,a111671a,a111672a,a111676a,a111677a,a111680a,a111683a,a111684a,a111685a,a111688a,a111691a,a111692a,a111695a,a111698a,a111699a,a111700a,a111704a,a111705a,a111708a,a111711a,a111712a,a111713a,a111716a,a111719a,a111720a,a111723a,a111726a,a111727a,a111728a,a111732a,a111733a,a111736a,a111739a,a111740a,a111741a,a111744a,a111747a,a111748a,a111751a,a111754a,a111755a,a111756a,a111760a,a111761a,a111764a,a111767a,a111768a,a111769a,a111772a,a111775a,a111776a,a111779a,a111782a,a111783a,a111784a,a111788a,a111789a,a111792a,a111795a,a111796a,a111797a,a111800a,a111803a,a111804a,a111807a,a111810a,a111811a,a111812a,a111816a,a111817a,a111820a,a111823a,a111824a,a111825a,a111828a,a111831a,a111832a,a111835a,a111838a,a111839a,a111840a,a111844a,a111845a,a111848a,a111851a,a111852a,a111853a,a111856a,a111859a,a111860a,a111863a,a111866a,a111867a,a111868a,a111872a,a111873a,a111876a,a111879a,a111880a,a111881a,a111884a,a111887a,a111888a,a111891a,a111894a,a111895a,a111896a,a111900a,a111901a,a111904a,a111907a,a111908a,a111909a,a111912a,a111915a,a111916a,a111919a,a111922a,a111923a,a111924a,a111928a,a111929a,a111932a,a111935a,a111936a,a111937a,a111940a,a111943a,a111944a,a111947a,a111950a,a111951a,a111952a,a111956a,a111957a,a111960a,a111963a,a111964a,a111965a,a111968a,a111971a,a111972a,a111975a,a111978a,a111979a,a111980a,a111984a,a111985a,a111988a,a111991a,a111992a,a111993a,a111996a,a111999a,a112000a,a112003a,a112006a,a112007a,a112008a,a112012a,a112013a,a112016a,a112019a,a112020a,a112021a,a112024a,a112027a,a112028a,a112031a,a112034a,a112035a,a112036a,a112040a,a112041a,a112044a,a112047a,a112048a,a112049a,a112052a,a112055a,a112056a,a112059a,a112062a,a112063a,a112064a,a112068a,a112069a,a112072a,a112075a,a112076a,a112077a,a112080a,a112083a,a112084a,a112087a,a112090a,a112091a,a112092a,a112096a,a112097a,a112100a,a112103a,a112104a,a112105a,a112108a,a112111a,a112112a,a112115a,a112118a,a112119a,a112120a,a112124a,a112125a,a112128a,a112131a,a112132a,a112133a,a112136a,a112139a,a112140a,a112143a,a112146a,a112147a,a112148a,a112152a,a112153a,a112156a,a112159a,a112160a,a112161a,a112164a,a112167a,a112168a,a112171a,a112174a,a112175a,a112176a,a112180a,a112181a,a112184a,a112187a,a112188a,a112189a,a112192a,a112195a,a112196a,a112199a,a112202a,a112203a,a112204a,a112208a,a112209a,a112212a,a112215a,a112216a,a112217a,a112220a,a112223a,a112224a,a112227a,a112230a,a112231a,a112232a,a112236a,a112237a,a112240a,a112243a,a112244a,a112245a,a112248a,a112251a,a112252a,a112255a,a112258a,a112259a,a112260a,a112264a,a112265a,a112268a,a112271a,a112272a,a112273a,a112276a,a112279a,a112280a,a112283a,a112286a,a112287a,a112288a,a112292a,a112293a,a112296a,a112299a,a112300a,a112301a,a112304a,a112307a,a112308a,a112311a,a112314a,a112315a,a112316a,a112320a,a112321a,a112324a,a112327a,a112328a,a112329a,a112332a,a112335a,a112336a,a112339a,a112342a,a112343a,a112344a,a112348a,a112349a,a112352a,a112355a,a112356a,a112357a,a112360a,a112363a,a112364a,a112367a,a112370a,a112371a,a112372a,a112376a,a112377a,a112380a,a112383a,a112384a,a112385a,a112388a,a112391a,a112392a,a112395a,a112398a,a112399a,a112400a,a112404a,a112405a,a112408a,a112411a,a112412a,a112413a,a112416a,a112419a,a112420a,a112423a,a112426a,a112427a,a112428a,a112432a,a112433a,a112436a,a112439a,a112440a,a112441a,a112444a,a112447a,a112448a,a112451a,a112454a,a112455a,a112456a,a112460a,a112461a,a112464a,a112467a,a112468a,a112469a,a112472a,a112475a,a112476a,a112479a,a112482a,a112483a,a112484a,a112488a,a112489a,a112492a,a112495a,a112496a,a112497a,a112500a,a112503a,a112504a,a112507a,a112510a,a112511a,a112512a,a112516a,a112517a,a112520a,a112523a,a112524a,a112525a,a112528a,a112531a,a112532a,a112535a,a112538a,a112539a,a112540a,a112544a,a112545a,a112548a,a112551a,a112552a,a112553a,a112556a,a112559a,a112560a,a112563a,a112566a,a112567a,a112568a,a112572a,a112573a,a112576a,a112579a,a112580a,a112581a,a112584a,a112587a,a112588a,a112591a,a112594a,a112595a,a112596a,a112600a,a112601a,a112604a,a112607a,a112608a,a112609a,a112612a,a112615a,a112616a,a112619a,a112622a,a112623a,a112624a,a112628a,a112629a,a112632a,a112635a,a112636a,a112637a,a112640a,a112643a,a112644a,a112647a,a112650a,a112651a,a112652a,a112656a,a112657a,a112660a,a112663a,a112664a,a112665a,a112668a,a112671a,a112672a,a112675a,a112678a,a112679a,a112680a,a112684a,a112685a,a112688a,a112691a,a112692a,a112693a,a112696a,a112699a,a112700a,a112703a,a112706a,a112707a,a112708a,a112712a,a112713a,a112716a,a112719a,a112720a,a112721a,a112724a,a112727a,a112728a,a112731a,a112734a,a112735a,a112736a,a112740a,a112741a,a112744a,a112747a,a112748a,a112749a,a112752a,a112755a,a112756a,a112759a,a112762a,a112763a,a112764a,a112768a,a112769a,a112772a,a112775a,a112776a,a112777a,a112780a,a112783a,a112784a,a112787a,a112790a,a112791a,a112792a,a112796a,a112797a,a112800a,a112803a,a112804a,a112805a,a112808a,a112811a,a112812a,a112815a,a112818a,a112819a,a112820a,a112824a,a112825a,a112828a,a112831a,a112832a,a112833a,a112836a,a112839a,a112840a,a112843a,a112846a,a112847a,a112848a,a112852a,a112853a,a112856a,a112859a,a112860a,a112861a,a112864a,a112867a,a112868a,a112871a,a112874a,a112875a,a112876a,a112880a,a112881a,a112884a,a112887a,a112888a,a112889a,a112892a,a112895a,a112896a,a112899a,a112902a,a112903a,a112904a,a112908a,a112909a,a112912a,a112915a,a112916a,a112917a,a112920a,a112923a,a112924a,a112927a,a112930a,a112931a,a112932a,a112936a,a112937a,a112940a,a112943a,a112944a,a112945a,a112948a,a112951a,a112952a,a112955a,a112958a,a112959a,a112960a,a112964a,a112965a,a112968a,a112971a,a112972a,a112973a,a112976a,a112979a,a112980a,a112983a,a112986a,a112987a,a112988a,a112992a,a112993a,a112996a,a112999a,a113000a,a113001a,a113004a,a113007a,a113008a,a113011a,a113014a,a113015a,a113016a,a113020a,a113021a,a113024a,a113027a,a113028a,a113029a,a113032a,a113035a,a113036a,a113039a,a113042a,a113043a,a113044a,a113048a,a113049a,a113052a,a113055a,a113056a,a113057a,a113060a,a113063a,a113064a,a113067a,a113070a,a113071a,a113072a,a113076a,a113077a,a113080a,a113083a,a113084a,a113085a,a113088a,a113091a,a113092a,a113095a,a113098a,a113099a,a113100a,a113104a,a113105a,a113108a,a113111a,a113112a,a113113a,a113116a,a113119a,a113120a,a113123a,a113126a,a113127a,a113128a,a113132a,a113133a,a113136a,a113139a,a113140a,a113141a,a113144a,a113147a,a113148a,a113151a,a113154a,a113155a,a113156a,a113160a,a113161a,a113164a,a113167a,a113168a,a113169a,a113172a,a113175a,a113176a,a113179a,a113182a,a113183a,a113184a,a113188a,a113189a,a113192a,a113195a,a113196a,a113197a,a113200a,a113203a,a113204a,a113207a,a113210a,a113211a,a113212a,a113216a,a113217a,a113220a,a113223a,a113224a,a113225a,a113228a,a113231a,a113232a,a113235a,a113238a,a113239a,a113240a,a113244a,a113245a,a113248a,a113251a,a113252a,a113253a,a113256a,a113259a,a113260a,a113263a,a113266a,a113267a,a113268a,a113272a,a113273a,a113276a,a113279a,a113280a,a113281a,a113284a,a113287a,a113288a,a113291a,a113294a,a113295a,a113296a,a113300a,a113301a,a113304a,a113307a,a113308a,a113309a,a113312a,a113315a,a113316a,a113319a,a113322a,a113323a,a113324a,a113328a,a113329a,a113332a,a113335a,a113336a,a113337a,a113340a,a113343a,a113344a,a113347a,a113350a,a113351a,a113352a,a113356a,a113357a,a113360a,a113363a,a113364a,a113365a,a113368a,a113371a,a113372a,a113375a,a113378a,a113379a,a113380a,a113384a,a113385a,a113388a,a113391a,a113392a,a113393a,a113396a,a113399a,a113400a,a113403a,a113406a,a113407a,a113408a,a113412a,a113413a,a113416a,a113419a,a113420a,a113421a,a113424a,a113427a,a113428a,a113431a,a113434a,a113435a,a113436a,a113440a,a113441a,a113444a,a113447a,a113448a,a113449a,a113452a,a113455a,a113456a,a113459a,a113462a,a113463a,a113464a,a113468a,a113469a,a113472a,a113475a,a113476a,a113477a,a113480a,a113483a,a113484a,a113487a,a113490a,a113491a,a113492a,a113496a,a113497a,a113500a,a113503a,a113504a,a113505a,a113508a,a113511a,a113512a,a113515a,a113518a,a113519a,a113520a,a113524a,a113525a,a113528a,a113531a,a113532a,a113533a,a113536a,a113539a,a113540a,a113543a,a113546a,a113547a,a113548a,a113552a,a113553a,a113556a,a113559a,a113560a,a113561a,a113564a,a113567a,a113568a,a113571a,a113574a,a113575a,a113576a,a113580a,a113581a,a113584a,a113587a,a113588a,a113589a,a113592a,a113595a,a113596a,a113599a,a113602a,a113603a,a113604a,a113608a,a113609a,a113612a,a113615a,a113616a,a113617a,a113620a,a113623a,a113624a,a113627a,a113630a,a113631a,a113632a,a113636a,a113637a,a113640a,a113643a,a113644a,a113645a,a113648a,a113651a,a113652a,a113655a,a113658a,a113659a,a113660a,a113664a,a113665a,a113668a,a113671a,a113672a,a113673a,a113676a,a113679a,a113680a,a113683a,a113686a,a113687a,a113688a,a113692a,a113693a,a113696a,a113699a,a113700a,a113701a,a113704a,a113707a,a113708a,a113711a,a113714a,a113715a,a113716a,a113720a,a113721a,a113724a,a113727a,a113728a,a113729a,a113732a,a113735a,a113736a,a113739a,a113742a,a113743a,a113744a,a113748a,a113749a,a113752a,a113755a,a113756a,a113757a,a113760a,a113763a,a113764a,a113767a,a113770a,a113771a,a113772a,a113776a,a113777a,a113780a,a113783a,a113784a,a113785a,a113788a,a113791a,a113792a,a113795a,a113798a,a113799a,a113800a,a113804a,a113805a,a113808a,a113811a,a113812a,a113813a,a113816a,a113819a,a113820a,a113823a,a113826a,a113827a,a113828a,a113832a,a113833a,a113836a,a113839a,a113840a,a113841a,a113844a,a113847a,a113848a,a113851a,a113854a,a113855a,a113856a,a113860a,a113861a,a113864a,a113867a,a113868a,a113869a,a113872a,a113875a,a113876a,a113879a,a113882a,a113883a,a113884a,a113888a,a113889a,a113892a,a113895a,a113896a,a113897a,a113900a,a113903a,a113904a,a113907a,a113910a,a113911a,a113912a,a113916a,a113917a,a113920a,a113923a,a113924a,a113925a,a113928a,a113931a,a113932a,a113935a,a113938a,a113939a,a113940a,a113944a,a113945a,a113948a,a113951a,a113952a,a113953a,a113956a,a113959a,a113960a,a113963a,a113966a,a113967a,a113968a,a113972a,a113973a,a113976a,a113979a,a113980a,a113981a,a113984a,a113987a,a113988a,a113991a,a113994a,a113995a,a113996a,a114000a,a114001a,a114004a,a114007a,a114008a,a114009a,a114012a,a114015a,a114016a,a114019a,a114022a,a114023a,a114024a,a114028a,a114029a,a114032a,a114035a,a114036a,a114037a,a114040a,a114043a,a114044a,a114047a,a114050a,a114051a,a114052a,a114056a,a114057a,a114060a,a114063a,a114064a,a114065a,a114068a,a114071a,a114072a,a114075a,a114078a,a114079a,a114080a,a114084a,a114085a,a114088a,a114091a,a114092a,a114093a,a114096a,a114099a,a114100a,a114103a,a114106a,a114107a,a114108a,a114112a,a114113a,a114116a,a114119a,a114120a,a114121a,a114124a,a114127a,a114128a,a114131a,a114134a,a114135a,a114136a,a114140a,a114141a,a114144a,a114147a,a114148a,a114149a,a114152a,a114155a,a114156a,a114159a,a114162a,a114163a,a114164a,a114168a,a114169a,a114172a,a114175a,a114176a,a114177a,a114180a,a114183a,a114184a,a114187a,a114190a,a114191a,a114192a,a114196a,a114197a,a114200a,a114203a,a114204a,a114205a,a114208a,a114211a,a114212a,a114215a,a114218a,a114219a,a114220a,a114224a,a114225a,a114228a,a114231a,a114232a,a114233a,a114236a,a114239a,a114240a,a114243a,a114246a,a114247a,a114248a,a114252a,a114253a,a114256a,a114259a,a114260a,a114261a,a114264a,a114267a,a114268a,a114271a,a114274a,a114275a,a114276a,a114280a,a114281a,a114284a,a114287a,a114288a,a114289a,a114292a,a114295a,a114296a,a114299a,a114302a,a114303a,a114304a,a114308a,a114309a,a114312a,a114315a,a114316a,a114317a,a114320a,a114323a,a114324a,a114327a,a114330a,a114331a,a114332a,a114336a,a114337a,a114340a,a114343a,a114344a,a114345a,a114348a,a114351a,a114352a,a114355a,a114358a,a114359a,a114360a,a114364a,a114365a,a114368a,a114371a,a114372a,a114373a,a114376a,a114379a,a114380a,a114383a,a114386a,a114387a,a114388a,a114392a,a114393a,a114396a,a114399a,a114400a,a114401a,a114404a,a114407a,a114408a,a114411a,a114414a,a114415a,a114416a,a114420a,a114421a,a114424a,a114427a,a114428a,a114429a,a114432a,a114435a,a114436a,a114439a,a114442a,a114443a,a114444a,a114448a,a114449a,a114452a,a114455a,a114456a,a114457a,a114460a,a114463a,a114464a,a114467a,a114470a,a114471a,a114472a,a114476a,a114477a,a114480a,a114483a,a114484a,a114485a,a114488a,a114491a,a114492a,a114495a,a114498a,a114499a,a114500a,a114504a,a114505a,a114508a,a114511a,a114512a,a114513a,a114516a,a114519a,a114520a,a114523a,a114526a,a114527a,a114528a,a114532a,a114533a,a114536a,a114539a,a114540a,a114541a,a114544a,a114547a,a114548a,a114551a,a114554a,a114555a,a114556a,a114560a,a114561a,a114564a,a114567a,a114568a,a114569a,a114572a,a114575a,a114576a,a114579a,a114582a,a114583a,a114584a,a114588a,a114589a,a114592a,a114595a,a114596a,a114597a,a114600a,a114603a,a114604a,a114607a,a114610a,a114611a,a114612a,a114616a,a114617a,a114620a,a114623a,a114624a,a114625a,a114628a,a114631a,a114632a,a114635a,a114638a,a114639a,a114640a,a114644a,a114645a,a114648a,a114651a,a114652a,a114653a,a114656a,a114659a,a114660a,a114663a,a114666a,a114667a,a114668a,a114672a,a114673a,a114676a,a114679a,a114680a,a114681a,a114684a,a114687a,a114688a,a114691a,a114694a,a114695a,a114696a,a114700a,a114701a,a114704a,a114707a,a114708a,a114709a,a114712a,a114715a,a114716a,a114719a,a114722a,a114723a,a114724a,a114728a,a114729a,a114732a,a114735a,a114736a,a114737a,a114740a,a114743a,a114744a,a114747a,a114750a,a114751a,a114752a,a114756a,a114757a,a114760a,a114763a,a114764a,a114765a,a114768a,a114771a,a114772a,a114775a,a114778a,a114779a,a114780a,a114784a,a114785a,a114788a,a114791a,a114792a,a114793a,a114796a,a114799a,a114800a,a114803a,a114806a,a114807a,a114808a,a114812a,a114813a,a114816a,a114819a,a114820a,a114821a,a114824a,a114827a,a114828a,a114831a,a114834a,a114835a,a114836a,a114840a,a114841a,a114844a,a114847a,a114848a,a114849a,a114852a,a114855a,a114856a,a114859a,a114862a,a114863a,a114864a,a114868a,a114869a,a114872a,a114875a,a114876a,a114877a,a114880a,a114883a,a114884a,a114887a,a114890a,a114891a,a114892a,a114896a,a114897a,a114900a,a114903a,a114904a,a114905a,a114908a,a114911a,a114912a,a114915a,a114918a,a114919a,a114920a,a114924a,a114925a,a114928a,a114931a,a114932a,a114933a,a114936a,a114939a,a114940a,a114943a,a114946a,a114947a,a114948a,a114952a,a114953a,a114956a,a114959a,a114960a,a114961a,a114964a,a114967a,a114968a,a114971a,a114974a,a114975a,a114976a,a114980a,a114981a,a114984a,a114987a,a114988a,a114989a,a114992a,a114995a,a114996a,a114999a,a115002a,a115003a,a115004a,a115008a,a115009a,a115012a,a115015a,a115016a,a115017a,a115020a,a115023a,a115024a,a115027a,a115030a,a115031a,a115032a,a115036a,a115037a,a115040a,a115043a,a115044a,a115045a,a115048a,a115051a,a115052a,a115055a,a115058a,a115059a,a115060a,a115064a,a115065a,a115068a,a115071a,a115072a,a115073a,a115076a,a115079a,a115080a,a115083a,a115086a,a115087a,a115088a,a115092a,a115093a,a115096a,a115099a,a115100a,a115101a,a115104a,a115107a,a115108a,a115111a,a115114a,a115115a,a115116a,a115120a,a115121a,a115124a,a115127a,a115128a,a115129a,a115132a,a115135a,a115136a,a115139a,a115142a,a115143a,a115144a,a115148a,a115149a,a115152a,a115155a,a115156a,a115157a,a115160a,a115163a,a115164a,a115167a,a115170a,a115171a,a115172a,a115176a,a115177a,a115180a,a115183a,a115184a,a115185a,a115188a,a115191a,a115192a,a115195a,a115198a,a115199a,a115200a,a115204a,a115205a,a115208a,a115211a,a115212a,a115213a,a115216a,a115219a,a115220a,a115223a,a115226a,a115227a,a115228a,a115232a,a115233a,a115236a,a115239a,a115240a,a115241a,a115244a,a115247a,a115248a,a115251a,a115254a,a115255a,a115256a,a115260a,a115261a,a115264a,a115267a,a115268a,a115269a,a115272a,a115275a,a115276a,a115279a,a115282a,a115283a,a115284a,a115288a,a115289a,a115292a,a115295a,a115296a,a115297a,a115300a,a115303a,a115304a,a115307a,a115310a,a115311a,a115312a,a115316a,a115317a,a115320a,a115323a,a115324a,a115325a,a115328a,a115331a,a115332a,a115335a,a115338a,a115339a,a115340a,a115344a,a115345a,a115348a,a115351a,a115352a,a115353a,a115356a,a115359a,a115360a,a115363a,a115366a,a115367a,a115368a,a115372a,a115373a,a115376a,a115379a,a115380a,a115381a,a115384a,a115387a,a115388a,a115391a,a115394a,a115395a,a115396a,a115400a,a115401a,a115404a,a115407a,a115408a,a115409a,a115412a,a115415a,a115416a,a115419a,a115422a,a115423a,a115424a,a115428a,a115429a,a115432a,a115435a,a115436a,a115437a,a115440a,a115443a,a115444a,a115447a,a115450a,a115451a,a115452a,a115456a,a115457a,a115460a,a115463a,a115464a,a115465a,a115468a,a115471a,a115472a,a115475a,a115478a,a115479a,a115480a,a115484a,a115485a,a115488a,a115491a,a115492a,a115493a,a115496a,a115499a,a115500a,a115503a,a115506a,a115507a,a115508a,a115512a,a115513a,a115516a,a115519a,a115520a,a115521a,a115524a,a115527a,a115528a,a115531a,a115534a,a115535a,a115536a,a115540a,a115541a,a115544a,a115547a,a115548a,a115549a,a115552a,a115555a,a115556a,a115559a,a115562a,a115563a,a115564a,a115568a,a115569a,a115572a,a115575a,a115576a,a115577a,a115580a,a115583a,a115584a,a115587a,a115590a,a115591a,a115592a,a115596a,a115597a,a115600a,a115603a,a115604a,a115605a,a115608a,a115611a,a115612a,a115615a,a115618a,a115619a,a115620a,a115624a,a115625a,a115628a,a115631a,a115632a,a115633a,a115636a,a115639a,a115640a,a115643a,a115646a,a115647a,a115648a,a115652a,a115653a,a115656a,a115659a,a115660a,a115661a,a115664a,a115667a,a115668a,a115671a,a115674a,a115675a,a115676a,a115680a,a115681a,a115684a,a115687a,a115688a,a115689a,a115692a,a115695a,a115696a,a115699a,a115702a,a115703a,a115704a,a115708a,a115709a,a115712a,a115715a,a115716a,a115717a,a115720a,a115723a,a115724a,a115727a,a115730a,a115731a,a115732a,a115736a,a115737a,a115740a,a115743a,a115744a,a115745a,a115748a,a115751a,a115752a,a115755a,a115758a,a115759a,a115760a,a115764a,a115765a,a115768a,a115771a,a115772a,a115773a,a115776a,a115779a,a115780a,a115783a,a115786a,a115787a,a115788a,a115792a,a115793a,a115796a,a115799a,a115800a,a115801a,a115804a,a115807a,a115808a,a115811a,a115814a,a115815a,a115816a,a115820a,a115821a,a115824a,a115827a,a115828a,a115829a,a115832a,a115835a,a115836a,a115839a,a115842a,a115843a,a115844a,a115848a,a115849a,a115852a,a115855a,a115856a,a115857a,a115860a,a115863a,a115864a,a115867a,a115870a,a115871a,a115872a,a115876a,a115877a,a115880a,a115883a,a115884a,a115885a,a115888a,a115891a,a115892a,a115895a,a115898a,a115899a,a115900a,a115904a,a115905a,a115908a,a115911a,a115912a,a115913a,a115916a,a115919a,a115920a,a115923a,a115926a,a115927a,a115928a,a115932a,a115933a,a115936a,a115939a,a115940a,a115941a,a115944a,a115947a,a115948a,a115951a,a115954a,a115955a,a115956a,a115960a,a115961a,a115964a,a115967a,a115968a,a115969a,a115972a,a115975a,a115976a,a115979a,a115982a,a115983a,a115984a,a115988a,a115989a,a115992a,a115995a,a115996a,a115997a,a116000a,a116003a,a116004a,a116007a,a116010a,a116011a,a116012a,a116016a,a116017a,a116020a,a116023a,a116024a,a116025a,a116028a,a116031a,a116032a,a116035a,a116038a,a116039a,a116040a,a116044a,a116045a,a116048a,a116051a,a116052a,a116053a,a116056a,a116059a,a116060a,a116063a,a116066a,a116067a,a116068a,a116072a,a116073a,a116076a,a116079a,a116080a,a116081a,a116084a,a116087a,a116088a,a116091a,a116094a,a116095a,a116096a,a116100a,a116101a,a116104a,a116107a,a116108a,a116109a,a116112a,a116115a,a116116a,a116119a,a116122a,a116123a,a116124a,a116128a,a116129a,a116132a,a116135a,a116136a,a116137a,a116140a,a116143a,a116144a,a116147a,a116150a,a116151a,a116152a,a116156a,a116157a,a116160a,a116163a,a116164a,a116165a,a116168a,a116171a,a116172a,a116175a,a116178a,a116179a,a116180a,a116184a,a116185a,a116188a,a116191a,a116192a,a116193a,a116196a,a116199a,a116200a,a116203a,a116206a,a116207a,a116208a,a116212a,a116213a,a116216a,a116219a,a116220a,a116221a,a116224a,a116227a,a116228a,a116231a,a116234a,a116235a,a116236a,a116240a,a116241a,a116244a,a116247a,a116248a,a116249a,a116252a,a116255a,a116256a,a116259a,a116262a,a116263a,a116264a,a116268a,a116269a,a116272a,a116275a,a116276a,a116277a,a116280a,a116283a,a116284a,a116287a,a116290a,a116291a,a116292a,a116296a,a116297a,a116300a,a116303a,a116304a,a116305a,a116308a,a116311a,a116312a,a116315a,a116318a,a116319a,a116320a,a116324a,a116325a,a116328a,a116331a,a116332a,a116333a,a116336a,a116339a,a116340a,a116343a,a116346a,a116347a,a116348a,a116352a,a116353a,a116356a,a116359a,a116360a,a116361a,a116364a,a116367a,a116368a,a116371a,a116374a,a116375a,a116376a,a116380a,a116381a,a116384a,a116387a,a116388a,a116389a,a116392a,a116395a,a116396a,a116399a,a116402a,a116403a,a116404a,a116408a,a116409a,a116412a,a116415a,a116416a,a116417a,a116420a,a116423a,a116424a,a116427a,a116430a,a116431a,a116432a,a116436a,a116437a,a116440a,a116443a,a116444a,a116445a,a116448a,a116451a,a116452a,a116455a,a116458a,a116459a,a116460a,a116464a,a116465a,a116468a,a116471a,a116472a,a116473a,a116476a,a116479a,a116480a,a116483a,a116486a,a116487a,a116488a,a116492a,a116493a,a116496a,a116499a,a116500a,a116501a,a116504a,a116507a,a116508a,a116511a,a116514a,a116515a,a116516a,a116520a,a116521a,a116524a,a116527a,a116528a,a116529a,a116532a,a116535a,a116536a,a116539a,a116542a,a116543a,a116544a,a116548a,a116549a,a116552a,a116555a,a116556a,a116557a,a116560a,a116563a,a116564a,a116567a,a116570a,a116571a,a116572a,a116576a,a116577a,a116580a,a116583a,a116584a,a116585a,a116588a,a116591a,a116592a,a116595a,a116598a,a116599a,a116600a,a116604a,a116605a,a116608a,a116611a,a116612a,a116613a,a116616a,a116619a,a116620a,a116623a,a116626a,a116627a,a116628a,a116632a,a116633a,a116636a,a116639a,a116640a,a116641a,a116644a,a116647a,a116648a,a116651a,a116654a,a116655a,a116656a,a116660a,a116661a,a116664a,a116667a,a116668a,a116669a,a116672a,a116675a,a116676a,a116679a,a116682a,a116683a,a116684a,a116688a,a116689a,a116692a,a116695a,a116696a,a116697a,a116700a,a116703a,a116704a,a116707a,a116710a,a116711a,a116712a,a116716a,a116717a,a116720a,a116723a,a116724a,a116725a,a116728a,a116731a,a116732a,a116735a,a116738a,a116739a,a116740a,a116744a,a116745a,a116748a,a116751a,a116752a,a116753a,a116756a,a116759a,a116760a,a116763a,a116766a,a116767a,a116768a,a116772a,a116773a,a116776a,a116779a,a116780a,a116781a,a116784a,a116787a,a116788a,a116791a,a116794a,a116795a,a116796a,a116800a,a116801a,a116804a,a116807a,a116808a,a116809a,a116812a,a116815a,a116816a,a116819a,a116822a,a116823a,a116824a,a116828a,a116829a,a116832a,a116835a,a116836a,a116837a,a116840a,a116843a,a116844a,a116847a,a116850a,a116851a,a116852a,a116855a,a116858a,a116859a,a116862a,a116865a,a116866a,a116867a,a116870a,a116873a,a116874a,a116877a,a116880a,a116881a,a116882a,a116885a,a116888a,a116889a,a116892a,a116895a,a116896a,a116897a,a116900a,a116903a,a116904a,a116907a,a116910a,a116911a,a116912a,a116915a,a116918a,a116919a,a116922a,a116925a,a116926a,a116927a,a116930a,a116933a,a116934a,a116937a,a116940a,a116941a,a116942a,a116945a,a116948a,a116949a,a116952a,a116955a,a116956a,a116957a,a116960a,a116963a,a116964a,a116967a,a116970a,a116971a,a116972a,a116975a,a116978a,a116979a,a116982a,a116985a,a116986a,a116987a,a116990a,a116993a,a116994a,a116997a,a117000a,a117001a,a117002a,a117005a,a117008a,a117009a,a117012a,a117015a,a117016a,a117017a,a117020a,a117023a,a117024a,a117027a,a117030a,a117031a,a117032a,a117035a,a117038a,a117039a,a117042a,a117045a,a117046a,a117047a,a117050a,a117053a,a117054a,a117057a,a117060a,a117061a,a117062a,a117065a,a117068a,a117069a,a117072a,a117075a,a117076a,a117077a,a117080a,a117083a,a117084a,a117087a,a117090a,a117091a,a117092a,a117095a,a117098a,a117099a,a117102a,a117105a,a117106a,a117107a,a117110a,a117113a,a117114a,a117117a,a117120a,a117121a,a117122a,a117125a,a117128a,a117129a,a117132a,a117135a,a117136a,a117137a,a117140a,a117143a,a117144a,a117147a,a117150a,a117151a,a117152a,a117155a,a117158a,a117159a,a117162a,a117165a,a117166a,a117167a,a117170a,a117173a,a117174a,a117177a,a117180a,a117181a,a117182a,a117185a,a117188a,a117189a,a117192a,a117195a,a117196a,a117197a,a117200a,a117203a,a117204a,a117207a,a117210a,a117211a,a117212a,a117215a,a117218a,a117219a,a117222a,a117225a,a117226a,a117227a,a117230a,a117233a,a117234a,a117237a,a117240a,a117241a,a117242a,a117245a,a117248a,a117249a,a117252a,a117255a,a117256a,a117257a,a117260a,a117263a,a117264a,a117267a,a117270a,a117271a,a117272a,a117275a,a117278a,a117279a,a117282a,a117285a,a117286a,a117287a,a117290a,a117293a,a117294a,a117297a,a117300a,a117301a,a117302a,a117305a,a117308a,a117309a,a117312a,a117315a,a117316a,a117317a,a117320a,a117323a,a117324a,a117327a,a117330a,a117331a,a117332a,a117335a,a117338a,a117339a,a117342a,a117345a,a117346a,a117347a,a117350a,a117353a,a117354a,a117357a,a117360a,a117361a,a117362a,a117365a,a117368a,a117369a,a117372a,a117375a,a117376a,a117377a,a117380a,a117383a,a117384a,a117387a,a117390a,a117391a,a117392a,a117395a,a117398a,a117399a,a117402a,a117405a,a117406a,a117407a,a117410a,a117413a,a117414a,a117417a,a117420a,a117421a,a117422a,a117425a,a117428a,a117429a,a117432a,a117435a,a117436a,a117437a,a117440a,a117443a,a117444a,a117447a,a117450a,a117451a,a117452a,a117455a,a117458a,a117459a,a117462a,a117465a,a117466a,a117467a,a117470a,a117473a,a117474a,a117477a,a117480a,a117481a,a117482a,a117485a,a117488a,a117489a,a117492a,a117495a,a117496a,a117497a,a117500a,a117503a,a117504a,a117507a,a117510a,a117511a,a117512a,a117515a,a117518a,a117519a,a117522a,a117525a,a117526a,a117527a,a117530a,a117533a,a117534a,a117537a,a117540a,a117541a,a117542a,a117545a,a117548a,a117549a,a117552a,a117555a,a117556a,a117557a,a117560a,a117563a,a117564a,a117567a,a117570a,a117571a,a117572a,a117575a,a117578a,a117579a,a117582a,a117585a,a117586a,a117587a,a117590a,a117593a,a117594a,a117597a,a117600a,a117601a,a117602a,a117605a,a117608a,a117609a,a117612a,a117615a,a117616a,a117617a,a117620a,a117623a,a117624a,a117627a,a117630a,a117631a,a117632a,a117635a,a117638a,a117639a,a117642a,a117645a,a117646a,a117647a,a117650a,a117653a,a117654a,a117657a,a117660a,a117661a,a117662a,a117665a,a117668a,a117669a,a117672a,a117675a,a117676a,a117677a,a117680a,a117683a,a117684a,a117687a,a117690a,a117691a,a117692a,a117695a,a117698a,a117699a,a117702a,a117705a,a117706a,a117707a,a117710a,a117713a,a117714a,a117717a,a117720a,a117721a,a117722a,a117725a,a117728a,a117729a,a117732a,a117735a,a117736a,a117737a,a117740a,a117743a,a117744a,a117747a,a117750a,a117751a,a117752a,a117755a,a117758a,a117759a,a117762a,a117765a,a117766a,a117767a,a117770a,a117773a,a117774a,a117777a,a117780a,a117781a,a117782a,a117785a,a117788a,a117789a,a117792a,a117795a,a117796a,a117797a,a117800a,a117803a,a117804a,a117807a,a117810a,a117811a,a117812a,a117815a,a117818a,a117819a,a117822a,a117825a,a117826a,a117827a,a117830a,a117833a,a117834a,a117837a,a117840a,a117841a,a117842a,a117845a,a117848a,a117849a,a117852a,a117855a,a117856a,a117857a,a117860a,a117863a,a117864a,a117867a,a117870a,a117871a,a117872a,a117875a,a117878a,a117879a,a117882a,a117885a,a117886a,a117887a,a117890a,a117893a,a117894a,a117897a,a117900a,a117901a,a117902a,a117905a,a117908a,a117909a,a117912a,a117915a,a117916a,a117917a,a117920a,a117923a,a117924a,a117927a,a117930a,a117931a,a117932a,a117935a,a117938a,a117939a,a117942a,a117945a,a117946a,a117947a,a117950a,a117953a,a117954a,a117957a,a117960a,a117961a,a117962a,a117965a,a117968a,a117969a,a117972a,a117975a,a117976a,a117977a,a117980a,a117983a,a117984a,a117987a,a117990a,a117991a,a117992a,a117995a,a117998a,a117999a,a118002a,a118005a,a118006a,a118007a,a118010a,a118013a,a118014a,a118017a,a118020a,a118021a,a118022a,a118025a,a118028a,a118029a,a118032a,a118035a,a118036a,a118037a,a118040a,a118043a,a118044a,a118047a,a118050a,a118051a,a118052a,a118055a,a118058a,a118059a,a118062a,a118065a,a118066a,a118067a,a118070a,a118073a,a118074a,a118077a,a118080a,a118081a,a118082a,a118085a,a118088a,a118089a,a118092a,a118095a,a118096a,a118097a,a118100a,a118103a,a118104a,a118107a,a118110a,a118111a,a118112a,a118115a,a118118a,a118119a,a118122a,a118125a,a118126a,a118127a,a118130a,a118133a,a118134a,a118137a,a118140a,a118141a,a118142a,a118145a,a118148a,a118149a,a118152a,a118155a,a118156a,a118157a,a118160a,a118163a,a118164a,a118167a,a118170a,a118171a,a118172a,a118175a,a118178a,a118179a,a118182a,a118185a,a118186a,a118187a,a118190a,a118193a,a118194a,a118197a,a118200a,a118201a,a118202a,a118205a,a118208a,a118209a,a118212a,a118215a,a118216a,a118217a,a118220a,a118223a,a118224a,a118227a,a118230a,a118231a,a118232a,a118235a,a118238a,a118239a,a118242a,a118245a,a118246a,a118247a,a118250a,a118253a,a118254a,a118257a,a118260a,a118261a,a118262a,a118265a,a118268a,a118269a,a118272a,a118275a,a118276a,a118277a,a118280a,a118283a,a118284a,a118287a,a118290a,a118291a,a118292a,a118295a,a118298a,a118299a,a118302a,a118305a,a118306a,a118307a,a118310a,a118313a,a118314a,a118317a,a118320a,a118321a,a118322a,a118325a,a118328a,a118329a,a118332a,a118335a,a118336a,a118337a,a118340a,a118343a,a118344a,a118347a,a118350a,a118351a,a118352a,a118355a,a118358a,a118359a,a118362a,a118365a,a118366a,a118367a,a118370a,a118373a,a118374a,a118377a,a118380a,a118381a,a118382a,a118385a,a118388a,a118389a,a118392a,a118395a,a118396a,a118397a,a118400a,a118403a,a118404a,a118407a,a118410a,a118411a,a118412a,a118415a,a118418a,a118419a,a118422a,a118425a,a118426a,a118427a,a118430a,a118433a,a118434a,a118437a,a118440a,a118441a,a118442a,a118445a,a118448a,a118449a,a118452a,a118455a,a118456a,a118457a,a118460a,a118463a,a118464a,a118467a,a118470a,a118471a,a118472a,a118475a,a118478a,a118479a,a118482a,a118485a,a118486a,a118487a,a118490a,a118493a,a118494a,a118497a,a118500a,a118501a,a118502a,a118505a,a118508a,a118509a,a118512a,a118515a,a118516a,a118517a,a118520a,a118523a,a118524a,a118527a,a118530a,a118531a,a118532a,a118535a,a118538a,a118539a,a118542a,a118545a,a118546a,a118547a,a118550a,a118553a,a118554a,a118557a,a118560a,a118561a,a118562a,a118565a,a118568a,a118569a,a118572a,a118575a,a118576a,a118577a,a118580a,a118583a,a118584a,a118587a,a118590a,a118591a,a118592a,a118595a,a118598a,a118599a,a118602a,a118605a,a118606a,a118607a,a118610a,a118613a,a118614a,a118617a,a118620a,a118621a,a118622a,a118625a,a118628a,a118629a,a118632a,a118635a,a118636a,a118637a,a118640a,a118643a,a118644a,a118647a,a118650a,a118651a,a118652a,a118655a,a118658a,a118659a,a118662a,a118665a,a118666a,a118667a,a118670a,a118673a,a118674a,a118677a,a118680a,a118681a,a118682a,a118685a,a118688a,a118689a,a118692a,a118695a,a118696a,a118697a,a118700a,a118703a,a118704a,a118707a,a118710a,a118711a,a118712a,a118715a,a118718a,a118719a,a118722a,a118725a,a118726a,a118727a,a118730a,a118733a,a118734a,a118737a,a118740a,a118741a,a118742a,a118745a,a118748a,a118749a,a118752a,a118755a,a118756a,a118757a,a118760a,a118763a,a118764a,a118767a,a118770a,a118771a,a118772a,a118775a,a118778a,a118779a,a118782a,a118785a,a118786a,a118787a,a118790a,a118793a,a118794a,a118797a,a118800a,a118801a,a118802a,a118805a,a118808a,a118809a,a118812a,a118815a,a118816a,a118817a,a118820a,a118823a,a118824a,a118827a,a118830a,a118831a,a118832a,a118835a,a118838a,a118839a,a118842a,a118845a,a118846a,a118847a,a118850a,a118853a,a118854a,a118857a,a118860a,a118861a,a118862a,a118865a,a118868a,a118869a,a118872a,a118875a,a118876a,a118877a,a118880a,a118883a,a118884a,a118887a,a118890a,a118891a,a118892a,a118895a,a118898a,a118899a,a118902a,a118905a,a118906a,a118907a,a118910a,a118913a,a118914a,a118917a,a118920a,a118921a,a118922a,a118925a,a118928a,a118929a,a118932a,a118935a,a118936a,a118937a,a118940a,a118943a,a118944a,a118947a,a118950a,a118951a,a118952a,a118955a,a118958a,a118959a,a118962a,a118965a,a118966a,a118967a,a118970a,a118973a,a118974a,a118977a,a118980a,a118981a,a118982a,a118985a,a118988a,a118989a,a118992a,a118995a,a118996a,a118997a,a119000a,a119003a,a119004a,a119007a,a119010a,a119011a,a119012a,a119015a,a119018a,a119019a,a119022a,a119025a,a119026a,a119027a,a119030a,a119033a,a119034a,a119037a,a119040a,a119041a,a119042a,a119045a,a119048a,a119049a,a119052a,a119055a,a119056a,a119057a,a119060a,a119063a,a119064a,a119067a,a119070a,a119071a,a119072a,a119075a,a119078a,a119079a,a119082a,a119085a,a119086a,a119087a,a119090a,a119093a,a119094a,a119097a,a119100a,a119101a,a119102a,a119105a,a119108a,a119109a,a119112a,a119115a,a119116a,a119117a,a119120a,a119123a,a119124a,a119127a,a119130a,a119131a,a119132a,a119135a,a119138a,a119139a,a119142a,a119145a,a119146a,a119147a,a119150a,a119153a,a119154a,a119157a,a119160a,a119161a,a119162a,a119165a,a119168a,a119169a,a119172a,a119175a,a119176a,a119177a,a119180a,a119183a,a119184a,a119187a,a119190a,a119191a,a119192a,a119195a,a119198a,a119199a,a119202a,a119205a,a119206a,a119207a,a119210a,a119213a,a119214a,a119217a,a119220a,a119221a,a119222a,a119225a,a119228a,a119229a,a119232a,a119235a,a119236a,a119237a,a119240a,a119243a,a119244a,a119247a,a119250a,a119251a,a119252a,a119255a,a119258a,a119259a,a119262a,a119265a,a119266a,a119267a,a119270a,a119273a,a119274a,a119277a,a119280a,a119281a,a119282a,a119285a,a119288a,a119289a,a119292a,a119295a,a119296a,a119297a,a119300a,a119303a,a119304a,a119307a,a119310a,a119311a,a119312a,a119315a,a119318a,a119319a,a119322a,a119325a,a119326a,a119327a,a119330a,a119333a,a119334a,a119337a,a119340a,a119341a,a119342a,a119345a,a119348a,a119349a,a119352a,a119355a,a119356a,a119357a,a119360a,a119363a,a119364a,a119367a,a119370a,a119371a,a119372a,a119375a,a119378a,a119379a,a119382a,a119385a,a119386a,a119387a,a119390a,a119393a,a119394a,a119397a,a119400a,a119401a,a119402a,a119405a,a119408a,a119409a,a119412a,a119415a,a119416a,a119417a,a119420a,a119423a,a119424a,a119427a,a119430a,a119431a,a119432a,a119435a,a119438a,a119439a,a119442a,a119445a,a119446a,a119447a,a119450a,a119453a,a119454a,a119457a,a119460a,a119461a,a119462a,a119465a,a119468a,a119469a,a119472a,a119475a,a119476a,a119477a,a119480a,a119483a,a119484a,a119487a,a119490a,a119491a,a119492a,a119495a,a119498a,a119499a,a119502a,a119505a,a119506a,a119507a,a119510a,a119513a,a119514a,a119517a,a119520a,a119521a,a119522a,a119525a,a119528a,a119529a,a119532a,a119535a,a119536a,a119537a,a119540a,a119543a,a119544a,a119547a,a119550a,a119551a,a119552a,a119555a,a119558a,a119559a,a119562a,a119565a,a119566a,a119567a,a119570a,a119573a,a119574a,a119577a,a119580a,a119581a,a119582a,a119585a,a119588a,a119589a,a119592a,a119595a,a119596a,a119597a,a119600a,a119603a,a119604a,a119607a,a119610a,a119611a,a119612a,a119615a,a119618a,a119619a,a119622a,a119625a,a119626a,a119627a,a119630a,a119633a,a119634a,a119637a,a119640a,a119641a,a119642a,a119645a,a119648a,a119649a,a119652a,a119655a,a119656a,a119657a,a119660a,a119663a,a119664a,a119667a,a119670a,a119671a,a119672a,a119675a,a119678a,a119679a,a119682a,a119685a,a119686a,a119687a,a119690a,a119693a,a119694a,a119697a,a119700a,a119701a,a119702a,a119705a,a119708a,a119709a,a119712a,a119715a,a119716a,a119717a,a119720a,a119723a,a119724a,a119727a,a119730a,a119731a,a119732a,a119735a,a119738a,a119739a,a119742a,a119745a,a119746a,a119747a,a119750a,a119753a,a119754a,a119757a,a119760a,a119761a,a119762a,a119765a,a119768a,a119769a,a119772a,a119775a,a119776a,a119777a,a119780a,a119783a,a119784a,a119787a,a119790a,a119791a,a119792a,a119795a,a119798a,a119799a,a119802a,a119805a,a119806a,a119807a,a119810a,a119813a,a119814a,a119817a,a119820a,a119821a,a119822a,a119825a,a119828a,a119829a,a119832a,a119835a,a119836a,a119837a,a119840a,a119843a,a119844a,a119847a,a119850a,a119851a,a119852a,a119855a,a119858a,a119859a,a119862a,a119865a,a119866a,a119867a,a119870a,a119873a,a119874a,a119877a,a119880a,a119881a,a119882a,a119885a,a119888a,a119889a,a119892a,a119895a,a119896a,a119897a,a119900a,a119903a,a119904a,a119907a,a119910a,a119911a,a119912a,a119915a,a119918a,a119919a,a119922a,a119925a,a119926a,a119927a,a119930a,a119933a,a119934a,a119937a,a119940a,a119941a,a119942a,a119945a,a119948a,a119949a,a119952a,a119955a,a119956a,a119957a,a119960a,a119963a,a119964a,a119967a,a119970a,a119971a,a119972a,a119975a,a119978a,a119979a,a119982a,a119985a,a119986a,a119987a,a119990a,a119993a,a119994a,a119997a,a120000a,a120001a,a120002a,a120005a,a120008a,a120009a,a120012a,a120015a,a120016a,a120017a,a120020a,a120023a,a120024a,a120027a,a120030a,a120031a,a120032a,a120035a,a120038a,a120039a,a120042a,a120045a,a120046a,a120047a,a120050a,a120053a,a120054a,a120057a,a120060a,a120061a,a120062a,a120065a,a120068a,a120069a,a120072a,a120075a,a120076a,a120077a,a120080a,a120083a,a120084a,a120087a,a120090a,a120091a,a120092a,a120095a,a120098a,a120099a,a120102a,a120105a,a120106a,a120107a,a120110a,a120113a,a120114a,a120117a,a120120a,a120121a,a120122a,a120125a,a120128a,a120129a,a120132a,a120135a,a120136a,a120137a,a120140a,a120143a,a120144a,a120147a,a120150a,a120151a,a120152a,a120155a,a120158a,a120159a,a120162a,a120165a,a120166a,a120167a,a120170a,a120173a,a120174a,a120177a,a120180a,a120181a,a120182a,a120185a,a120188a,a120189a,a120192a,a120195a,a120196a,a120197a,a120200a,a120203a,a120204a,a120207a,a120210a,a120211a,a120212a,a120215a,a120218a,a120219a,a120222a,a120225a,a120226a,a120227a,a120230a,a120233a,a120234a,a120237a,a120240a,a120241a,a120242a,a120245a,a120248a,a120249a,a120252a,a120255a,a120256a,a120257a,a120260a,a120263a,a120264a,a120267a,a120270a,a120271a,a120272a,a120275a,a120278a,a120279a,a120282a,a120285a,a120286a,a120287a,a120290a,a120293a,a120294a,a120297a,a120300a,a120301a,a120302a,a120305a,a120308a,a120309a,a120312a,a120315a,a120316a,a120317a,a120320a,a120323a,a120324a,a120327a,a120330a,a120331a,a120332a,a120335a,a120338a,a120339a,a120342a,a120345a,a120346a,a120347a,a120350a,a120353a,a120354a,a120357a,a120360a,a120361a,a120362a,a120365a,a120368a,a120369a,a120372a,a120375a,a120376a,a120377a,a120380a,a120383a,a120384a,a120387a,a120390a,a120391a,a120392a,a120395a,a120398a,a120399a,a120402a,a120405a,a120406a,a120407a,a120410a,a120413a,a120414a,a120417a,a120420a,a120421a,a120422a,a120425a,a120428a,a120429a,a120432a,a120435a,a120436a,a120437a,a120440a,a120443a,a120444a,a120447a,a120450a,a120451a,a120452a,a120455a,a120458a,a120459a,a120462a,a120465a,a120466a,a120467a,a120470a,a120473a,a120474a,a120477a,a120480a,a120481a,a120482a,a120485a,a120488a,a120489a,a120492a,a120495a,a120496a,a120497a,a120500a,a120503a,a120504a,a120507a,a120510a,a120511a,a120512a,a120515a,a120518a,a120519a,a120522a,a120525a,a120526a,a120527a,a120530a,a120533a,a120534a,a120537a,a120540a,a120541a,a120542a,a120545a,a120548a,a120549a,a120552a,a120555a,a120556a,a120557a,a120560a,a120563a,a120564a,a120567a,a120570a,a120571a,a120572a,a120575a,a120578a,a120579a,a120582a,a120585a,a120586a,a120587a,a120590a,a120593a,a120594a,a120597a,a120600a,a120601a,a120602a,a120605a,a120608a,a120609a,a120612a,a120615a,a120616a,a120617a,a120620a,a120623a,a120624a,a120627a,a120630a,a120631a,a120632a,a120635a,a120638a,a120639a,a120642a,a120645a,a120646a,a120647a,a120650a,a120653a,a120654a,a120657a,a120660a,a120661a,a120662a,a120665a,a120668a,a120669a,a120672a,a120675a,a120676a,a120677a,a120680a,a120683a,a120684a,a120687a,a120690a,a120691a,a120692a,a120695a,a120698a,a120699a,a120702a,a120705a,a120706a,a120707a,a120710a,a120713a,a120714a,a120717a,a120720a,a120721a,a120722a,a120725a,a120728a,a120729a,a120732a,a120735a,a120736a,a120737a,a120740a,a120743a,a120744a,a120747a,a120750a,a120751a,a120752a,a120755a,a120758a,a120759a,a120762a,a120765a,a120766a,a120767a,a120770a,a120773a,a120774a,a120777a,a120780a,a120781a,a120782a,a120785a,a120788a,a120789a,a120792a,a120795a,a120796a,a120797a,a120800a,a120803a,a120804a,a120807a,a120810a,a120811a,a120812a,a120815a,a120818a,a120819a,a120822a,a120825a,a120826a,a120827a,a120830a,a120833a,a120834a,a120837a,a120840a,a120841a,a120842a,a120845a,a120848a,a120849a,a120852a,a120855a,a120856a,a120857a,a120860a,a120863a,a120864a,a120867a,a120870a,a120871a,a120872a,a120875a,a120878a,a120879a,a120882a,a120885a,a120886a,a120887a,a120890a,a120893a,a120894a,a120897a,a120900a,a120901a,a120902a,a120905a,a120908a,a120909a,a120912a,a120915a,a120916a,a120917a,a120920a,a120923a,a120924a,a120927a,a120930a,a120931a,a120932a,a120935a,a120938a,a120939a,a120942a,a120945a,a120946a,a120947a,a120950a,a120953a,a120954a,a120957a,a120960a,a120961a,a120962a,a120965a,a120968a,a120969a,a120972a,a120975a,a120976a,a120977a,a120980a,a120983a,a120984a,a120987a,a120990a,a120991a,a120992a,a120995a,a120998a,a120999a,a121002a,a121005a,a121006a,a121007a,a121010a,a121013a,a121014a,a121017a,a121020a,a121021a,a121022a,a121025a,a121028a,a121029a,a121032a,a121035a,a121036a,a121037a,a121040a,a121043a,a121044a,a121047a,a121050a,a121051a,a121052a,a121055a,a121058a,a121059a,a121062a,a121065a,a121066a,a121067a,a121070a,a121073a,a121074a,a121077a,a121080a,a121081a,a121082a,a121085a,a121088a,a121089a,a121092a,a121095a,a121096a,a121097a,a121100a,a121103a,a121104a,a121107a,a121110a,a121111a,a121112a,a121115a,a121118a,a121119a,a121122a,a121125a,a121126a,a121127a,a121130a,a121133a,a121134a,a121137a,a121140a,a121141a,a121142a,a121145a,a121148a,a121149a,a121152a,a121155a,a121156a,a121157a,a121160a,a121163a,a121164a,a121167a,a121170a,a121171a,a121172a,a121175a,a121178a,a121179a,a121182a,a121185a,a121186a,a121187a,a121190a,a121193a,a121194a,a121197a,a121200a,a121201a,a121202a,a121205a,a121208a,a121209a,a121212a,a121215a,a121216a,a121217a,a121220a,a121223a,a121224a,a121227a,a121230a,a121231a,a121232a,a121235a,a121238a,a121239a,a121242a,a121245a,a121246a,a121247a,a121250a,a121253a,a121254a,a121257a,a121260a,a121261a,a121262a,a121265a,a121268a,a121269a,a121272a,a121275a,a121276a,a121277a,a121280a,a121283a,a121284a,a121287a,a121290a,a121291a,a121292a,a121295a,a121298a,a121299a,a121302a,a121305a,a121306a,a121307a,a121310a,a121313a,a121314a,a121317a,a121320a,a121321a,a121322a,a121325a,a121328a,a121329a,a121332a,a121335a,a121336a,a121337a,a121340a,a121343a,a121344a,a121347a,a121350a,a121351a,a121352a,a121355a,a121358a,a121359a,a121362a,a121365a,a121366a,a121367a,a121370a,a121373a,a121374a,a121377a,a121380a,a121381a,a121382a,a121385a,a121388a,a121389a,a121392a,a121395a,a121396a,a121397a,a121400a,a121403a,a121404a,a121407a,a121410a,a121411a,a121412a,a121415a,a121418a,a121419a,a121422a,a121425a,a121426a,a121427a,a121430a,a121433a,a121434a,a121437a,a121440a,a121441a,a121442a,a121445a,a121448a,a121449a,a121452a,a121455a,a121456a,a121457a,a121460a,a121463a,a121464a,a121467a,a121470a,a121471a,a121472a,a121475a,a121478a,a121479a,a121482a,a121485a,a121486a,a121487a,a121490a,a121493a,a121494a,a121497a,a121500a,a121501a,a121502a,a121505a,a121508a,a121509a,a121512a,a121515a,a121516a,a121517a,a121520a,a121523a,a121524a,a121527a,a121530a,a121531a,a121532a,a121535a,a121538a,a121539a,a121542a,a121545a,a121546a,a121547a,a121550a,a121553a,a121554a,a121557a,a121560a,a121561a,a121562a,a121565a,a121568a,a121569a,a121572a,a121575a,a121576a,a121577a,a121580a,a121583a,a121584a,a121587a,a121590a,a121591a,a121592a,a121595a,a121598a,a121599a,a121602a,a121605a,a121606a,a121607a,a121610a,a121613a,a121614a,a121617a,a121620a,a121621a,a121622a,a121625a,a121628a,a121629a,a121632a,a121635a,a121636a,a121637a,a121640a,a121643a,a121644a,a121647a,a121650a,a121651a,a121652a,a121655a,a121658a,a121659a,a121662a,a121665a,a121666a,a121667a,a121670a,a121673a,a121674a,a121677a,a121680a,a121681a,a121682a,a121685a,a121688a,a121689a,a121692a,a121695a,a121696a,a121697a,a121700a,a121703a,a121704a,a121707a,a121710a,a121711a,a121712a,a121715a,a121718a,a121719a,a121722a,a121725a,a121726a,a121727a,a121730a,a121733a,a121734a,a121737a,a121740a,a121741a,a121742a,a121745a,a121748a,a121749a,a121752a,a121755a,a121756a,a121757a,a121760a,a121763a,a121764a,a121767a,a121770a,a121771a,a121772a,a121775a,a121778a,a121779a,a121782a,a121785a,a121786a,a121787a,a121790a,a121793a,a121794a,a121797a,a121800a,a121801a,a121802a,a121805a,a121808a,a121809a,a121812a,a121815a,a121816a,a121817a,a121820a,a121823a,a121824a,a121827a,a121830a,a121831a,a121832a,a121835a,a121838a,a121839a,a121842a,a121845a,a121846a,a121847a,a121850a,a121853a,a121854a,a121857a,a121860a,a121861a,a121862a,a121865a,a121868a,a121869a,a121872a,a121875a,a121876a,a121877a,a121880a,a121883a,a121884a,a121887a,a121890a,a121891a,a121892a,a121895a,a121898a,a121899a,a121902a,a121905a,a121906a,a121907a,a121910a,a121913a,a121914a,a121917a,a121920a,a121921a,a121922a,a121925a,a121928a,a121929a,a121932a,a121935a,a121936a,a121937a,a121940a,a121943a,a121944a,a121947a,a121950a,a121951a,a121952a,a121955a,a121958a,a121959a,a121962a,a121965a,a121966a,a121967a,a121970a,a121973a,a121974a,a121977a,a121980a,a121981a,a121982a,a121985a,a121988a,a121989a,a121992a,a121995a,a121996a,a121997a,a122000a,a122003a,a122004a,a122007a,a122010a,a122011a,a122012a,a122015a,a122018a,a122019a,a122022a,a122025a,a122026a,a122027a,a122030a,a122033a,a122034a,a122037a,a122040a,a122041a,a122042a,a122045a,a122048a,a122049a,a122052a,a122055a,a122056a,a122057a,a122060a,a122063a,a122064a,a122067a,a122070a,a122071a,a122072a,a122075a,a122078a,a122079a,a122082a,a122085a,a122086a,a122087a,a122090a,a122093a,a122094a,a122097a,a122100a,a122101a,a122102a,a122105a,a122108a,a122109a,a122112a,a122115a,a122116a,a122117a,a122120a,a122123a,a122124a,a122127a,a122130a,a122131a,a122132a,a122135a,a122138a,a122139a,a122142a,a122145a,a122146a,a122147a,a122150a,a122153a,a122154a,a122157a,a122160a,a122161a,a122162a,a122165a,a122168a,a122169a,a122172a,a122175a,a122176a,a122177a,a122180a,a122183a,a122184a,a122187a,a122190a,a122191a,a122192a,a122195a,a122198a,a122199a,a122202a,a122205a,a122206a,a122207a,a122210a,a122213a,a122214a,a122217a,a122220a,a122221a,a122222a,a122225a,a122228a,a122229a,a122232a,a122235a,a122236a,a122237a,a122240a,a122243a,a122244a,a122247a,a122250a,a122251a,a122252a,a122255a,a122258a,a122259a,a122262a,a122265a,a122266a,a122267a,a122270a,a122273a,a122274a,a122277a,a122280a,a122281a,a122282a,a122285a,a122288a,a122289a,a122292a,a122295a,a122296a,a122297a,a122300a,a122303a,a122304a,a122307a,a122310a,a122311a,a122312a,a122315a,a122318a,a122319a,a122322a,a122325a,a122326a,a122327a,a122330a,a122333a,a122334a,a122337a,a122340a,a122341a,a122342a,a122345a,a122348a,a122349a,a122352a,a122355a,a122356a,a122357a,a122360a,a122363a,a122364a,a122367a,a122370a,a122371a,a122372a,a122375a,a122378a,a122379a,a122382a,a122385a,a122386a,a122387a,a122390a,a122393a,a122394a,a122397a,a122400a,a122401a,a122402a,a122405a,a122408a,a122409a,a122412a,a122415a,a122416a,a122417a,a122420a,a122423a,a122424a,a122427a,a122430a,a122431a,a122432a,a122435a,a122438a,a122439a,a122442a,a122445a,a122446a,a122447a,a122450a,a122453a,a122454a,a122457a,a122460a,a122461a,a122462a,a122465a,a122468a,a122469a,a122472a,a122475a,a122476a,a122477a,a122480a,a122483a,a122484a,a122487a,a122490a,a122491a,a122492a,a122495a,a122498a,a122499a,a122502a,a122505a,a122506a,a122507a,a122510a,a122513a,a122514a,a122517a,a122520a,a122521a,a122522a,a122525a,a122528a,a122529a,a122532a,a122535a,a122536a,a122537a,a122540a,a122543a,a122544a,a122547a,a122550a,a122551a,a122552a,a122555a,a122558a,a122559a,a122562a,a122565a,a122566a,a122567a,a122570a,a122573a,a122574a,a122577a,a122580a,a122581a,a122582a,a122585a,a122588a,a122589a,a122592a,a122595a,a122596a,a122597a,a122600a,a122603a,a122604a,a122607a,a122610a,a122611a,a122612a,a122615a,a122618a,a122619a,a122622a,a122625a,a122626a,a122627a,a122630a,a122633a,a122634a,a122637a,a122640a,a122641a,a122642a,a122645a,a122648a,a122649a,a122652a,a122655a,a122656a,a122657a,a122660a,a122663a,a122664a,a122667a,a122670a,a122671a,a122672a,a122675a,a122678a,a122679a,a122682a,a122685a,a122686a,a122687a,a122690a,a122693a,a122694a,a122697a,a122700a,a122701a,a122702a,a122705a,a122708a,a122709a,a122712a,a122715a,a122716a,a122717a,a122720a,a122723a,a122724a,a122727a,a122730a,a122731a,a122732a,a122735a,a122738a,a122739a,a122742a,a122745a,a122746a,a122747a,a122750a,a122753a,a122754a,a122757a,a122760a,a122761a,a122762a,a122765a,a122768a,a122769a,a122772a,a122775a,a122776a,a122777a,a122780a,a122783a,a122784a,a122787a,a122790a,a122791a,a122792a,a122795a,a122798a,a122799a,a122802a,a122805a,a122806a,a122807a,a122810a,a122813a,a122814a,a122817a,a122820a,a122821a,a122822a,a122825a,a122828a,a122829a,a122832a,a122835a,a122836a,a122837a,a122840a,a122843a,a122844a,a122847a,a122850a,a122851a,a122852a,a122855a,a122858a,a122859a,a122862a,a122865a,a122866a,a122867a,a122870a,a122873a,a122874a,a122877a,a122880a,a122881a,a122882a,a122885a,a122888a,a122889a,a122892a,a122895a,a122896a,a122897a,a122900a,a122903a,a122904a,a122907a,a122910a,a122911a,a122912a,a122915a,a122918a,a122919a,a122922a,a122925a,a122926a,a122927a,a122930a,a122933a,a122934a,a122937a,a122940a,a122941a,a122942a,a122945a,a122948a,a122949a,a122952a,a122955a,a122956a,a122957a,a122960a,a122963a,a122964a,a122967a,a122970a,a122971a,a122972a,a122975a,a122978a,a122979a,a122982a,a122985a,a122986a,a122987a,a122990a,a122993a,a122994a,a122997a,a123000a,a123001a,a123002a,a123005a,a123008a,a123009a,a123012a,a123015a,a123016a,a123017a,a123020a,a123023a,a123024a,a123027a,a123030a,a123031a,a123032a,a123035a,a123038a,a123039a,a123042a,a123045a,a123046a,a123047a,a123050a,a123053a,a123054a,a123057a,a123060a,a123061a,a123062a,a123065a,a123068a,a123069a,a123072a,a123075a,a123076a,a123077a,a123080a,a123083a,a123084a,a123087a,a123090a,a123091a,a123092a,a123095a,a123098a,a123099a,a123102a,a123105a,a123106a,a123107a,a123110a,a123113a,a123114a,a123117a,a123120a,a123121a,a123122a,a123125a,a123128a,a123129a,a123132a,a123135a,a123136a,a123137a,a123140a,a123143a,a123144a,a123147a,a123150a,a123151a,a123152a,a123155a,a123158a,a123159a,a123162a,a123165a,a123166a,a123167a,a123170a,a123173a,a123174a,a123177a,a123180a,a123181a,a123182a,a123185a,a123188a,a123189a,a123192a,a123195a,a123196a,a123197a,a123200a,a123203a,a123204a,a123207a,a123210a,a123211a,a123212a,a123215a,a123218a,a123219a,a123222a,a123225a,a123226a,a123227a,a123230a,a123233a,a123234a,a123237a,a123240a,a123241a,a123242a,a123245a,a123248a,a123249a,a123252a,a123255a,a123256a,a123257a,a123260a,a123263a,a123264a,a123267a,a123270a,a123271a,a123272a,a123275a,a123278a,a123279a,a123282a,a123285a,a123286a,a123287a,a123290a,a123293a,a123294a,a123297a,a123300a,a123301a,a123302a,a123305a,a123308a,a123309a,a123312a,a123315a,a123316a,a123317a,a123320a,a123323a,a123324a,a123327a,a123330a,a123331a,a123332a,a123335a,a123338a,a123339a,a123342a,a123345a,a123346a,a123347a,a123350a,a123353a,a123354a,a123357a,a123360a,a123361a,a123362a,a123365a,a123368a,a123369a,a123372a,a123375a,a123376a,a123377a,a123380a,a123383a,a123384a,a123387a,a123390a,a123391a,a123392a,a123395a,a123398a,a123399a,a123402a,a123405a,a123406a,a123407a,a123410a,a123413a,a123414a,a123417a,a123420a,a123421a,a123422a,a123425a,a123428a,a123429a,a123432a,a123435a,a123436a,a123437a,a123440a,a123443a,a123444a,a123447a,a123450a,a123451a,a123452a,a123455a,a123458a,a123459a,a123462a,a123465a,a123466a,a123467a,a123470a,a123473a,a123474a,a123477a,a123480a,a123481a,a123482a,a123485a,a123488a,a123489a,a123492a,a123495a,a123496a,a123497a,a123500a,a123503a,a123504a,a123507a,a123510a,a123511a,a123512a,a123515a,a123518a,a123519a,a123522a,a123525a,a123526a,a123527a,a123530a,a123533a,a123534a,a123537a,a123540a,a123541a,a123542a,a123545a,a123548a,a123549a,a123552a,a123555a,a123556a,a123557a,a123560a,a123563a,a123564a,a123567a,a123570a,a123571a,a123572a,a123575a,a123578a,a123579a,a123582a,a123585a,a123586a,a123587a,a123590a,a123593a,a123594a,a123597a,a123600a,a123601a,a123602a,a123605a,a123608a,a123609a,a123612a,a123615a,a123616a,a123617a,a123620a,a123623a,a123624a,a123627a,a123630a,a123631a,a123632a,a123635a,a123638a,a123639a,a123642a,a123645a,a123646a,a123647a,a123650a,a123653a,a123654a,a123657a,a123660a,a123661a,a123662a,a123665a,a123668a,a123669a,a123672a,a123675a,a123676a,a123677a,a123680a,a123683a,a123684a,a123687a,a123690a,a123691a,a123692a,a123695a,a123698a,a123699a,a123702a,a123705a,a123706a,a123707a,a123710a,a123713a,a123714a,a123717a,a123720a,a123721a,a123722a,a123725a,a123728a,a123729a,a123732a,a123735a,a123736a,a123737a,a123740a,a123743a,a123744a,a123747a,a123750a,a123751a,a123752a,a123755a,a123758a,a123759a,a123762a,a123765a,a123766a,a123767a,a123770a,a123773a,a123774a,a123777a,a123780a,a123781a,a123782a,a123785a,a123788a,a123789a,a123792a,a123795a,a123796a,a123797a,a123800a,a123803a,a123804a,a123807a,a123810a,a123811a,a123812a,a123815a,a123818a,a123819a,a123822a,a123825a,a123826a,a123827a,a123830a,a123833a,a123834a,a123837a,a123840a,a123841a,a123842a,a123845a,a123848a,a123849a,a123852a,a123855a,a123856a,a123857a,a123860a,a123863a,a123864a,a123867a,a123870a,a123871a,a123872a,a123875a,a123878a,a123879a,a123882a,a123885a,a123886a,a123887a,a123890a,a123893a,a123894a,a123897a,a123900a,a123901a,a123902a,a123905a,a123908a,a123909a,a123912a,a123915a,a123916a,a123917a,a123920a,a123923a,a123924a,a123927a,a123930a,a123931a,a123932a,a123935a,a123938a,a123939a,a123942a,a123945a,a123946a,a123947a,a123950a,a123953a,a123954a,a123957a,a123960a,a123961a,a123962a,a123965a,a123968a,a123969a,a123972a,a123975a,a123976a,a123977a,a123980a,a123983a,a123984a,a123987a,a123990a,a123991a,a123992a,a123995a,a123998a,a123999a,a124002a,a124005a,a124006a,a124007a,a124010a,a124013a,a124014a,a124017a,a124020a,a124021a,a124022a,a124025a,a124028a,a124029a,a124032a,a124035a,a124036a,a124037a,a124040a,a124043a,a124044a,a124047a,a124050a,a124051a,a124052a,a124055a,a124058a,a124059a,a124062a,a124065a,a124066a,a124067a,a124070a,a124073a,a124074a,a124077a,a124080a,a124081a,a124082a,a124085a,a124088a,a124089a,a124092a,a124095a,a124096a,a124097a,a124100a,a124103a,a124104a,a124107a,a124110a,a124111a,a124112a,a124115a,a124118a,a124119a,a124122a,a124125a,a124126a,a124127a,a124130a,a124133a,a124134a,a124137a,a124140a,a124141a,a124142a,a124145a,a124148a,a124149a,a124152a,a124155a,a124156a,a124157a,a124160a,a124163a,a124164a,a124167a,a124170a,a124171a,a124172a,a124175a,a124178a,a124179a,a124182a,a124185a,a124186a,a124187a,a124190a,a124193a,a124194a,a124197a,a124200a,a124201a,a124202a,a124205a,a124208a,a124209a,a124212a,a124215a,a124216a,a124217a,a124220a,a124223a,a124224a,a124227a,a124230a,a124231a,a124232a,a124235a,a124238a,a124239a,a124242a,a124245a,a124246a,a124247a,a124250a,a124253a,a124254a,a124257a,a124260a,a124261a,a124262a,a124265a,a124268a,a124269a,a124272a,a124275a,a124276a,a124277a,a124280a,a124283a,a124284a,a124287a,a124290a,a124291a,a124292a,a124295a,a124298a,a124299a,a124302a,a124305a,a124306a,a124307a,a124310a,a124313a,a124314a,a124317a,a124320a,a124321a,a124322a,a124325a,a124328a,a124329a,a124332a,a124335a,a124336a,a124337a,a124340a,a124343a,a124344a,a124347a,a124350a,a124351a,a124352a,a124355a,a124358a,a124359a,a124362a,a124365a,a124366a,a124367a,a124370a,a124373a,a124374a,a124377a,a124380a,a124381a,a124382a,a124385a,a124388a,a124389a,a124392a,a124395a,a124396a,a124397a,a124400a,a124403a,a124404a,a124407a,a124410a,a124411a,a124412a,a124415a,a124418a,a124419a,a124422a,a124425a,a124426a,a124427a,a124430a,a124433a,a124434a,a124437a,a124440a,a124441a,a124442a,a124445a,a124448a,a124449a,a124452a,a124455a,a124456a,a124457a,a124460a,a124463a,a124464a,a124467a,a124470a,a124471a,a124472a,a124475a,a124478a,a124479a,a124482a,a124485a,a124486a,a124487a,a124490a,a124493a,a124494a,a124497a,a124500a,a124501a,a124502a,a124505a,a124508a,a124509a,a124512a,a124515a,a124516a,a124517a,a124520a,a124523a,a124524a,a124527a,a124530a,a124531a,a124532a,a124535a,a124538a,a124539a,a124542a,a124545a,a124546a,a124547a,a124550a,a124553a,a124554a,a124557a,a124560a,a124561a,a124562a,a124565a,a124568a,a124569a,a124572a,a124575a,a124576a,a124577a,a124580a,a124583a,a124584a,a124587a,a124590a,a124591a,a124592a,a124595a,a124598a,a124599a,a124602a,a124605a,a124606a,a124607a,a124610a,a124613a,a124614a,a124617a,a124620a,a124621a,a124622a,a124625a,a124628a,a124629a,a124632a,a124635a,a124636a,a124637a,a124640a,a124643a,a124644a,a124647a,a124650a,a124651a,a124652a,a124655a,a124658a,a124659a,a124662a,a124665a,a124666a,a124667a,a124670a,a124673a,a124674a,a124677a,a124680a,a124681a,a124682a,a124685a,a124688a,a124689a,a124692a,a124695a,a124696a,a124697a,a124700a,a124703a,a124704a,a124707a,a124710a,a124711a,a124712a,a124715a,a124718a,a124719a,a124722a,a124725a,a124726a,a124727a,a124730a,a124733a,a124734a,a124737a,a124740a,a124741a,a124742a,a124745a,a124748a,a124749a,a124752a,a124755a,a124756a,a124757a,a124760a,a124763a,a124764a,a124767a,a124770a,a124771a,a124772a,a124775a,a124778a,a124779a,a124782a,a124785a,a124786a,a124787a,a124790a,a124793a,a124794a,a124797a,a124800a,a124801a,a124802a,a124805a,a124808a,a124809a,a124812a,a124815a,a124816a,a124817a,a124820a,a124823a,a124824a,a124827a,a124830a,a124831a,a124832a,a124835a,a124838a,a124839a,a124842a,a124845a,a124846a,a124847a,a124850a,a124853a,a124854a,a124857a,a124860a,a124861a,a124862a,a124865a,a124868a,a124869a,a124872a,a124875a,a124876a,a124877a,a124880a,a124883a,a124884a,a124887a,a124890a,a124891a,a124892a,a124895a,a124898a,a124899a,a124902a,a124905a,a124906a,a124907a,a124910a,a124913a,a124914a,a124917a,a124920a,a124921a,a124922a,a124925a,a124928a,a124929a,a124932a,a124935a,a124936a,a124937a,a124940a,a124943a,a124944a,a124947a,a124950a,a124951a,a124952a,a124955a,a124958a,a124959a,a124962a,a124965a,a124966a,a124967a,a124970a,a124973a,a124974a,a124977a,a124980a,a124981a,a124982a,a124985a,a124988a,a124989a,a124992a,a124995a,a124996a,a124997a,a125000a,a125003a,a125004a,a125007a,a125010a,a125011a,a125012a,a125015a,a125018a,a125019a,a125022a,a125025a,a125026a,a125027a,a125030a,a125033a,a125034a,a125037a,a125040a,a125041a,a125042a,a125045a,a125048a,a125049a,a125052a,a125055a,a125056a,a125057a,a125060a,a125063a,a125064a,a125067a,a125070a,a125071a,a125072a,a125075a,a125078a,a125079a,a125082a,a125085a,a125086a,a125087a,a125090a,a125093a,a125094a,a125097a,a125100a,a125101a,a125102a,a125105a,a125108a,a125109a,a125112a,a125115a,a125116a,a125117a,a125120a,a125123a,a125124a,a125127a,a125130a,a125131a,a125132a,a125135a,a125138a,a125139a,a125142a,a125145a,a125146a,a125147a,a125150a,a125153a,a125154a,a125157a,a125160a,a125161a,a125162a,a125165a,a125168a,a125169a,a125172a,a125175a,a125176a,a125177a,a125180a,a125183a,a125184a,a125187a,a125190a,a125191a,a125192a,a125195a,a125198a,a125199a,a125202a,a125205a,a125206a,a125207a,a125210a,a125213a,a125214a,a125217a,a125220a,a125221a,a125222a,a125225a,a125228a,a125229a,a125232a,a125235a,a125236a,a125237a,a125240a,a125243a,a125244a,a125247a,a125250a,a125251a,a125252a,a125255a,a125258a,a125259a,a125262a,a125265a,a125266a,a125267a,a125270a,a125273a,a125274a,a125277a,a125280a,a125281a,a125282a,a125285a,a125288a,a125289a,a125292a,a125295a,a125296a,a125297a,a125300a,a125303a,a125304a,a125307a,a125310a,a125311a,a125312a,a125315a,a125318a,a125319a,a125322a,a125325a,a125326a,a125327a,a125330a,a125333a,a125334a,a125337a,a125340a,a125341a,a125342a,a125345a,a125348a,a125349a,a125352a,a125355a,a125356a,a125357a,a125360a,a125363a,a125364a,a125367a,a125370a,a125371a,a125372a,a125375a,a125378a,a125379a,a125382a,a125385a,a125386a,a125387a,a125390a,a125393a,a125394a,a125397a,a125400a,a125401a,a125402a,a125405a,a125408a,a125409a,a125412a,a125415a,a125416a,a125417a,a125420a,a125423a,a125424a,a125427a,a125430a,a125431a,a125432a,a125435a,a125438a,a125439a,a125442a,a125445a,a125446a,a125447a,a125450a,a125453a,a125454a,a125457a,a125460a,a125461a,a125462a,a125465a,a125468a,a125469a,a125472a,a125475a,a125476a,a125477a,a125480a,a125483a,a125484a,a125487a,a125490a,a125491a,a125492a,a125495a,a125498a,a125499a,a125502a,a125505a,a125506a,a125507a,a125510a,a125513a,a125514a,a125517a,a125520a,a125521a,a125522a,a125525a,a125528a,a125529a,a125532a,a125535a,a125536a,a125537a,a125540a,a125543a,a125544a,a125547a,a125550a,a125551a,a125552a,a125555a,a125558a,a125559a,a125562a,a125565a,a125566a,a125567a,a125570a,a125573a,a125574a,a125577a,a125580a,a125581a,a125582a,a125585a,a125588a,a125589a,a125592a,a125595a,a125596a,a125597a,a125600a,a125603a,a125604a,a125607a,a125610a,a125611a,a125612a,a125615a,a125618a,a125619a,a125622a,a125625a,a125626a,a125627a,a125630a,a125633a,a125634a,a125637a,a125640a,a125641a,a125642a,a125645a,a125648a,a125649a,a125652a,a125655a,a125656a,a125657a,a125660a,a125663a,a125664a,a125667a,a125670a,a125671a,a125672a,a125675a,a125678a,a125679a,a125682a,a125685a,a125686a,a125687a,a125690a,a125693a,a125694a,a125697a,a125700a,a125701a,a125702a,a125705a,a125708a,a125709a,a125712a,a125715a,a125716a,a125717a,a125720a,a125723a,a125724a,a125727a,a125730a,a125731a,a125732a,a125735a,a125738a,a125739a,a125742a,a125745a,a125746a,a125747a,a125750a,a125753a,a125754a,a125757a,a125760a,a125761a,a125762a,a125765a,a125768a,a125769a,a125772a,a125775a,a125776a,a125777a,a125780a,a125783a,a125784a,a125787a,a125790a,a125791a,a125792a,a125795a,a125798a,a125799a,a125802a,a125805a,a125806a,a125807a,a125810a,a125813a,a125814a,a125817a,a125820a,a125821a,a125822a,a125825a,a125828a,a125829a,a125832a,a125835a,a125836a,a125837a,a125840a,a125843a,a125844a,a125847a,a125850a,a125851a,a125852a,a125855a,a125858a,a125859a,a125862a,a125865a,a125866a,a125867a,a125870a,a125873a,a125874a,a125877a,a125880a,a125881a,a125882a,a125885a,a125888a,a125889a,a125892a,a125895a,a125896a,a125897a,a125900a,a125903a,a125904a,a125907a,a125910a,a125911a,a125912a,a125915a,a125918a,a125919a,a125922a,a125925a,a125926a,a125927a,a125930a,a125933a,a125934a,a125937a,a125940a,a125941a,a125942a,a125945a,a125948a,a125949a,a125952a,a125955a,a125956a,a125957a,a125960a,a125963a,a125964a,a125967a,a125970a,a125971a,a125972a,a125975a,a125978a,a125979a,a125982a,a125985a,a125986a,a125987a,a125990a,a125993a,a125994a,a125997a,a126000a,a126001a,a126002a,a126005a,a126008a,a126009a,a126012a,a126015a,a126016a,a126017a,a126020a,a126023a,a126024a,a126027a,a126030a,a126031a,a126032a,a126035a,a126038a,a126039a,a126042a,a126045a,a126046a,a126047a,a126050a,a126053a,a126054a,a126057a,a126060a,a126061a,a126062a,a126065a,a126068a,a126069a,a126072a,a126075a,a126076a,a126077a,a126080a,a126083a,a126084a,a126087a,a126090a,a126091a,a126092a,a126095a,a126098a,a126099a,a126102a,a126105a,a126106a,a126107a,a126110a,a126113a,a126114a,a126117a,a126120a,a126121a,a126122a,a126125a,a126128a,a126129a,a126132a,a126135a,a126136a,a126137a,a126140a,a126143a,a126144a,a126147a,a126150a,a126151a,a126152a,a126155a,a126158a,a126159a,a126162a,a126165a,a126166a,a126167a,a126170a,a126173a,a126174a,a126177a,a126180a,a126181a,a126182a,a126185a,a126188a,a126189a,a126192a,a126195a,a126196a,a126197a,a126200a,a126203a,a126204a,a126207a,a126210a,a126211a,a126212a,a126215a,a126218a,a126219a,a126222a,a126225a,a126226a,a126227a,a126230a,a126233a,a126234a,a126237a,a126240a,a126241a,a126242a,a126245a,a126248a,a126249a,a126252a,a126255a,a126256a,a126257a,a126260a,a126263a,a126264a,a126267a,a126270a,a126271a,a126272a,a126275a,a126278a,a126279a,a126282a,a126285a,a126286a,a126287a,a126290a,a126293a,a126294a,a126297a,a126300a,a126301a,a126302a,a126305a,a126308a,a126309a,a126312a,a126315a,a126316a,a126317a,a126320a,a126323a,a126324a,a126327a,a126330a,a126331a,a126332a,a126335a,a126338a,a126339a,a126342a,a126345a,a126346a,a126347a,a126350a,a126353a,a126354a,a126357a,a126360a,a126361a,a126362a,a126365a,a126368a,a126369a,a126372a,a126375a,a126376a,a126377a,a126380a,a126383a,a126384a,a126387a,a126390a,a126391a,a126392a,a126395a,a126398a,a126399a,a126402a,a126405a,a126406a,a126407a,a126410a,a126413a,a126414a,a126417a,a126420a,a126421a,a126422a,a126425a,a126428a,a126429a,a126432a,a126435a,a126436a,a126437a,a126440a,a126443a,a126444a,a126447a,a126450a,a126451a,a126452a,a126455a,a126458a,a126459a,a126462a,a126465a,a126466a,a126467a,a126470a,a126473a,a126474a,a126477a,a126480a,a126481a,a126482a,a126485a,a126488a,a126489a,a126492a,a126495a,a126496a,a126497a,a126500a,a126503a,a126504a,a126507a,a126510a,a126511a,a126512a,a126515a,a126518a,a126519a,a126522a,a126525a,a126526a,a126527a,a126530a,a126533a,a126534a,a126537a,a126540a,a126541a,a126542a,a126545a,a126548a,a126549a,a126552a,a126555a,a126556a,a126557a,a126560a,a126563a,a126564a,a126567a,a126570a,a126571a,a126572a,a126575a,a126578a,a126579a,a126582a,a126585a,a126586a,a126587a,a126590a,a126593a,a126594a,a126597a,a126600a,a126601a,a126602a,a126605a,a126608a,a126609a,a126612a,a126615a,a126616a,a126617a,a126620a,a126623a,a126624a,a126627a,a126630a,a126631a,a126632a,a126635a,a126638a,a126639a,a126642a,a126645a,a126646a,a126647a,a126650a,a126653a,a126654a,a126657a,a126660a,a126661a,a126662a,a126665a,a126668a,a126669a,a126672a,a126675a,a126676a,a126677a,a126680a,a126683a,a126684a,a126687a,a126690a,a126691a,a126692a,a126695a,a126698a,a126699a,a126702a,a126705a,a126706a,a126707a,a126710a,a126713a,a126714a,a126717a,a126720a,a126721a,a126722a,a126725a,a126728a,a126729a,a126732a,a126735a,a126736a,a126737a,a126740a,a126743a,a126744a,a126747a,a126750a,a126751a,a126752a,a126755a,a126758a,a126759a,a126762a,a126765a,a126766a,a126767a,a126770a,a126773a,a126774a,a126777a,a126780a,a126781a,a126782a,a126785a,a126788a,a126789a,a126792a,a126795a,a126796a,a126797a,a126800a,a126803a,a126804a,a126807a,a126810a,a126811a,a126812a,a126815a,a126818a,a126819a,a126822a,a126825a,a126826a,a126827a,a126830a,a126833a,a126834a,a126837a,a126840a,a126841a,a126842a,a126845a,a126848a,a126849a,a126852a,a126855a,a126856a,a126857a,a126860a,a126863a,a126864a,a126867a,a126870a,a126871a,a126872a,a126875a,a126878a,a126879a,a126882a,a126885a,a126886a,a126887a,a126890a,a126893a,a126894a,a126897a,a126900a,a126901a,a126902a,a126905a,a126908a,a126909a,a126912a,a126915a,a126916a,a126917a,a126920a,a126923a,a126924a,a126927a,a126930a,a126931a,a126932a,a126935a,a126938a,a126939a,a126942a,a126945a,a126946a,a126947a,a126950a,a126953a,a126954a,a126957a,a126960a,a126961a,a126962a,a126965a,a126968a,a126969a,a126972a,a126975a,a126976a,a126977a,a126980a,a126983a,a126984a,a126987a,a126990a,a126991a,a126992a,a126995a,a126998a,a126999a,a127002a,a127005a,a127006a,a127007a,a127010a,a127013a,a127014a,a127017a,a127020a,a127021a,a127022a,a127025a,a127028a,a127029a,a127032a,a127035a,a127036a,a127037a,a127040a,a127043a,a127044a,a127047a,a127050a,a127051a,a127052a,a127055a,a127058a,a127059a,a127062a,a127065a,a127066a,a127067a,a127070a,a127073a,a127074a,a127077a,a127080a,a127081a,a127082a,a127085a,a127088a,a127089a,a127092a,a127095a,a127096a,a127097a,a127100a,a127103a,a127104a,a127107a,a127110a,a127111a,a127112a,a127115a,a127118a,a127119a,a127122a,a127125a,a127126a,a127127a,a127130a,a127133a,a127134a,a127137a,a127140a,a127141a,a127142a,a127145a,a127148a,a127149a,a127152a,a127155a,a127156a,a127157a,a127160a,a127163a,a127164a,a127167a,a127170a,a127171a,a127172a,a127175a,a127178a,a127179a,a127182a,a127185a,a127186a,a127187a,a127190a,a127193a,a127194a,a127197a,a127200a,a127201a,a127202a,a127205a,a127208a,a127209a,a127212a,a127215a,a127216a,a127217a,a127220a,a127223a,a127224a,a127227a,a127230a,a127231a,a127232a,a127235a,a127238a,a127239a,a127242a,a127245a,a127246a,a127247a,a127250a,a127253a,a127254a,a127257a,a127260a,a127261a,a127262a,a127265a,a127268a,a127269a,a127272a,a127275a,a127276a,a127277a,a127280a,a127283a,a127284a,a127287a,a127290a,a127291a,a127292a,a127295a,a127298a,a127299a,a127302a,a127305a,a127306a,a127307a,a127310a,a127313a,a127314a,a127317a,a127320a,a127321a,a127322a,a127325a,a127328a,a127329a,a127332a,a127335a,a127336a,a127337a,a127340a,a127343a,a127344a,a127347a,a127350a,a127351a,a127352a,a127355a,a127358a,a127359a,a127362a,a127365a,a127366a,a127367a,a127370a,a127373a,a127374a,a127377a,a127380a,a127381a,a127382a,a127385a,a127388a,a127389a,a127392a,a127395a,a127396a,a127397a,a127400a,a127403a,a127404a,a127407a,a127410a,a127411a,a127412a,a127415a,a127418a,a127419a,a127422a,a127425a,a127426a,a127427a,a127430a,a127433a,a127434a,a127437a,a127440a,a127441a,a127442a,a127445a,a127448a,a127449a,a127452a,a127455a,a127456a,a127457a,a127460a,a127463a,a127464a,a127467a,a127470a,a127471a,a127472a,a127475a,a127478a,a127479a,a127482a,a127485a,a127486a,a127487a,a127490a,a127493a,a127494a,a127497a,a127500a,a127501a,a127502a,a127505a,a127508a,a127509a,a127512a,a127515a,a127516a,a127517a,a127520a,a127523a,a127524a,a127527a,a127530a,a127531a,a127532a,a127535a,a127538a,a127539a,a127542a,a127545a,a127546a,a127547a,a127550a,a127553a,a127554a,a127557a,a127560a,a127561a,a127562a,a127565a,a127568a,a127569a,a127572a,a127575a,a127576a,a127577a,a127580a,a127583a,a127584a,a127587a,a127590a,a127591a,a127592a,a127595a,a127598a,a127599a,a127602a,a127605a,a127606a,a127607a,a127610a,a127613a,a127614a,a127617a,a127620a,a127621a,a127622a,a127625a,a127628a,a127629a,a127632a,a127635a,a127636a,a127637a,a127640a,a127643a,a127644a,a127647a,a127650a,a127651a,a127652a,a127655a,a127658a,a127659a,a127662a,a127665a,a127666a,a127667a,a127670a,a127673a,a127674a,a127677a,a127680a,a127681a,a127682a,a127685a,a127688a,a127689a,a127692a,a127695a,a127696a,a127697a,a127700a,a127703a,a127704a,a127707a,a127710a,a127711a,a127712a,a127715a,a127718a,a127719a,a127722a,a127725a,a127726a,a127727a,a127730a,a127733a,a127734a,a127737a,a127740a,a127741a,a127742a,a127745a,a127748a,a127749a,a127752a,a127755a,a127756a,a127757a,a127760a,a127763a,a127764a,a127767a,a127770a,a127771a,a127772a,a127775a,a127778a,a127779a,a127782a,a127785a,a127786a,a127787a,a127790a,a127793a,a127794a,a127797a,a127800a,a127801a,a127802a,a127805a,a127808a,a127809a,a127812a,a127815a,a127816a,a127817a,a127820a,a127823a,a127824a,a127827a,a127830a,a127831a,a127832a,a127835a,a127838a,a127839a,a127842a,a127845a,a127846a,a127847a,a127850a,a127853a,a127854a,a127857a,a127860a,a127861a,a127862a,a127865a,a127868a,a127869a,a127872a,a127875a,a127876a,a127877a,a127880a,a127883a,a127884a,a127887a,a127890a,a127891a,a127892a,a127895a,a127898a,a127899a,a127902a,a127905a,a127906a,a127907a,a127910a,a127913a,a127914a,a127917a,a127920a,a127921a,a127922a,a127925a,a127928a,a127929a,a127932a,a127935a,a127936a,a127937a,a127940a,a127943a,a127944a,a127947a,a127950a,a127951a,a127952a,a127955a,a127958a,a127959a,a127962a,a127965a,a127966a,a127967a,a127970a,a127973a,a127974a,a127977a,a127980a,a127981a,a127982a,a127985a,a127988a,a127989a,a127992a,a127995a,a127996a,a127997a,a128000a,a128003a,a128004a,a128007a,a128010a,a128011a,a128012a,a128015a,a128018a,a128019a,a128022a,a128025a,a128026a,a128027a,a128030a,a128033a,a128034a,a128037a,a128040a,a128041a,a128042a,a128045a,a128048a,a128049a,a128052a,a128055a,a128056a,a128057a,a128060a,a128063a,a128064a,a128067a,a128070a,a128071a,a128072a,a128075a,a128078a,a128079a,a128082a,a128085a,a128086a,a128087a,a128090a,a128093a,a128094a,a128097a,a128100a,a128101a,a128102a,a128105a,a128108a,a128109a,a128112a,a128115a,a128116a,a128117a,a128120a,a128123a,a128124a,a128127a,a128130a,a128131a,a128132a,a128135a,a128138a,a128139a,a128142a,a128145a,a128146a,a128147a,a128150a,a128153a,a128154a,a128157a,a128160a,a128161a,a128162a,a128165a,a128168a,a128169a,a128172a,a128175a,a128176a,a128177a,a128180a,a128183a,a128184a,a128187a,a128190a,a128191a,a128192a,a128195a,a128198a,a128199a,a128202a,a128205a,a128206a,a128207a,a128210a,a128213a,a128214a,a128217a,a128220a,a128221a,a128222a,a128225a,a128228a,a128229a,a128232a,a128235a,a128236a,a128237a,a128240a,a128243a,a128244a,a128247a,a128250a,a128251a,a128252a,a128255a,a128258a,a128259a,a128262a,a128265a,a128266a,a128267a,a128270a,a128273a,a128274a,a128277a,a128280a,a128281a,a128282a,a128285a,a128288a,a128289a,a128292a,a128295a,a128296a,a128297a,a128300a,a128303a,a128304a,a128307a,a128310a,a128311a,a128312a,a128315a,a128318a,a128319a,a128322a,a128325a,a128326a,a128327a,a128330a,a128333a,a128334a,a128337a,a128340a,a128341a,a128342a,a128345a,a128348a,a128349a,a128352a,a128355a,a128356a,a128357a,a128360a,a128363a,a128364a,a128367a,a128370a,a128371a,a128372a,a128375a,a128378a,a128379a,a128382a,a128385a,a128386a,a128387a,a128390a,a128393a,a128394a,a128397a,a128400a,a128401a,a128402a,a128405a,a128408a,a128409a,a128412a,a128415a,a128416a,a128417a,a128420a,a128423a,a128424a,a128427a,a128430a,a128431a,a128432a,a128435a,a128438a,a128439a,a128442a,a128445a,a128446a,a128447a,a128450a,a128453a,a128454a,a128457a,a128460a,a128461a,a128462a,a128465a,a128468a,a128469a,a128472a,a128475a,a128476a,a128477a,a128480a,a128483a,a128484a,a128487a,a128490a,a128491a,a128492a,a128495a,a128498a,a128499a,a128502a,a128505a,a128506a,a128507a,a128510a,a128513a,a128514a,a128517a,a128520a,a128521a,a128522a,a128525a,a128528a,a128529a,a128532a,a128535a,a128536a,a128537a,a128540a,a128543a,a128544a,a128547a,a128550a,a128551a,a128552a,a128555a,a128558a,a128559a,a128562a,a128565a,a128566a,a128567a,a128570a,a128573a,a128574a,a128577a,a128580a,a128581a,a128582a,a128585a,a128588a,a128589a,a128592a,a128595a,a128596a,a128597a,a128600a,a128603a,a128604a,a128607a,a128610a,a128611a,a128612a,a128615a,a128618a,a128619a,a128622a,a128625a,a128626a,a128627a,a128630a,a128633a,a128634a,a128637a,a128640a,a128641a,a128642a,a128645a,a128648a,a128649a,a128652a,a128655a,a128656a,a128657a,a128660a,a128663a,a128664a,a128667a,a128670a,a128671a,a128672a,a128675a,a128678a,a128679a,a128682a,a128685a,a128686a,a128687a,a128690a,a128693a,a128694a,a128697a,a128700a,a128701a,a128702a,a128705a,a128708a,a128709a,a128712a,a128715a,a128716a,a128717a,a128720a,a128723a,a128724a,a128727a,a128730a,a128731a,a128732a,a128735a,a128738a,a128739a,a128742a,a128745a,a128746a,a128747a,a128750a,a128753a,a128754a,a128757a,a128760a,a128761a,a128762a,a128765a,a128768a,a128769a,a128772a,a128775a,a128776a,a128777a,a128780a,a128783a,a128784a,a128787a,a128790a,a128791a,a128792a,a128795a,a128798a,a128799a,a128802a,a128805a,a128806a,a128807a,a128810a,a128813a,a128814a,a128817a,a128820a,a128821a,a128822a,a128825a,a128828a,a128829a,a128832a,a128835a,a128836a,a128837a,a128840a,a128843a,a128844a,a128847a,a128850a,a128851a,a128852a,a128855a,a128858a,a128859a,a128862a,a128865a,a128866a,a128867a,a128870a,a128873a,a128874a,a128877a,a128880a,a128881a,a128882a,a128885a,a128888a,a128889a,a128892a,a128895a,a128896a,a128897a,a128900a,a128903a,a128904a,a128907a,a128910a,a128911a,a128912a,a128915a,a128918a,a128919a,a128922a,a128925a,a128926a,a128927a,a128930a,a128933a,a128934a,a128937a,a128940a,a128941a,a128942a,a128945a,a128948a,a128949a,a128952a,a128955a,a128956a,a128957a,a128960a,a128963a,a128964a,a128967a,a128970a,a128971a,a128972a,a128975a,a128978a,a128979a,a128982a,a128985a,a128986a,a128987a,a128990a,a128993a,a128994a,a128997a,a129000a,a129001a,a129002a,a129005a,a129008a,a129009a,a129012a,a129015a,a129016a,a129017a,a129020a,a129023a,a129024a,a129027a,a129030a,a129031a,a129032a,a129035a,a129038a,a129039a,a129042a,a129045a,a129046a,a129047a,a129050a,a129053a,a129054a,a129057a,a129060a,a129061a,a129062a,a129065a,a129068a,a129069a,a129072a,a129075a,a129076a,a129077a,a129080a,a129083a,a129084a,a129087a,a129090a,a129091a,a129092a,a129095a,a129098a,a129099a,a129102a,a129105a,a129106a,a129107a,a129110a,a129113a,a129114a,a129117a,a129120a,a129121a,a129122a,a129125a,a129128a,a129129a,a129132a,a129135a,a129136a,a129137a,a129140a,a129143a,a129144a,a129147a,a129150a,a129151a,a129152a,a129155a,a129158a,a129159a,a129162a,a129165a,a129166a,a129167a,a129170a,a129173a,a129174a,a129177a,a129180a,a129181a,a129182a,a129185a,a129188a,a129189a,a129192a,a129195a,a129196a,a129197a,a129200a,a129203a,a129204a,a129207a,a129210a,a129211a,a129212a,a129215a,a129218a,a129219a,a129222a,a129225a,a129226a,a129227a,a129230a,a129233a,a129234a,a129237a,a129240a,a129241a,a129242a,a129245a,a129248a,a129249a,a129252a,a129255a,a129256a,a129257a,a129260a,a129263a,a129264a,a129267a,a129270a,a129271a,a129272a,a129275a,a129278a,a129279a,a129282a,a129285a,a129286a,a129287a,a129290a,a129293a,a129294a,a129297a,a129300a,a129301a,a129302a,a129305a,a129308a,a129309a,a129312a,a129315a,a129316a,a129317a,a129320a,a129323a,a129324a,a129327a,a129330a,a129331a,a129332a,a129335a,a129338a,a129339a,a129342a,a129345a,a129346a,a129347a,a129350a,a129353a,a129354a,a129357a,a129360a,a129361a,a129362a,a129365a,a129368a,a129369a,a129372a,a129375a,a129376a,a129377a,a129380a,a129383a,a129384a,a129387a,a129390a,a129391a,a129392a,a129395a,a129398a,a129399a,a129402a,a129405a,a129406a,a129407a,a129410a,a129413a,a129414a,a129417a,a129420a,a129421a,a129422a,a129425a,a129428a,a129429a,a129432a,a129435a,a129436a,a129437a,a129440a,a129443a,a129444a,a129447a,a129450a,a129451a,a129452a,a129455a,a129458a,a129459a,a129462a,a129465a,a129466a,a129467a,a129470a,a129473a,a129474a,a129477a,a129480a,a129481a,a129482a,a129485a,a129488a,a129489a,a129492a,a129495a,a129496a,a129497a,a129500a,a129503a,a129504a,a129507a,a129510a,a129511a,a129512a,a129515a,a129518a,a129519a,a129522a,a129525a,a129526a,a129527a,a129530a,a129533a,a129534a,a129537a,a129540a,a129541a,a129542a,a129545a,a129548a,a129549a,a129552a,a129555a,a129556a,a129557a,a129560a,a129563a,a129564a,a129567a,a129570a,a129571a,a129572a,a129575a,a129578a,a129579a,a129582a,a129585a,a129586a,a129587a,a129590a,a129593a,a129594a,a129597a,a129600a,a129601a,a129602a,a129605a,a129608a,a129609a,a129612a,a129615a,a129616a,a129617a,a129620a,a129623a,a129624a,a129627a,a129630a,a129631a,a129632a,a129635a,a129638a,a129639a,a129642a,a129645a,a129646a,a129647a,a129650a,a129653a,a129654a,a129657a,a129660a,a129661a,a129662a,a129665a,a129668a,a129669a,a129672a,a129675a,a129676a,a129677a,a129680a,a129683a,a129684a,a129687a,a129690a,a129691a,a129692a,a129695a,a129698a,a129699a,a129702a,a129705a,a129706a,a129707a,a129710a,a129713a,a129714a,a129717a,a129720a,a129721a,a129722a,a129725a,a129728a,a129729a,a129732a,a129735a,a129736a,a129737a,a129740a,a129743a,a129744a,a129747a,a129750a,a129751a,a129752a,a129755a,a129758a,a129759a,a129762a,a129765a,a129766a,a129767a,a129770a,a129773a,a129774a,a129777a,a129780a,a129781a,a129782a,a129785a,a129788a,a129789a,a129792a,a129795a,a129796a,a129797a,a129800a,a129803a,a129804a,a129807a,a129810a,a129811a,a129812a,a129815a,a129818a,a129819a,a129822a,a129825a,a129826a,a129827a,a129830a,a129833a,a129834a,a129837a,a129840a,a129841a,a129842a,a129845a,a129848a,a129849a,a129852a,a129855a,a129856a,a129857a,a129860a,a129863a,a129864a,a129867a,a129870a,a129871a,a129872a,a129875a,a129878a,a129879a,a129882a,a129885a,a129886a,a129887a,a129890a,a129893a,a129894a,a129897a,a129900a,a129901a,a129902a,a129905a,a129908a,a129909a,a129912a,a129915a,a129916a,a129917a,a129920a,a129923a,a129924a,a129927a,a129930a,a129931a,a129932a,a129935a,a129938a,a129939a,a129942a,a129945a,a129946a,a129947a,a129950a,a129953a,a129954a,a129957a,a129960a,a129961a,a129962a,a129965a,a129968a,a129969a,a129972a,a129975a,a129976a,a129977a,a129980a,a129983a,a129984a,a129987a,a129990a,a129991a,a129992a,a129995a,a129998a,a129999a,a130002a,a130005a,a130006a,a130007a,a130010a,a130013a,a130014a,a130017a,a130020a,a130021a,a130022a,a130025a,a130028a,a130029a,a130032a,a130035a,a130036a,a130037a,a130040a,a130043a,a130044a,a130047a,a130050a,a130051a,a130052a,a130055a,a130058a,a130059a,a130062a,a130065a,a130066a,a130067a,a130070a,a130073a,a130074a,a130077a,a130080a,a130081a,a130082a,a130085a,a130088a,a130089a,a130092a,a130095a,a130096a,a130097a,a130100a,a130103a,a130104a,a130107a,a130110a,a130111a,a130112a,a130115a,a130118a,a130119a,a130122a,a130125a,a130126a,a130127a,a130130a,a130133a,a130134a,a130137a,a130140a,a130141a,a130142a,a130145a,a130148a,a130149a,a130152a,a130155a,a130156a,a130157a,a130160a,a130163a,a130164a,a130167a,a130170a,a130171a,a130172a,a130175a,a130178a,a130179a,a130182a,a130185a,a130186a,a130187a,a130190a,a130193a,a130194a,a130197a,a130200a,a130201a,a130202a,a130205a,a130208a,a130209a,a130212a,a130215a,a130216a,a130217a,a130220a,a130223a,a130224a,a130227a,a130230a,a130231a,a130232a,a130235a,a130238a,a130239a,a130242a,a130245a,a130246a,a130247a,a130250a,a130253a,a130254a,a130257a,a130260a,a130261a,a130262a,a130265a,a130268a,a130269a,a130272a,a130275a,a130276a,a130277a,a130280a,a130283a,a130284a,a130287a,a130290a,a130291a,a130292a,a130295a,a130298a,a130299a,a130302a,a130305a,a130306a,a130307a,a130310a,a130313a,a130314a,a130317a,a130320a,a130321a,a130322a,a130325a,a130328a,a130329a,a130332a,a130335a,a130336a,a130337a,a130340a,a130343a,a130344a,a130347a,a130350a,a130351a,a130352a,a130355a,a130358a,a130359a,a130362a,a130365a,a130366a,a130367a,a130370a,a130373a,a130374a,a130377a,a130380a,a130381a,a130382a,a130385a,a130388a,a130389a,a130392a,a130395a,a130396a,a130397a,a130400a,a130403a,a130404a,a130407a,a130410a,a130411a,a130412a,a130415a,a130418a,a130419a,a130422a,a130425a,a130426a,a130427a,a130430a,a130433a,a130434a,a130437a,a130440a,a130441a,a130442a,a130445a,a130448a,a130449a,a130452a,a130455a,a130456a,a130457a,a130460a,a130463a,a130464a,a130467a,a130470a,a130471a,a130472a,a130475a,a130478a,a130479a,a130482a,a130485a,a130486a,a130487a,a130490a,a130493a,a130494a,a130497a,a130500a,a130501a,a130502a,a130505a,a130508a,a130509a,a130512a,a130515a,a130516a,a130517a,a130520a,a130523a,a130524a,a130527a,a130530a,a130531a,a130532a,a130535a,a130538a,a130539a,a130542a,a130545a,a130546a,a130547a,a130550a,a130553a,a130554a,a130557a,a130560a,a130561a,a130562a,a130565a,a130568a,a130569a,a130572a,a130575a,a130576a,a130577a,a130580a,a130583a,a130584a,a130587a,a130590a,a130591a,a130592a,a130595a,a130598a,a130599a,a130602a,a130605a,a130606a,a130607a,a130610a,a130613a,a130614a,a130617a,a130620a,a130621a,a130622a,a130625a,a130628a,a130629a,a130632a,a130635a,a130636a,a130637a,a130640a,a130643a,a130644a,a130647a,a130650a,a130651a,a130652a,a130655a,a130658a,a130659a,a130662a,a130665a,a130666a,a130667a,a130670a,a130673a,a130674a,a130677a,a130680a,a130681a,a130682a,a130685a,a130688a,a130689a,a130692a,a130695a,a130696a,a130697a,a130700a,a130703a,a130704a,a130707a,a130710a,a130711a,a130712a,a130715a,a130718a,a130719a,a130722a,a130725a,a130726a,a130727a,a130730a,a130733a,a130734a,a130737a,a130740a,a130741a,a130742a,a130745a,a130748a,a130749a,a130752a,a130755a,a130756a,a130757a,a130760a,a130763a,a130764a,a130767a,a130770a,a130771a,a130772a,a130775a,a130778a,a130779a,a130782a,a130785a,a130786a,a130787a,a130790a,a130793a,a130794a,a130797a,a130800a,a130801a,a130802a,a130805a,a130808a,a130809a,a130812a,a130815a,a130816a,a130817a,a130820a,a130823a,a130824a,a130827a,a130830a,a130831a,a130832a,a130835a,a130838a,a130839a,a130842a,a130845a,a130846a,a130847a,a130850a,a130853a,a130854a,a130857a,a130860a,a130861a,a130862a,a130865a,a130868a,a130869a,a130872a,a130875a,a130876a,a130877a,a130880a,a130883a,a130884a,a130887a,a130890a,a130891a,a130892a,a130895a,a130898a,a130899a,a130902a,a130905a,a130906a,a130907a,a130910a,a130913a,a130914a,a130917a,a130920a,a130921a,a130922a,a130925a,a130928a,a130929a,a130932a,a130935a,a130936a,a130937a,a130940a,a130943a,a130944a,a130947a,a130950a,a130951a,a130952a,a130955a,a130958a,a130959a,a130962a,a130965a,a130966a,a130967a,a130970a,a130973a,a130974a,a130977a,a130980a,a130981a,a130982a,a130985a,a130988a,a130989a,a130992a,a130995a,a130996a,a130997a,a131000a,a131003a,a131004a,a131007a,a131010a,a131011a,a131012a,a131015a,a131018a,a131019a,a131022a,a131025a,a131026a,a131027a,a131030a,a131033a,a131034a,a131037a,a131040a,a131041a,a131042a,a131045a,a131048a,a131049a,a131052a,a131055a,a131056a,a131057a,a131060a,a131063a,a131064a,a131067a,a131070a,a131071a,a131072a,a131075a,a131078a,a131079a,a131082a,a131085a,a131086a,a131087a,a131090a,a131093a,a131094a,a131097a,a131100a,a131101a,a131102a,a131105a,a131108a,a131109a,a131112a,a131115a,a131116a,a131117a,a131120a,a131123a,a131124a,a131127a,a131130a,a131131a,a131132a,a131135a,a131138a,a131139a,a131142a,a131145a,a131146a,a131147a,a131150a,a131153a,a131154a,a131157a,a131160a,a131161a,a131162a,a131165a,a131168a,a131169a,a131172a,a131175a,a131176a,a131177a,a131180a,a131183a,a131184a,a131187a,a131190a,a131191a,a131192a,a131195a,a131198a,a131199a,a131202a,a131205a,a131206a,a131207a,a131210a,a131213a,a131214a,a131217a,a131220a,a131221a,a131222a,a131225a,a131228a,a131229a,a131232a,a131235a,a131236a,a131237a,a131240a,a131243a,a131244a,a131247a,a131250a,a131251a,a131252a: std_logic;
begin

A40 <=( a14272a ) or ( a9515a );
 a1a <=( a131252a  and  a131237a );
 a2a <=( a131222a  and  a131207a );
 a3a <=( a131192a  and  a131177a );
 a4a <=( a131162a  and  a131147a );
 a5a <=( a131132a  and  a131117a );
 a6a <=( a131102a  and  a131087a );
 a7a <=( a131072a  and  a131057a );
 a8a <=( a131042a  and  a131027a );
 a9a <=( a131012a  and  a130997a );
 a10a <=( a130982a  and  a130967a );
 a11a <=( a130952a  and  a130937a );
 a12a <=( a130922a  and  a130907a );
 a13a <=( a130892a  and  a130877a );
 a14a <=( a130862a  and  a130847a );
 a15a <=( a130832a  and  a130817a );
 a16a <=( a130802a  and  a130787a );
 a17a <=( a130772a  and  a130757a );
 a18a <=( a130742a  and  a130727a );
 a19a <=( a130712a  and  a130697a );
 a20a <=( a130682a  and  a130667a );
 a21a <=( a130652a  and  a130637a );
 a22a <=( a130622a  and  a130607a );
 a23a <=( a130592a  and  a130577a );
 a24a <=( a130562a  and  a130547a );
 a25a <=( a130532a  and  a130517a );
 a26a <=( a130502a  and  a130487a );
 a27a <=( a130472a  and  a130457a );
 a28a <=( a130442a  and  a130427a );
 a29a <=( a130412a  and  a130397a );
 a30a <=( a130382a  and  a130367a );
 a31a <=( a130352a  and  a130337a );
 a32a <=( a130322a  and  a130307a );
 a33a <=( a130292a  and  a130277a );
 a34a <=( a130262a  and  a130247a );
 a35a <=( a130232a  and  a130217a );
 a36a <=( a130202a  and  a130187a );
 a37a <=( a130172a  and  a130157a );
 a38a <=( a130142a  and  a130127a );
 a39a <=( a130112a  and  a130097a );
 a40a <=( a130082a  and  a130067a );
 a41a <=( a130052a  and  a130037a );
 a42a <=( a130022a  and  a130007a );
 a43a <=( a129992a  and  a129977a );
 a44a <=( a129962a  and  a129947a );
 a45a <=( a129932a  and  a129917a );
 a46a <=( a129902a  and  a129887a );
 a47a <=( a129872a  and  a129857a );
 a48a <=( a129842a  and  a129827a );
 a49a <=( a129812a  and  a129797a );
 a50a <=( a129782a  and  a129767a );
 a51a <=( a129752a  and  a129737a );
 a52a <=( a129722a  and  a129707a );
 a53a <=( a129692a  and  a129677a );
 a54a <=( a129662a  and  a129647a );
 a55a <=( a129632a  and  a129617a );
 a56a <=( a129602a  and  a129587a );
 a57a <=( a129572a  and  a129557a );
 a58a <=( a129542a  and  a129527a );
 a59a <=( a129512a  and  a129497a );
 a60a <=( a129482a  and  a129467a );
 a61a <=( a129452a  and  a129437a );
 a62a <=( a129422a  and  a129407a );
 a63a <=( a129392a  and  a129377a );
 a64a <=( a129362a  and  a129347a );
 a65a <=( a129332a  and  a129317a );
 a66a <=( a129302a  and  a129287a );
 a67a <=( a129272a  and  a129257a );
 a68a <=( a129242a  and  a129227a );
 a69a <=( a129212a  and  a129197a );
 a70a <=( a129182a  and  a129167a );
 a71a <=( a129152a  and  a129137a );
 a72a <=( a129122a  and  a129107a );
 a73a <=( a129092a  and  a129077a );
 a74a <=( a129062a  and  a129047a );
 a75a <=( a129032a  and  a129017a );
 a76a <=( a129002a  and  a128987a );
 a77a <=( a128972a  and  a128957a );
 a78a <=( a128942a  and  a128927a );
 a79a <=( a128912a  and  a128897a );
 a80a <=( a128882a  and  a128867a );
 a81a <=( a128852a  and  a128837a );
 a82a <=( a128822a  and  a128807a );
 a83a <=( a128792a  and  a128777a );
 a84a <=( a128762a  and  a128747a );
 a85a <=( a128732a  and  a128717a );
 a86a <=( a128702a  and  a128687a );
 a87a <=( a128672a  and  a128657a );
 a88a <=( a128642a  and  a128627a );
 a89a <=( a128612a  and  a128597a );
 a90a <=( a128582a  and  a128567a );
 a91a <=( a128552a  and  a128537a );
 a92a <=( a128522a  and  a128507a );
 a93a <=( a128492a  and  a128477a );
 a94a <=( a128462a  and  a128447a );
 a95a <=( a128432a  and  a128417a );
 a96a <=( a128402a  and  a128387a );
 a97a <=( a128372a  and  a128357a );
 a98a <=( a128342a  and  a128327a );
 a99a <=( a128312a  and  a128297a );
 a100a <=( a128282a  and  a128267a );
 a101a <=( a128252a  and  a128237a );
 a102a <=( a128222a  and  a128207a );
 a103a <=( a128192a  and  a128177a );
 a104a <=( a128162a  and  a128147a );
 a105a <=( a128132a  and  a128117a );
 a106a <=( a128102a  and  a128087a );
 a107a <=( a128072a  and  a128057a );
 a108a <=( a128042a  and  a128027a );
 a109a <=( a128012a  and  a127997a );
 a110a <=( a127982a  and  a127967a );
 a111a <=( a127952a  and  a127937a );
 a112a <=( a127922a  and  a127907a );
 a113a <=( a127892a  and  a127877a );
 a114a <=( a127862a  and  a127847a );
 a115a <=( a127832a  and  a127817a );
 a116a <=( a127802a  and  a127787a );
 a117a <=( a127772a  and  a127757a );
 a118a <=( a127742a  and  a127727a );
 a119a <=( a127712a  and  a127697a );
 a120a <=( a127682a  and  a127667a );
 a121a <=( a127652a  and  a127637a );
 a122a <=( a127622a  and  a127607a );
 a123a <=( a127592a  and  a127577a );
 a124a <=( a127562a  and  a127547a );
 a125a <=( a127532a  and  a127517a );
 a126a <=( a127502a  and  a127487a );
 a127a <=( a127472a  and  a127457a );
 a128a <=( a127442a  and  a127427a );
 a129a <=( a127412a  and  a127397a );
 a130a <=( a127382a  and  a127367a );
 a131a <=( a127352a  and  a127337a );
 a132a <=( a127322a  and  a127307a );
 a133a <=( a127292a  and  a127277a );
 a134a <=( a127262a  and  a127247a );
 a135a <=( a127232a  and  a127217a );
 a136a <=( a127202a  and  a127187a );
 a137a <=( a127172a  and  a127157a );
 a138a <=( a127142a  and  a127127a );
 a139a <=( a127112a  and  a127097a );
 a140a <=( a127082a  and  a127067a );
 a141a <=( a127052a  and  a127037a );
 a142a <=( a127022a  and  a127007a );
 a143a <=( a126992a  and  a126977a );
 a144a <=( a126962a  and  a126947a );
 a145a <=( a126932a  and  a126917a );
 a146a <=( a126902a  and  a126887a );
 a147a <=( a126872a  and  a126857a );
 a148a <=( a126842a  and  a126827a );
 a149a <=( a126812a  and  a126797a );
 a150a <=( a126782a  and  a126767a );
 a151a <=( a126752a  and  a126737a );
 a152a <=( a126722a  and  a126707a );
 a153a <=( a126692a  and  a126677a );
 a154a <=( a126662a  and  a126647a );
 a155a <=( a126632a  and  a126617a );
 a156a <=( a126602a  and  a126587a );
 a157a <=( a126572a  and  a126557a );
 a158a <=( a126542a  and  a126527a );
 a159a <=( a126512a  and  a126497a );
 a160a <=( a126482a  and  a126467a );
 a161a <=( a126452a  and  a126437a );
 a162a <=( a126422a  and  a126407a );
 a163a <=( a126392a  and  a126377a );
 a164a <=( a126362a  and  a126347a );
 a165a <=( a126332a  and  a126317a );
 a166a <=( a126302a  and  a126287a );
 a167a <=( a126272a  and  a126257a );
 a168a <=( a126242a  and  a126227a );
 a169a <=( a126212a  and  a126197a );
 a170a <=( a126182a  and  a126167a );
 a171a <=( a126152a  and  a126137a );
 a172a <=( a126122a  and  a126107a );
 a173a <=( a126092a  and  a126077a );
 a174a <=( a126062a  and  a126047a );
 a175a <=( a126032a  and  a126017a );
 a176a <=( a126002a  and  a125987a );
 a177a <=( a125972a  and  a125957a );
 a178a <=( a125942a  and  a125927a );
 a179a <=( a125912a  and  a125897a );
 a180a <=( a125882a  and  a125867a );
 a181a <=( a125852a  and  a125837a );
 a182a <=( a125822a  and  a125807a );
 a183a <=( a125792a  and  a125777a );
 a184a <=( a125762a  and  a125747a );
 a185a <=( a125732a  and  a125717a );
 a186a <=( a125702a  and  a125687a );
 a187a <=( a125672a  and  a125657a );
 a188a <=( a125642a  and  a125627a );
 a189a <=( a125612a  and  a125597a );
 a190a <=( a125582a  and  a125567a );
 a191a <=( a125552a  and  a125537a );
 a192a <=( a125522a  and  a125507a );
 a193a <=( a125492a  and  a125477a );
 a194a <=( a125462a  and  a125447a );
 a195a <=( a125432a  and  a125417a );
 a196a <=( a125402a  and  a125387a );
 a197a <=( a125372a  and  a125357a );
 a198a <=( a125342a  and  a125327a );
 a199a <=( a125312a  and  a125297a );
 a200a <=( a125282a  and  a125267a );
 a201a <=( a125252a  and  a125237a );
 a202a <=( a125222a  and  a125207a );
 a203a <=( a125192a  and  a125177a );
 a204a <=( a125162a  and  a125147a );
 a205a <=( a125132a  and  a125117a );
 a206a <=( a125102a  and  a125087a );
 a207a <=( a125072a  and  a125057a );
 a208a <=( a125042a  and  a125027a );
 a209a <=( a125012a  and  a124997a );
 a210a <=( a124982a  and  a124967a );
 a211a <=( a124952a  and  a124937a );
 a212a <=( a124922a  and  a124907a );
 a213a <=( a124892a  and  a124877a );
 a214a <=( a124862a  and  a124847a );
 a215a <=( a124832a  and  a124817a );
 a216a <=( a124802a  and  a124787a );
 a217a <=( a124772a  and  a124757a );
 a218a <=( a124742a  and  a124727a );
 a219a <=( a124712a  and  a124697a );
 a220a <=( a124682a  and  a124667a );
 a221a <=( a124652a  and  a124637a );
 a222a <=( a124622a  and  a124607a );
 a223a <=( a124592a  and  a124577a );
 a224a <=( a124562a  and  a124547a );
 a225a <=( a124532a  and  a124517a );
 a226a <=( a124502a  and  a124487a );
 a227a <=( a124472a  and  a124457a );
 a228a <=( a124442a  and  a124427a );
 a229a <=( a124412a  and  a124397a );
 a230a <=( a124382a  and  a124367a );
 a231a <=( a124352a  and  a124337a );
 a232a <=( a124322a  and  a124307a );
 a233a <=( a124292a  and  a124277a );
 a234a <=( a124262a  and  a124247a );
 a235a <=( a124232a  and  a124217a );
 a236a <=( a124202a  and  a124187a );
 a237a <=( a124172a  and  a124157a );
 a238a <=( a124142a  and  a124127a );
 a239a <=( a124112a  and  a124097a );
 a240a <=( a124082a  and  a124067a );
 a241a <=( a124052a  and  a124037a );
 a242a <=( a124022a  and  a124007a );
 a243a <=( a123992a  and  a123977a );
 a244a <=( a123962a  and  a123947a );
 a245a <=( a123932a  and  a123917a );
 a246a <=( a123902a  and  a123887a );
 a247a <=( a123872a  and  a123857a );
 a248a <=( a123842a  and  a123827a );
 a249a <=( a123812a  and  a123797a );
 a250a <=( a123782a  and  a123767a );
 a251a <=( a123752a  and  a123737a );
 a252a <=( a123722a  and  a123707a );
 a253a <=( a123692a  and  a123677a );
 a254a <=( a123662a  and  a123647a );
 a255a <=( a123632a  and  a123617a );
 a256a <=( a123602a  and  a123587a );
 a257a <=( a123572a  and  a123557a );
 a258a <=( a123542a  and  a123527a );
 a259a <=( a123512a  and  a123497a );
 a260a <=( a123482a  and  a123467a );
 a261a <=( a123452a  and  a123437a );
 a262a <=( a123422a  and  a123407a );
 a263a <=( a123392a  and  a123377a );
 a264a <=( a123362a  and  a123347a );
 a265a <=( a123332a  and  a123317a );
 a266a <=( a123302a  and  a123287a );
 a267a <=( a123272a  and  a123257a );
 a268a <=( a123242a  and  a123227a );
 a269a <=( a123212a  and  a123197a );
 a270a <=( a123182a  and  a123167a );
 a271a <=( a123152a  and  a123137a );
 a272a <=( a123122a  and  a123107a );
 a273a <=( a123092a  and  a123077a );
 a274a <=( a123062a  and  a123047a );
 a275a <=( a123032a  and  a123017a );
 a276a <=( a123002a  and  a122987a );
 a277a <=( a122972a  and  a122957a );
 a278a <=( a122942a  and  a122927a );
 a279a <=( a122912a  and  a122897a );
 a280a <=( a122882a  and  a122867a );
 a281a <=( a122852a  and  a122837a );
 a282a <=( a122822a  and  a122807a );
 a283a <=( a122792a  and  a122777a );
 a284a <=( a122762a  and  a122747a );
 a285a <=( a122732a  and  a122717a );
 a286a <=( a122702a  and  a122687a );
 a287a <=( a122672a  and  a122657a );
 a288a <=( a122642a  and  a122627a );
 a289a <=( a122612a  and  a122597a );
 a290a <=( a122582a  and  a122567a );
 a291a <=( a122552a  and  a122537a );
 a292a <=( a122522a  and  a122507a );
 a293a <=( a122492a  and  a122477a );
 a294a <=( a122462a  and  a122447a );
 a295a <=( a122432a  and  a122417a );
 a296a <=( a122402a  and  a122387a );
 a297a <=( a122372a  and  a122357a );
 a298a <=( a122342a  and  a122327a );
 a299a <=( a122312a  and  a122297a );
 a300a <=( a122282a  and  a122267a );
 a301a <=( a122252a  and  a122237a );
 a302a <=( a122222a  and  a122207a );
 a303a <=( a122192a  and  a122177a );
 a304a <=( a122162a  and  a122147a );
 a305a <=( a122132a  and  a122117a );
 a306a <=( a122102a  and  a122087a );
 a307a <=( a122072a  and  a122057a );
 a308a <=( a122042a  and  a122027a );
 a309a <=( a122012a  and  a121997a );
 a310a <=( a121982a  and  a121967a );
 a311a <=( a121952a  and  a121937a );
 a312a <=( a121922a  and  a121907a );
 a313a <=( a121892a  and  a121877a );
 a314a <=( a121862a  and  a121847a );
 a315a <=( a121832a  and  a121817a );
 a316a <=( a121802a  and  a121787a );
 a317a <=( a121772a  and  a121757a );
 a318a <=( a121742a  and  a121727a );
 a319a <=( a121712a  and  a121697a );
 a320a <=( a121682a  and  a121667a );
 a321a <=( a121652a  and  a121637a );
 a322a <=( a121622a  and  a121607a );
 a323a <=( a121592a  and  a121577a );
 a324a <=( a121562a  and  a121547a );
 a325a <=( a121532a  and  a121517a );
 a326a <=( a121502a  and  a121487a );
 a327a <=( a121472a  and  a121457a );
 a328a <=( a121442a  and  a121427a );
 a329a <=( a121412a  and  a121397a );
 a330a <=( a121382a  and  a121367a );
 a331a <=( a121352a  and  a121337a );
 a332a <=( a121322a  and  a121307a );
 a333a <=( a121292a  and  a121277a );
 a334a <=( a121262a  and  a121247a );
 a335a <=( a121232a  and  a121217a );
 a336a <=( a121202a  and  a121187a );
 a337a <=( a121172a  and  a121157a );
 a338a <=( a121142a  and  a121127a );
 a339a <=( a121112a  and  a121097a );
 a340a <=( a121082a  and  a121067a );
 a341a <=( a121052a  and  a121037a );
 a342a <=( a121022a  and  a121007a );
 a343a <=( a120992a  and  a120977a );
 a344a <=( a120962a  and  a120947a );
 a345a <=( a120932a  and  a120917a );
 a346a <=( a120902a  and  a120887a );
 a347a <=( a120872a  and  a120857a );
 a348a <=( a120842a  and  a120827a );
 a349a <=( a120812a  and  a120797a );
 a350a <=( a120782a  and  a120767a );
 a351a <=( a120752a  and  a120737a );
 a352a <=( a120722a  and  a120707a );
 a353a <=( a120692a  and  a120677a );
 a354a <=( a120662a  and  a120647a );
 a355a <=( a120632a  and  a120617a );
 a356a <=( a120602a  and  a120587a );
 a357a <=( a120572a  and  a120557a );
 a358a <=( a120542a  and  a120527a );
 a359a <=( a120512a  and  a120497a );
 a360a <=( a120482a  and  a120467a );
 a361a <=( a120452a  and  a120437a );
 a362a <=( a120422a  and  a120407a );
 a363a <=( a120392a  and  a120377a );
 a364a <=( a120362a  and  a120347a );
 a365a <=( a120332a  and  a120317a );
 a366a <=( a120302a  and  a120287a );
 a367a <=( a120272a  and  a120257a );
 a368a <=( a120242a  and  a120227a );
 a369a <=( a120212a  and  a120197a );
 a370a <=( a120182a  and  a120167a );
 a371a <=( a120152a  and  a120137a );
 a372a <=( a120122a  and  a120107a );
 a373a <=( a120092a  and  a120077a );
 a374a <=( a120062a  and  a120047a );
 a375a <=( a120032a  and  a120017a );
 a376a <=( a120002a  and  a119987a );
 a377a <=( a119972a  and  a119957a );
 a378a <=( a119942a  and  a119927a );
 a379a <=( a119912a  and  a119897a );
 a380a <=( a119882a  and  a119867a );
 a381a <=( a119852a  and  a119837a );
 a382a <=( a119822a  and  a119807a );
 a383a <=( a119792a  and  a119777a );
 a384a <=( a119762a  and  a119747a );
 a385a <=( a119732a  and  a119717a );
 a386a <=( a119702a  and  a119687a );
 a387a <=( a119672a  and  a119657a );
 a388a <=( a119642a  and  a119627a );
 a389a <=( a119612a  and  a119597a );
 a390a <=( a119582a  and  a119567a );
 a391a <=( a119552a  and  a119537a );
 a392a <=( a119522a  and  a119507a );
 a393a <=( a119492a  and  a119477a );
 a394a <=( a119462a  and  a119447a );
 a395a <=( a119432a  and  a119417a );
 a396a <=( a119402a  and  a119387a );
 a397a <=( a119372a  and  a119357a );
 a398a <=( a119342a  and  a119327a );
 a399a <=( a119312a  and  a119297a );
 a400a <=( a119282a  and  a119267a );
 a401a <=( a119252a  and  a119237a );
 a402a <=( a119222a  and  a119207a );
 a403a <=( a119192a  and  a119177a );
 a404a <=( a119162a  and  a119147a );
 a405a <=( a119132a  and  a119117a );
 a406a <=( a119102a  and  a119087a );
 a407a <=( a119072a  and  a119057a );
 a408a <=( a119042a  and  a119027a );
 a409a <=( a119012a  and  a118997a );
 a410a <=( a118982a  and  a118967a );
 a411a <=( a118952a  and  a118937a );
 a412a <=( a118922a  and  a118907a );
 a413a <=( a118892a  and  a118877a );
 a414a <=( a118862a  and  a118847a );
 a415a <=( a118832a  and  a118817a );
 a416a <=( a118802a  and  a118787a );
 a417a <=( a118772a  and  a118757a );
 a418a <=( a118742a  and  a118727a );
 a419a <=( a118712a  and  a118697a );
 a420a <=( a118682a  and  a118667a );
 a421a <=( a118652a  and  a118637a );
 a422a <=( a118622a  and  a118607a );
 a423a <=( a118592a  and  a118577a );
 a424a <=( a118562a  and  a118547a );
 a425a <=( a118532a  and  a118517a );
 a426a <=( a118502a  and  a118487a );
 a427a <=( a118472a  and  a118457a );
 a428a <=( a118442a  and  a118427a );
 a429a <=( a118412a  and  a118397a );
 a430a <=( a118382a  and  a118367a );
 a431a <=( a118352a  and  a118337a );
 a432a <=( a118322a  and  a118307a );
 a433a <=( a118292a  and  a118277a );
 a434a <=( a118262a  and  a118247a );
 a435a <=( a118232a  and  a118217a );
 a436a <=( a118202a  and  a118187a );
 a437a <=( a118172a  and  a118157a );
 a438a <=( a118142a  and  a118127a );
 a439a <=( a118112a  and  a118097a );
 a440a <=( a118082a  and  a118067a );
 a441a <=( a118052a  and  a118037a );
 a442a <=( a118022a  and  a118007a );
 a443a <=( a117992a  and  a117977a );
 a444a <=( a117962a  and  a117947a );
 a445a <=( a117932a  and  a117917a );
 a446a <=( a117902a  and  a117887a );
 a447a <=( a117872a  and  a117857a );
 a448a <=( a117842a  and  a117827a );
 a449a <=( a117812a  and  a117797a );
 a450a <=( a117782a  and  a117767a );
 a451a <=( a117752a  and  a117737a );
 a452a <=( a117722a  and  a117707a );
 a453a <=( a117692a  and  a117677a );
 a454a <=( a117662a  and  a117647a );
 a455a <=( a117632a  and  a117617a );
 a456a <=( a117602a  and  a117587a );
 a457a <=( a117572a  and  a117557a );
 a458a <=( a117542a  and  a117527a );
 a459a <=( a117512a  and  a117497a );
 a460a <=( a117482a  and  a117467a );
 a461a <=( a117452a  and  a117437a );
 a462a <=( a117422a  and  a117407a );
 a463a <=( a117392a  and  a117377a );
 a464a <=( a117362a  and  a117347a );
 a465a <=( a117332a  and  a117317a );
 a466a <=( a117302a  and  a117287a );
 a467a <=( a117272a  and  a117257a );
 a468a <=( a117242a  and  a117227a );
 a469a <=( a117212a  and  a117197a );
 a470a <=( a117182a  and  a117167a );
 a471a <=( a117152a  and  a117137a );
 a472a <=( a117122a  and  a117107a );
 a473a <=( a117092a  and  a117077a );
 a474a <=( a117062a  and  a117047a );
 a475a <=( a117032a  and  a117017a );
 a476a <=( a117002a  and  a116987a );
 a477a <=( a116972a  and  a116957a );
 a478a <=( a116942a  and  a116927a );
 a479a <=( a116912a  and  a116897a );
 a480a <=( a116882a  and  a116867a );
 a481a <=( a116852a  and  a116837a );
 a482a <=( a116824a  and  a116809a );
 a483a <=( a116796a  and  a116781a );
 a484a <=( a116768a  and  a116753a );
 a485a <=( a116740a  and  a116725a );
 a486a <=( a116712a  and  a116697a );
 a487a <=( a116684a  and  a116669a );
 a488a <=( a116656a  and  a116641a );
 a489a <=( a116628a  and  a116613a );
 a490a <=( a116600a  and  a116585a );
 a491a <=( a116572a  and  a116557a );
 a492a <=( a116544a  and  a116529a );
 a493a <=( a116516a  and  a116501a );
 a494a <=( a116488a  and  a116473a );
 a495a <=( a116460a  and  a116445a );
 a496a <=( a116432a  and  a116417a );
 a497a <=( a116404a  and  a116389a );
 a498a <=( a116376a  and  a116361a );
 a499a <=( a116348a  and  a116333a );
 a500a <=( a116320a  and  a116305a );
 a501a <=( a116292a  and  a116277a );
 a502a <=( a116264a  and  a116249a );
 a503a <=( a116236a  and  a116221a );
 a504a <=( a116208a  and  a116193a );
 a505a <=( a116180a  and  a116165a );
 a506a <=( a116152a  and  a116137a );
 a507a <=( a116124a  and  a116109a );
 a508a <=( a116096a  and  a116081a );
 a509a <=( a116068a  and  a116053a );
 a510a <=( a116040a  and  a116025a );
 a511a <=( a116012a  and  a115997a );
 a512a <=( a115984a  and  a115969a );
 a513a <=( a115956a  and  a115941a );
 a514a <=( a115928a  and  a115913a );
 a515a <=( a115900a  and  a115885a );
 a516a <=( a115872a  and  a115857a );
 a517a <=( a115844a  and  a115829a );
 a518a <=( a115816a  and  a115801a );
 a519a <=( a115788a  and  a115773a );
 a520a <=( a115760a  and  a115745a );
 a521a <=( a115732a  and  a115717a );
 a522a <=( a115704a  and  a115689a );
 a523a <=( a115676a  and  a115661a );
 a524a <=( a115648a  and  a115633a );
 a525a <=( a115620a  and  a115605a );
 a526a <=( a115592a  and  a115577a );
 a527a <=( a115564a  and  a115549a );
 a528a <=( a115536a  and  a115521a );
 a529a <=( a115508a  and  a115493a );
 a530a <=( a115480a  and  a115465a );
 a531a <=( a115452a  and  a115437a );
 a532a <=( a115424a  and  a115409a );
 a533a <=( a115396a  and  a115381a );
 a534a <=( a115368a  and  a115353a );
 a535a <=( a115340a  and  a115325a );
 a536a <=( a115312a  and  a115297a );
 a537a <=( a115284a  and  a115269a );
 a538a <=( a115256a  and  a115241a );
 a539a <=( a115228a  and  a115213a );
 a540a <=( a115200a  and  a115185a );
 a541a <=( a115172a  and  a115157a );
 a542a <=( a115144a  and  a115129a );
 a543a <=( a115116a  and  a115101a );
 a544a <=( a115088a  and  a115073a );
 a545a <=( a115060a  and  a115045a );
 a546a <=( a115032a  and  a115017a );
 a547a <=( a115004a  and  a114989a );
 a548a <=( a114976a  and  a114961a );
 a549a <=( a114948a  and  a114933a );
 a550a <=( a114920a  and  a114905a );
 a551a <=( a114892a  and  a114877a );
 a552a <=( a114864a  and  a114849a );
 a553a <=( a114836a  and  a114821a );
 a554a <=( a114808a  and  a114793a );
 a555a <=( a114780a  and  a114765a );
 a556a <=( a114752a  and  a114737a );
 a557a <=( a114724a  and  a114709a );
 a558a <=( a114696a  and  a114681a );
 a559a <=( a114668a  and  a114653a );
 a560a <=( a114640a  and  a114625a );
 a561a <=( a114612a  and  a114597a );
 a562a <=( a114584a  and  a114569a );
 a563a <=( a114556a  and  a114541a );
 a564a <=( a114528a  and  a114513a );
 a565a <=( a114500a  and  a114485a );
 a566a <=( a114472a  and  a114457a );
 a567a <=( a114444a  and  a114429a );
 a568a <=( a114416a  and  a114401a );
 a569a <=( a114388a  and  a114373a );
 a570a <=( a114360a  and  a114345a );
 a571a <=( a114332a  and  a114317a );
 a572a <=( a114304a  and  a114289a );
 a573a <=( a114276a  and  a114261a );
 a574a <=( a114248a  and  a114233a );
 a575a <=( a114220a  and  a114205a );
 a576a <=( a114192a  and  a114177a );
 a577a <=( a114164a  and  a114149a );
 a578a <=( a114136a  and  a114121a );
 a579a <=( a114108a  and  a114093a );
 a580a <=( a114080a  and  a114065a );
 a581a <=( a114052a  and  a114037a );
 a582a <=( a114024a  and  a114009a );
 a583a <=( a113996a  and  a113981a );
 a584a <=( a113968a  and  a113953a );
 a585a <=( a113940a  and  a113925a );
 a586a <=( a113912a  and  a113897a );
 a587a <=( a113884a  and  a113869a );
 a588a <=( a113856a  and  a113841a );
 a589a <=( a113828a  and  a113813a );
 a590a <=( a113800a  and  a113785a );
 a591a <=( a113772a  and  a113757a );
 a592a <=( a113744a  and  a113729a );
 a593a <=( a113716a  and  a113701a );
 a594a <=( a113688a  and  a113673a );
 a595a <=( a113660a  and  a113645a );
 a596a <=( a113632a  and  a113617a );
 a597a <=( a113604a  and  a113589a );
 a598a <=( a113576a  and  a113561a );
 a599a <=( a113548a  and  a113533a );
 a600a <=( a113520a  and  a113505a );
 a601a <=( a113492a  and  a113477a );
 a602a <=( a113464a  and  a113449a );
 a603a <=( a113436a  and  a113421a );
 a604a <=( a113408a  and  a113393a );
 a605a <=( a113380a  and  a113365a );
 a606a <=( a113352a  and  a113337a );
 a607a <=( a113324a  and  a113309a );
 a608a <=( a113296a  and  a113281a );
 a609a <=( a113268a  and  a113253a );
 a610a <=( a113240a  and  a113225a );
 a611a <=( a113212a  and  a113197a );
 a612a <=( a113184a  and  a113169a );
 a613a <=( a113156a  and  a113141a );
 a614a <=( a113128a  and  a113113a );
 a615a <=( a113100a  and  a113085a );
 a616a <=( a113072a  and  a113057a );
 a617a <=( a113044a  and  a113029a );
 a618a <=( a113016a  and  a113001a );
 a619a <=( a112988a  and  a112973a );
 a620a <=( a112960a  and  a112945a );
 a621a <=( a112932a  and  a112917a );
 a622a <=( a112904a  and  a112889a );
 a623a <=( a112876a  and  a112861a );
 a624a <=( a112848a  and  a112833a );
 a625a <=( a112820a  and  a112805a );
 a626a <=( a112792a  and  a112777a );
 a627a <=( a112764a  and  a112749a );
 a628a <=( a112736a  and  a112721a );
 a629a <=( a112708a  and  a112693a );
 a630a <=( a112680a  and  a112665a );
 a631a <=( a112652a  and  a112637a );
 a632a <=( a112624a  and  a112609a );
 a633a <=( a112596a  and  a112581a );
 a634a <=( a112568a  and  a112553a );
 a635a <=( a112540a  and  a112525a );
 a636a <=( a112512a  and  a112497a );
 a637a <=( a112484a  and  a112469a );
 a638a <=( a112456a  and  a112441a );
 a639a <=( a112428a  and  a112413a );
 a640a <=( a112400a  and  a112385a );
 a641a <=( a112372a  and  a112357a );
 a642a <=( a112344a  and  a112329a );
 a643a <=( a112316a  and  a112301a );
 a644a <=( a112288a  and  a112273a );
 a645a <=( a112260a  and  a112245a );
 a646a <=( a112232a  and  a112217a );
 a647a <=( a112204a  and  a112189a );
 a648a <=( a112176a  and  a112161a );
 a649a <=( a112148a  and  a112133a );
 a650a <=( a112120a  and  a112105a );
 a651a <=( a112092a  and  a112077a );
 a652a <=( a112064a  and  a112049a );
 a653a <=( a112036a  and  a112021a );
 a654a <=( a112008a  and  a111993a );
 a655a <=( a111980a  and  a111965a );
 a656a <=( a111952a  and  a111937a );
 a657a <=( a111924a  and  a111909a );
 a658a <=( a111896a  and  a111881a );
 a659a <=( a111868a  and  a111853a );
 a660a <=( a111840a  and  a111825a );
 a661a <=( a111812a  and  a111797a );
 a662a <=( a111784a  and  a111769a );
 a663a <=( a111756a  and  a111741a );
 a664a <=( a111728a  and  a111713a );
 a665a <=( a111700a  and  a111685a );
 a666a <=( a111672a  and  a111657a );
 a667a <=( a111644a  and  a111629a );
 a668a <=( a111616a  and  a111601a );
 a669a <=( a111588a  and  a111573a );
 a670a <=( a111560a  and  a111545a );
 a671a <=( a111532a  and  a111517a );
 a672a <=( a111504a  and  a111489a );
 a673a <=( a111476a  and  a111461a );
 a674a <=( a111448a  and  a111433a );
 a675a <=( a111420a  and  a111405a );
 a676a <=( a111392a  and  a111377a );
 a677a <=( a111364a  and  a111349a );
 a678a <=( a111336a  and  a111321a );
 a679a <=( a111308a  and  a111293a );
 a680a <=( a111280a  and  a111265a );
 a681a <=( a111252a  and  a111237a );
 a682a <=( a111224a  and  a111209a );
 a683a <=( a111196a  and  a111181a );
 a684a <=( a111168a  and  a111153a );
 a685a <=( a111140a  and  a111125a );
 a686a <=( a111112a  and  a111097a );
 a687a <=( a111084a  and  a111069a );
 a688a <=( a111056a  and  a111041a );
 a689a <=( a111028a  and  a111013a );
 a690a <=( a111000a  and  a110985a );
 a691a <=( a110972a  and  a110957a );
 a692a <=( a110944a  and  a110929a );
 a693a <=( a110916a  and  a110901a );
 a694a <=( a110888a  and  a110873a );
 a695a <=( a110860a  and  a110845a );
 a696a <=( a110832a  and  a110817a );
 a697a <=( a110804a  and  a110789a );
 a698a <=( a110776a  and  a110761a );
 a699a <=( a110748a  and  a110733a );
 a700a <=( a110720a  and  a110705a );
 a701a <=( a110692a  and  a110677a );
 a702a <=( a110664a  and  a110649a );
 a703a <=( a110636a  and  a110621a );
 a704a <=( a110608a  and  a110593a );
 a705a <=( a110580a  and  a110565a );
 a706a <=( a110552a  and  a110537a );
 a707a <=( a110524a  and  a110509a );
 a708a <=( a110496a  and  a110481a );
 a709a <=( a110468a  and  a110453a );
 a710a <=( a110440a  and  a110425a );
 a711a <=( a110412a  and  a110397a );
 a712a <=( a110384a  and  a110369a );
 a713a <=( a110356a  and  a110341a );
 a714a <=( a110328a  and  a110313a );
 a715a <=( a110300a  and  a110285a );
 a716a <=( a110272a  and  a110257a );
 a717a <=( a110244a  and  a110229a );
 a718a <=( a110216a  and  a110201a );
 a719a <=( a110188a  and  a110173a );
 a720a <=( a110160a  and  a110145a );
 a721a <=( a110132a  and  a110117a );
 a722a <=( a110104a  and  a110089a );
 a723a <=( a110076a  and  a110061a );
 a724a <=( a110048a  and  a110033a );
 a725a <=( a110020a  and  a110005a );
 a726a <=( a109992a  and  a109977a );
 a727a <=( a109964a  and  a109949a );
 a728a <=( a109936a  and  a109921a );
 a729a <=( a109908a  and  a109893a );
 a730a <=( a109880a  and  a109865a );
 a731a <=( a109852a  and  a109837a );
 a732a <=( a109824a  and  a109809a );
 a733a <=( a109796a  and  a109781a );
 a734a <=( a109768a  and  a109753a );
 a735a <=( a109740a  and  a109725a );
 a736a <=( a109712a  and  a109697a );
 a737a <=( a109684a  and  a109669a );
 a738a <=( a109656a  and  a109641a );
 a739a <=( a109628a  and  a109613a );
 a740a <=( a109600a  and  a109585a );
 a741a <=( a109572a  and  a109557a );
 a742a <=( a109544a  and  a109529a );
 a743a <=( a109516a  and  a109501a );
 a744a <=( a109488a  and  a109473a );
 a745a <=( a109460a  and  a109445a );
 a746a <=( a109432a  and  a109417a );
 a747a <=( a109404a  and  a109389a );
 a748a <=( a109376a  and  a109361a );
 a749a <=( a109348a  and  a109333a );
 a750a <=( a109320a  and  a109305a );
 a751a <=( a109292a  and  a109277a );
 a752a <=( a109264a  and  a109249a );
 a753a <=( a109236a  and  a109221a );
 a754a <=( a109208a  and  a109193a );
 a755a <=( a109180a  and  a109165a );
 a756a <=( a109152a  and  a109137a );
 a757a <=( a109124a  and  a109109a );
 a758a <=( a109096a  and  a109081a );
 a759a <=( a109068a  and  a109053a );
 a760a <=( a109040a  and  a109025a );
 a761a <=( a109012a  and  a108997a );
 a762a <=( a108984a  and  a108969a );
 a763a <=( a108956a  and  a108941a );
 a764a <=( a108928a  and  a108913a );
 a765a <=( a108900a  and  a108885a );
 a766a <=( a108872a  and  a108857a );
 a767a <=( a108844a  and  a108829a );
 a768a <=( a108816a  and  a108801a );
 a769a <=( a108788a  and  a108773a );
 a770a <=( a108760a  and  a108745a );
 a771a <=( a108732a  and  a108717a );
 a772a <=( a108704a  and  a108689a );
 a773a <=( a108676a  and  a108661a );
 a774a <=( a108648a  and  a108633a );
 a775a <=( a108620a  and  a108605a );
 a776a <=( a108592a  and  a108577a );
 a777a <=( a108564a  and  a108549a );
 a778a <=( a108536a  and  a108521a );
 a779a <=( a108508a  and  a108493a );
 a780a <=( a108480a  and  a108465a );
 a781a <=( a108452a  and  a108437a );
 a782a <=( a108424a  and  a108409a );
 a783a <=( a108396a  and  a108381a );
 a784a <=( a108368a  and  a108353a );
 a785a <=( a108340a  and  a108325a );
 a786a <=( a108312a  and  a108297a );
 a787a <=( a108284a  and  a108269a );
 a788a <=( a108256a  and  a108241a );
 a789a <=( a108228a  and  a108213a );
 a790a <=( a108200a  and  a108185a );
 a791a <=( a108172a  and  a108157a );
 a792a <=( a108144a  and  a108129a );
 a793a <=( a108116a  and  a108101a );
 a794a <=( a108088a  and  a108073a );
 a795a <=( a108060a  and  a108045a );
 a796a <=( a108032a  and  a108017a );
 a797a <=( a108004a  and  a107989a );
 a798a <=( a107976a  and  a107961a );
 a799a <=( a107948a  and  a107933a );
 a800a <=( a107920a  and  a107905a );
 a801a <=( a107892a  and  a107877a );
 a802a <=( a107864a  and  a107849a );
 a803a <=( a107836a  and  a107821a );
 a804a <=( a107808a  and  a107793a );
 a805a <=( a107780a  and  a107765a );
 a806a <=( a107752a  and  a107737a );
 a807a <=( a107724a  and  a107709a );
 a808a <=( a107696a  and  a107681a );
 a809a <=( a107668a  and  a107653a );
 a810a <=( a107640a  and  a107625a );
 a811a <=( a107612a  and  a107597a );
 a812a <=( a107584a  and  a107569a );
 a813a <=( a107556a  and  a107541a );
 a814a <=( a107528a  and  a107513a );
 a815a <=( a107500a  and  a107485a );
 a816a <=( a107472a  and  a107457a );
 a817a <=( a107444a  and  a107429a );
 a818a <=( a107416a  and  a107401a );
 a819a <=( a107388a  and  a107373a );
 a820a <=( a107360a  and  a107345a );
 a821a <=( a107332a  and  a107317a );
 a822a <=( a107304a  and  a107289a );
 a823a <=( a107276a  and  a107261a );
 a824a <=( a107248a  and  a107233a );
 a825a <=( a107220a  and  a107205a );
 a826a <=( a107192a  and  a107177a );
 a827a <=( a107164a  and  a107149a );
 a828a <=( a107136a  and  a107121a );
 a829a <=( a107108a  and  a107093a );
 a830a <=( a107080a  and  a107065a );
 a831a <=( a107052a  and  a107037a );
 a832a <=( a107024a  and  a107009a );
 a833a <=( a106996a  and  a106981a );
 a834a <=( a106968a  and  a106953a );
 a835a <=( a106940a  and  a106925a );
 a836a <=( a106912a  and  a106897a );
 a837a <=( a106884a  and  a106869a );
 a838a <=( a106856a  and  a106841a );
 a839a <=( a106828a  and  a106813a );
 a840a <=( a106800a  and  a106785a );
 a841a <=( a106772a  and  a106757a );
 a842a <=( a106744a  and  a106729a );
 a843a <=( a106716a  and  a106701a );
 a844a <=( a106688a  and  a106673a );
 a845a <=( a106660a  and  a106645a );
 a846a <=( a106632a  and  a106617a );
 a847a <=( a106604a  and  a106589a );
 a848a <=( a106576a  and  a106561a );
 a849a <=( a106548a  and  a106533a );
 a850a <=( a106520a  and  a106505a );
 a851a <=( a106492a  and  a106477a );
 a852a <=( a106464a  and  a106449a );
 a853a <=( a106436a  and  a106421a );
 a854a <=( a106408a  and  a106393a );
 a855a <=( a106380a  and  a106365a );
 a856a <=( a106352a  and  a106337a );
 a857a <=( a106324a  and  a106309a );
 a858a <=( a106296a  and  a106281a );
 a859a <=( a106268a  and  a106253a );
 a860a <=( a106240a  and  a106225a );
 a861a <=( a106212a  and  a106197a );
 a862a <=( a106184a  and  a106169a );
 a863a <=( a106156a  and  a106141a );
 a864a <=( a106128a  and  a106113a );
 a865a <=( a106100a  and  a106085a );
 a866a <=( a106072a  and  a106057a );
 a867a <=( a106044a  and  a106029a );
 a868a <=( a106016a  and  a106001a );
 a869a <=( a105988a  and  a105973a );
 a870a <=( a105960a  and  a105945a );
 a871a <=( a105932a  and  a105917a );
 a872a <=( a105904a  and  a105889a );
 a873a <=( a105876a  and  a105861a );
 a874a <=( a105848a  and  a105833a );
 a875a <=( a105820a  and  a105805a );
 a876a <=( a105792a  and  a105777a );
 a877a <=( a105764a  and  a105749a );
 a878a <=( a105736a  and  a105721a );
 a879a <=( a105708a  and  a105693a );
 a880a <=( a105680a  and  a105665a );
 a881a <=( a105652a  and  a105637a );
 a882a <=( a105624a  and  a105609a );
 a883a <=( a105596a  and  a105581a );
 a884a <=( a105568a  and  a105553a );
 a885a <=( a105540a  and  a105525a );
 a886a <=( a105512a  and  a105497a );
 a887a <=( a105484a  and  a105469a );
 a888a <=( a105456a  and  a105441a );
 a889a <=( a105428a  and  a105413a );
 a890a <=( a105400a  and  a105385a );
 a891a <=( a105372a  and  a105357a );
 a892a <=( a105344a  and  a105329a );
 a893a <=( a105316a  and  a105301a );
 a894a <=( a105288a  and  a105273a );
 a895a <=( a105260a  and  a105245a );
 a896a <=( a105232a  and  a105217a );
 a897a <=( a105204a  and  a105189a );
 a898a <=( a105176a  and  a105161a );
 a899a <=( a105148a  and  a105133a );
 a900a <=( a105120a  and  a105105a );
 a901a <=( a105092a  and  a105077a );
 a902a <=( a105064a  and  a105049a );
 a903a <=( a105036a  and  a105021a );
 a904a <=( a105008a  and  a104993a );
 a905a <=( a104980a  and  a104965a );
 a906a <=( a104952a  and  a104937a );
 a907a <=( a104924a  and  a104909a );
 a908a <=( a104896a  and  a104881a );
 a909a <=( a104868a  and  a104853a );
 a910a <=( a104840a  and  a104825a );
 a911a <=( a104812a  and  a104797a );
 a912a <=( a104784a  and  a104769a );
 a913a <=( a104756a  and  a104741a );
 a914a <=( a104728a  and  a104713a );
 a915a <=( a104700a  and  a104685a );
 a916a <=( a104672a  and  a104657a );
 a917a <=( a104644a  and  a104629a );
 a918a <=( a104616a  and  a104601a );
 a919a <=( a104588a  and  a104573a );
 a920a <=( a104560a  and  a104545a );
 a921a <=( a104532a  and  a104517a );
 a922a <=( a104504a  and  a104489a );
 a923a <=( a104476a  and  a104461a );
 a924a <=( a104448a  and  a104433a );
 a925a <=( a104420a  and  a104405a );
 a926a <=( a104392a  and  a104377a );
 a927a <=( a104364a  and  a104349a );
 a928a <=( a104336a  and  a104321a );
 a929a <=( a104308a  and  a104293a );
 a930a <=( a104280a  and  a104265a );
 a931a <=( a104252a  and  a104237a );
 a932a <=( a104224a  and  a104209a );
 a933a <=( a104196a  and  a104181a );
 a934a <=( a104168a  and  a104153a );
 a935a <=( a104140a  and  a104125a );
 a936a <=( a104112a  and  a104097a );
 a937a <=( a104084a  and  a104069a );
 a938a <=( a104056a  and  a104041a );
 a939a <=( a104028a  and  a104013a );
 a940a <=( a104000a  and  a103985a );
 a941a <=( a103972a  and  a103957a );
 a942a <=( a103944a  and  a103929a );
 a943a <=( a103916a  and  a103901a );
 a944a <=( a103888a  and  a103873a );
 a945a <=( a103860a  and  a103845a );
 a946a <=( a103832a  and  a103817a );
 a947a <=( a103804a  and  a103789a );
 a948a <=( a103776a  and  a103761a );
 a949a <=( a103748a  and  a103733a );
 a950a <=( a103720a  and  a103705a );
 a951a <=( a103692a  and  a103677a );
 a952a <=( a103664a  and  a103649a );
 a953a <=( a103636a  and  a103621a );
 a954a <=( a103608a  and  a103593a );
 a955a <=( a103580a  and  a103565a );
 a956a <=( a103552a  and  a103537a );
 a957a <=( a103524a  and  a103509a );
 a958a <=( a103496a  and  a103481a );
 a959a <=( a103468a  and  a103453a );
 a960a <=( a103440a  and  a103425a );
 a961a <=( a103412a  and  a103397a );
 a962a <=( a103384a  and  a103369a );
 a963a <=( a103356a  and  a103341a );
 a964a <=( a103328a  and  a103313a );
 a965a <=( a103300a  and  a103285a );
 a966a <=( a103272a  and  a103257a );
 a967a <=( a103244a  and  a103229a );
 a968a <=( a103216a  and  a103201a );
 a969a <=( a103188a  and  a103173a );
 a970a <=( a103160a  and  a103145a );
 a971a <=( a103132a  and  a103117a );
 a972a <=( a103104a  and  a103089a );
 a973a <=( a103076a  and  a103061a );
 a974a <=( a103048a  and  a103033a );
 a975a <=( a103020a  and  a103005a );
 a976a <=( a102992a  and  a102977a );
 a977a <=( a102964a  and  a102951a );
 a978a <=( a102938a  and  a102925a );
 a979a <=( a102912a  and  a102899a );
 a980a <=( a102886a  and  a102873a );
 a981a <=( a102860a  and  a102847a );
 a982a <=( a102834a  and  a102821a );
 a983a <=( a102808a  and  a102795a );
 a984a <=( a102782a  and  a102769a );
 a985a <=( a102756a  and  a102743a );
 a986a <=( a102730a  and  a102717a );
 a987a <=( a102704a  and  a102691a );
 a988a <=( a102678a  and  a102665a );
 a989a <=( a102652a  and  a102639a );
 a990a <=( a102626a  and  a102613a );
 a991a <=( a102600a  and  a102587a );
 a992a <=( a102574a  and  a102561a );
 a993a <=( a102548a  and  a102535a );
 a994a <=( a102522a  and  a102509a );
 a995a <=( a102496a  and  a102483a );
 a996a <=( a102470a  and  a102457a );
 a997a <=( a102444a  and  a102431a );
 a998a <=( a102418a  and  a102405a );
 a999a <=( a102392a  and  a102379a );
 a1000a <=( a102366a  and  a102353a );
 a1001a <=( a102340a  and  a102327a );
 a1002a <=( a102314a  and  a102301a );
 a1003a <=( a102288a  and  a102275a );
 a1004a <=( a102262a  and  a102249a );
 a1005a <=( a102236a  and  a102223a );
 a1006a <=( a102210a  and  a102197a );
 a1007a <=( a102184a  and  a102171a );
 a1008a <=( a102158a  and  a102145a );
 a1009a <=( a102132a  and  a102119a );
 a1010a <=( a102106a  and  a102093a );
 a1011a <=( a102080a  and  a102067a );
 a1012a <=( a102054a  and  a102041a );
 a1013a <=( a102028a  and  a102015a );
 a1014a <=( a102002a  and  a101989a );
 a1015a <=( a101976a  and  a101963a );
 a1016a <=( a101950a  and  a101937a );
 a1017a <=( a101924a  and  a101911a );
 a1018a <=( a101898a  and  a101885a );
 a1019a <=( a101872a  and  a101859a );
 a1020a <=( a101846a  and  a101833a );
 a1021a <=( a101820a  and  a101807a );
 a1022a <=( a101794a  and  a101781a );
 a1023a <=( a101768a  and  a101755a );
 a1024a <=( a101742a  and  a101729a );
 a1025a <=( a101716a  and  a101703a );
 a1026a <=( a101690a  and  a101677a );
 a1027a <=( a101664a  and  a101651a );
 a1028a <=( a101638a  and  a101625a );
 a1029a <=( a101612a  and  a101599a );
 a1030a <=( a101586a  and  a101573a );
 a1031a <=( a101560a  and  a101547a );
 a1032a <=( a101534a  and  a101521a );
 a1033a <=( a101508a  and  a101495a );
 a1034a <=( a101482a  and  a101469a );
 a1035a <=( a101456a  and  a101443a );
 a1036a <=( a101430a  and  a101417a );
 a1037a <=( a101404a  and  a101391a );
 a1038a <=( a101378a  and  a101365a );
 a1039a <=( a101352a  and  a101339a );
 a1040a <=( a101326a  and  a101313a );
 a1041a <=( a101300a  and  a101287a );
 a1042a <=( a101274a  and  a101261a );
 a1043a <=( a101248a  and  a101235a );
 a1044a <=( a101222a  and  a101209a );
 a1045a <=( a101196a  and  a101183a );
 a1046a <=( a101170a  and  a101157a );
 a1047a <=( a101144a  and  a101131a );
 a1048a <=( a101118a  and  a101105a );
 a1049a <=( a101092a  and  a101079a );
 a1050a <=( a101066a  and  a101053a );
 a1051a <=( a101040a  and  a101027a );
 a1052a <=( a101014a  and  a101001a );
 a1053a <=( a100988a  and  a100975a );
 a1054a <=( a100962a  and  a100949a );
 a1055a <=( a100936a  and  a100923a );
 a1056a <=( a100910a  and  a100897a );
 a1057a <=( a100884a  and  a100871a );
 a1058a <=( a100858a  and  a100845a );
 a1059a <=( a100832a  and  a100819a );
 a1060a <=( a100806a  and  a100793a );
 a1061a <=( a100780a  and  a100767a );
 a1062a <=( a100754a  and  a100741a );
 a1063a <=( a100728a  and  a100715a );
 a1064a <=( a100702a  and  a100689a );
 a1065a <=( a100676a  and  a100663a );
 a1066a <=( a100650a  and  a100637a );
 a1067a <=( a100624a  and  a100611a );
 a1068a <=( a100598a  and  a100585a );
 a1069a <=( a100572a  and  a100559a );
 a1070a <=( a100546a  and  a100533a );
 a1071a <=( a100520a  and  a100507a );
 a1072a <=( a100494a  and  a100481a );
 a1073a <=( a100468a  and  a100455a );
 a1074a <=( a100442a  and  a100429a );
 a1075a <=( a100416a  and  a100403a );
 a1076a <=( a100390a  and  a100377a );
 a1077a <=( a100364a  and  a100351a );
 a1078a <=( a100338a  and  a100325a );
 a1079a <=( a100312a  and  a100299a );
 a1080a <=( a100286a  and  a100273a );
 a1081a <=( a100260a  and  a100247a );
 a1082a <=( a100234a  and  a100221a );
 a1083a <=( a100208a  and  a100195a );
 a1084a <=( a100182a  and  a100169a );
 a1085a <=( a100156a  and  a100143a );
 a1086a <=( a100130a  and  a100117a );
 a1087a <=( a100104a  and  a100091a );
 a1088a <=( a100078a  and  a100065a );
 a1089a <=( a100052a  and  a100039a );
 a1090a <=( a100026a  and  a100013a );
 a1091a <=( a100000a  and  a99987a );
 a1092a <=( a99974a  and  a99961a );
 a1093a <=( a99948a  and  a99935a );
 a1094a <=( a99922a  and  a99909a );
 a1095a <=( a99896a  and  a99883a );
 a1096a <=( a99870a  and  a99857a );
 a1097a <=( a99844a  and  a99831a );
 a1098a <=( a99818a  and  a99805a );
 a1099a <=( a99792a  and  a99779a );
 a1100a <=( a99766a  and  a99753a );
 a1101a <=( a99740a  and  a99727a );
 a1102a <=( a99714a  and  a99701a );
 a1103a <=( a99688a  and  a99675a );
 a1104a <=( a99662a  and  a99649a );
 a1105a <=( a99636a  and  a99623a );
 a1106a <=( a99610a  and  a99597a );
 a1107a <=( a99584a  and  a99571a );
 a1108a <=( a99558a  and  a99545a );
 a1109a <=( a99532a  and  a99519a );
 a1110a <=( a99506a  and  a99493a );
 a1111a <=( a99480a  and  a99467a );
 a1112a <=( a99454a  and  a99441a );
 a1113a <=( a99428a  and  a99415a );
 a1114a <=( a99402a  and  a99389a );
 a1115a <=( a99376a  and  a99363a );
 a1116a <=( a99350a  and  a99337a );
 a1117a <=( a99324a  and  a99311a );
 a1118a <=( a99298a  and  a99285a );
 a1119a <=( a99272a  and  a99259a );
 a1120a <=( a99246a  and  a99233a );
 a1121a <=( a99220a  and  a99207a );
 a1122a <=( a99194a  and  a99181a );
 a1123a <=( a99168a  and  a99155a );
 a1124a <=( a99142a  and  a99129a );
 a1125a <=( a99116a  and  a99103a );
 a1126a <=( a99090a  and  a99077a );
 a1127a <=( a99064a  and  a99051a );
 a1128a <=( a99038a  and  a99025a );
 a1129a <=( a99012a  and  a98999a );
 a1130a <=( a98986a  and  a98973a );
 a1131a <=( a98960a  and  a98947a );
 a1132a <=( a98934a  and  a98921a );
 a1133a <=( a98908a  and  a98895a );
 a1134a <=( a98882a  and  a98869a );
 a1135a <=( a98856a  and  a98843a );
 a1136a <=( a98830a  and  a98817a );
 a1137a <=( a98804a  and  a98791a );
 a1138a <=( a98778a  and  a98765a );
 a1139a <=( a98752a  and  a98739a );
 a1140a <=( a98726a  and  a98713a );
 a1141a <=( a98700a  and  a98687a );
 a1142a <=( a98674a  and  a98661a );
 a1143a <=( a98648a  and  a98635a );
 a1144a <=( a98622a  and  a98609a );
 a1145a <=( a98596a  and  a98583a );
 a1146a <=( a98570a  and  a98557a );
 a1147a <=( a98544a  and  a98531a );
 a1148a <=( a98518a  and  a98505a );
 a1149a <=( a98492a  and  a98479a );
 a1150a <=( a98466a  and  a98453a );
 a1151a <=( a98440a  and  a98427a );
 a1152a <=( a98414a  and  a98401a );
 a1153a <=( a98388a  and  a98375a );
 a1154a <=( a98362a  and  a98349a );
 a1155a <=( a98336a  and  a98323a );
 a1156a <=( a98310a  and  a98297a );
 a1157a <=( a98284a  and  a98271a );
 a1158a <=( a98258a  and  a98245a );
 a1159a <=( a98232a  and  a98219a );
 a1160a <=( a98206a  and  a98193a );
 a1161a <=( a98180a  and  a98167a );
 a1162a <=( a98154a  and  a98141a );
 a1163a <=( a98128a  and  a98115a );
 a1164a <=( a98102a  and  a98089a );
 a1165a <=( a98076a  and  a98063a );
 a1166a <=( a98050a  and  a98037a );
 a1167a <=( a98024a  and  a98011a );
 a1168a <=( a97998a  and  a97985a );
 a1169a <=( a97972a  and  a97959a );
 a1170a <=( a97946a  and  a97933a );
 a1171a <=( a97920a  and  a97907a );
 a1172a <=( a97894a  and  a97881a );
 a1173a <=( a97868a  and  a97855a );
 a1174a <=( a97842a  and  a97829a );
 a1175a <=( a97816a  and  a97803a );
 a1176a <=( a97790a  and  a97777a );
 a1177a <=( a97764a  and  a97751a );
 a1178a <=( a97738a  and  a97725a );
 a1179a <=( a97712a  and  a97699a );
 a1180a <=( a97686a  and  a97673a );
 a1181a <=( a97660a  and  a97647a );
 a1182a <=( a97634a  and  a97621a );
 a1183a <=( a97608a  and  a97595a );
 a1184a <=( a97582a  and  a97569a );
 a1185a <=( a97556a  and  a97543a );
 a1186a <=( a97530a  and  a97517a );
 a1187a <=( a97504a  and  a97491a );
 a1188a <=( a97478a  and  a97465a );
 a1189a <=( a97452a  and  a97439a );
 a1190a <=( a97426a  and  a97413a );
 a1191a <=( a97400a  and  a97387a );
 a1192a <=( a97374a  and  a97361a );
 a1193a <=( a97348a  and  a97335a );
 a1194a <=( a97322a  and  a97309a );
 a1195a <=( a97296a  and  a97283a );
 a1196a <=( a97270a  and  a97257a );
 a1197a <=( a97244a  and  a97231a );
 a1198a <=( a97218a  and  a97205a );
 a1199a <=( a97192a  and  a97179a );
 a1200a <=( a97166a  and  a97153a );
 a1201a <=( a97140a  and  a97127a );
 a1202a <=( a97114a  and  a97101a );
 a1203a <=( a97088a  and  a97075a );
 a1204a <=( a97062a  and  a97049a );
 a1205a <=( a97036a  and  a97023a );
 a1206a <=( a97010a  and  a96997a );
 a1207a <=( a96984a  and  a96971a );
 a1208a <=( a96958a  and  a96945a );
 a1209a <=( a96932a  and  a96919a );
 a1210a <=( a96906a  and  a96893a );
 a1211a <=( a96880a  and  a96867a );
 a1212a <=( a96854a  and  a96841a );
 a1213a <=( a96828a  and  a96815a );
 a1214a <=( a96802a  and  a96789a );
 a1215a <=( a96776a  and  a96763a );
 a1216a <=( a96750a  and  a96737a );
 a1217a <=( a96724a  and  a96711a );
 a1218a <=( a96698a  and  a96685a );
 a1219a <=( a96672a  and  a96659a );
 a1220a <=( a96646a  and  a96633a );
 a1221a <=( a96620a  and  a96607a );
 a1222a <=( a96594a  and  a96581a );
 a1223a <=( a96568a  and  a96555a );
 a1224a <=( a96542a  and  a96529a );
 a1225a <=( a96516a  and  a96503a );
 a1226a <=( a96490a  and  a96477a );
 a1227a <=( a96464a  and  a96451a );
 a1228a <=( a96438a  and  a96425a );
 a1229a <=( a96412a  and  a96399a );
 a1230a <=( a96386a  and  a96373a );
 a1231a <=( a96360a  and  a96347a );
 a1232a <=( a96334a  and  a96321a );
 a1233a <=( a96308a  and  a96295a );
 a1234a <=( a96282a  and  a96269a );
 a1235a <=( a96256a  and  a96243a );
 a1236a <=( a96230a  and  a96217a );
 a1237a <=( a96204a  and  a96191a );
 a1238a <=( a96178a  and  a96165a );
 a1239a <=( a96152a  and  a96139a );
 a1240a <=( a96126a  and  a96113a );
 a1241a <=( a96100a  and  a96087a );
 a1242a <=( a96074a  and  a96061a );
 a1243a <=( a96048a  and  a96035a );
 a1244a <=( a96022a  and  a96009a );
 a1245a <=( a95996a  and  a95983a );
 a1246a <=( a95970a  and  a95957a );
 a1247a <=( a95944a  and  a95931a );
 a1248a <=( a95918a  and  a95905a );
 a1249a <=( a95892a  and  a95879a );
 a1250a <=( a95866a  and  a95853a );
 a1251a <=( a95840a  and  a95827a );
 a1252a <=( a95814a  and  a95801a );
 a1253a <=( a95788a  and  a95775a );
 a1254a <=( a95762a  and  a95749a );
 a1255a <=( a95736a  and  a95723a );
 a1256a <=( a95710a  and  a95697a );
 a1257a <=( a95684a  and  a95671a );
 a1258a <=( a95658a  and  a95645a );
 a1259a <=( a95632a  and  a95619a );
 a1260a <=( a95606a  and  a95593a );
 a1261a <=( a95580a  and  a95567a );
 a1262a <=( a95554a  and  a95541a );
 a1263a <=( a95528a  and  a95515a );
 a1264a <=( a95502a  and  a95489a );
 a1265a <=( a95476a  and  a95463a );
 a1266a <=( a95450a  and  a95437a );
 a1267a <=( a95424a  and  a95411a );
 a1268a <=( a95398a  and  a95385a );
 a1269a <=( a95372a  and  a95359a );
 a1270a <=( a95346a  and  a95333a );
 a1271a <=( a95320a  and  a95307a );
 a1272a <=( a95294a  and  a95281a );
 a1273a <=( a95268a  and  a95255a );
 a1274a <=( a95242a  and  a95229a );
 a1275a <=( a95216a  and  a95203a );
 a1276a <=( a95190a  and  a95177a );
 a1277a <=( a95164a  and  a95151a );
 a1278a <=( a95138a  and  a95125a );
 a1279a <=( a95112a  and  a95099a );
 a1280a <=( a95086a  and  a95073a );
 a1281a <=( a95060a  and  a95047a );
 a1282a <=( a95034a  and  a95021a );
 a1283a <=( a95008a  and  a94995a );
 a1284a <=( a94982a  and  a94969a );
 a1285a <=( a94956a  and  a94943a );
 a1286a <=( a94930a  and  a94917a );
 a1287a <=( a94904a  and  a94891a );
 a1288a <=( a94878a  and  a94865a );
 a1289a <=( a94852a  and  a94839a );
 a1290a <=( a94826a  and  a94813a );
 a1291a <=( a94800a  and  a94787a );
 a1292a <=( a94774a  and  a94761a );
 a1293a <=( a94748a  and  a94735a );
 a1294a <=( a94722a  and  a94709a );
 a1295a <=( a94696a  and  a94683a );
 a1296a <=( a94670a  and  a94657a );
 a1297a <=( a94644a  and  a94631a );
 a1298a <=( a94618a  and  a94605a );
 a1299a <=( a94592a  and  a94579a );
 a1300a <=( a94566a  and  a94553a );
 a1301a <=( a94540a  and  a94527a );
 a1302a <=( a94514a  and  a94501a );
 a1303a <=( a94488a  and  a94475a );
 a1304a <=( a94462a  and  a94449a );
 a1305a <=( a94436a  and  a94423a );
 a1306a <=( a94410a  and  a94397a );
 a1307a <=( a94384a  and  a94371a );
 a1308a <=( a94358a  and  a94345a );
 a1309a <=( a94332a  and  a94319a );
 a1310a <=( a94306a  and  a94293a );
 a1311a <=( a94280a  and  a94267a );
 a1312a <=( a94254a  and  a94241a );
 a1313a <=( a94228a  and  a94215a );
 a1314a <=( a94202a  and  a94189a );
 a1315a <=( a94176a  and  a94163a );
 a1316a <=( a94150a  and  a94137a );
 a1317a <=( a94124a  and  a94111a );
 a1318a <=( a94098a  and  a94085a );
 a1319a <=( a94072a  and  a94059a );
 a1320a <=( a94046a  and  a94033a );
 a1321a <=( a94020a  and  a94007a );
 a1322a <=( a93994a  and  a93981a );
 a1323a <=( a93968a  and  a93955a );
 a1324a <=( a93942a  and  a93929a );
 a1325a <=( a93916a  and  a93903a );
 a1326a <=( a93890a  and  a93877a );
 a1327a <=( a93864a  and  a93851a );
 a1328a <=( a93838a  and  a93825a );
 a1329a <=( a93812a  and  a93799a );
 a1330a <=( a93786a  and  a93773a );
 a1331a <=( a93760a  and  a93747a );
 a1332a <=( a93734a  and  a93721a );
 a1333a <=( a93708a  and  a93695a );
 a1334a <=( a93682a  and  a93669a );
 a1335a <=( a93656a  and  a93643a );
 a1336a <=( a93630a  and  a93617a );
 a1337a <=( a93604a  and  a93591a );
 a1338a <=( a93578a  and  a93565a );
 a1339a <=( a93552a  and  a93539a );
 a1340a <=( a93526a  and  a93513a );
 a1341a <=( a93500a  and  a93487a );
 a1342a <=( a93474a  and  a93461a );
 a1343a <=( a93448a  and  a93435a );
 a1344a <=( a93422a  and  a93409a );
 a1345a <=( a93396a  and  a93383a );
 a1346a <=( a93370a  and  a93357a );
 a1347a <=( a93344a  and  a93331a );
 a1348a <=( a93318a  and  a93305a );
 a1349a <=( a93292a  and  a93279a );
 a1350a <=( a93266a  and  a93253a );
 a1351a <=( a93240a  and  a93227a );
 a1352a <=( a93214a  and  a93201a );
 a1353a <=( a93188a  and  a93175a );
 a1354a <=( a93162a  and  a93149a );
 a1355a <=( a93136a  and  a93123a );
 a1356a <=( a93110a  and  a93097a );
 a1357a <=( a93084a  and  a93071a );
 a1358a <=( a93058a  and  a93045a );
 a1359a <=( a93032a  and  a93019a );
 a1360a <=( a93006a  and  a92993a );
 a1361a <=( a92980a  and  a92967a );
 a1362a <=( a92954a  and  a92941a );
 a1363a <=( a92928a  and  a92915a );
 a1364a <=( a92902a  and  a92889a );
 a1365a <=( a92876a  and  a92863a );
 a1366a <=( a92850a  and  a92837a );
 a1367a <=( a92824a  and  a92811a );
 a1368a <=( a92798a  and  a92785a );
 a1369a <=( a92772a  and  a92759a );
 a1370a <=( a92746a  and  a92733a );
 a1371a <=( a92720a  and  a92707a );
 a1372a <=( a92694a  and  a92681a );
 a1373a <=( a92668a  and  a92655a );
 a1374a <=( a92642a  and  a92629a );
 a1375a <=( a92616a  and  a92603a );
 a1376a <=( a92590a  and  a92577a );
 a1377a <=( a92564a  and  a92551a );
 a1378a <=( a92538a  and  a92525a );
 a1379a <=( a92512a  and  a92499a );
 a1380a <=( a92486a  and  a92473a );
 a1381a <=( a92460a  and  a92447a );
 a1382a <=( a92434a  and  a92421a );
 a1383a <=( a92408a  and  a92395a );
 a1384a <=( a92382a  and  a92369a );
 a1385a <=( a92356a  and  a92343a );
 a1386a <=( a92330a  and  a92317a );
 a1387a <=( a92304a  and  a92291a );
 a1388a <=( a92278a  and  a92265a );
 a1389a <=( a92252a  and  a92239a );
 a1390a <=( a92226a  and  a92213a );
 a1391a <=( a92200a  and  a92187a );
 a1392a <=( a92174a  and  a92161a );
 a1393a <=( a92148a  and  a92135a );
 a1394a <=( a92122a  and  a92109a );
 a1395a <=( a92096a  and  a92083a );
 a1396a <=( a92070a  and  a92057a );
 a1397a <=( a92044a  and  a92031a );
 a1398a <=( a92018a  and  a92005a );
 a1399a <=( a91992a  and  a91979a );
 a1400a <=( a91966a  and  a91953a );
 a1401a <=( a91940a  and  a91927a );
 a1402a <=( a91914a  and  a91901a );
 a1403a <=( a91888a  and  a91875a );
 a1404a <=( a91862a  and  a91849a );
 a1405a <=( a91836a  and  a91823a );
 a1406a <=( a91810a  and  a91797a );
 a1407a <=( a91784a  and  a91771a );
 a1408a <=( a91758a  and  a91745a );
 a1409a <=( a91732a  and  a91719a );
 a1410a <=( a91706a  and  a91693a );
 a1411a <=( a91680a  and  a91667a );
 a1412a <=( a91654a  and  a91641a );
 a1413a <=( a91628a  and  a91615a );
 a1414a <=( a91602a  and  a91589a );
 a1415a <=( a91576a  and  a91563a );
 a1416a <=( a91550a  and  a91537a );
 a1417a <=( a91524a  and  a91511a );
 a1418a <=( a91498a  and  a91485a );
 a1419a <=( a91472a  and  a91459a );
 a1420a <=( a91446a  and  a91433a );
 a1421a <=( a91420a  and  a91407a );
 a1422a <=( a91394a  and  a91381a );
 a1423a <=( a91368a  and  a91355a );
 a1424a <=( a91342a  and  a91329a );
 a1425a <=( a91316a  and  a91303a );
 a1426a <=( a91290a  and  a91277a );
 a1427a <=( a91264a  and  a91251a );
 a1428a <=( a91238a  and  a91225a );
 a1429a <=( a91212a  and  a91199a );
 a1430a <=( a91186a  and  a91173a );
 a1431a <=( a91160a  and  a91147a );
 a1432a <=( a91134a  and  a91121a );
 a1433a <=( a91108a  and  a91095a );
 a1434a <=( a91082a  and  a91069a );
 a1435a <=( a91056a  and  a91043a );
 a1436a <=( a91030a  and  a91017a );
 a1437a <=( a91004a  and  a90991a );
 a1438a <=( a90978a  and  a90965a );
 a1439a <=( a90952a  and  a90939a );
 a1440a <=( a90926a  and  a90913a );
 a1441a <=( a90900a  and  a90887a );
 a1442a <=( a90874a  and  a90861a );
 a1443a <=( a90848a  and  a90835a );
 a1444a <=( a90822a  and  a90809a );
 a1445a <=( a90796a  and  a90783a );
 a1446a <=( a90770a  and  a90757a );
 a1447a <=( a90744a  and  a90731a );
 a1448a <=( a90718a  and  a90705a );
 a1449a <=( a90692a  and  a90679a );
 a1450a <=( a90666a  and  a90653a );
 a1451a <=( a90640a  and  a90627a );
 a1452a <=( a90614a  and  a90601a );
 a1453a <=( a90588a  and  a90575a );
 a1454a <=( a90562a  and  a90549a );
 a1455a <=( a90536a  and  a90523a );
 a1456a <=( a90510a  and  a90497a );
 a1457a <=( a90484a  and  a90471a );
 a1458a <=( a90458a  and  a90445a );
 a1459a <=( a90432a  and  a90419a );
 a1460a <=( a90406a  and  a90393a );
 a1461a <=( a90380a  and  a90367a );
 a1462a <=( a90354a  and  a90341a );
 a1463a <=( a90328a  and  a90315a );
 a1464a <=( a90302a  and  a90289a );
 a1465a <=( a90276a  and  a90263a );
 a1466a <=( a90250a  and  a90237a );
 a1467a <=( a90224a  and  a90211a );
 a1468a <=( a90198a  and  a90185a );
 a1469a <=( a90172a  and  a90159a );
 a1470a <=( a90146a  and  a90133a );
 a1471a <=( a90120a  and  a90107a );
 a1472a <=( a90094a  and  a90081a );
 a1473a <=( a90068a  and  a90055a );
 a1474a <=( a90042a  and  a90029a );
 a1475a <=( a90016a  and  a90003a );
 a1476a <=( a89990a  and  a89977a );
 a1477a <=( a89964a  and  a89951a );
 a1478a <=( a89938a  and  a89925a );
 a1479a <=( a89912a  and  a89899a );
 a1480a <=( a89886a  and  a89873a );
 a1481a <=( a89860a  and  a89847a );
 a1482a <=( a89834a  and  a89821a );
 a1483a <=( a89808a  and  a89795a );
 a1484a <=( a89782a  and  a89769a );
 a1485a <=( a89756a  and  a89743a );
 a1486a <=( a89730a  and  a89717a );
 a1487a <=( a89704a  and  a89691a );
 a1488a <=( a89678a  and  a89665a );
 a1489a <=( a89652a  and  a89639a );
 a1490a <=( a89626a  and  a89613a );
 a1491a <=( a89600a  and  a89587a );
 a1492a <=( a89574a  and  a89561a );
 a1493a <=( a89548a  and  a89535a );
 a1494a <=( a89522a  and  a89509a );
 a1495a <=( a89496a  and  a89483a );
 a1496a <=( a89470a  and  a89457a );
 a1497a <=( a89444a  and  a89431a );
 a1498a <=( a89418a  and  a89405a );
 a1499a <=( a89392a  and  a89379a );
 a1500a <=( a89366a  and  a89353a );
 a1501a <=( a89340a  and  a89327a );
 a1502a <=( a89314a  and  a89301a );
 a1503a <=( a89288a  and  a89275a );
 a1504a <=( a89262a  and  a89249a );
 a1505a <=( a89236a  and  a89223a );
 a1506a <=( a89210a  and  a89197a );
 a1507a <=( a89184a  and  a89171a );
 a1508a <=( a89158a  and  a89145a );
 a1509a <=( a89132a  and  a89119a );
 a1510a <=( a89106a  and  a89093a );
 a1511a <=( a89080a  and  a89067a );
 a1512a <=( a89054a  and  a89041a );
 a1513a <=( a89028a  and  a89015a );
 a1514a <=( a89002a  and  a88989a );
 a1515a <=( a88976a  and  a88963a );
 a1516a <=( a88950a  and  a88937a );
 a1517a <=( a88924a  and  a88911a );
 a1518a <=( a88898a  and  a88885a );
 a1519a <=( a88872a  and  a88859a );
 a1520a <=( a88846a  and  a88833a );
 a1521a <=( a88820a  and  a88807a );
 a1522a <=( a88794a  and  a88781a );
 a1523a <=( a88768a  and  a88755a );
 a1524a <=( a88742a  and  a88729a );
 a1525a <=( a88716a  and  a88703a );
 a1526a <=( a88690a  and  a88677a );
 a1527a <=( a88664a  and  a88651a );
 a1528a <=( a88638a  and  a88625a );
 a1529a <=( a88612a  and  a88599a );
 a1530a <=( a88586a  and  a88573a );
 a1531a <=( a88560a  and  a88547a );
 a1532a <=( a88534a  and  a88521a );
 a1533a <=( a88508a  and  a88495a );
 a1534a <=( a88482a  and  a88469a );
 a1535a <=( a88456a  and  a88443a );
 a1536a <=( a88430a  and  a88417a );
 a1537a <=( a88404a  and  a88391a );
 a1538a <=( a88378a  and  a88365a );
 a1539a <=( a88352a  and  a88339a );
 a1540a <=( a88326a  and  a88313a );
 a1541a <=( a88300a  and  a88287a );
 a1542a <=( a88274a  and  a88261a );
 a1543a <=( a88248a  and  a88235a );
 a1544a <=( a88222a  and  a88209a );
 a1545a <=( a88196a  and  a88183a );
 a1546a <=( a88170a  and  a88157a );
 a1547a <=( a88144a  and  a88131a );
 a1548a <=( a88118a  and  a88105a );
 a1549a <=( a88092a  and  a88079a );
 a1550a <=( a88066a  and  a88053a );
 a1551a <=( a88040a  and  a88027a );
 a1552a <=( a88014a  and  a88001a );
 a1553a <=( a87988a  and  a87975a );
 a1554a <=( a87962a  and  a87949a );
 a1555a <=( a87936a  and  a87923a );
 a1556a <=( a87910a  and  a87897a );
 a1557a <=( a87884a  and  a87871a );
 a1558a <=( a87858a  and  a87845a );
 a1559a <=( a87832a  and  a87819a );
 a1560a <=( a87806a  and  a87793a );
 a1561a <=( a87780a  and  a87767a );
 a1562a <=( a87754a  and  a87741a );
 a1563a <=( a87728a  and  a87715a );
 a1564a <=( a87702a  and  a87689a );
 a1565a <=( a87676a  and  a87663a );
 a1566a <=( a87650a  and  a87637a );
 a1567a <=( a87624a  and  a87611a );
 a1568a <=( a87598a  and  a87585a );
 a1569a <=( a87572a  and  a87559a );
 a1570a <=( a87546a  and  a87533a );
 a1571a <=( a87520a  and  a87507a );
 a1572a <=( a87494a  and  a87481a );
 a1573a <=( a87468a  and  a87455a );
 a1574a <=( a87442a  and  a87429a );
 a1575a <=( a87416a  and  a87403a );
 a1576a <=( a87390a  and  a87377a );
 a1577a <=( a87364a  and  a87351a );
 a1578a <=( a87338a  and  a87325a );
 a1579a <=( a87312a  and  a87299a );
 a1580a <=( a87286a  and  a87273a );
 a1581a <=( a87260a  and  a87247a );
 a1582a <=( a87234a  and  a87221a );
 a1583a <=( a87208a  and  a87195a );
 a1584a <=( a87182a  and  a87169a );
 a1585a <=( a87156a  and  a87143a );
 a1586a <=( a87130a  and  a87117a );
 a1587a <=( a87104a  and  a87091a );
 a1588a <=( a87078a  and  a87065a );
 a1589a <=( a87052a  and  a87039a );
 a1590a <=( a87026a  and  a87013a );
 a1591a <=( a87000a  and  a86987a );
 a1592a <=( a86974a  and  a86961a );
 a1593a <=( a86948a  and  a86935a );
 a1594a <=( a86922a  and  a86909a );
 a1595a <=( a86896a  and  a86883a );
 a1596a <=( a86870a  and  a86857a );
 a1597a <=( a86844a  and  a86831a );
 a1598a <=( a86818a  and  a86805a );
 a1599a <=( a86792a  and  a86779a );
 a1600a <=( a86766a  and  a86753a );
 a1601a <=( a86740a  and  a86727a );
 a1602a <=( a86714a  and  a86701a );
 a1603a <=( a86688a  and  a86675a );
 a1604a <=( a86662a  and  a86649a );
 a1605a <=( a86636a  and  a86623a );
 a1606a <=( a86610a  and  a86597a );
 a1607a <=( a86584a  and  a86571a );
 a1608a <=( a86558a  and  a86545a );
 a1609a <=( a86532a  and  a86519a );
 a1610a <=( a86506a  and  a86493a );
 a1611a <=( a86480a  and  a86467a );
 a1612a <=( a86454a  and  a86441a );
 a1613a <=( a86428a  and  a86415a );
 a1614a <=( a86402a  and  a86389a );
 a1615a <=( a86376a  and  a86363a );
 a1616a <=( a86350a  and  a86337a );
 a1617a <=( a86324a  and  a86311a );
 a1618a <=( a86298a  and  a86285a );
 a1619a <=( a86272a  and  a86259a );
 a1620a <=( a86246a  and  a86233a );
 a1621a <=( a86220a  and  a86207a );
 a1622a <=( a86194a  and  a86181a );
 a1623a <=( a86168a  and  a86155a );
 a1624a <=( a86142a  and  a86129a );
 a1625a <=( a86116a  and  a86103a );
 a1626a <=( a86090a  and  a86077a );
 a1627a <=( a86064a  and  a86051a );
 a1628a <=( a86038a  and  a86025a );
 a1629a <=( a86012a  and  a85999a );
 a1630a <=( a85986a  and  a85973a );
 a1631a <=( a85960a  and  a85947a );
 a1632a <=( a85934a  and  a85921a );
 a1633a <=( a85908a  and  a85895a );
 a1634a <=( a85882a  and  a85869a );
 a1635a <=( a85856a  and  a85843a );
 a1636a <=( a85830a  and  a85817a );
 a1637a <=( a85804a  and  a85791a );
 a1638a <=( a85778a  and  a85765a );
 a1639a <=( a85752a  and  a85739a );
 a1640a <=( a85726a  and  a85713a );
 a1641a <=( a85700a  and  a85687a );
 a1642a <=( a85674a  and  a85661a );
 a1643a <=( a85648a  and  a85635a );
 a1644a <=( a85622a  and  a85609a );
 a1645a <=( a85596a  and  a85583a );
 a1646a <=( a85570a  and  a85557a );
 a1647a <=( a85544a  and  a85531a );
 a1648a <=( a85518a  and  a85505a );
 a1649a <=( a85492a  and  a85479a );
 a1650a <=( a85466a  and  a85453a );
 a1651a <=( a85440a  and  a85427a );
 a1652a <=( a85414a  and  a85401a );
 a1653a <=( a85388a  and  a85375a );
 a1654a <=( a85362a  and  a85349a );
 a1655a <=( a85336a  and  a85323a );
 a1656a <=( a85310a  and  a85297a );
 a1657a <=( a85284a  and  a85271a );
 a1658a <=( a85258a  and  a85245a );
 a1659a <=( a85232a  and  a85219a );
 a1660a <=( a85206a  and  a85193a );
 a1661a <=( a85180a  and  a85167a );
 a1662a <=( a85154a  and  a85141a );
 a1663a <=( a85128a  and  a85115a );
 a1664a <=( a85102a  and  a85089a );
 a1665a <=( a85076a  and  a85063a );
 a1666a <=( a85050a  and  a85037a );
 a1667a <=( a85024a  and  a85011a );
 a1668a <=( a84998a  and  a84985a );
 a1669a <=( a84972a  and  a84959a );
 a1670a <=( a84946a  and  a84933a );
 a1671a <=( a84920a  and  a84907a );
 a1672a <=( a84894a  and  a84881a );
 a1673a <=( a84868a  and  a84855a );
 a1674a <=( a84842a  and  a84829a );
 a1675a <=( a84816a  and  a84803a );
 a1676a <=( a84790a  and  a84777a );
 a1677a <=( a84764a  and  a84751a );
 a1678a <=( a84738a  and  a84725a );
 a1679a <=( a84712a  and  a84699a );
 a1680a <=( a84686a  and  a84673a );
 a1681a <=( a84660a  and  a84647a );
 a1682a <=( a84634a  and  a84621a );
 a1683a <=( a84608a  and  a84595a );
 a1684a <=( a84582a  and  a84569a );
 a1685a <=( a84556a  and  a84543a );
 a1686a <=( a84530a  and  a84517a );
 a1687a <=( a84504a  and  a84491a );
 a1688a <=( a84478a  and  a84465a );
 a1689a <=( a84452a  and  a84439a );
 a1690a <=( a84426a  and  a84413a );
 a1691a <=( a84400a  and  a84387a );
 a1692a <=( a84374a  and  a84361a );
 a1693a <=( a84348a  and  a84335a );
 a1694a <=( a84322a  and  a84309a );
 a1695a <=( a84296a  and  a84283a );
 a1696a <=( a84270a  and  a84257a );
 a1697a <=( a84244a  and  a84231a );
 a1698a <=( a84218a  and  a84205a );
 a1699a <=( a84192a  and  a84179a );
 a1700a <=( a84166a  and  a84153a );
 a1701a <=( a84140a  and  a84127a );
 a1702a <=( a84114a  and  a84101a );
 a1703a <=( a84088a  and  a84075a );
 a1704a <=( a84062a  and  a84049a );
 a1705a <=( a84036a  and  a84023a );
 a1706a <=( a84010a  and  a83997a );
 a1707a <=( a83984a  and  a83971a );
 a1708a <=( a83958a  and  a83945a );
 a1709a <=( a83932a  and  a83919a );
 a1710a <=( a83906a  and  a83893a );
 a1711a <=( a83880a  and  a83867a );
 a1712a <=( a83854a  and  a83841a );
 a1713a <=( a83828a  and  a83815a );
 a1714a <=( a83802a  and  a83789a );
 a1715a <=( a83776a  and  a83763a );
 a1716a <=( a83750a  and  a83737a );
 a1717a <=( a83724a  and  a83711a );
 a1718a <=( a83698a  and  a83685a );
 a1719a <=( a83672a  and  a83659a );
 a1720a <=( a83646a  and  a83633a );
 a1721a <=( a83620a  and  a83607a );
 a1722a <=( a83594a  and  a83581a );
 a1723a <=( a83568a  and  a83555a );
 a1724a <=( a83542a  and  a83529a );
 a1725a <=( a83516a  and  a83503a );
 a1726a <=( a83490a  and  a83477a );
 a1727a <=( a83464a  and  a83451a );
 a1728a <=( a83438a  and  a83425a );
 a1729a <=( a83412a  and  a83399a );
 a1730a <=( a83386a  and  a83373a );
 a1731a <=( a83360a  and  a83347a );
 a1732a <=( a83334a  and  a83321a );
 a1733a <=( a83308a  and  a83295a );
 a1734a <=( a83282a  and  a83269a );
 a1735a <=( a83256a  and  a83243a );
 a1736a <=( a83230a  and  a83217a );
 a1737a <=( a83204a  and  a83191a );
 a1738a <=( a83178a  and  a83165a );
 a1739a <=( a83152a  and  a83139a );
 a1740a <=( a83126a  and  a83113a );
 a1741a <=( a83100a  and  a83087a );
 a1742a <=( a83074a  and  a83061a );
 a1743a <=( a83048a  and  a83035a );
 a1744a <=( a83022a  and  a83009a );
 a1745a <=( a82996a  and  a82983a );
 a1746a <=( a82970a  and  a82957a );
 a1747a <=( a82944a  and  a82931a );
 a1748a <=( a82918a  and  a82905a );
 a1749a <=( a82892a  and  a82879a );
 a1750a <=( a82866a  and  a82853a );
 a1751a <=( a82840a  and  a82827a );
 a1752a <=( a82814a  and  a82801a );
 a1753a <=( a82788a  and  a82775a );
 a1754a <=( a82762a  and  a82749a );
 a1755a <=( a82736a  and  a82723a );
 a1756a <=( a82710a  and  a82697a );
 a1757a <=( a82684a  and  a82671a );
 a1758a <=( a82658a  and  a82645a );
 a1759a <=( a82632a  and  a82619a );
 a1760a <=( a82606a  and  a82593a );
 a1761a <=( a82580a  and  a82567a );
 a1762a <=( a82554a  and  a82541a );
 a1763a <=( a82528a  and  a82515a );
 a1764a <=( a82502a  and  a82489a );
 a1765a <=( a82476a  and  a82463a );
 a1766a <=( a82450a  and  a82437a );
 a1767a <=( a82424a  and  a82411a );
 a1768a <=( a82398a  and  a82385a );
 a1769a <=( a82372a  and  a82359a );
 a1770a <=( a82346a  and  a82333a );
 a1771a <=( a82320a  and  a82307a );
 a1772a <=( a82294a  and  a82281a );
 a1773a <=( a82268a  and  a82255a );
 a1774a <=( a82242a  and  a82229a );
 a1775a <=( a82216a  and  a82203a );
 a1776a <=( a82190a  and  a82177a );
 a1777a <=( a82164a  and  a82151a );
 a1778a <=( a82138a  and  a82125a );
 a1779a <=( a82112a  and  a82099a );
 a1780a <=( a82086a  and  a82073a );
 a1781a <=( a82060a  and  a82047a );
 a1782a <=( a82034a  and  a82021a );
 a1783a <=( a82008a  and  a81995a );
 a1784a <=( a81982a  and  a81969a );
 a1785a <=( a81956a  and  a81943a );
 a1786a <=( a81930a  and  a81917a );
 a1787a <=( a81904a  and  a81891a );
 a1788a <=( a81878a  and  a81865a );
 a1789a <=( a81852a  and  a81839a );
 a1790a <=( a81826a  and  a81813a );
 a1791a <=( a81800a  and  a81787a );
 a1792a <=( a81774a  and  a81761a );
 a1793a <=( a81748a  and  a81735a );
 a1794a <=( a81722a  and  a81709a );
 a1795a <=( a81696a  and  a81683a );
 a1796a <=( a81670a  and  a81657a );
 a1797a <=( a81644a  and  a81631a );
 a1798a <=( a81618a  and  a81605a );
 a1799a <=( a81592a  and  a81579a );
 a1800a <=( a81566a  and  a81553a );
 a1801a <=( a81540a  and  a81527a );
 a1802a <=( a81514a  and  a81501a );
 a1803a <=( a81488a  and  a81475a );
 a1804a <=( a81462a  and  a81449a );
 a1805a <=( a81436a  and  a81423a );
 a1806a <=( a81410a  and  a81397a );
 a1807a <=( a81384a  and  a81371a );
 a1808a <=( a81358a  and  a81345a );
 a1809a <=( a81332a  and  a81319a );
 a1810a <=( a81306a  and  a81293a );
 a1811a <=( a81280a  and  a81267a );
 a1812a <=( a81254a  and  a81241a );
 a1813a <=( a81228a  and  a81215a );
 a1814a <=( a81202a  and  a81189a );
 a1815a <=( a81176a  and  a81163a );
 a1816a <=( a81150a  and  a81137a );
 a1817a <=( a81124a  and  a81111a );
 a1818a <=( a81098a  and  a81085a );
 a1819a <=( a81072a  and  a81059a );
 a1820a <=( a81046a  and  a81033a );
 a1821a <=( a81020a  and  a81007a );
 a1822a <=( a80994a  and  a80981a );
 a1823a <=( a80968a  and  a80955a );
 a1824a <=( a80942a  and  a80929a );
 a1825a <=( a80916a  and  a80903a );
 a1826a <=( a80890a  and  a80877a );
 a1827a <=( a80864a  and  a80851a );
 a1828a <=( a80838a  and  a80825a );
 a1829a <=( a80812a  and  a80799a );
 a1830a <=( a80786a  and  a80773a );
 a1831a <=( a80760a  and  a80747a );
 a1832a <=( a80734a  and  a80721a );
 a1833a <=( a80708a  and  a80695a );
 a1834a <=( a80682a  and  a80669a );
 a1835a <=( a80656a  and  a80643a );
 a1836a <=( a80630a  and  a80617a );
 a1837a <=( a80604a  and  a80591a );
 a1838a <=( a80578a  and  a80565a );
 a1839a <=( a80552a  and  a80539a );
 a1840a <=( a80526a  and  a80513a );
 a1841a <=( a80500a  and  a80487a );
 a1842a <=( a80474a  and  a80461a );
 a1843a <=( a80448a  and  a80435a );
 a1844a <=( a80422a  and  a80409a );
 a1845a <=( a80396a  and  a80383a );
 a1846a <=( a80370a  and  a80357a );
 a1847a <=( a80344a  and  a80331a );
 a1848a <=( a80318a  and  a80305a );
 a1849a <=( a80292a  and  a80279a );
 a1850a <=( a80266a  and  a80253a );
 a1851a <=( a80240a  and  a80227a );
 a1852a <=( a80214a  and  a80201a );
 a1853a <=( a80188a  and  a80175a );
 a1854a <=( a80162a  and  a80149a );
 a1855a <=( a80136a  and  a80123a );
 a1856a <=( a80110a  and  a80097a );
 a1857a <=( a80084a  and  a80071a );
 a1858a <=( a80058a  and  a80045a );
 a1859a <=( a80032a  and  a80019a );
 a1860a <=( a80006a  and  a79993a );
 a1861a <=( a79980a  and  a79967a );
 a1862a <=( a79954a  and  a79941a );
 a1863a <=( a79928a  and  a79915a );
 a1864a <=( a79902a  and  a79889a );
 a1865a <=( a79876a  and  a79863a );
 a1866a <=( a79850a  and  a79837a );
 a1867a <=( a79824a  and  a79811a );
 a1868a <=( a79798a  and  a79785a );
 a1869a <=( a79772a  and  a79759a );
 a1870a <=( a79746a  and  a79733a );
 a1871a <=( a79720a  and  a79707a );
 a1872a <=( a79694a  and  a79681a );
 a1873a <=( a79668a  and  a79655a );
 a1874a <=( a79642a  and  a79629a );
 a1875a <=( a79616a  and  a79603a );
 a1876a <=( a79590a  and  a79577a );
 a1877a <=( a79564a  and  a79551a );
 a1878a <=( a79538a  and  a79525a );
 a1879a <=( a79512a  and  a79499a );
 a1880a <=( a79486a  and  a79473a );
 a1881a <=( a79460a  and  a79447a );
 a1882a <=( a79434a  and  a79421a );
 a1883a <=( a79408a  and  a79395a );
 a1884a <=( a79382a  and  a79369a );
 a1885a <=( a79356a  and  a79343a );
 a1886a <=( a79330a  and  a79317a );
 a1887a <=( a79304a  and  a79291a );
 a1888a <=( a79278a  and  a79265a );
 a1889a <=( a79252a  and  a79239a );
 a1890a <=( a79226a  and  a79213a );
 a1891a <=( a79200a  and  a79187a );
 a1892a <=( a79174a  and  a79161a );
 a1893a <=( a79148a  and  a79135a );
 a1894a <=( a79122a  and  a79109a );
 a1895a <=( a79096a  and  a79083a );
 a1896a <=( a79070a  and  a79057a );
 a1897a <=( a79044a  and  a79031a );
 a1898a <=( a79018a  and  a79005a );
 a1899a <=( a78992a  and  a78979a );
 a1900a <=( a78966a  and  a78953a );
 a1901a <=( a78940a  and  a78927a );
 a1902a <=( a78914a  and  a78901a );
 a1903a <=( a78888a  and  a78875a );
 a1904a <=( a78862a  and  a78849a );
 a1905a <=( a78836a  and  a78823a );
 a1906a <=( a78810a  and  a78797a );
 a1907a <=( a78784a  and  a78771a );
 a1908a <=( a78758a  and  a78745a );
 a1909a <=( a78732a  and  a78719a );
 a1910a <=( a78706a  and  a78693a );
 a1911a <=( a78680a  and  a78667a );
 a1912a <=( a78654a  and  a78641a );
 a1913a <=( a78628a  and  a78615a );
 a1914a <=( a78602a  and  a78589a );
 a1915a <=( a78576a  and  a78563a );
 a1916a <=( a78550a  and  a78537a );
 a1917a <=( a78524a  and  a78511a );
 a1918a <=( a78498a  and  a78485a );
 a1919a <=( a78472a  and  a78459a );
 a1920a <=( a78446a  and  a78433a );
 a1921a <=( a78420a  and  a78407a );
 a1922a <=( a78394a  and  a78381a );
 a1923a <=( a78368a  and  a78355a );
 a1924a <=( a78342a  and  a78329a );
 a1925a <=( a78316a  and  a78303a );
 a1926a <=( a78290a  and  a78277a );
 a1927a <=( a78264a  and  a78251a );
 a1928a <=( a78238a  and  a78225a );
 a1929a <=( a78212a  and  a78199a );
 a1930a <=( a78186a  and  a78173a );
 a1931a <=( a78160a  and  a78147a );
 a1932a <=( a78134a  and  a78121a );
 a1933a <=( a78108a  and  a78095a );
 a1934a <=( a78082a  and  a78069a );
 a1935a <=( a78056a  and  a78043a );
 a1936a <=( a78030a  and  a78017a );
 a1937a <=( a78004a  and  a77991a );
 a1938a <=( a77978a  and  a77965a );
 a1939a <=( a77952a  and  a77939a );
 a1940a <=( a77926a  and  a77913a );
 a1941a <=( a77900a  and  a77887a );
 a1942a <=( a77874a  and  a77861a );
 a1943a <=( a77848a  and  a77835a );
 a1944a <=( a77822a  and  a77809a );
 a1945a <=( a77796a  and  a77783a );
 a1946a <=( a77770a  and  a77757a );
 a1947a <=( a77744a  and  a77731a );
 a1948a <=( a77718a  and  a77705a );
 a1949a <=( a77692a  and  a77679a );
 a1950a <=( a77666a  and  a77653a );
 a1951a <=( a77640a  and  a77627a );
 a1952a <=( a77614a  and  a77601a );
 a1953a <=( a77588a  and  a77575a );
 a1954a <=( a77562a  and  a77549a );
 a1955a <=( a77536a  and  a77523a );
 a1956a <=( a77510a  and  a77497a );
 a1957a <=( a77484a  and  a77471a );
 a1958a <=( a77458a  and  a77445a );
 a1959a <=( a77432a  and  a77419a );
 a1960a <=( a77406a  and  a77393a );
 a1961a <=( a77380a  and  a77367a );
 a1962a <=( a77354a  and  a77341a );
 a1963a <=( a77328a  and  a77315a );
 a1964a <=( a77302a  and  a77289a );
 a1965a <=( a77276a  and  a77263a );
 a1966a <=( a77250a  and  a77237a );
 a1967a <=( a77224a  and  a77211a );
 a1968a <=( a77198a  and  a77185a );
 a1969a <=( a77172a  and  a77159a );
 a1970a <=( a77146a  and  a77133a );
 a1971a <=( a77120a  and  a77107a );
 a1972a <=( a77094a  and  a77081a );
 a1973a <=( a77068a  and  a77055a );
 a1974a <=( a77042a  and  a77029a );
 a1975a <=( a77016a  and  a77003a );
 a1976a <=( a76990a  and  a76977a );
 a1977a <=( a76964a  and  a76951a );
 a1978a <=( a76938a  and  a76925a );
 a1979a <=( a76912a  and  a76899a );
 a1980a <=( a76886a  and  a76873a );
 a1981a <=( a76860a  and  a76847a );
 a1982a <=( a76834a  and  a76821a );
 a1983a <=( a76808a  and  a76795a );
 a1984a <=( a76782a  and  a76769a );
 a1985a <=( a76756a  and  a76743a );
 a1986a <=( a76730a  and  a76717a );
 a1987a <=( a76704a  and  a76691a );
 a1988a <=( a76678a  and  a76665a );
 a1989a <=( a76652a  and  a76639a );
 a1990a <=( a76626a  and  a76613a );
 a1991a <=( a76600a  and  a76587a );
 a1992a <=( a76574a  and  a76561a );
 a1993a <=( a76548a  and  a76535a );
 a1994a <=( a76522a  and  a76509a );
 a1995a <=( a76496a  and  a76483a );
 a1996a <=( a76470a  and  a76457a );
 a1997a <=( a76444a  and  a76431a );
 a1998a <=( a76418a  and  a76405a );
 a1999a <=( a76392a  and  a76379a );
 a2000a <=( a76366a  and  a76353a );
 a2001a <=( a76340a  and  a76327a );
 a2002a <=( a76314a  and  a76301a );
 a2003a <=( a76288a  and  a76275a );
 a2004a <=( a76262a  and  a76249a );
 a2005a <=( a76236a  and  a76223a );
 a2006a <=( a76210a  and  a76197a );
 a2007a <=( a76184a  and  a76171a );
 a2008a <=( a76158a  and  a76145a );
 a2009a <=( a76132a  and  a76119a );
 a2010a <=( a76106a  and  a76093a );
 a2011a <=( a76080a  and  a76067a );
 a2012a <=( a76054a  and  a76041a );
 a2013a <=( a76028a  and  a76015a );
 a2014a <=( a76002a  and  a75989a );
 a2015a <=( a75976a  and  a75963a );
 a2016a <=( a75950a  and  a75937a );
 a2017a <=( a75924a  and  a75911a );
 a2018a <=( a75898a  and  a75885a );
 a2019a <=( a75872a  and  a75859a );
 a2020a <=( a75846a  and  a75833a );
 a2021a <=( a75820a  and  a75807a );
 a2022a <=( a75794a  and  a75781a );
 a2023a <=( a75768a  and  a75755a );
 a2024a <=( a75742a  and  a75729a );
 a2025a <=( a75716a  and  a75703a );
 a2026a <=( a75690a  and  a75677a );
 a2027a <=( a75664a  and  a75651a );
 a2028a <=( a75638a  and  a75625a );
 a2029a <=( a75612a  and  a75599a );
 a2030a <=( a75586a  and  a75573a );
 a2031a <=( a75560a  and  a75547a );
 a2032a <=( a75534a  and  a75521a );
 a2033a <=( a75508a  and  a75495a );
 a2034a <=( a75482a  and  a75469a );
 a2035a <=( a75456a  and  a75443a );
 a2036a <=( a75430a  and  a75417a );
 a2037a <=( a75404a  and  a75391a );
 a2038a <=( a75378a  and  a75365a );
 a2039a <=( a75352a  and  a75339a );
 a2040a <=( a75326a  and  a75313a );
 a2041a <=( a75300a  and  a75287a );
 a2042a <=( a75274a  and  a75261a );
 a2043a <=( a75248a  and  a75235a );
 a2044a <=( a75222a  and  a75209a );
 a2045a <=( a75196a  and  a75183a );
 a2046a <=( a75170a  and  a75157a );
 a2047a <=( a75144a  and  a75131a );
 a2048a <=( a75118a  and  a75105a );
 a2049a <=( a75092a  and  a75079a );
 a2050a <=( a75066a  and  a75053a );
 a2051a <=( a75040a  and  a75027a );
 a2052a <=( a75014a  and  a75001a );
 a2053a <=( a74988a  and  a74975a );
 a2054a <=( a74962a  and  a74949a );
 a2055a <=( a74936a  and  a74923a );
 a2056a <=( a74910a  and  a74897a );
 a2057a <=( a74884a  and  a74871a );
 a2058a <=( a74858a  and  a74845a );
 a2059a <=( a74832a  and  a74819a );
 a2060a <=( a74806a  and  a74793a );
 a2061a <=( a74780a  and  a74767a );
 a2062a <=( a74754a  and  a74741a );
 a2063a <=( a74728a  and  a74715a );
 a2064a <=( a74702a  and  a74689a );
 a2065a <=( a74676a  and  a74663a );
 a2066a <=( a74650a  and  a74637a );
 a2067a <=( a74624a  and  a74611a );
 a2068a <=( a74598a  and  a74585a );
 a2069a <=( a74572a  and  a74559a );
 a2070a <=( a74546a  and  a74533a );
 a2071a <=( a74520a  and  a74507a );
 a2072a <=( a74494a  and  a74481a );
 a2073a <=( a74468a  and  a74455a );
 a2074a <=( a74442a  and  a74429a );
 a2075a <=( a74416a  and  a74403a );
 a2076a <=( a74390a  and  a74377a );
 a2077a <=( a74364a  and  a74351a );
 a2078a <=( a74338a  and  a74325a );
 a2079a <=( a74312a  and  a74299a );
 a2080a <=( a74286a  and  a74273a );
 a2081a <=( a74260a  and  a74247a );
 a2082a <=( a74234a  and  a74221a );
 a2083a <=( a74208a  and  a74195a );
 a2084a <=( a74182a  and  a74169a );
 a2085a <=( a74156a  and  a74143a );
 a2086a <=( a74130a  and  a74117a );
 a2087a <=( a74104a  and  a74091a );
 a2088a <=( a74078a  and  a74065a );
 a2089a <=( a74052a  and  a74039a );
 a2090a <=( a74026a  and  a74013a );
 a2091a <=( a74000a  and  a73987a );
 a2092a <=( a73974a  and  a73961a );
 a2093a <=( a73948a  and  a73935a );
 a2094a <=( a73922a  and  a73909a );
 a2095a <=( a73896a  and  a73883a );
 a2096a <=( a73870a  and  a73857a );
 a2097a <=( a73844a  and  a73831a );
 a2098a <=( a73818a  and  a73805a );
 a2099a <=( a73792a  and  a73779a );
 a2100a <=( a73766a  and  a73753a );
 a2101a <=( a73740a  and  a73727a );
 a2102a <=( a73714a  and  a73701a );
 a2103a <=( a73688a  and  a73675a );
 a2104a <=( a73662a  and  a73649a );
 a2105a <=( a73636a  and  a73623a );
 a2106a <=( a73610a  and  a73597a );
 a2107a <=( a73584a  and  a73571a );
 a2108a <=( a73558a  and  a73545a );
 a2109a <=( a73532a  and  a73519a );
 a2110a <=( a73506a  and  a73493a );
 a2111a <=( a73480a  and  a73467a );
 a2112a <=( a73454a  and  a73441a );
 a2113a <=( a73428a  and  a73415a );
 a2114a <=( a73402a  and  a73389a );
 a2115a <=( a73376a  and  a73363a );
 a2116a <=( a73350a  and  a73337a );
 a2117a <=( a73324a  and  a73311a );
 a2118a <=( a73298a  and  a73285a );
 a2119a <=( a73272a  and  a73259a );
 a2120a <=( a73246a  and  a73233a );
 a2121a <=( a73220a  and  a73207a );
 a2122a <=( a73194a  and  a73181a );
 a2123a <=( a73168a  and  a73155a );
 a2124a <=( a73142a  and  a73129a );
 a2125a <=( a73116a  and  a73103a );
 a2126a <=( a73090a  and  a73077a );
 a2127a <=( a73064a  and  a73051a );
 a2128a <=( a73038a  and  a73025a );
 a2129a <=( a73012a  and  a72999a );
 a2130a <=( a72986a  and  a72973a );
 a2131a <=( a72960a  and  a72947a );
 a2132a <=( a72934a  and  a72921a );
 a2133a <=( a72908a  and  a72895a );
 a2134a <=( a72882a  and  a72869a );
 a2135a <=( a72856a  and  a72843a );
 a2136a <=( a72830a  and  a72817a );
 a2137a <=( a72804a  and  a72791a );
 a2138a <=( a72778a  and  a72765a );
 a2139a <=( a72752a  and  a72739a );
 a2140a <=( a72726a  and  a72713a );
 a2141a <=( a72700a  and  a72687a );
 a2142a <=( a72674a  and  a72661a );
 a2143a <=( a72648a  and  a72635a );
 a2144a <=( a72622a  and  a72609a );
 a2145a <=( a72596a  and  a72583a );
 a2146a <=( a72570a  and  a72557a );
 a2147a <=( a72544a  and  a72531a );
 a2148a <=( a72518a  and  a72505a );
 a2149a <=( a72492a  and  a72479a );
 a2150a <=( a72466a  and  a72453a );
 a2151a <=( a72440a  and  a72427a );
 a2152a <=( a72414a  and  a72401a );
 a2153a <=( a72388a  and  a72375a );
 a2154a <=( a72362a  and  a72349a );
 a2155a <=( a72336a  and  a72323a );
 a2156a <=( a72310a  and  a72297a );
 a2157a <=( a72284a  and  a72271a );
 a2158a <=( a72258a  and  a72245a );
 a2159a <=( a72232a  and  a72219a );
 a2160a <=( a72206a  and  a72193a );
 a2161a <=( a72180a  and  a72167a );
 a2162a <=( a72154a  and  a72141a );
 a2163a <=( a72128a  and  a72115a );
 a2164a <=( a72102a  and  a72089a );
 a2165a <=( a72076a  and  a72063a );
 a2166a <=( a72050a  and  a72037a );
 a2167a <=( a72024a  and  a72011a );
 a2168a <=( a71998a  and  a71985a );
 a2169a <=( a71972a  and  a71959a );
 a2170a <=( a71946a  and  a71933a );
 a2171a <=( a71920a  and  a71907a );
 a2172a <=( a71894a  and  a71881a );
 a2173a <=( a71868a  and  a71855a );
 a2174a <=( a71842a  and  a71829a );
 a2175a <=( a71816a  and  a71803a );
 a2176a <=( a71790a  and  a71777a );
 a2177a <=( a71764a  and  a71751a );
 a2178a <=( a71738a  and  a71725a );
 a2179a <=( a71712a  and  a71699a );
 a2180a <=( a71686a  and  a71673a );
 a2181a <=( a71660a  and  a71647a );
 a2182a <=( a71634a  and  a71621a );
 a2183a <=( a71608a  and  a71595a );
 a2184a <=( a71582a  and  a71569a );
 a2185a <=( a71556a  and  a71543a );
 a2186a <=( a71530a  and  a71517a );
 a2187a <=( a71504a  and  a71491a );
 a2188a <=( a71478a  and  a71465a );
 a2189a <=( a71452a  and  a71439a );
 a2190a <=( a71426a  and  a71413a );
 a2191a <=( a71400a  and  a71387a );
 a2192a <=( a71374a  and  a71361a );
 a2193a <=( a71348a  and  a71335a );
 a2194a <=( a71322a  and  a71309a );
 a2195a <=( a71296a  and  a71283a );
 a2196a <=( a71270a  and  a71257a );
 a2197a <=( a71244a  and  a71231a );
 a2198a <=( a71218a  and  a71205a );
 a2199a <=( a71192a  and  a71179a );
 a2200a <=( a71166a  and  a71153a );
 a2201a <=( a71140a  and  a71127a );
 a2202a <=( a71114a  and  a71101a );
 a2203a <=( a71088a  and  a71075a );
 a2204a <=( a71062a  and  a71049a );
 a2205a <=( a71036a  and  a71023a );
 a2206a <=( a71010a  and  a70997a );
 a2207a <=( a70984a  and  a70971a );
 a2208a <=( a70958a  and  a70945a );
 a2209a <=( a70932a  and  a70919a );
 a2210a <=( a70906a  and  a70893a );
 a2211a <=( a70880a  and  a70867a );
 a2212a <=( a70854a  and  a70841a );
 a2213a <=( a70828a  and  a70815a );
 a2214a <=( a70802a  and  a70789a );
 a2215a <=( a70776a  and  a70763a );
 a2216a <=( a70750a  and  a70737a );
 a2217a <=( a70724a  and  a70711a );
 a2218a <=( a70698a  and  a70685a );
 a2219a <=( a70672a  and  a70659a );
 a2220a <=( a70646a  and  a70633a );
 a2221a <=( a70620a  and  a70607a );
 a2222a <=( a70594a  and  a70581a );
 a2223a <=( a70568a  and  a70555a );
 a2224a <=( a70542a  and  a70529a );
 a2225a <=( a70516a  and  a70503a );
 a2226a <=( a70490a  and  a70477a );
 a2227a <=( a70464a  and  a70451a );
 a2228a <=( a70438a  and  a70425a );
 a2229a <=( a70412a  and  a70399a );
 a2230a <=( a70386a  and  a70373a );
 a2231a <=( a70360a  and  a70347a );
 a2232a <=( a70334a  and  a70321a );
 a2233a <=( a70308a  and  a70295a );
 a2234a <=( a70282a  and  a70269a );
 a2235a <=( a70256a  and  a70243a );
 a2236a <=( a70230a  and  a70217a );
 a2237a <=( a70204a  and  a70191a );
 a2238a <=( a70178a  and  a70165a );
 a2239a <=( a70152a  and  a70139a );
 a2240a <=( a70126a  and  a70113a );
 a2241a <=( a70100a  and  a70087a );
 a2242a <=( a70074a  and  a70061a );
 a2243a <=( a70048a  and  a70035a );
 a2244a <=( a70022a  and  a70009a );
 a2245a <=( a69996a  and  a69983a );
 a2246a <=( a69970a  and  a69957a );
 a2247a <=( a69944a  and  a69931a );
 a2248a <=( a69918a  and  a69905a );
 a2249a <=( a69892a  and  a69879a );
 a2250a <=( a69866a  and  a69853a );
 a2251a <=( a69840a  and  a69827a );
 a2252a <=( a69814a  and  a69801a );
 a2253a <=( a69788a  and  a69775a );
 a2254a <=( a69762a  and  a69749a );
 a2255a <=( a69736a  and  a69723a );
 a2256a <=( a69710a  and  a69697a );
 a2257a <=( a69684a  and  a69671a );
 a2258a <=( a69658a  and  a69645a );
 a2259a <=( a69632a  and  a69619a );
 a2260a <=( a69606a  and  a69593a );
 a2261a <=( a69580a  and  a69567a );
 a2262a <=( a69554a  and  a69541a );
 a2263a <=( a69528a  and  a69515a );
 a2264a <=( a69502a  and  a69489a );
 a2265a <=( a69476a  and  a69463a );
 a2266a <=( a69450a  and  a69437a );
 a2267a <=( a69424a  and  a69411a );
 a2268a <=( a69398a  and  a69385a );
 a2269a <=( a69372a  and  a69359a );
 a2270a <=( a69346a  and  a69333a );
 a2271a <=( a69320a  and  a69307a );
 a2272a <=( a69294a  and  a69281a );
 a2273a <=( a69268a  and  a69255a );
 a2274a <=( a69242a  and  a69229a );
 a2275a <=( a69216a  and  a69203a );
 a2276a <=( a69190a  and  a69177a );
 a2277a <=( a69164a  and  a69151a );
 a2278a <=( a69138a  and  a69125a );
 a2279a <=( a69112a  and  a69099a );
 a2280a <=( a69086a  and  a69073a );
 a2281a <=( a69060a  and  a69047a );
 a2282a <=( a69034a  and  a69021a );
 a2283a <=( a69008a  and  a68995a );
 a2284a <=( a68982a  and  a68969a );
 a2285a <=( a68956a  and  a68943a );
 a2286a <=( a68930a  and  a68917a );
 a2287a <=( a68904a  and  a68891a );
 a2288a <=( a68878a  and  a68865a );
 a2289a <=( a68852a  and  a68839a );
 a2290a <=( a68826a  and  a68813a );
 a2291a <=( a68800a  and  a68787a );
 a2292a <=( a68774a  and  a68761a );
 a2293a <=( a68748a  and  a68735a );
 a2294a <=( a68722a  and  a68709a );
 a2295a <=( a68696a  and  a68683a );
 a2296a <=( a68670a  and  a68657a );
 a2297a <=( a68644a  and  a68631a );
 a2298a <=( a68618a  and  a68605a );
 a2299a <=( a68592a  and  a68579a );
 a2300a <=( a68566a  and  a68553a );
 a2301a <=( a68540a  and  a68527a );
 a2302a <=( a68514a  and  a68501a );
 a2303a <=( a68488a  and  a68475a );
 a2304a <=( a68462a  and  a68449a );
 a2305a <=( a68436a  and  a68423a );
 a2306a <=( a68410a  and  a68397a );
 a2307a <=( a68384a  and  a68371a );
 a2308a <=( a68358a  and  a68345a );
 a2309a <=( a68332a  and  a68319a );
 a2310a <=( a68306a  and  a68293a );
 a2311a <=( a68280a  and  a68267a );
 a2312a <=( a68254a  and  a68241a );
 a2313a <=( a68228a  and  a68215a );
 a2314a <=( a68202a  and  a68189a );
 a2315a <=( a68176a  and  a68163a );
 a2316a <=( a68150a  and  a68137a );
 a2317a <=( a68124a  and  a68111a );
 a2318a <=( a68098a  and  a68085a );
 a2319a <=( a68072a  and  a68059a );
 a2320a <=( a68046a  and  a68033a );
 a2321a <=( a68020a  and  a68007a );
 a2322a <=( a67994a  and  a67981a );
 a2323a <=( a67968a  and  a67955a );
 a2324a <=( a67942a  and  a67929a );
 a2325a <=( a67916a  and  a67903a );
 a2326a <=( a67890a  and  a67877a );
 a2327a <=( a67864a  and  a67851a );
 a2328a <=( a67838a  and  a67825a );
 a2329a <=( a67812a  and  a67799a );
 a2330a <=( a67786a  and  a67773a );
 a2331a <=( a67760a  and  a67747a );
 a2332a <=( a67734a  and  a67721a );
 a2333a <=( a67708a  and  a67695a );
 a2334a <=( a67682a  and  a67669a );
 a2335a <=( a67656a  and  a67643a );
 a2336a <=( a67630a  and  a67617a );
 a2337a <=( a67604a  and  a67591a );
 a2338a <=( a67578a  and  a67565a );
 a2339a <=( a67552a  and  a67539a );
 a2340a <=( a67526a  and  a67513a );
 a2341a <=( a67500a  and  a67487a );
 a2342a <=( a67474a  and  a67461a );
 a2343a <=( a67448a  and  a67435a );
 a2344a <=( a67422a  and  a67409a );
 a2345a <=( a67396a  and  a67383a );
 a2346a <=( a67370a  and  a67357a );
 a2347a <=( a67344a  and  a67331a );
 a2348a <=( a67318a  and  a67305a );
 a2349a <=( a67292a  and  a67279a );
 a2350a <=( a67266a  and  a67253a );
 a2351a <=( a67240a  and  a67227a );
 a2352a <=( a67214a  and  a67201a );
 a2353a <=( a67188a  and  a67175a );
 a2354a <=( a67162a  and  a67149a );
 a2355a <=( a67136a  and  a67123a );
 a2356a <=( a67110a  and  a67097a );
 a2357a <=( a67084a  and  a67071a );
 a2358a <=( a67058a  and  a67045a );
 a2359a <=( a67032a  and  a67019a );
 a2360a <=( a67006a  and  a66993a );
 a2361a <=( a66980a  and  a66967a );
 a2362a <=( a66954a  and  a66941a );
 a2363a <=( a66928a  and  a66915a );
 a2364a <=( a66902a  and  a66889a );
 a2365a <=( a66876a  and  a66863a );
 a2366a <=( a66850a  and  a66837a );
 a2367a <=( a66824a  and  a66811a );
 a2368a <=( a66798a  and  a66785a );
 a2369a <=( a66772a  and  a66759a );
 a2370a <=( a66746a  and  a66733a );
 a2371a <=( a66720a  and  a66707a );
 a2372a <=( a66694a  and  a66681a );
 a2373a <=( a66668a  and  a66655a );
 a2374a <=( a66642a  and  a66629a );
 a2375a <=( a66616a  and  a66603a );
 a2376a <=( a66590a  and  a66577a );
 a2377a <=( a66564a  and  a66551a );
 a2378a <=( a66538a  and  a66525a );
 a2379a <=( a66512a  and  a66499a );
 a2380a <=( a66486a  and  a66473a );
 a2381a <=( a66460a  and  a66447a );
 a2382a <=( a66434a  and  a66421a );
 a2383a <=( a66408a  and  a66395a );
 a2384a <=( a66382a  and  a66369a );
 a2385a <=( a66356a  and  a66343a );
 a2386a <=( a66330a  and  a66317a );
 a2387a <=( a66304a  and  a66291a );
 a2388a <=( a66278a  and  a66265a );
 a2389a <=( a66252a  and  a66239a );
 a2390a <=( a66226a  and  a66213a );
 a2391a <=( a66200a  and  a66187a );
 a2392a <=( a66174a  and  a66161a );
 a2393a <=( a66148a  and  a66135a );
 a2394a <=( a66122a  and  a66109a );
 a2395a <=( a66096a  and  a66083a );
 a2396a <=( a66070a  and  a66057a );
 a2397a <=( a66044a  and  a66031a );
 a2398a <=( a66018a  and  a66005a );
 a2399a <=( a65992a  and  a65979a );
 a2400a <=( a65966a  and  a65953a );
 a2401a <=( a65940a  and  a65927a );
 a2402a <=( a65914a  and  a65901a );
 a2403a <=( a65888a  and  a65875a );
 a2404a <=( a65862a  and  a65849a );
 a2405a <=( a65836a  and  a65823a );
 a2406a <=( a65810a  and  a65797a );
 a2407a <=( a65784a  and  a65771a );
 a2408a <=( a65758a  and  a65745a );
 a2409a <=( a65732a  and  a65719a );
 a2410a <=( a65706a  and  a65693a );
 a2411a <=( a65680a  and  a65667a );
 a2412a <=( a65654a  and  a65641a );
 a2413a <=( a65628a  and  a65615a );
 a2414a <=( a65602a  and  a65589a );
 a2415a <=( a65576a  and  a65563a );
 a2416a <=( a65550a  and  a65537a );
 a2417a <=( a65524a  and  a65511a );
 a2418a <=( a65498a  and  a65485a );
 a2419a <=( a65472a  and  a65459a );
 a2420a <=( a65446a  and  a65433a );
 a2421a <=( a65420a  and  a65407a );
 a2422a <=( a65394a  and  a65381a );
 a2423a <=( a65368a  and  a65355a );
 a2424a <=( a65342a  and  a65329a );
 a2425a <=( a65316a  and  a65303a );
 a2426a <=( a65290a  and  a65277a );
 a2427a <=( a65264a  and  a65251a );
 a2428a <=( a65238a  and  a65225a );
 a2429a <=( a65212a  and  a65199a );
 a2430a <=( a65186a  and  a65173a );
 a2431a <=( a65160a  and  a65147a );
 a2432a <=( a65134a  and  a65121a );
 a2433a <=( a65108a  and  a65095a );
 a2434a <=( a65084a  and  a65071a );
 a2435a <=( a65060a  and  a65047a );
 a2436a <=( a65036a  and  a65023a );
 a2437a <=( a65012a  and  a64999a );
 a2438a <=( a64988a  and  a64975a );
 a2439a <=( a64964a  and  a64951a );
 a2440a <=( a64940a  and  a64927a );
 a2441a <=( a64916a  and  a64903a );
 a2442a <=( a64892a  and  a64879a );
 a2443a <=( a64868a  and  a64855a );
 a2444a <=( a64844a  and  a64831a );
 a2445a <=( a64820a  and  a64807a );
 a2446a <=( a64796a  and  a64783a );
 a2447a <=( a64772a  and  a64759a );
 a2448a <=( a64748a  and  a64735a );
 a2449a <=( a64724a  and  a64711a );
 a2450a <=( a64700a  and  a64687a );
 a2451a <=( a64676a  and  a64663a );
 a2452a <=( a64652a  and  a64639a );
 a2453a <=( a64628a  and  a64615a );
 a2454a <=( a64604a  and  a64591a );
 a2455a <=( a64580a  and  a64567a );
 a2456a <=( a64556a  and  a64543a );
 a2457a <=( a64532a  and  a64519a );
 a2458a <=( a64508a  and  a64495a );
 a2459a <=( a64484a  and  a64471a );
 a2460a <=( a64460a  and  a64447a );
 a2461a <=( a64436a  and  a64423a );
 a2462a <=( a64412a  and  a64399a );
 a2463a <=( a64388a  and  a64375a );
 a2464a <=( a64364a  and  a64351a );
 a2465a <=( a64340a  and  a64327a );
 a2466a <=( a64316a  and  a64303a );
 a2467a <=( a64292a  and  a64279a );
 a2468a <=( a64268a  and  a64255a );
 a2469a <=( a64244a  and  a64231a );
 a2470a <=( a64220a  and  a64207a );
 a2471a <=( a64196a  and  a64183a );
 a2472a <=( a64172a  and  a64159a );
 a2473a <=( a64148a  and  a64135a );
 a2474a <=( a64124a  and  a64111a );
 a2475a <=( a64100a  and  a64087a );
 a2476a <=( a64076a  and  a64063a );
 a2477a <=( a64052a  and  a64039a );
 a2478a <=( a64028a  and  a64015a );
 a2479a <=( a64004a  and  a63991a );
 a2480a <=( a63980a  and  a63967a );
 a2481a <=( a63956a  and  a63943a );
 a2482a <=( a63932a  and  a63919a );
 a2483a <=( a63908a  and  a63895a );
 a2484a <=( a63884a  and  a63871a );
 a2485a <=( a63860a  and  a63847a );
 a2486a <=( a63836a  and  a63823a );
 a2487a <=( a63812a  and  a63799a );
 a2488a <=( a63788a  and  a63775a );
 a2489a <=( a63764a  and  a63751a );
 a2490a <=( a63740a  and  a63727a );
 a2491a <=( a63716a  and  a63703a );
 a2492a <=( a63692a  and  a63679a );
 a2493a <=( a63668a  and  a63655a );
 a2494a <=( a63644a  and  a63631a );
 a2495a <=( a63620a  and  a63607a );
 a2496a <=( a63596a  and  a63583a );
 a2497a <=( a63572a  and  a63559a );
 a2498a <=( a63548a  and  a63535a );
 a2499a <=( a63524a  and  a63511a );
 a2500a <=( a63500a  and  a63487a );
 a2501a <=( a63476a  and  a63463a );
 a2502a <=( a63452a  and  a63439a );
 a2503a <=( a63428a  and  a63415a );
 a2504a <=( a63404a  and  a63391a );
 a2505a <=( a63380a  and  a63367a );
 a2506a <=( a63356a  and  a63343a );
 a2507a <=( a63332a  and  a63319a );
 a2508a <=( a63308a  and  a63295a );
 a2509a <=( a63284a  and  a63271a );
 a2510a <=( a63260a  and  a63247a );
 a2511a <=( a63236a  and  a63223a );
 a2512a <=( a63212a  and  a63199a );
 a2513a <=( a63188a  and  a63175a );
 a2514a <=( a63164a  and  a63151a );
 a2515a <=( a63140a  and  a63127a );
 a2516a <=( a63116a  and  a63103a );
 a2517a <=( a63092a  and  a63079a );
 a2518a <=( a63068a  and  a63055a );
 a2519a <=( a63044a  and  a63031a );
 a2520a <=( a63020a  and  a63007a );
 a2521a <=( a62996a  and  a62983a );
 a2522a <=( a62972a  and  a62959a );
 a2523a <=( a62948a  and  a62935a );
 a2524a <=( a62924a  and  a62911a );
 a2525a <=( a62900a  and  a62887a );
 a2526a <=( a62876a  and  a62863a );
 a2527a <=( a62852a  and  a62839a );
 a2528a <=( a62828a  and  a62815a );
 a2529a <=( a62804a  and  a62791a );
 a2530a <=( a62780a  and  a62767a );
 a2531a <=( a62756a  and  a62743a );
 a2532a <=( a62732a  and  a62719a );
 a2533a <=( a62708a  and  a62695a );
 a2534a <=( a62684a  and  a62671a );
 a2535a <=( a62660a  and  a62647a );
 a2536a <=( a62636a  and  a62623a );
 a2537a <=( a62612a  and  a62599a );
 a2538a <=( a62588a  and  a62575a );
 a2539a <=( a62564a  and  a62551a );
 a2540a <=( a62540a  and  a62527a );
 a2541a <=( a62516a  and  a62503a );
 a2542a <=( a62492a  and  a62479a );
 a2543a <=( a62468a  and  a62455a );
 a2544a <=( a62444a  and  a62431a );
 a2545a <=( a62420a  and  a62407a );
 a2546a <=( a62396a  and  a62383a );
 a2547a <=( a62372a  and  a62359a );
 a2548a <=( a62348a  and  a62335a );
 a2549a <=( a62324a  and  a62311a );
 a2550a <=( a62300a  and  a62287a );
 a2551a <=( a62276a  and  a62263a );
 a2552a <=( a62252a  and  a62239a );
 a2553a <=( a62228a  and  a62215a );
 a2554a <=( a62204a  and  a62191a );
 a2555a <=( a62180a  and  a62167a );
 a2556a <=( a62156a  and  a62143a );
 a2557a <=( a62132a  and  a62119a );
 a2558a <=( a62108a  and  a62095a );
 a2559a <=( a62084a  and  a62071a );
 a2560a <=( a62060a  and  a62047a );
 a2561a <=( a62036a  and  a62023a );
 a2562a <=( a62012a  and  a61999a );
 a2563a <=( a61988a  and  a61975a );
 a2564a <=( a61964a  and  a61951a );
 a2565a <=( a61940a  and  a61927a );
 a2566a <=( a61916a  and  a61903a );
 a2567a <=( a61892a  and  a61879a );
 a2568a <=( a61868a  and  a61855a );
 a2569a <=( a61844a  and  a61831a );
 a2570a <=( a61820a  and  a61807a );
 a2571a <=( a61796a  and  a61783a );
 a2572a <=( a61772a  and  a61759a );
 a2573a <=( a61748a  and  a61735a );
 a2574a <=( a61724a  and  a61711a );
 a2575a <=( a61700a  and  a61687a );
 a2576a <=( a61676a  and  a61663a );
 a2577a <=( a61652a  and  a61639a );
 a2578a <=( a61628a  and  a61615a );
 a2579a <=( a61604a  and  a61591a );
 a2580a <=( a61580a  and  a61567a );
 a2581a <=( a61556a  and  a61543a );
 a2582a <=( a61532a  and  a61519a );
 a2583a <=( a61508a  and  a61495a );
 a2584a <=( a61484a  and  a61471a );
 a2585a <=( a61460a  and  a61447a );
 a2586a <=( a61436a  and  a61423a );
 a2587a <=( a61412a  and  a61399a );
 a2588a <=( a61388a  and  a61375a );
 a2589a <=( a61364a  and  a61351a );
 a2590a <=( a61340a  and  a61327a );
 a2591a <=( a61316a  and  a61303a );
 a2592a <=( a61292a  and  a61279a );
 a2593a <=( a61268a  and  a61255a );
 a2594a <=( a61244a  and  a61231a );
 a2595a <=( a61220a  and  a61207a );
 a2596a <=( a61196a  and  a61183a );
 a2597a <=( a61172a  and  a61159a );
 a2598a <=( a61148a  and  a61135a );
 a2599a <=( a61124a  and  a61111a );
 a2600a <=( a61100a  and  a61087a );
 a2601a <=( a61076a  and  a61063a );
 a2602a <=( a61052a  and  a61039a );
 a2603a <=( a61028a  and  a61015a );
 a2604a <=( a61004a  and  a60991a );
 a2605a <=( a60980a  and  a60967a );
 a2606a <=( a60956a  and  a60943a );
 a2607a <=( a60932a  and  a60919a );
 a2608a <=( a60908a  and  a60895a );
 a2609a <=( a60884a  and  a60871a );
 a2610a <=( a60860a  and  a60847a );
 a2611a <=( a60836a  and  a60823a );
 a2612a <=( a60812a  and  a60799a );
 a2613a <=( a60788a  and  a60775a );
 a2614a <=( a60764a  and  a60751a );
 a2615a <=( a60740a  and  a60727a );
 a2616a <=( a60716a  and  a60703a );
 a2617a <=( a60692a  and  a60679a );
 a2618a <=( a60668a  and  a60655a );
 a2619a <=( a60644a  and  a60631a );
 a2620a <=( a60620a  and  a60607a );
 a2621a <=( a60596a  and  a60583a );
 a2622a <=( a60572a  and  a60559a );
 a2623a <=( a60548a  and  a60535a );
 a2624a <=( a60524a  and  a60511a );
 a2625a <=( a60500a  and  a60487a );
 a2626a <=( a60476a  and  a60463a );
 a2627a <=( a60452a  and  a60439a );
 a2628a <=( a60428a  and  a60415a );
 a2629a <=( a60404a  and  a60391a );
 a2630a <=( a60380a  and  a60367a );
 a2631a <=( a60356a  and  a60343a );
 a2632a <=( a60332a  and  a60319a );
 a2633a <=( a60308a  and  a60295a );
 a2634a <=( a60284a  and  a60271a );
 a2635a <=( a60260a  and  a60247a );
 a2636a <=( a60236a  and  a60223a );
 a2637a <=( a60212a  and  a60199a );
 a2638a <=( a60188a  and  a60175a );
 a2639a <=( a60164a  and  a60151a );
 a2640a <=( a60140a  and  a60127a );
 a2641a <=( a60116a  and  a60103a );
 a2642a <=( a60092a  and  a60079a );
 a2643a <=( a60068a  and  a60055a );
 a2644a <=( a60044a  and  a60031a );
 a2645a <=( a60020a  and  a60007a );
 a2646a <=( a59996a  and  a59983a );
 a2647a <=( a59972a  and  a59959a );
 a2648a <=( a59948a  and  a59935a );
 a2649a <=( a59924a  and  a59911a );
 a2650a <=( a59900a  and  a59887a );
 a2651a <=( a59876a  and  a59863a );
 a2652a <=( a59852a  and  a59839a );
 a2653a <=( a59828a  and  a59815a );
 a2654a <=( a59804a  and  a59791a );
 a2655a <=( a59780a  and  a59767a );
 a2656a <=( a59756a  and  a59743a );
 a2657a <=( a59732a  and  a59719a );
 a2658a <=( a59708a  and  a59695a );
 a2659a <=( a59684a  and  a59671a );
 a2660a <=( a59660a  and  a59647a );
 a2661a <=( a59636a  and  a59623a );
 a2662a <=( a59612a  and  a59599a );
 a2663a <=( a59588a  and  a59575a );
 a2664a <=( a59564a  and  a59551a );
 a2665a <=( a59540a  and  a59527a );
 a2666a <=( a59516a  and  a59503a );
 a2667a <=( a59492a  and  a59479a );
 a2668a <=( a59468a  and  a59455a );
 a2669a <=( a59444a  and  a59431a );
 a2670a <=( a59420a  and  a59407a );
 a2671a <=( a59396a  and  a59383a );
 a2672a <=( a59372a  and  a59359a );
 a2673a <=( a59348a  and  a59335a );
 a2674a <=( a59324a  and  a59311a );
 a2675a <=( a59300a  and  a59287a );
 a2676a <=( a59276a  and  a59263a );
 a2677a <=( a59252a  and  a59239a );
 a2678a <=( a59228a  and  a59215a );
 a2679a <=( a59204a  and  a59191a );
 a2680a <=( a59180a  and  a59167a );
 a2681a <=( a59156a  and  a59143a );
 a2682a <=( a59132a  and  a59119a );
 a2683a <=( a59108a  and  a59095a );
 a2684a <=( a59084a  and  a59071a );
 a2685a <=( a59060a  and  a59047a );
 a2686a <=( a59036a  and  a59023a );
 a2687a <=( a59012a  and  a58999a );
 a2688a <=( a58988a  and  a58975a );
 a2689a <=( a58964a  and  a58951a );
 a2690a <=( a58940a  and  a58927a );
 a2691a <=( a58916a  and  a58903a );
 a2692a <=( a58892a  and  a58879a );
 a2693a <=( a58868a  and  a58855a );
 a2694a <=( a58844a  and  a58831a );
 a2695a <=( a58820a  and  a58807a );
 a2696a <=( a58796a  and  a58783a );
 a2697a <=( a58772a  and  a58759a );
 a2698a <=( a58748a  and  a58735a );
 a2699a <=( a58724a  and  a58711a );
 a2700a <=( a58700a  and  a58687a );
 a2701a <=( a58676a  and  a58663a );
 a2702a <=( a58652a  and  a58639a );
 a2703a <=( a58628a  and  a58615a );
 a2704a <=( a58604a  and  a58591a );
 a2705a <=( a58580a  and  a58567a );
 a2706a <=( a58556a  and  a58543a );
 a2707a <=( a58532a  and  a58519a );
 a2708a <=( a58508a  and  a58495a );
 a2709a <=( a58484a  and  a58471a );
 a2710a <=( a58460a  and  a58447a );
 a2711a <=( a58436a  and  a58423a );
 a2712a <=( a58412a  and  a58399a );
 a2713a <=( a58388a  and  a58375a );
 a2714a <=( a58364a  and  a58351a );
 a2715a <=( a58340a  and  a58327a );
 a2716a <=( a58316a  and  a58303a );
 a2717a <=( a58292a  and  a58279a );
 a2718a <=( a58268a  and  a58255a );
 a2719a <=( a58244a  and  a58231a );
 a2720a <=( a58220a  and  a58207a );
 a2721a <=( a58196a  and  a58183a );
 a2722a <=( a58172a  and  a58159a );
 a2723a <=( a58148a  and  a58135a );
 a2724a <=( a58124a  and  a58111a );
 a2725a <=( a58100a  and  a58087a );
 a2726a <=( a58076a  and  a58063a );
 a2727a <=( a58052a  and  a58039a );
 a2728a <=( a58028a  and  a58015a );
 a2729a <=( a58004a  and  a57991a );
 a2730a <=( a57980a  and  a57967a );
 a2731a <=( a57956a  and  a57943a );
 a2732a <=( a57932a  and  a57919a );
 a2733a <=( a57908a  and  a57895a );
 a2734a <=( a57884a  and  a57871a );
 a2735a <=( a57860a  and  a57847a );
 a2736a <=( a57836a  and  a57823a );
 a2737a <=( a57812a  and  a57799a );
 a2738a <=( a57788a  and  a57775a );
 a2739a <=( a57764a  and  a57751a );
 a2740a <=( a57740a  and  a57727a );
 a2741a <=( a57716a  and  a57703a );
 a2742a <=( a57692a  and  a57679a );
 a2743a <=( a57668a  and  a57655a );
 a2744a <=( a57644a  and  a57631a );
 a2745a <=( a57620a  and  a57607a );
 a2746a <=( a57596a  and  a57583a );
 a2747a <=( a57572a  and  a57559a );
 a2748a <=( a57548a  and  a57535a );
 a2749a <=( a57524a  and  a57511a );
 a2750a <=( a57500a  and  a57487a );
 a2751a <=( a57476a  and  a57463a );
 a2752a <=( a57452a  and  a57439a );
 a2753a <=( a57428a  and  a57415a );
 a2754a <=( a57404a  and  a57391a );
 a2755a <=( a57380a  and  a57367a );
 a2756a <=( a57356a  and  a57343a );
 a2757a <=( a57332a  and  a57319a );
 a2758a <=( a57308a  and  a57295a );
 a2759a <=( a57284a  and  a57271a );
 a2760a <=( a57260a  and  a57247a );
 a2761a <=( a57236a  and  a57223a );
 a2762a <=( a57212a  and  a57199a );
 a2763a <=( a57188a  and  a57175a );
 a2764a <=( a57164a  and  a57151a );
 a2765a <=( a57140a  and  a57127a );
 a2766a <=( a57116a  and  a57103a );
 a2767a <=( a57092a  and  a57079a );
 a2768a <=( a57068a  and  a57055a );
 a2769a <=( a57044a  and  a57031a );
 a2770a <=( a57020a  and  a57007a );
 a2771a <=( a56996a  and  a56983a );
 a2772a <=( a56972a  and  a56959a );
 a2773a <=( a56948a  and  a56935a );
 a2774a <=( a56924a  and  a56911a );
 a2775a <=( a56900a  and  a56887a );
 a2776a <=( a56876a  and  a56863a );
 a2777a <=( a56852a  and  a56839a );
 a2778a <=( a56828a  and  a56815a );
 a2779a <=( a56804a  and  a56791a );
 a2780a <=( a56780a  and  a56767a );
 a2781a <=( a56756a  and  a56743a );
 a2782a <=( a56732a  and  a56719a );
 a2783a <=( a56708a  and  a56695a );
 a2784a <=( a56684a  and  a56671a );
 a2785a <=( a56660a  and  a56647a );
 a2786a <=( a56636a  and  a56623a );
 a2787a <=( a56612a  and  a56599a );
 a2788a <=( a56588a  and  a56575a );
 a2789a <=( a56564a  and  a56551a );
 a2790a <=( a56540a  and  a56527a );
 a2791a <=( a56516a  and  a56503a );
 a2792a <=( a56492a  and  a56479a );
 a2793a <=( a56468a  and  a56455a );
 a2794a <=( a56444a  and  a56431a );
 a2795a <=( a56420a  and  a56407a );
 a2796a <=( a56396a  and  a56383a );
 a2797a <=( a56372a  and  a56359a );
 a2798a <=( a56348a  and  a56335a );
 a2799a <=( a56324a  and  a56311a );
 a2800a <=( a56300a  and  a56287a );
 a2801a <=( a56276a  and  a56263a );
 a2802a <=( a56252a  and  a56239a );
 a2803a <=( a56228a  and  a56215a );
 a2804a <=( a56204a  and  a56191a );
 a2805a <=( a56180a  and  a56167a );
 a2806a <=( a56156a  and  a56143a );
 a2807a <=( a56132a  and  a56119a );
 a2808a <=( a56108a  and  a56095a );
 a2809a <=( a56084a  and  a56071a );
 a2810a <=( a56060a  and  a56047a );
 a2811a <=( a56036a  and  a56023a );
 a2812a <=( a56012a  and  a55999a );
 a2813a <=( a55988a  and  a55975a );
 a2814a <=( a55964a  and  a55951a );
 a2815a <=( a55940a  and  a55927a );
 a2816a <=( a55916a  and  a55903a );
 a2817a <=( a55892a  and  a55879a );
 a2818a <=( a55868a  and  a55855a );
 a2819a <=( a55844a  and  a55831a );
 a2820a <=( a55820a  and  a55807a );
 a2821a <=( a55796a  and  a55783a );
 a2822a <=( a55772a  and  a55759a );
 a2823a <=( a55748a  and  a55735a );
 a2824a <=( a55724a  and  a55711a );
 a2825a <=( a55700a  and  a55687a );
 a2826a <=( a55676a  and  a55663a );
 a2827a <=( a55652a  and  a55639a );
 a2828a <=( a55628a  and  a55615a );
 a2829a <=( a55604a  and  a55591a );
 a2830a <=( a55580a  and  a55567a );
 a2831a <=( a55556a  and  a55543a );
 a2832a <=( a55532a  and  a55519a );
 a2833a <=( a55508a  and  a55495a );
 a2834a <=( a55484a  and  a55471a );
 a2835a <=( a55460a  and  a55447a );
 a2836a <=( a55436a  and  a55423a );
 a2837a <=( a55412a  and  a55399a );
 a2838a <=( a55388a  and  a55375a );
 a2839a <=( a55364a  and  a55351a );
 a2840a <=( a55340a  and  a55327a );
 a2841a <=( a55316a  and  a55303a );
 a2842a <=( a55292a  and  a55279a );
 a2843a <=( a55268a  and  a55255a );
 a2844a <=( a55244a  and  a55231a );
 a2845a <=( a55220a  and  a55207a );
 a2846a <=( a55196a  and  a55183a );
 a2847a <=( a55172a  and  a55159a );
 a2848a <=( a55148a  and  a55135a );
 a2849a <=( a55124a  and  a55111a );
 a2850a <=( a55100a  and  a55087a );
 a2851a <=( a55076a  and  a55063a );
 a2852a <=( a55052a  and  a55039a );
 a2853a <=( a55028a  and  a55015a );
 a2854a <=( a55004a  and  a54991a );
 a2855a <=( a54980a  and  a54967a );
 a2856a <=( a54956a  and  a54943a );
 a2857a <=( a54932a  and  a54919a );
 a2858a <=( a54908a  and  a54895a );
 a2859a <=( a54884a  and  a54871a );
 a2860a <=( a54860a  and  a54847a );
 a2861a <=( a54836a  and  a54823a );
 a2862a <=( a54812a  and  a54799a );
 a2863a <=( a54788a  and  a54775a );
 a2864a <=( a54764a  and  a54751a );
 a2865a <=( a54740a  and  a54727a );
 a2866a <=( a54716a  and  a54703a );
 a2867a <=( a54692a  and  a54679a );
 a2868a <=( a54668a  and  a54655a );
 a2869a <=( a54644a  and  a54631a );
 a2870a <=( a54620a  and  a54607a );
 a2871a <=( a54596a  and  a54583a );
 a2872a <=( a54572a  and  a54559a );
 a2873a <=( a54548a  and  a54535a );
 a2874a <=( a54524a  and  a54511a );
 a2875a <=( a54500a  and  a54487a );
 a2876a <=( a54476a  and  a54463a );
 a2877a <=( a54452a  and  a54439a );
 a2878a <=( a54428a  and  a54415a );
 a2879a <=( a54404a  and  a54391a );
 a2880a <=( a54380a  and  a54367a );
 a2881a <=( a54356a  and  a54343a );
 a2882a <=( a54332a  and  a54319a );
 a2883a <=( a54308a  and  a54295a );
 a2884a <=( a54284a  and  a54271a );
 a2885a <=( a54260a  and  a54247a );
 a2886a <=( a54236a  and  a54223a );
 a2887a <=( a54212a  and  a54199a );
 a2888a <=( a54188a  and  a54175a );
 a2889a <=( a54164a  and  a54151a );
 a2890a <=( a54140a  and  a54127a );
 a2891a <=( a54116a  and  a54103a );
 a2892a <=( a54092a  and  a54079a );
 a2893a <=( a54068a  and  a54055a );
 a2894a <=( a54044a  and  a54031a );
 a2895a <=( a54020a  and  a54007a );
 a2896a <=( a53996a  and  a53983a );
 a2897a <=( a53972a  and  a53959a );
 a2898a <=( a53948a  and  a53935a );
 a2899a <=( a53924a  and  a53911a );
 a2900a <=( a53900a  and  a53887a );
 a2901a <=( a53876a  and  a53863a );
 a2902a <=( a53852a  and  a53839a );
 a2903a <=( a53828a  and  a53815a );
 a2904a <=( a53804a  and  a53791a );
 a2905a <=( a53780a  and  a53767a );
 a2906a <=( a53756a  and  a53743a );
 a2907a <=( a53732a  and  a53719a );
 a2908a <=( a53708a  and  a53695a );
 a2909a <=( a53684a  and  a53671a );
 a2910a <=( a53660a  and  a53647a );
 a2911a <=( a53636a  and  a53623a );
 a2912a <=( a53612a  and  a53599a );
 a2913a <=( a53588a  and  a53575a );
 a2914a <=( a53564a  and  a53551a );
 a2915a <=( a53540a  and  a53527a );
 a2916a <=( a53516a  and  a53503a );
 a2917a <=( a53492a  and  a53479a );
 a2918a <=( a53468a  and  a53455a );
 a2919a <=( a53444a  and  a53431a );
 a2920a <=( a53420a  and  a53407a );
 a2921a <=( a53396a  and  a53383a );
 a2922a <=( a53372a  and  a53359a );
 a2923a <=( a53348a  and  a53335a );
 a2924a <=( a53324a  and  a53311a );
 a2925a <=( a53300a  and  a53287a );
 a2926a <=( a53276a  and  a53263a );
 a2927a <=( a53252a  and  a53239a );
 a2928a <=( a53228a  and  a53215a );
 a2929a <=( a53204a  and  a53191a );
 a2930a <=( a53180a  and  a53167a );
 a2931a <=( a53156a  and  a53143a );
 a2932a <=( a53132a  and  a53119a );
 a2933a <=( a53108a  and  a53095a );
 a2934a <=( a53084a  and  a53071a );
 a2935a <=( a53060a  and  a53047a );
 a2936a <=( a53036a  and  a53023a );
 a2937a <=( a53012a  and  a52999a );
 a2938a <=( a52988a  and  a52975a );
 a2939a <=( a52964a  and  a52951a );
 a2940a <=( a52940a  and  a52927a );
 a2941a <=( a52916a  and  a52903a );
 a2942a <=( a52892a  and  a52879a );
 a2943a <=( a52868a  and  a52855a );
 a2944a <=( a52844a  and  a52831a );
 a2945a <=( a52820a  and  a52807a );
 a2946a <=( a52796a  and  a52783a );
 a2947a <=( a52772a  and  a52759a );
 a2948a <=( a52748a  and  a52735a );
 a2949a <=( a52724a  and  a52711a );
 a2950a <=( a52700a  and  a52687a );
 a2951a <=( a52676a  and  a52663a );
 a2952a <=( a52652a  and  a52639a );
 a2953a <=( a52628a  and  a52615a );
 a2954a <=( a52604a  and  a52591a );
 a2955a <=( a52580a  and  a52567a );
 a2956a <=( a52556a  and  a52543a );
 a2957a <=( a52532a  and  a52519a );
 a2958a <=( a52508a  and  a52495a );
 a2959a <=( a52484a  and  a52471a );
 a2960a <=( a52460a  and  a52447a );
 a2961a <=( a52436a  and  a52423a );
 a2962a <=( a52412a  and  a52399a );
 a2963a <=( a52388a  and  a52375a );
 a2964a <=( a52364a  and  a52351a );
 a2965a <=( a52340a  and  a52327a );
 a2966a <=( a52316a  and  a52303a );
 a2967a <=( a52292a  and  a52279a );
 a2968a <=( a52268a  and  a52255a );
 a2969a <=( a52244a  and  a52231a );
 a2970a <=( a52220a  and  a52207a );
 a2971a <=( a52196a  and  a52183a );
 a2972a <=( a52172a  and  a52159a );
 a2973a <=( a52148a  and  a52135a );
 a2974a <=( a52124a  and  a52111a );
 a2975a <=( a52100a  and  a52087a );
 a2976a <=( a52076a  and  a52063a );
 a2977a <=( a52052a  and  a52039a );
 a2978a <=( a52028a  and  a52015a );
 a2979a <=( a52004a  and  a51991a );
 a2980a <=( a51980a  and  a51967a );
 a2981a <=( a51956a  and  a51943a );
 a2982a <=( a51932a  and  a51919a );
 a2983a <=( a51908a  and  a51895a );
 a2984a <=( a51884a  and  a51871a );
 a2985a <=( a51860a  and  a51847a );
 a2986a <=( a51836a  and  a51823a );
 a2987a <=( a51812a  and  a51799a );
 a2988a <=( a51788a  and  a51775a );
 a2989a <=( a51764a  and  a51751a );
 a2990a <=( a51740a  and  a51727a );
 a2991a <=( a51716a  and  a51703a );
 a2992a <=( a51692a  and  a51679a );
 a2993a <=( a51668a  and  a51655a );
 a2994a <=( a51644a  and  a51631a );
 a2995a <=( a51620a  and  a51607a );
 a2996a <=( a51596a  and  a51583a );
 a2997a <=( a51572a  and  a51559a );
 a2998a <=( a51548a  and  a51535a );
 a2999a <=( a51524a  and  a51511a );
 a3000a <=( a51500a  and  a51487a );
 a3001a <=( a51476a  and  a51463a );
 a3002a <=( a51452a  and  a51439a );
 a3003a <=( a51428a  and  a51415a );
 a3004a <=( a51404a  and  a51391a );
 a3005a <=( a51380a  and  a51367a );
 a3006a <=( a51356a  and  a51343a );
 a3007a <=( a51332a  and  a51319a );
 a3008a <=( a51308a  and  a51295a );
 a3009a <=( a51284a  and  a51271a );
 a3010a <=( a51260a  and  a51247a );
 a3011a <=( a51236a  and  a51223a );
 a3012a <=( a51212a  and  a51199a );
 a3013a <=( a51188a  and  a51175a );
 a3014a <=( a51164a  and  a51151a );
 a3015a <=( a51140a  and  a51127a );
 a3016a <=( a51116a  and  a51103a );
 a3017a <=( a51092a  and  a51079a );
 a3018a <=( a51068a  and  a51055a );
 a3019a <=( a51044a  and  a51031a );
 a3020a <=( a51020a  and  a51007a );
 a3021a <=( a50996a  and  a50983a );
 a3022a <=( a50972a  and  a50959a );
 a3023a <=( a50948a  and  a50935a );
 a3024a <=( a50924a  and  a50911a );
 a3025a <=( a50900a  and  a50887a );
 a3026a <=( a50876a  and  a50863a );
 a3027a <=( a50852a  and  a50839a );
 a3028a <=( a50828a  and  a50815a );
 a3029a <=( a50804a  and  a50791a );
 a3030a <=( a50780a  and  a50767a );
 a3031a <=( a50756a  and  a50743a );
 a3032a <=( a50732a  and  a50719a );
 a3033a <=( a50708a  and  a50695a );
 a3034a <=( a50684a  and  a50671a );
 a3035a <=( a50660a  and  a50647a );
 a3036a <=( a50636a  and  a50623a );
 a3037a <=( a50612a  and  a50599a );
 a3038a <=( a50588a  and  a50575a );
 a3039a <=( a50564a  and  a50551a );
 a3040a <=( a50540a  and  a50527a );
 a3041a <=( a50516a  and  a50503a );
 a3042a <=( a50492a  and  a50479a );
 a3043a <=( a50468a  and  a50455a );
 a3044a <=( a50444a  and  a50431a );
 a3045a <=( a50420a  and  a50407a );
 a3046a <=( a50396a  and  a50383a );
 a3047a <=( a50372a  and  a50359a );
 a3048a <=( a50348a  and  a50335a );
 a3049a <=( a50324a  and  a50311a );
 a3050a <=( a50300a  and  a50287a );
 a3051a <=( a50276a  and  a50263a );
 a3052a <=( a50252a  and  a50239a );
 a3053a <=( a50228a  and  a50215a );
 a3054a <=( a50204a  and  a50191a );
 a3055a <=( a50180a  and  a50167a );
 a3056a <=( a50156a  and  a50143a );
 a3057a <=( a50132a  and  a50119a );
 a3058a <=( a50108a  and  a50095a );
 a3059a <=( a50084a  and  a50071a );
 a3060a <=( a50060a  and  a50047a );
 a3061a <=( a50036a  and  a50023a );
 a3062a <=( a50012a  and  a49999a );
 a3063a <=( a49988a  and  a49975a );
 a3064a <=( a49964a  and  a49951a );
 a3065a <=( a49940a  and  a49927a );
 a3066a <=( a49916a  and  a49903a );
 a3067a <=( a49892a  and  a49879a );
 a3068a <=( a49868a  and  a49855a );
 a3069a <=( a49844a  and  a49831a );
 a3070a <=( a49820a  and  a49807a );
 a3071a <=( a49796a  and  a49783a );
 a3072a <=( a49772a  and  a49759a );
 a3073a <=( a49748a  and  a49735a );
 a3074a <=( a49724a  and  a49711a );
 a3075a <=( a49700a  and  a49687a );
 a3076a <=( a49676a  and  a49663a );
 a3077a <=( a49652a  and  a49639a );
 a3078a <=( a49628a  and  a49615a );
 a3079a <=( a49604a  and  a49591a );
 a3080a <=( a49580a  and  a49567a );
 a3081a <=( a49556a  and  a49543a );
 a3082a <=( a49532a  and  a49519a );
 a3083a <=( a49508a  and  a49495a );
 a3084a <=( a49484a  and  a49471a );
 a3085a <=( a49460a  and  a49447a );
 a3086a <=( a49436a  and  a49423a );
 a3087a <=( a49412a  and  a49399a );
 a3088a <=( a49388a  and  a49375a );
 a3089a <=( a49364a  and  a49351a );
 a3090a <=( a49340a  and  a49327a );
 a3091a <=( a49316a  and  a49303a );
 a3092a <=( a49292a  and  a49279a );
 a3093a <=( a49268a  and  a49255a );
 a3094a <=( a49244a  and  a49231a );
 a3095a <=( a49220a  and  a49207a );
 a3096a <=( a49196a  and  a49183a );
 a3097a <=( a49172a  and  a49159a );
 a3098a <=( a49148a  and  a49135a );
 a3099a <=( a49124a  and  a49111a );
 a3100a <=( a49100a  and  a49087a );
 a3101a <=( a49076a  and  a49063a );
 a3102a <=( a49052a  and  a49039a );
 a3103a <=( a49028a  and  a49015a );
 a3104a <=( a49004a  and  a48991a );
 a3105a <=( a48980a  and  a48967a );
 a3106a <=( a48956a  and  a48943a );
 a3107a <=( a48932a  and  a48919a );
 a3108a <=( a48908a  and  a48895a );
 a3109a <=( a48884a  and  a48871a );
 a3110a <=( a48860a  and  a48847a );
 a3111a <=( a48836a  and  a48823a );
 a3112a <=( a48812a  and  a48799a );
 a3113a <=( a48788a  and  a48775a );
 a3114a <=( a48764a  and  a48751a );
 a3115a <=( a48740a  and  a48727a );
 a3116a <=( a48716a  and  a48703a );
 a3117a <=( a48692a  and  a48679a );
 a3118a <=( a48668a  and  a48655a );
 a3119a <=( a48644a  and  a48631a );
 a3120a <=( a48620a  and  a48607a );
 a3121a <=( a48596a  and  a48583a );
 a3122a <=( a48572a  and  a48559a );
 a3123a <=( a48548a  and  a48535a );
 a3124a <=( a48524a  and  a48511a );
 a3125a <=( a48500a  and  a48487a );
 a3126a <=( a48476a  and  a48463a );
 a3127a <=( a48452a  and  a48439a );
 a3128a <=( a48428a  and  a48415a );
 a3129a <=( a48404a  and  a48391a );
 a3130a <=( a48380a  and  a48367a );
 a3131a <=( a48356a  and  a48343a );
 a3132a <=( a48332a  and  a48319a );
 a3133a <=( a48308a  and  a48295a );
 a3134a <=( a48284a  and  a48271a );
 a3135a <=( a48260a  and  a48247a );
 a3136a <=( a48236a  and  a48223a );
 a3137a <=( a48212a  and  a48199a );
 a3138a <=( a48188a  and  a48175a );
 a3139a <=( a48164a  and  a48151a );
 a3140a <=( a48140a  and  a48127a );
 a3141a <=( a48116a  and  a48103a );
 a3142a <=( a48092a  and  a48079a );
 a3143a <=( a48068a  and  a48055a );
 a3144a <=( a48044a  and  a48031a );
 a3145a <=( a48020a  and  a48007a );
 a3146a <=( a47996a  and  a47983a );
 a3147a <=( a47972a  and  a47959a );
 a3148a <=( a47948a  and  a47935a );
 a3149a <=( a47924a  and  a47911a );
 a3150a <=( a47900a  and  a47887a );
 a3151a <=( a47876a  and  a47863a );
 a3152a <=( a47852a  and  a47839a );
 a3153a <=( a47828a  and  a47815a );
 a3154a <=( a47804a  and  a47791a );
 a3155a <=( a47780a  and  a47767a );
 a3156a <=( a47756a  and  a47743a );
 a3157a <=( a47732a  and  a47719a );
 a3158a <=( a47708a  and  a47695a );
 a3159a <=( a47684a  and  a47671a );
 a3160a <=( a47660a  and  a47647a );
 a3161a <=( a47636a  and  a47623a );
 a3162a <=( a47612a  and  a47599a );
 a3163a <=( a47588a  and  a47575a );
 a3164a <=( a47564a  and  a47551a );
 a3165a <=( a47540a  and  a47527a );
 a3166a <=( a47516a  and  a47503a );
 a3167a <=( a47492a  and  a47479a );
 a3168a <=( a47468a  and  a47455a );
 a3169a <=( a47444a  and  a47431a );
 a3170a <=( a47420a  and  a47407a );
 a3171a <=( a47396a  and  a47383a );
 a3172a <=( a47372a  and  a47359a );
 a3173a <=( a47348a  and  a47335a );
 a3174a <=( a47324a  and  a47311a );
 a3175a <=( a47300a  and  a47287a );
 a3176a <=( a47276a  and  a47263a );
 a3177a <=( a47252a  and  a47239a );
 a3178a <=( a47228a  and  a47215a );
 a3179a <=( a47204a  and  a47191a );
 a3180a <=( a47180a  and  a47167a );
 a3181a <=( a47156a  and  a47143a );
 a3182a <=( a47132a  and  a47119a );
 a3183a <=( a47108a  and  a47095a );
 a3184a <=( a47084a  and  a47071a );
 a3185a <=( a47060a  and  a47047a );
 a3186a <=( a47036a  and  a47023a );
 a3187a <=( a47012a  and  a46999a );
 a3188a <=( a46988a  and  a46975a );
 a3189a <=( a46964a  and  a46951a );
 a3190a <=( a46940a  and  a46927a );
 a3191a <=( a46916a  and  a46903a );
 a3192a <=( a46892a  and  a46879a );
 a3193a <=( a46868a  and  a46855a );
 a3194a <=( a46844a  and  a46831a );
 a3195a <=( a46820a  and  a46807a );
 a3196a <=( a46796a  and  a46783a );
 a3197a <=( a46772a  and  a46759a );
 a3198a <=( a46748a  and  a46735a );
 a3199a <=( a46724a  and  a46711a );
 a3200a <=( a46700a  and  a46687a );
 a3201a <=( a46676a  and  a46663a );
 a3202a <=( a46652a  and  a46639a );
 a3203a <=( a46628a  and  a46615a );
 a3204a <=( a46604a  and  a46591a );
 a3205a <=( a46580a  and  a46567a );
 a3206a <=( a46556a  and  a46543a );
 a3207a <=( a46532a  and  a46519a );
 a3208a <=( a46508a  and  a46495a );
 a3209a <=( a46484a  and  a46471a );
 a3210a <=( a46460a  and  a46447a );
 a3211a <=( a46436a  and  a46423a );
 a3212a <=( a46412a  and  a46399a );
 a3213a <=( a46388a  and  a46375a );
 a3214a <=( a46364a  and  a46351a );
 a3215a <=( a46340a  and  a46327a );
 a3216a <=( a46316a  and  a46303a );
 a3217a <=( a46292a  and  a46279a );
 a3218a <=( a46268a  and  a46255a );
 a3219a <=( a46244a  and  a46231a );
 a3220a <=( a46220a  and  a46207a );
 a3221a <=( a46196a  and  a46183a );
 a3222a <=( a46172a  and  a46159a );
 a3223a <=( a46148a  and  a46135a );
 a3224a <=( a46124a  and  a46111a );
 a3225a <=( a46100a  and  a46087a );
 a3226a <=( a46076a  and  a46063a );
 a3227a <=( a46052a  and  a46039a );
 a3228a <=( a46028a  and  a46015a );
 a3229a <=( a46004a  and  a45991a );
 a3230a <=( a45980a  and  a45967a );
 a3231a <=( a45956a  and  a45943a );
 a3232a <=( a45932a  and  a45919a );
 a3233a <=( a45908a  and  a45895a );
 a3234a <=( a45884a  and  a45871a );
 a3235a <=( a45860a  and  a45847a );
 a3236a <=( a45836a  and  a45823a );
 a3237a <=( a45812a  and  a45799a );
 a3238a <=( a45788a  and  a45775a );
 a3239a <=( a45764a  and  a45751a );
 a3240a <=( a45740a  and  a45727a );
 a3241a <=( a45716a  and  a45703a );
 a3242a <=( a45692a  and  a45679a );
 a3243a <=( a45668a  and  a45655a );
 a3244a <=( a45644a  and  a45631a );
 a3245a <=( a45620a  and  a45607a );
 a3246a <=( a45596a  and  a45583a );
 a3247a <=( a45572a  and  a45559a );
 a3248a <=( a45548a  and  a45535a );
 a3249a <=( a45524a  and  a45511a );
 a3250a <=( a45500a  and  a45487a );
 a3251a <=( a45476a  and  a45463a );
 a3252a <=( a45452a  and  a45439a );
 a3253a <=( a45428a  and  a45415a );
 a3254a <=( a45404a  and  a45391a );
 a3255a <=( a45380a  and  a45367a );
 a3256a <=( a45356a  and  a45343a );
 a3257a <=( a45332a  and  a45319a );
 a3258a <=( a45308a  and  a45295a );
 a3259a <=( a45284a  and  a45271a );
 a3260a <=( a45260a  and  a45247a );
 a3261a <=( a45236a  and  a45223a );
 a3262a <=( a45212a  and  a45199a );
 a3263a <=( a45188a  and  a45175a );
 a3264a <=( a45164a  and  a45151a );
 a3265a <=( a45140a  and  a45127a );
 a3266a <=( a45116a  and  a45103a );
 a3267a <=( a45092a  and  a45079a );
 a3268a <=( a45068a  and  a45055a );
 a3269a <=( a45044a  and  a45031a );
 a3270a <=( a45020a  and  a45007a );
 a3271a <=( a44996a  and  a44983a );
 a3272a <=( a44972a  and  a44959a );
 a3273a <=( a44948a  and  a44935a );
 a3274a <=( a44924a  and  a44911a );
 a3275a <=( a44900a  and  a44887a );
 a3276a <=( a44876a  and  a44863a );
 a3277a <=( a44852a  and  a44839a );
 a3278a <=( a44828a  and  a44815a );
 a3279a <=( a44804a  and  a44791a );
 a3280a <=( a44780a  and  a44767a );
 a3281a <=( a44756a  and  a44743a );
 a3282a <=( a44732a  and  a44719a );
 a3283a <=( a44708a  and  a44695a );
 a3284a <=( a44684a  and  a44671a );
 a3285a <=( a44660a  and  a44647a );
 a3286a <=( a44636a  and  a44623a );
 a3287a <=( a44612a  and  a44599a );
 a3288a <=( a44588a  and  a44575a );
 a3289a <=( a44564a  and  a44553a );
 a3290a <=( a44542a  and  a44531a );
 a3291a <=( a44520a  and  a44509a );
 a3292a <=( a44498a  and  a44487a );
 a3293a <=( a44476a  and  a44465a );
 a3294a <=( a44454a  and  a44443a );
 a3295a <=( a44432a  and  a44421a );
 a3296a <=( a44410a  and  a44399a );
 a3297a <=( a44388a  and  a44377a );
 a3298a <=( a44366a  and  a44355a );
 a3299a <=( a44344a  and  a44333a );
 a3300a <=( a44322a  and  a44311a );
 a3301a <=( a44300a  and  a44289a );
 a3302a <=( a44278a  and  a44267a );
 a3303a <=( a44256a  and  a44245a );
 a3304a <=( a44234a  and  a44223a );
 a3305a <=( a44212a  and  a44201a );
 a3306a <=( a44190a  and  a44179a );
 a3307a <=( a44168a  and  a44157a );
 a3308a <=( a44146a  and  a44135a );
 a3309a <=( a44124a  and  a44113a );
 a3310a <=( a44102a  and  a44091a );
 a3311a <=( a44080a  and  a44069a );
 a3312a <=( a44058a  and  a44047a );
 a3313a <=( a44036a  and  a44025a );
 a3314a <=( a44014a  and  a44003a );
 a3315a <=( a43992a  and  a43981a );
 a3316a <=( a43970a  and  a43959a );
 a3317a <=( a43948a  and  a43937a );
 a3318a <=( a43926a  and  a43915a );
 a3319a <=( a43904a  and  a43893a );
 a3320a <=( a43882a  and  a43871a );
 a3321a <=( a43860a  and  a43849a );
 a3322a <=( a43838a  and  a43827a );
 a3323a <=( a43816a  and  a43805a );
 a3324a <=( a43794a  and  a43783a );
 a3325a <=( a43772a  and  a43761a );
 a3326a <=( a43750a  and  a43739a );
 a3327a <=( a43728a  and  a43717a );
 a3328a <=( a43706a  and  a43695a );
 a3329a <=( a43684a  and  a43673a );
 a3330a <=( a43662a  and  a43651a );
 a3331a <=( a43640a  and  a43629a );
 a3332a <=( a43618a  and  a43607a );
 a3333a <=( a43596a  and  a43585a );
 a3334a <=( a43574a  and  a43563a );
 a3335a <=( a43552a  and  a43541a );
 a3336a <=( a43530a  and  a43519a );
 a3337a <=( a43508a  and  a43497a );
 a3338a <=( a43486a  and  a43475a );
 a3339a <=( a43464a  and  a43453a );
 a3340a <=( a43442a  and  a43431a );
 a3341a <=( a43420a  and  a43409a );
 a3342a <=( a43398a  and  a43387a );
 a3343a <=( a43376a  and  a43365a );
 a3344a <=( a43354a  and  a43343a );
 a3345a <=( a43332a  and  a43321a );
 a3346a <=( a43310a  and  a43299a );
 a3347a <=( a43288a  and  a43277a );
 a3348a <=( a43266a  and  a43255a );
 a3349a <=( a43244a  and  a43233a );
 a3350a <=( a43222a  and  a43211a );
 a3351a <=( a43200a  and  a43189a );
 a3352a <=( a43178a  and  a43167a );
 a3353a <=( a43156a  and  a43145a );
 a3354a <=( a43134a  and  a43123a );
 a3355a <=( a43112a  and  a43101a );
 a3356a <=( a43090a  and  a43079a );
 a3357a <=( a43068a  and  a43057a );
 a3358a <=( a43046a  and  a43035a );
 a3359a <=( a43024a  and  a43013a );
 a3360a <=( a43002a  and  a42991a );
 a3361a <=( a42980a  and  a42969a );
 a3362a <=( a42958a  and  a42947a );
 a3363a <=( a42936a  and  a42925a );
 a3364a <=( a42914a  and  a42903a );
 a3365a <=( a42892a  and  a42881a );
 a3366a <=( a42870a  and  a42859a );
 a3367a <=( a42848a  and  a42837a );
 a3368a <=( a42826a  and  a42815a );
 a3369a <=( a42804a  and  a42793a );
 a3370a <=( a42782a  and  a42771a );
 a3371a <=( a42760a  and  a42749a );
 a3372a <=( a42738a  and  a42727a );
 a3373a <=( a42716a  and  a42705a );
 a3374a <=( a42694a  and  a42683a );
 a3375a <=( a42672a  and  a42661a );
 a3376a <=( a42650a  and  a42639a );
 a3377a <=( a42628a  and  a42617a );
 a3378a <=( a42606a  and  a42595a );
 a3379a <=( a42584a  and  a42573a );
 a3380a <=( a42562a  and  a42551a );
 a3381a <=( a42540a  and  a42529a );
 a3382a <=( a42518a  and  a42507a );
 a3383a <=( a42496a  and  a42485a );
 a3384a <=( a42474a  and  a42463a );
 a3385a <=( a42452a  and  a42441a );
 a3386a <=( a42430a  and  a42419a );
 a3387a <=( a42408a  and  a42397a );
 a3388a <=( a42386a  and  a42375a );
 a3389a <=( a42364a  and  a42353a );
 a3390a <=( a42342a  and  a42331a );
 a3391a <=( a42320a  and  a42309a );
 a3392a <=( a42298a  and  a42287a );
 a3393a <=( a42276a  and  a42265a );
 a3394a <=( a42254a  and  a42243a );
 a3395a <=( a42232a  and  a42221a );
 a3396a <=( a42210a  and  a42199a );
 a3397a <=( a42188a  and  a42177a );
 a3398a <=( a42166a  and  a42155a );
 a3399a <=( a42144a  and  a42133a );
 a3400a <=( a42122a  and  a42111a );
 a3401a <=( a42100a  and  a42089a );
 a3402a <=( a42078a  and  a42067a );
 a3403a <=( a42056a  and  a42045a );
 a3404a <=( a42034a  and  a42023a );
 a3405a <=( a42012a  and  a42001a );
 a3406a <=( a41990a  and  a41979a );
 a3407a <=( a41968a  and  a41957a );
 a3408a <=( a41946a  and  a41935a );
 a3409a <=( a41924a  and  a41913a );
 a3410a <=( a41902a  and  a41891a );
 a3411a <=( a41880a  and  a41869a );
 a3412a <=( a41858a  and  a41847a );
 a3413a <=( a41836a  and  a41825a );
 a3414a <=( a41814a  and  a41803a );
 a3415a <=( a41792a  and  a41781a );
 a3416a <=( a41770a  and  a41759a );
 a3417a <=( a41748a  and  a41737a );
 a3418a <=( a41726a  and  a41715a );
 a3419a <=( a41704a  and  a41693a );
 a3420a <=( a41682a  and  a41671a );
 a3421a <=( a41660a  and  a41649a );
 a3422a <=( a41638a  and  a41627a );
 a3423a <=( a41616a  and  a41605a );
 a3424a <=( a41594a  and  a41583a );
 a3425a <=( a41572a  and  a41561a );
 a3426a <=( a41550a  and  a41539a );
 a3427a <=( a41528a  and  a41517a );
 a3428a <=( a41506a  and  a41495a );
 a3429a <=( a41484a  and  a41473a );
 a3430a <=( a41462a  and  a41451a );
 a3431a <=( a41440a  and  a41429a );
 a3432a <=( a41418a  and  a41407a );
 a3433a <=( a41396a  and  a41385a );
 a3434a <=( a41374a  and  a41363a );
 a3435a <=( a41352a  and  a41341a );
 a3436a <=( a41330a  and  a41319a );
 a3437a <=( a41308a  and  a41297a );
 a3438a <=( a41286a  and  a41275a );
 a3439a <=( a41264a  and  a41253a );
 a3440a <=( a41242a  and  a41231a );
 a3441a <=( a41220a  and  a41209a );
 a3442a <=( a41198a  and  a41187a );
 a3443a <=( a41176a  and  a41165a );
 a3444a <=( a41154a  and  a41143a );
 a3445a <=( a41132a  and  a41121a );
 a3446a <=( a41110a  and  a41099a );
 a3447a <=( a41088a  and  a41077a );
 a3448a <=( a41066a  and  a41055a );
 a3449a <=( a41044a  and  a41033a );
 a3450a <=( a41022a  and  a41011a );
 a3451a <=( a41000a  and  a40989a );
 a3452a <=( a40978a  and  a40967a );
 a3453a <=( a40956a  and  a40945a );
 a3454a <=( a40934a  and  a40923a );
 a3455a <=( a40912a  and  a40901a );
 a3456a <=( a40890a  and  a40879a );
 a3457a <=( a40868a  and  a40857a );
 a3458a <=( a40846a  and  a40835a );
 a3459a <=( a40824a  and  a40813a );
 a3460a <=( a40802a  and  a40791a );
 a3461a <=( a40780a  and  a40769a );
 a3462a <=( a40758a  and  a40747a );
 a3463a <=( a40736a  and  a40725a );
 a3464a <=( a40714a  and  a40703a );
 a3465a <=( a40692a  and  a40681a );
 a3466a <=( a40670a  and  a40659a );
 a3467a <=( a40648a  and  a40637a );
 a3468a <=( a40626a  and  a40615a );
 a3469a <=( a40604a  and  a40593a );
 a3470a <=( a40582a  and  a40571a );
 a3471a <=( a40560a  and  a40549a );
 a3472a <=( a40538a  and  a40527a );
 a3473a <=( a40516a  and  a40505a );
 a3474a <=( a40494a  and  a40483a );
 a3475a <=( a40472a  and  a40461a );
 a3476a <=( a40450a  and  a40439a );
 a3477a <=( a40428a  and  a40417a );
 a3478a <=( a40406a  and  a40395a );
 a3479a <=( a40384a  and  a40373a );
 a3480a <=( a40362a  and  a40351a );
 a3481a <=( a40340a  and  a40329a );
 a3482a <=( a40318a  and  a40307a );
 a3483a <=( a40296a  and  a40285a );
 a3484a <=( a40274a  and  a40263a );
 a3485a <=( a40252a  and  a40241a );
 a3486a <=( a40230a  and  a40219a );
 a3487a <=( a40208a  and  a40197a );
 a3488a <=( a40186a  and  a40175a );
 a3489a <=( a40164a  and  a40153a );
 a3490a <=( a40142a  and  a40131a );
 a3491a <=( a40120a  and  a40109a );
 a3492a <=( a40098a  and  a40087a );
 a3493a <=( a40076a  and  a40065a );
 a3494a <=( a40054a  and  a40043a );
 a3495a <=( a40032a  and  a40021a );
 a3496a <=( a40010a  and  a39999a );
 a3497a <=( a39988a  and  a39977a );
 a3498a <=( a39966a  and  a39955a );
 a3499a <=( a39944a  and  a39933a );
 a3500a <=( a39922a  and  a39911a );
 a3501a <=( a39900a  and  a39889a );
 a3502a <=( a39878a  and  a39867a );
 a3503a <=( a39856a  and  a39845a );
 a3504a <=( a39834a  and  a39823a );
 a3505a <=( a39812a  and  a39801a );
 a3506a <=( a39790a  and  a39779a );
 a3507a <=( a39768a  and  a39757a );
 a3508a <=( a39746a  and  a39735a );
 a3509a <=( a39724a  and  a39713a );
 a3510a <=( a39702a  and  a39691a );
 a3511a <=( a39680a  and  a39669a );
 a3512a <=( a39658a  and  a39647a );
 a3513a <=( a39636a  and  a39625a );
 a3514a <=( a39614a  and  a39603a );
 a3515a <=( a39592a  and  a39581a );
 a3516a <=( a39570a  and  a39559a );
 a3517a <=( a39548a  and  a39537a );
 a3518a <=( a39526a  and  a39515a );
 a3519a <=( a39504a  and  a39493a );
 a3520a <=( a39482a  and  a39471a );
 a3521a <=( a39460a  and  a39449a );
 a3522a <=( a39438a  and  a39427a );
 a3523a <=( a39416a  and  a39405a );
 a3524a <=( a39394a  and  a39383a );
 a3525a <=( a39372a  and  a39361a );
 a3526a <=( a39350a  and  a39339a );
 a3527a <=( a39328a  and  a39317a );
 a3528a <=( a39306a  and  a39295a );
 a3529a <=( a39284a  and  a39273a );
 a3530a <=( a39262a  and  a39251a );
 a3531a <=( a39240a  and  a39229a );
 a3532a <=( a39218a  and  a39207a );
 a3533a <=( a39196a  and  a39185a );
 a3534a <=( a39174a  and  a39163a );
 a3535a <=( a39152a  and  a39141a );
 a3536a <=( a39130a  and  a39119a );
 a3537a <=( a39108a  and  a39097a );
 a3538a <=( a39086a  and  a39075a );
 a3539a <=( a39064a  and  a39053a );
 a3540a <=( a39042a  and  a39031a );
 a3541a <=( a39020a  and  a39009a );
 a3542a <=( a38998a  and  a38987a );
 a3543a <=( a38976a  and  a38965a );
 a3544a <=( a38954a  and  a38943a );
 a3545a <=( a38932a  and  a38921a );
 a3546a <=( a38910a  and  a38899a );
 a3547a <=( a38888a  and  a38877a );
 a3548a <=( a38866a  and  a38855a );
 a3549a <=( a38844a  and  a38833a );
 a3550a <=( a38822a  and  a38811a );
 a3551a <=( a38800a  and  a38789a );
 a3552a <=( a38778a  and  a38767a );
 a3553a <=( a38756a  and  a38745a );
 a3554a <=( a38734a  and  a38723a );
 a3555a <=( a38712a  and  a38701a );
 a3556a <=( a38690a  and  a38679a );
 a3557a <=( a38668a  and  a38657a );
 a3558a <=( a38646a  and  a38635a );
 a3559a <=( a38624a  and  a38613a );
 a3560a <=( a38602a  and  a38591a );
 a3561a <=( a38580a  and  a38569a );
 a3562a <=( a38558a  and  a38547a );
 a3563a <=( a38536a  and  a38525a );
 a3564a <=( a38514a  and  a38503a );
 a3565a <=( a38492a  and  a38481a );
 a3566a <=( a38470a  and  a38459a );
 a3567a <=( a38448a  and  a38437a );
 a3568a <=( a38426a  and  a38415a );
 a3569a <=( a38404a  and  a38393a );
 a3570a <=( a38382a  and  a38371a );
 a3571a <=( a38360a  and  a38349a );
 a3572a <=( a38338a  and  a38327a );
 a3573a <=( a38316a  and  a38305a );
 a3574a <=( a38294a  and  a38283a );
 a3575a <=( a38272a  and  a38261a );
 a3576a <=( a38250a  and  a38239a );
 a3577a <=( a38228a  and  a38217a );
 a3578a <=( a38206a  and  a38195a );
 a3579a <=( a38184a  and  a38173a );
 a3580a <=( a38162a  and  a38151a );
 a3581a <=( a38140a  and  a38129a );
 a3582a <=( a38118a  and  a38107a );
 a3583a <=( a38096a  and  a38085a );
 a3584a <=( a38074a  and  a38063a );
 a3585a <=( a38052a  and  a38041a );
 a3586a <=( a38030a  and  a38019a );
 a3587a <=( a38008a  and  a37997a );
 a3588a <=( a37986a  and  a37975a );
 a3589a <=( a37964a  and  a37953a );
 a3590a <=( a37942a  and  a37931a );
 a3591a <=( a37920a  and  a37909a );
 a3592a <=( a37898a  and  a37887a );
 a3593a <=( a37876a  and  a37865a );
 a3594a <=( a37854a  and  a37843a );
 a3595a <=( a37832a  and  a37821a );
 a3596a <=( a37810a  and  a37799a );
 a3597a <=( a37788a  and  a37777a );
 a3598a <=( a37766a  and  a37755a );
 a3599a <=( a37744a  and  a37733a );
 a3600a <=( a37722a  and  a37711a );
 a3601a <=( a37700a  and  a37689a );
 a3602a <=( a37678a  and  a37667a );
 a3603a <=( a37656a  and  a37645a );
 a3604a <=( a37634a  and  a37623a );
 a3605a <=( a37612a  and  a37601a );
 a3606a <=( a37590a  and  a37579a );
 a3607a <=( a37568a  and  a37557a );
 a3608a <=( a37546a  and  a37535a );
 a3609a <=( a37524a  and  a37513a );
 a3610a <=( a37502a  and  a37491a );
 a3611a <=( a37480a  and  a37469a );
 a3612a <=( a37458a  and  a37447a );
 a3613a <=( a37436a  and  a37425a );
 a3614a <=( a37414a  and  a37403a );
 a3615a <=( a37392a  and  a37381a );
 a3616a <=( a37370a  and  a37359a );
 a3617a <=( a37348a  and  a37337a );
 a3618a <=( a37326a  and  a37315a );
 a3619a <=( a37304a  and  a37293a );
 a3620a <=( a37282a  and  a37271a );
 a3621a <=( a37260a  and  a37249a );
 a3622a <=( a37238a  and  a37227a );
 a3623a <=( a37216a  and  a37205a );
 a3624a <=( a37194a  and  a37183a );
 a3625a <=( a37172a  and  a37161a );
 a3626a <=( a37150a  and  a37139a );
 a3627a <=( a37128a  and  a37117a );
 a3628a <=( a37106a  and  a37095a );
 a3629a <=( a37084a  and  a37073a );
 a3630a <=( a37062a  and  a37051a );
 a3631a <=( a37040a  and  a37029a );
 a3632a <=( a37018a  and  a37007a );
 a3633a <=( a36996a  and  a36985a );
 a3634a <=( a36974a  and  a36963a );
 a3635a <=( a36952a  and  a36941a );
 a3636a <=( a36930a  and  a36919a );
 a3637a <=( a36908a  and  a36897a );
 a3638a <=( a36886a  and  a36875a );
 a3639a <=( a36864a  and  a36853a );
 a3640a <=( a36842a  and  a36831a );
 a3641a <=( a36820a  and  a36809a );
 a3642a <=( a36798a  and  a36787a );
 a3643a <=( a36776a  and  a36765a );
 a3644a <=( a36754a  and  a36743a );
 a3645a <=( a36732a  and  a36721a );
 a3646a <=( a36710a  and  a36699a );
 a3647a <=( a36688a  and  a36677a );
 a3648a <=( a36666a  and  a36655a );
 a3649a <=( a36644a  and  a36633a );
 a3650a <=( a36622a  and  a36611a );
 a3651a <=( a36600a  and  a36589a );
 a3652a <=( a36578a  and  a36567a );
 a3653a <=( a36556a  and  a36545a );
 a3654a <=( a36534a  and  a36523a );
 a3655a <=( a36512a  and  a36501a );
 a3656a <=( a36490a  and  a36479a );
 a3657a <=( a36468a  and  a36457a );
 a3658a <=( a36446a  and  a36435a );
 a3659a <=( a36424a  and  a36413a );
 a3660a <=( a36402a  and  a36391a );
 a3661a <=( a36380a  and  a36369a );
 a3662a <=( a36358a  and  a36347a );
 a3663a <=( a36336a  and  a36325a );
 a3664a <=( a36314a  and  a36303a );
 a3665a <=( a36292a  and  a36281a );
 a3666a <=( a36270a  and  a36259a );
 a3667a <=( a36248a  and  a36237a );
 a3668a <=( a36226a  and  a36215a );
 a3669a <=( a36204a  and  a36193a );
 a3670a <=( a36182a  and  a36171a );
 a3671a <=( a36160a  and  a36149a );
 a3672a <=( a36138a  and  a36127a );
 a3673a <=( a36116a  and  a36105a );
 a3674a <=( a36094a  and  a36083a );
 a3675a <=( a36072a  and  a36061a );
 a3676a <=( a36050a  and  a36039a );
 a3677a <=( a36028a  and  a36017a );
 a3678a <=( a36006a  and  a35995a );
 a3679a <=( a35984a  and  a35973a );
 a3680a <=( a35962a  and  a35951a );
 a3681a <=( a35940a  and  a35929a );
 a3682a <=( a35918a  and  a35907a );
 a3683a <=( a35896a  and  a35885a );
 a3684a <=( a35874a  and  a35863a );
 a3685a <=( a35852a  and  a35841a );
 a3686a <=( a35830a  and  a35819a );
 a3687a <=( a35808a  and  a35797a );
 a3688a <=( a35786a  and  a35775a );
 a3689a <=( a35764a  and  a35753a );
 a3690a <=( a35742a  and  a35731a );
 a3691a <=( a35720a  and  a35709a );
 a3692a <=( a35698a  and  a35687a );
 a3693a <=( a35676a  and  a35665a );
 a3694a <=( a35654a  and  a35643a );
 a3695a <=( a35632a  and  a35621a );
 a3696a <=( a35610a  and  a35599a );
 a3697a <=( a35588a  and  a35577a );
 a3698a <=( a35566a  and  a35555a );
 a3699a <=( a35544a  and  a35533a );
 a3700a <=( a35522a  and  a35511a );
 a3701a <=( a35500a  and  a35489a );
 a3702a <=( a35478a  and  a35467a );
 a3703a <=( a35456a  and  a35445a );
 a3704a <=( a35434a  and  a35423a );
 a3705a <=( a35412a  and  a35401a );
 a3706a <=( a35390a  and  a35379a );
 a3707a <=( a35368a  and  a35357a );
 a3708a <=( a35346a  and  a35335a );
 a3709a <=( a35324a  and  a35313a );
 a3710a <=( a35302a  and  a35291a );
 a3711a <=( a35280a  and  a35269a );
 a3712a <=( a35258a  and  a35247a );
 a3713a <=( a35236a  and  a35225a );
 a3714a <=( a35214a  and  a35203a );
 a3715a <=( a35192a  and  a35181a );
 a3716a <=( a35170a  and  a35159a );
 a3717a <=( a35148a  and  a35137a );
 a3718a <=( a35126a  and  a35115a );
 a3719a <=( a35104a  and  a35093a );
 a3720a <=( a35082a  and  a35071a );
 a3721a <=( a35060a  and  a35049a );
 a3722a <=( a35038a  and  a35027a );
 a3723a <=( a35016a  and  a35005a );
 a3724a <=( a34994a  and  a34983a );
 a3725a <=( a34972a  and  a34961a );
 a3726a <=( a34950a  and  a34939a );
 a3727a <=( a34928a  and  a34917a );
 a3728a <=( a34906a  and  a34895a );
 a3729a <=( a34884a  and  a34873a );
 a3730a <=( a34862a  and  a34851a );
 a3731a <=( a34840a  and  a34829a );
 a3732a <=( a34818a  and  a34807a );
 a3733a <=( a34796a  and  a34785a );
 a3734a <=( a34774a  and  a34763a );
 a3735a <=( a34752a  and  a34741a );
 a3736a <=( a34730a  and  a34719a );
 a3737a <=( a34708a  and  a34697a );
 a3738a <=( a34686a  and  a34675a );
 a3739a <=( a34664a  and  a34653a );
 a3740a <=( a34642a  and  a34631a );
 a3741a <=( a34620a  and  a34609a );
 a3742a <=( a34598a  and  a34587a );
 a3743a <=( a34576a  and  a34565a );
 a3744a <=( a34554a  and  a34543a );
 a3745a <=( a34532a  and  a34521a );
 a3746a <=( a34510a  and  a34499a );
 a3747a <=( a34488a  and  a34477a );
 a3748a <=( a34466a  and  a34455a );
 a3749a <=( a34444a  and  a34433a );
 a3750a <=( a34422a  and  a34411a );
 a3751a <=( a34400a  and  a34389a );
 a3752a <=( a34378a  and  a34367a );
 a3753a <=( a34356a  and  a34345a );
 a3754a <=( a34334a  and  a34323a );
 a3755a <=( a34312a  and  a34301a );
 a3756a <=( a34290a  and  a34279a );
 a3757a <=( a34268a  and  a34257a );
 a3758a <=( a34246a  and  a34235a );
 a3759a <=( a34224a  and  a34213a );
 a3760a <=( a34202a  and  a34191a );
 a3761a <=( a34180a  and  a34169a );
 a3762a <=( a34158a  and  a34147a );
 a3763a <=( a34136a  and  a34125a );
 a3764a <=( a34114a  and  a34103a );
 a3765a <=( a34092a  and  a34081a );
 a3766a <=( a34070a  and  a34059a );
 a3767a <=( a34048a  and  a34037a );
 a3768a <=( a34026a  and  a34015a );
 a3769a <=( a34004a  and  a33993a );
 a3770a <=( a33982a  and  a33971a );
 a3771a <=( a33960a  and  a33949a );
 a3772a <=( a33938a  and  a33927a );
 a3773a <=( a33916a  and  a33905a );
 a3774a <=( a33894a  and  a33883a );
 a3775a <=( a33872a  and  a33861a );
 a3776a <=( a33850a  and  a33839a );
 a3777a <=( a33828a  and  a33817a );
 a3778a <=( a33806a  and  a33795a );
 a3779a <=( a33784a  and  a33773a );
 a3780a <=( a33762a  and  a33751a );
 a3781a <=( a33740a  and  a33729a );
 a3782a <=( a33718a  and  a33707a );
 a3783a <=( a33696a  and  a33685a );
 a3784a <=( a33674a  and  a33663a );
 a3785a <=( a33652a  and  a33641a );
 a3786a <=( a33630a  and  a33619a );
 a3787a <=( a33608a  and  a33597a );
 a3788a <=( a33586a  and  a33575a );
 a3789a <=( a33564a  and  a33553a );
 a3790a <=( a33542a  and  a33531a );
 a3791a <=( a33520a  and  a33509a );
 a3792a <=( a33498a  and  a33487a );
 a3793a <=( a33476a  and  a33465a );
 a3794a <=( a33454a  and  a33443a );
 a3795a <=( a33432a  and  a33421a );
 a3796a <=( a33410a  and  a33399a );
 a3797a <=( a33388a  and  a33377a );
 a3798a <=( a33366a  and  a33355a );
 a3799a <=( a33344a  and  a33333a );
 a3800a <=( a33322a  and  a33311a );
 a3801a <=( a33300a  and  a33289a );
 a3802a <=( a33278a  and  a33267a );
 a3803a <=( a33256a  and  a33245a );
 a3804a <=( a33234a  and  a33223a );
 a3805a <=( a33212a  and  a33201a );
 a3806a <=( a33190a  and  a33179a );
 a3807a <=( a33168a  and  a33157a );
 a3808a <=( a33146a  and  a33135a );
 a3809a <=( a33124a  and  a33113a );
 a3810a <=( a33102a  and  a33091a );
 a3811a <=( a33080a  and  a33069a );
 a3812a <=( a33058a  and  a33047a );
 a3813a <=( a33036a  and  a33025a );
 a3814a <=( a33014a  and  a33003a );
 a3815a <=( a32992a  and  a32981a );
 a3816a <=( a32970a  and  a32959a );
 a3817a <=( a32948a  and  a32937a );
 a3818a <=( a32926a  and  a32915a );
 a3819a <=( a32904a  and  a32893a );
 a3820a <=( a32882a  and  a32871a );
 a3821a <=( a32860a  and  a32849a );
 a3822a <=( a32838a  and  a32827a );
 a3823a <=( a32816a  and  a32805a );
 a3824a <=( a32794a  and  a32783a );
 a3825a <=( a32772a  and  a32761a );
 a3826a <=( a32750a  and  a32739a );
 a3827a <=( a32728a  and  a32717a );
 a3828a <=( a32706a  and  a32695a );
 a3829a <=( a32684a  and  a32673a );
 a3830a <=( a32662a  and  a32651a );
 a3831a <=( a32640a  and  a32629a );
 a3832a <=( a32618a  and  a32607a );
 a3833a <=( a32596a  and  a32585a );
 a3834a <=( a32574a  and  a32563a );
 a3835a <=( a32552a  and  a32541a );
 a3836a <=( a32530a  and  a32519a );
 a3837a <=( a32508a  and  a32497a );
 a3838a <=( a32486a  and  a32475a );
 a3839a <=( a32464a  and  a32453a );
 a3840a <=( a32442a  and  a32431a );
 a3841a <=( a32420a  and  a32409a );
 a3842a <=( a32398a  and  a32387a );
 a3843a <=( a32376a  and  a32365a );
 a3844a <=( a32354a  and  a32343a );
 a3845a <=( a32332a  and  a32321a );
 a3846a <=( a32310a  and  a32299a );
 a3847a <=( a32288a  and  a32277a );
 a3848a <=( a32266a  and  a32255a );
 a3849a <=( a32244a  and  a32233a );
 a3850a <=( a32222a  and  a32211a );
 a3851a <=( a32200a  and  a32189a );
 a3852a <=( a32178a  and  a32167a );
 a3853a <=( a32156a  and  a32145a );
 a3854a <=( a32134a  and  a32123a );
 a3855a <=( a32112a  and  a32101a );
 a3856a <=( a32090a  and  a32079a );
 a3857a <=( a32068a  and  a32057a );
 a3858a <=( a32046a  and  a32035a );
 a3859a <=( a32024a  and  a32013a );
 a3860a <=( a32002a  and  a31991a );
 a3861a <=( a31980a  and  a31969a );
 a3862a <=( a31958a  and  a31947a );
 a3863a <=( a31936a  and  a31925a );
 a3864a <=( a31914a  and  a31903a );
 a3865a <=( a31892a  and  a31881a );
 a3866a <=( a31870a  and  a31859a );
 a3867a <=( a31848a  and  a31837a );
 a3868a <=( a31826a  and  a31815a );
 a3869a <=( a31804a  and  a31793a );
 a3870a <=( a31782a  and  a31771a );
 a3871a <=( a31760a  and  a31749a );
 a3872a <=( a31738a  and  a31727a );
 a3873a <=( a31716a  and  a31705a );
 a3874a <=( a31694a  and  a31683a );
 a3875a <=( a31672a  and  a31661a );
 a3876a <=( a31650a  and  a31639a );
 a3877a <=( a31628a  and  a31617a );
 a3878a <=( a31606a  and  a31595a );
 a3879a <=( a31584a  and  a31573a );
 a3880a <=( a31562a  and  a31551a );
 a3881a <=( a31540a  and  a31529a );
 a3882a <=( a31518a  and  a31507a );
 a3883a <=( a31496a  and  a31485a );
 a3884a <=( a31474a  and  a31463a );
 a3885a <=( a31452a  and  a31441a );
 a3886a <=( a31430a  and  a31419a );
 a3887a <=( a31408a  and  a31397a );
 a3888a <=( a31386a  and  a31375a );
 a3889a <=( a31364a  and  a31353a );
 a3890a <=( a31342a  and  a31331a );
 a3891a <=( a31320a  and  a31309a );
 a3892a <=( a31298a  and  a31287a );
 a3893a <=( a31276a  and  a31265a );
 a3894a <=( a31254a  and  a31243a );
 a3895a <=( a31232a  and  a31221a );
 a3896a <=( a31210a  and  a31199a );
 a3897a <=( a31188a  and  a31177a );
 a3898a <=( a31166a  and  a31155a );
 a3899a <=( a31144a  and  a31133a );
 a3900a <=( a31122a  and  a31111a );
 a3901a <=( a31100a  and  a31089a );
 a3902a <=( a31078a  and  a31067a );
 a3903a <=( a31056a  and  a31045a );
 a3904a <=( a31034a  and  a31023a );
 a3905a <=( a31012a  and  a31001a );
 a3906a <=( a30990a  and  a30979a );
 a3907a <=( a30968a  and  a30957a );
 a3908a <=( a30946a  and  a30935a );
 a3909a <=( a30924a  and  a30913a );
 a3910a <=( a30902a  and  a30891a );
 a3911a <=( a30880a  and  a30869a );
 a3912a <=( a30858a  and  a30847a );
 a3913a <=( a30836a  and  a30825a );
 a3914a <=( a30814a  and  a30803a );
 a3915a <=( a30792a  and  a30781a );
 a3916a <=( a30770a  and  a30759a );
 a3917a <=( a30748a  and  a30737a );
 a3918a <=( a30726a  and  a30715a );
 a3919a <=( a30704a  and  a30693a );
 a3920a <=( a30682a  and  a30671a );
 a3921a <=( a30660a  and  a30649a );
 a3922a <=( a30638a  and  a30627a );
 a3923a <=( a30616a  and  a30605a );
 a3924a <=( a30594a  and  a30583a );
 a3925a <=( a30572a  and  a30561a );
 a3926a <=( a30550a  and  a30539a );
 a3927a <=( a30528a  and  a30517a );
 a3928a <=( a30506a  and  a30495a );
 a3929a <=( a30484a  and  a30473a );
 a3930a <=( a30462a  and  a30451a );
 a3931a <=( a30440a  and  a30429a );
 a3932a <=( a30418a  and  a30407a );
 a3933a <=( a30396a  and  a30385a );
 a3934a <=( a30374a  and  a30363a );
 a3935a <=( a30352a  and  a30341a );
 a3936a <=( a30330a  and  a30319a );
 a3937a <=( a30308a  and  a30297a );
 a3938a <=( a30286a  and  a30275a );
 a3939a <=( a30264a  and  a30253a );
 a3940a <=( a30242a  and  a30231a );
 a3941a <=( a30220a  and  a30209a );
 a3942a <=( a30198a  and  a30187a );
 a3943a <=( a30176a  and  a30165a );
 a3944a <=( a30154a  and  a30143a );
 a3945a <=( a30132a  and  a30121a );
 a3946a <=( a30110a  and  a30099a );
 a3947a <=( a30088a  and  a30077a );
 a3948a <=( a30066a  and  a30055a );
 a3949a <=( a30044a  and  a30033a );
 a3950a <=( a30022a  and  a30011a );
 a3951a <=( a30000a  and  a29989a );
 a3952a <=( a29978a  and  a29967a );
 a3953a <=( a29956a  and  a29945a );
 a3954a <=( a29934a  and  a29923a );
 a3955a <=( a29912a  and  a29901a );
 a3956a <=( a29890a  and  a29879a );
 a3957a <=( a29868a  and  a29857a );
 a3958a <=( a29846a  and  a29835a );
 a3959a <=( a29824a  and  a29813a );
 a3960a <=( a29802a  and  a29791a );
 a3961a <=( a29780a  and  a29769a );
 a3962a <=( a29758a  and  a29747a );
 a3963a <=( a29736a  and  a29725a );
 a3964a <=( a29714a  and  a29703a );
 a3965a <=( a29692a  and  a29681a );
 a3966a <=( a29670a  and  a29659a );
 a3967a <=( a29648a  and  a29637a );
 a3968a <=( a29626a  and  a29615a );
 a3969a <=( a29604a  and  a29593a );
 a3970a <=( a29582a  and  a29571a );
 a3971a <=( a29560a  and  a29549a );
 a3972a <=( a29538a  and  a29527a );
 a3973a <=( a29516a  and  a29505a );
 a3974a <=( a29494a  and  a29483a );
 a3975a <=( a29472a  and  a29461a );
 a3976a <=( a29450a  and  a29439a );
 a3977a <=( a29428a  and  a29417a );
 a3978a <=( a29406a  and  a29395a );
 a3979a <=( a29384a  and  a29373a );
 a3980a <=( a29362a  and  a29351a );
 a3981a <=( a29340a  and  a29329a );
 a3982a <=( a29318a  and  a29307a );
 a3983a <=( a29296a  and  a29285a );
 a3984a <=( a29274a  and  a29263a );
 a3985a <=( a29252a  and  a29241a );
 a3986a <=( a29230a  and  a29219a );
 a3987a <=( a29208a  and  a29197a );
 a3988a <=( a29186a  and  a29175a );
 a3989a <=( a29164a  and  a29153a );
 a3990a <=( a29142a  and  a29131a );
 a3991a <=( a29120a  and  a29109a );
 a3992a <=( a29098a  and  a29087a );
 a3993a <=( a29076a  and  a29065a );
 a3994a <=( a29054a  and  a29043a );
 a3995a <=( a29032a  and  a29021a );
 a3996a <=( a29010a  and  a28999a );
 a3997a <=( a28988a  and  a28977a );
 a3998a <=( a28966a  and  a28955a );
 a3999a <=( a28944a  and  a28933a );
 a4000a <=( a28922a  and  a28911a );
 a4001a <=( a28900a  and  a28889a );
 a4002a <=( a28878a  and  a28867a );
 a4003a <=( a28856a  and  a28845a );
 a4004a <=( a28834a  and  a28823a );
 a4005a <=( a28812a  and  a28801a );
 a4006a <=( a28790a  and  a28779a );
 a4007a <=( a28768a  and  a28757a );
 a4008a <=( a28746a  and  a28735a );
 a4009a <=( a28724a  and  a28713a );
 a4010a <=( a28702a  and  a28691a );
 a4011a <=( a28680a  and  a28669a );
 a4012a <=( a28658a  and  a28647a );
 a4013a <=( a28636a  and  a28625a );
 a4014a <=( a28614a  and  a28603a );
 a4015a <=( a28592a  and  a28581a );
 a4016a <=( a28570a  and  a28559a );
 a4017a <=( a28548a  and  a28537a );
 a4018a <=( a28526a  and  a28515a );
 a4019a <=( a28504a  and  a28493a );
 a4020a <=( a28482a  and  a28471a );
 a4021a <=( a28460a  and  a28449a );
 a4022a <=( a28438a  and  a28427a );
 a4023a <=( a28416a  and  a28405a );
 a4024a <=( a28394a  and  a28383a );
 a4025a <=( a28372a  and  a28361a );
 a4026a <=( a28350a  and  a28339a );
 a4027a <=( a28328a  and  a28317a );
 a4028a <=( a28306a  and  a28295a );
 a4029a <=( a28284a  and  a28273a );
 a4030a <=( a28262a  and  a28251a );
 a4031a <=( a28240a  and  a28229a );
 a4032a <=( a28218a  and  a28207a );
 a4033a <=( a28196a  and  a28185a );
 a4034a <=( a28174a  and  a28163a );
 a4035a <=( a28152a  and  a28141a );
 a4036a <=( a28130a  and  a28119a );
 a4037a <=( a28108a  and  a28097a );
 a4038a <=( a28086a  and  a28075a );
 a4039a <=( a28064a  and  a28053a );
 a4040a <=( a28042a  and  a28031a );
 a4041a <=( a28020a  and  a28009a );
 a4042a <=( a27998a  and  a27987a );
 a4043a <=( a27976a  and  a27965a );
 a4044a <=( a27954a  and  a27943a );
 a4045a <=( a27932a  and  a27921a );
 a4046a <=( a27910a  and  a27899a );
 a4047a <=( a27888a  and  a27877a );
 a4048a <=( a27866a  and  a27855a );
 a4049a <=( a27844a  and  a27833a );
 a4050a <=( a27822a  and  a27811a );
 a4051a <=( a27800a  and  a27789a );
 a4052a <=( a27778a  and  a27767a );
 a4053a <=( a27756a  and  a27745a );
 a4054a <=( a27734a  and  a27723a );
 a4055a <=( a27712a  and  a27701a );
 a4056a <=( a27690a  and  a27679a );
 a4057a <=( a27668a  and  a27657a );
 a4058a <=( a27646a  and  a27635a );
 a4059a <=( a27624a  and  a27613a );
 a4060a <=( a27602a  and  a27591a );
 a4061a <=( a27580a  and  a27569a );
 a4062a <=( a27558a  and  a27547a );
 a4063a <=( a27536a  and  a27525a );
 a4064a <=( a27514a  and  a27503a );
 a4065a <=( a27492a  and  a27481a );
 a4066a <=( a27470a  and  a27459a );
 a4067a <=( a27448a  and  a27437a );
 a4068a <=( a27426a  and  a27415a );
 a4069a <=( a27404a  and  a27393a );
 a4070a <=( a27382a  and  a27371a );
 a4071a <=( a27360a  and  a27349a );
 a4072a <=( a27338a  and  a27327a );
 a4073a <=( a27316a  and  a27305a );
 a4074a <=( a27294a  and  a27283a );
 a4075a <=( a27272a  and  a27261a );
 a4076a <=( a27250a  and  a27239a );
 a4077a <=( a27228a  and  a27217a );
 a4078a <=( a27206a  and  a27195a );
 a4079a <=( a27184a  and  a27173a );
 a4080a <=( a27162a  and  a27151a );
 a4081a <=( a27140a  and  a27129a );
 a4082a <=( a27118a  and  a27107a );
 a4083a <=( a27096a  and  a27085a );
 a4084a <=( a27074a  and  a27063a );
 a4085a <=( a27052a  and  a27041a );
 a4086a <=( a27030a  and  a27019a );
 a4087a <=( a27008a  and  a26997a );
 a4088a <=( a26986a  and  a26975a );
 a4089a <=( a26964a  and  a26953a );
 a4090a <=( a26942a  and  a26931a );
 a4091a <=( a26920a  and  a26909a );
 a4092a <=( a26898a  and  a26887a );
 a4093a <=( a26876a  and  a26865a );
 a4094a <=( a26854a  and  a26843a );
 a4095a <=( a26832a  and  a26821a );
 a4096a <=( a26810a  and  a26799a );
 a4097a <=( a26788a  and  a26777a );
 a4098a <=( a26766a  and  a26755a );
 a4099a <=( a26744a  and  a26733a );
 a4100a <=( a26722a  and  a26711a );
 a4101a <=( a26700a  and  a26689a );
 a4102a <=( a26678a  and  a26667a );
 a4103a <=( a26656a  and  a26645a );
 a4104a <=( a26634a  and  a26623a );
 a4105a <=( a26612a  and  a26601a );
 a4106a <=( a26590a  and  a26579a );
 a4107a <=( a26568a  and  a26557a );
 a4108a <=( a26546a  and  a26535a );
 a4109a <=( a26524a  and  a26513a );
 a4110a <=( a26502a  and  a26491a );
 a4111a <=( a26480a  and  a26469a );
 a4112a <=( a26458a  and  a26447a );
 a4113a <=( a26436a  and  a26425a );
 a4114a <=( a26414a  and  a26403a );
 a4115a <=( a26392a  and  a26381a );
 a4116a <=( a26370a  and  a26359a );
 a4117a <=( a26348a  and  a26337a );
 a4118a <=( a26326a  and  a26315a );
 a4119a <=( a26304a  and  a26293a );
 a4120a <=( a26282a  and  a26271a );
 a4121a <=( a26260a  and  a26249a );
 a4122a <=( a26238a  and  a26227a );
 a4123a <=( a26216a  and  a26205a );
 a4124a <=( a26194a  and  a26183a );
 a4125a <=( a26172a  and  a26161a );
 a4126a <=( a26150a  and  a26139a );
 a4127a <=( a26128a  and  a26117a );
 a4128a <=( a26106a  and  a26095a );
 a4129a <=( a26084a  and  a26073a );
 a4130a <=( a26062a  and  a26051a );
 a4131a <=( a26040a  and  a26029a );
 a4132a <=( a26018a  and  a26007a );
 a4133a <=( a25996a  and  a25985a );
 a4134a <=( a25974a  and  a25963a );
 a4135a <=( a25952a  and  a25941a );
 a4136a <=( a25930a  and  a25919a );
 a4137a <=( a25908a  and  a25897a );
 a4138a <=( a25886a  and  a25875a );
 a4139a <=( a25864a  and  a25853a );
 a4140a <=( a25842a  and  a25831a );
 a4141a <=( a25820a  and  a25809a );
 a4142a <=( a25798a  and  a25787a );
 a4143a <=( a25776a  and  a25765a );
 a4144a <=( a25754a  and  a25743a );
 a4145a <=( a25732a  and  a25721a );
 a4146a <=( a25710a  and  a25699a );
 a4147a <=( a25688a  and  a25677a );
 a4148a <=( a25666a  and  a25655a );
 a4149a <=( a25644a  and  a25633a );
 a4150a <=( a25622a  and  a25611a );
 a4151a <=( a25600a  and  a25589a );
 a4152a <=( a25578a  and  a25567a );
 a4153a <=( a25556a  and  a25545a );
 a4154a <=( a25534a  and  a25523a );
 a4155a <=( a25512a  and  a25501a );
 a4156a <=( a25490a  and  a25479a );
 a4157a <=( a25468a  and  a25457a );
 a4158a <=( a25446a  and  a25435a );
 a4159a <=( a25424a  and  a25413a );
 a4160a <=( a25402a  and  a25391a );
 a4161a <=( a25380a  and  a25369a );
 a4162a <=( a25358a  and  a25347a );
 a4163a <=( a25336a  and  a25325a );
 a4164a <=( a25314a  and  a25303a );
 a4165a <=( a25292a  and  a25281a );
 a4166a <=( a25270a  and  a25259a );
 a4167a <=( a25248a  and  a25237a );
 a4168a <=( a25226a  and  a25215a );
 a4169a <=( a25204a  and  a25193a );
 a4170a <=( a25184a  and  a25173a );
 a4171a <=( a25164a  and  a25153a );
 a4172a <=( a25144a  and  a25133a );
 a4173a <=( a25124a  and  a25113a );
 a4174a <=( a25104a  and  a25093a );
 a4175a <=( a25084a  and  a25073a );
 a4176a <=( a25064a  and  a25053a );
 a4177a <=( a25044a  and  a25033a );
 a4178a <=( a25024a  and  a25013a );
 a4179a <=( a25004a  and  a24993a );
 a4180a <=( a24984a  and  a24973a );
 a4181a <=( a24964a  and  a24953a );
 a4182a <=( a24944a  and  a24933a );
 a4183a <=( a24924a  and  a24913a );
 a4184a <=( a24904a  and  a24893a );
 a4185a <=( a24884a  and  a24873a );
 a4186a <=( a24864a  and  a24853a );
 a4187a <=( a24844a  and  a24833a );
 a4188a <=( a24824a  and  a24813a );
 a4189a <=( a24804a  and  a24793a );
 a4190a <=( a24784a  and  a24773a );
 a4191a <=( a24764a  and  a24753a );
 a4192a <=( a24744a  and  a24733a );
 a4193a <=( a24724a  and  a24713a );
 a4194a <=( a24704a  and  a24693a );
 a4195a <=( a24684a  and  a24673a );
 a4196a <=( a24664a  and  a24653a );
 a4197a <=( a24644a  and  a24633a );
 a4198a <=( a24624a  and  a24613a );
 a4199a <=( a24604a  and  a24593a );
 a4200a <=( a24584a  and  a24573a );
 a4201a <=( a24564a  and  a24553a );
 a4202a <=( a24544a  and  a24533a );
 a4203a <=( a24524a  and  a24513a );
 a4204a <=( a24504a  and  a24493a );
 a4205a <=( a24484a  and  a24473a );
 a4206a <=( a24464a  and  a24453a );
 a4207a <=( a24444a  and  a24433a );
 a4208a <=( a24424a  and  a24413a );
 a4209a <=( a24404a  and  a24393a );
 a4210a <=( a24384a  and  a24373a );
 a4211a <=( a24364a  and  a24353a );
 a4212a <=( a24344a  and  a24333a );
 a4213a <=( a24324a  and  a24313a );
 a4214a <=( a24304a  and  a24293a );
 a4215a <=( a24284a  and  a24273a );
 a4216a <=( a24264a  and  a24253a );
 a4217a <=( a24244a  and  a24233a );
 a4218a <=( a24224a  and  a24213a );
 a4219a <=( a24204a  and  a24193a );
 a4220a <=( a24184a  and  a24173a );
 a4221a <=( a24164a  and  a24153a );
 a4222a <=( a24144a  and  a24133a );
 a4223a <=( a24124a  and  a24113a );
 a4224a <=( a24104a  and  a24093a );
 a4225a <=( a24084a  and  a24073a );
 a4226a <=( a24064a  and  a24053a );
 a4227a <=( a24044a  and  a24033a );
 a4228a <=( a24024a  and  a24013a );
 a4229a <=( a24004a  and  a23993a );
 a4230a <=( a23984a  and  a23973a );
 a4231a <=( a23964a  and  a23953a );
 a4232a <=( a23944a  and  a23933a );
 a4233a <=( a23924a  and  a23913a );
 a4234a <=( a23904a  and  a23893a );
 a4235a <=( a23884a  and  a23873a );
 a4236a <=( a23864a  and  a23853a );
 a4237a <=( a23844a  and  a23833a );
 a4238a <=( a23824a  and  a23813a );
 a4239a <=( a23804a  and  a23793a );
 a4240a <=( a23784a  and  a23773a );
 a4241a <=( a23764a  and  a23753a );
 a4242a <=( a23744a  and  a23733a );
 a4243a <=( a23724a  and  a23713a );
 a4244a <=( a23704a  and  a23693a );
 a4245a <=( a23684a  and  a23673a );
 a4246a <=( a23664a  and  a23653a );
 a4247a <=( a23644a  and  a23633a );
 a4248a <=( a23624a  and  a23613a );
 a4249a <=( a23604a  and  a23593a );
 a4250a <=( a23584a  and  a23573a );
 a4251a <=( a23564a  and  a23553a );
 a4252a <=( a23544a  and  a23533a );
 a4253a <=( a23524a  and  a23513a );
 a4254a <=( a23504a  and  a23493a );
 a4255a <=( a23484a  and  a23473a );
 a4256a <=( a23464a  and  a23453a );
 a4257a <=( a23444a  and  a23433a );
 a4258a <=( a23424a  and  a23413a );
 a4259a <=( a23404a  and  a23393a );
 a4260a <=( a23384a  and  a23373a );
 a4261a <=( a23364a  and  a23353a );
 a4262a <=( a23344a  and  a23333a );
 a4263a <=( a23324a  and  a23313a );
 a4264a <=( a23304a  and  a23293a );
 a4265a <=( a23284a  and  a23273a );
 a4266a <=( a23264a  and  a23253a );
 a4267a <=( a23244a  and  a23233a );
 a4268a <=( a23224a  and  a23213a );
 a4269a <=( a23204a  and  a23193a );
 a4270a <=( a23184a  and  a23173a );
 a4271a <=( a23164a  and  a23153a );
 a4272a <=( a23144a  and  a23133a );
 a4273a <=( a23124a  and  a23113a );
 a4274a <=( a23104a  and  a23093a );
 a4275a <=( a23084a  and  a23073a );
 a4276a <=( a23064a  and  a23053a );
 a4277a <=( a23044a  and  a23033a );
 a4278a <=( a23024a  and  a23013a );
 a4279a <=( a23004a  and  a22993a );
 a4280a <=( a22984a  and  a22973a );
 a4281a <=( a22964a  and  a22953a );
 a4282a <=( a22944a  and  a22933a );
 a4283a <=( a22924a  and  a22913a );
 a4284a <=( a22904a  and  a22893a );
 a4285a <=( a22884a  and  a22873a );
 a4286a <=( a22864a  and  a22853a );
 a4287a <=( a22844a  and  a22833a );
 a4288a <=( a22824a  and  a22813a );
 a4289a <=( a22804a  and  a22793a );
 a4290a <=( a22784a  and  a22773a );
 a4291a <=( a22764a  and  a22753a );
 a4292a <=( a22744a  and  a22733a );
 a4293a <=( a22724a  and  a22713a );
 a4294a <=( a22704a  and  a22693a );
 a4295a <=( a22684a  and  a22673a );
 a4296a <=( a22664a  and  a22653a );
 a4297a <=( a22644a  and  a22633a );
 a4298a <=( a22624a  and  a22613a );
 a4299a <=( a22604a  and  a22593a );
 a4300a <=( a22584a  and  a22573a );
 a4301a <=( a22564a  and  a22553a );
 a4302a <=( a22544a  and  a22533a );
 a4303a <=( a22524a  and  a22513a );
 a4304a <=( a22504a  and  a22493a );
 a4305a <=( a22484a  and  a22473a );
 a4306a <=( a22464a  and  a22453a );
 a4307a <=( a22444a  and  a22433a );
 a4308a <=( a22424a  and  a22413a );
 a4309a <=( a22404a  and  a22393a );
 a4310a <=( a22384a  and  a22373a );
 a4311a <=( a22364a  and  a22353a );
 a4312a <=( a22344a  and  a22333a );
 a4313a <=( a22324a  and  a22313a );
 a4314a <=( a22304a  and  a22293a );
 a4315a <=( a22284a  and  a22273a );
 a4316a <=( a22264a  and  a22253a );
 a4317a <=( a22244a  and  a22233a );
 a4318a <=( a22224a  and  a22213a );
 a4319a <=( a22204a  and  a22193a );
 a4320a <=( a22184a  and  a22173a );
 a4321a <=( a22164a  and  a22153a );
 a4322a <=( a22144a  and  a22133a );
 a4323a <=( a22124a  and  a22113a );
 a4324a <=( a22104a  and  a22093a );
 a4325a <=( a22084a  and  a22073a );
 a4326a <=( a22064a  and  a22053a );
 a4327a <=( a22044a  and  a22033a );
 a4328a <=( a22024a  and  a22013a );
 a4329a <=( a22004a  and  a21993a );
 a4330a <=( a21984a  and  a21973a );
 a4331a <=( a21964a  and  a21953a );
 a4332a <=( a21944a  and  a21933a );
 a4333a <=( a21924a  and  a21913a );
 a4334a <=( a21904a  and  a21893a );
 a4335a <=( a21884a  and  a21873a );
 a4336a <=( a21864a  and  a21853a );
 a4337a <=( a21844a  and  a21833a );
 a4338a <=( a21824a  and  a21813a );
 a4339a <=( a21804a  and  a21793a );
 a4340a <=( a21784a  and  a21773a );
 a4341a <=( a21764a  and  a21753a );
 a4342a <=( a21744a  and  a21733a );
 a4343a <=( a21724a  and  a21713a );
 a4344a <=( a21704a  and  a21693a );
 a4345a <=( a21684a  and  a21673a );
 a4346a <=( a21664a  and  a21653a );
 a4347a <=( a21644a  and  a21633a );
 a4348a <=( a21624a  and  a21613a );
 a4349a <=( a21604a  and  a21593a );
 a4350a <=( a21584a  and  a21573a );
 a4351a <=( a21564a  and  a21553a );
 a4352a <=( a21544a  and  a21533a );
 a4353a <=( a21524a  and  a21513a );
 a4354a <=( a21504a  and  a21493a );
 a4355a <=( a21484a  and  a21473a );
 a4356a <=( a21464a  and  a21453a );
 a4357a <=( a21444a  and  a21433a );
 a4358a <=( a21424a  and  a21413a );
 a4359a <=( a21404a  and  a21393a );
 a4360a <=( a21384a  and  a21373a );
 a4361a <=( a21364a  and  a21353a );
 a4362a <=( a21344a  and  a21333a );
 a4363a <=( a21324a  and  a21313a );
 a4364a <=( a21304a  and  a21293a );
 a4365a <=( a21284a  and  a21273a );
 a4366a <=( a21264a  and  a21253a );
 a4367a <=( a21244a  and  a21233a );
 a4368a <=( a21224a  and  a21213a );
 a4369a <=( a21204a  and  a21193a );
 a4370a <=( a21184a  and  a21173a );
 a4371a <=( a21164a  and  a21153a );
 a4372a <=( a21144a  and  a21133a );
 a4373a <=( a21124a  and  a21113a );
 a4374a <=( a21104a  and  a21093a );
 a4375a <=( a21084a  and  a21073a );
 a4376a <=( a21064a  and  a21053a );
 a4377a <=( a21044a  and  a21033a );
 a4378a <=( a21024a  and  a21013a );
 a4379a <=( a21004a  and  a20993a );
 a4380a <=( a20984a  and  a20973a );
 a4381a <=( a20964a  and  a20953a );
 a4382a <=( a20944a  and  a20933a );
 a4383a <=( a20924a  and  a20913a );
 a4384a <=( a20904a  and  a20893a );
 a4385a <=( a20884a  and  a20873a );
 a4386a <=( a20864a  and  a20853a );
 a4387a <=( a20844a  and  a20833a );
 a4388a <=( a20824a  and  a20813a );
 a4389a <=( a20804a  and  a20793a );
 a4390a <=( a20784a  and  a20773a );
 a4391a <=( a20764a  and  a20753a );
 a4392a <=( a20744a  and  a20733a );
 a4393a <=( a20724a  and  a20713a );
 a4394a <=( a20704a  and  a20693a );
 a4395a <=( a20684a  and  a20673a );
 a4396a <=( a20664a  and  a20653a );
 a4397a <=( a20644a  and  a20633a );
 a4398a <=( a20624a  and  a20613a );
 a4399a <=( a20604a  and  a20593a );
 a4400a <=( a20584a  and  a20573a );
 a4401a <=( a20564a  and  a20553a );
 a4402a <=( a20544a  and  a20533a );
 a4403a <=( a20524a  and  a20513a );
 a4404a <=( a20504a  and  a20493a );
 a4405a <=( a20484a  and  a20473a );
 a4406a <=( a20464a  and  a20453a );
 a4407a <=( a20444a  and  a20433a );
 a4408a <=( a20424a  and  a20413a );
 a4409a <=( a20404a  and  a20393a );
 a4410a <=( a20384a  and  a20373a );
 a4411a <=( a20364a  and  a20353a );
 a4412a <=( a20344a  and  a20333a );
 a4413a <=( a20324a  and  a20313a );
 a4414a <=( a20304a  and  a20293a );
 a4415a <=( a20284a  and  a20273a );
 a4416a <=( a20264a  and  a20253a );
 a4417a <=( a20244a  and  a20233a );
 a4418a <=( a20224a  and  a20213a );
 a4419a <=( a20204a  and  a20193a );
 a4420a <=( a20184a  and  a20173a );
 a4421a <=( a20164a  and  a20153a );
 a4422a <=( a20144a  and  a20133a );
 a4423a <=( a20124a  and  a20113a );
 a4424a <=( a20104a  and  a20093a );
 a4425a <=( a20084a  and  a20073a );
 a4426a <=( a20064a  and  a20053a );
 a4427a <=( a20044a  and  a20033a );
 a4428a <=( a20024a  and  a20013a );
 a4429a <=( a20004a  and  a19993a );
 a4430a <=( a19984a  and  a19973a );
 a4431a <=( a19964a  and  a19953a );
 a4432a <=( a19944a  and  a19933a );
 a4433a <=( a19924a  and  a19913a );
 a4434a <=( a19904a  and  a19893a );
 a4435a <=( a19884a  and  a19873a );
 a4436a <=( a19864a  and  a19853a );
 a4437a <=( a19844a  and  a19833a );
 a4438a <=( a19824a  and  a19813a );
 a4439a <=( a19804a  and  a19793a );
 a4440a <=( a19784a  and  a19773a );
 a4441a <=( a19764a  and  a19753a );
 a4442a <=( a19744a  and  a19733a );
 a4443a <=( a19724a  and  a19713a );
 a4444a <=( a19704a  and  a19693a );
 a4445a <=( a19684a  and  a19673a );
 a4446a <=( a19664a  and  a19653a );
 a4447a <=( a19644a  and  a19633a );
 a4448a <=( a19624a  and  a19613a );
 a4449a <=( a19604a  and  a19593a );
 a4450a <=( a19584a  and  a19573a );
 a4451a <=( a19564a  and  a19553a );
 a4452a <=( a19544a  and  a19533a );
 a4453a <=( a19524a  and  a19513a );
 a4454a <=( a19504a  and  a19493a );
 a4455a <=( a19484a  and  a19473a );
 a4456a <=( a19464a  and  a19453a );
 a4457a <=( a19444a  and  a19433a );
 a4458a <=( a19424a  and  a19413a );
 a4459a <=( a19404a  and  a19393a );
 a4460a <=( a19384a  and  a19373a );
 a4461a <=( a19364a  and  a19353a );
 a4462a <=( a19344a  and  a19333a );
 a4463a <=( a19324a  and  a19313a );
 a4464a <=( a19304a  and  a19293a );
 a4465a <=( a19284a  and  a19273a );
 a4466a <=( a19264a  and  a19253a );
 a4467a <=( a19244a  and  a19233a );
 a4468a <=( a19224a  and  a19213a );
 a4469a <=( a19204a  and  a19193a );
 a4470a <=( a19184a  and  a19173a );
 a4471a <=( a19164a  and  a19153a );
 a4472a <=( a19144a  and  a19133a );
 a4473a <=( a19124a  and  a19113a );
 a4474a <=( a19104a  and  a19093a );
 a4475a <=( a19084a  and  a19073a );
 a4476a <=( a19064a  and  a19053a );
 a4477a <=( a19044a  and  a19033a );
 a4478a <=( a19024a  and  a19013a );
 a4479a <=( a19004a  and  a18993a );
 a4480a <=( a18984a  and  a18973a );
 a4481a <=( a18964a  and  a18953a );
 a4482a <=( a18944a  and  a18933a );
 a4483a <=( a18924a  and  a18913a );
 a4484a <=( a18904a  and  a18893a );
 a4485a <=( a18884a  and  a18873a );
 a4486a <=( a18864a  and  a18853a );
 a4487a <=( a18844a  and  a18833a );
 a4488a <=( a18824a  and  a18813a );
 a4489a <=( a18804a  and  a18793a );
 a4490a <=( a18784a  and  a18773a );
 a4491a <=( a18764a  and  a18753a );
 a4492a <=( a18744a  and  a18733a );
 a4493a <=( a18724a  and  a18713a );
 a4494a <=( a18704a  and  a18693a );
 a4495a <=( a18684a  and  a18673a );
 a4496a <=( a18664a  and  a18653a );
 a4497a <=( a18644a  and  a18633a );
 a4498a <=( a18624a  and  a18613a );
 a4499a <=( a18604a  and  a18593a );
 a4500a <=( a18584a  and  a18573a );
 a4501a <=( a18564a  and  a18553a );
 a4502a <=( a18544a  and  a18533a );
 a4503a <=( a18524a  and  a18513a );
 a4504a <=( a18504a  and  a18493a );
 a4505a <=( a18484a  and  a18473a );
 a4506a <=( a18464a  and  a18453a );
 a4507a <=( a18444a  and  a18433a );
 a4508a <=( a18424a  and  a18413a );
 a4509a <=( a18404a  and  a18393a );
 a4510a <=( a18384a  and  a18373a );
 a4511a <=( a18364a  and  a18353a );
 a4512a <=( a18344a  and  a18333a );
 a4513a <=( a18324a  and  a18313a );
 a4514a <=( a18304a  and  a18293a );
 a4515a <=( a18284a  and  a18273a );
 a4516a <=( a18264a  and  a18253a );
 a4517a <=( a18244a  and  a18233a );
 a4518a <=( a18224a  and  a18213a );
 a4519a <=( a18204a  and  a18193a );
 a4520a <=( a18184a  and  a18173a );
 a4521a <=( a18164a  and  a18153a );
 a4522a <=( a18144a  and  a18133a );
 a4523a <=( a18124a  and  a18113a );
 a4524a <=( a18104a  and  a18093a );
 a4525a <=( a18084a  and  a18073a );
 a4526a <=( a18064a  and  a18053a );
 a4527a <=( a18044a  and  a18033a );
 a4528a <=( a18024a  and  a18013a );
 a4529a <=( a18004a  and  a17993a );
 a4530a <=( a17984a  and  a17973a );
 a4531a <=( a17964a  and  a17953a );
 a4532a <=( a17944a  and  a17933a );
 a4533a <=( a17924a  and  a17913a );
 a4534a <=( a17904a  and  a17893a );
 a4535a <=( a17884a  and  a17873a );
 a4536a <=( a17864a  and  a17853a );
 a4537a <=( a17844a  and  a17835a );
 a4538a <=( a17826a  and  a17817a );
 a4539a <=( a17808a  and  a17799a );
 a4540a <=( a17790a  and  a17781a );
 a4541a <=( a17772a  and  a17763a );
 a4542a <=( a17754a  and  a17745a );
 a4543a <=( a17736a  and  a17727a );
 a4544a <=( a17718a  and  a17709a );
 a4545a <=( a17700a  and  a17691a );
 a4546a <=( a17682a  and  a17673a );
 a4547a <=( a17664a  and  a17655a );
 a4548a <=( a17646a  and  a17637a );
 a4549a <=( a17628a  and  a17619a );
 a4550a <=( a17610a  and  a17601a );
 a4551a <=( a17592a  and  a17583a );
 a4552a <=( a17574a  and  a17565a );
 a4553a <=( a17556a  and  a17547a );
 a4554a <=( a17538a  and  a17529a );
 a4555a <=( a17520a  and  a17511a );
 a4556a <=( a17502a  and  a17493a );
 a4557a <=( a17484a  and  a17475a );
 a4558a <=( a17466a  and  a17457a );
 a4559a <=( a17448a  and  a17439a );
 a4560a <=( a17430a  and  a17421a );
 a4561a <=( a17412a  and  a17403a );
 a4562a <=( a17394a  and  a17385a );
 a4563a <=( a17376a  and  a17367a );
 a4564a <=( a17358a  and  a17349a );
 a4565a <=( a17340a  and  a17331a );
 a4566a <=( a17322a  and  a17313a );
 a4567a <=( a17304a  and  a17295a );
 a4568a <=( a17286a  and  a17277a );
 a4569a <=( a17268a  and  a17259a );
 a4570a <=( a17250a  and  a17241a );
 a4571a <=( a17232a  and  a17223a );
 a4572a <=( a17214a  and  a17205a );
 a4573a <=( a17196a  and  a17187a );
 a4574a <=( a17178a  and  a17169a );
 a4575a <=( a17160a  and  a17151a );
 a4576a <=( a17142a  and  a17133a );
 a4577a <=( a17124a  and  a17115a );
 a4578a <=( a17106a  and  a17097a );
 a4579a <=( a17088a  and  a17079a );
 a4580a <=( a17070a  and  a17061a );
 a4581a <=( a17052a  and  a17043a );
 a4582a <=( a17034a  and  a17025a );
 a4583a <=( a17016a  and  a17007a );
 a4584a <=( a16998a  and  a16989a );
 a4585a <=( a16980a  and  a16971a );
 a4586a <=( a16962a  and  a16953a );
 a4587a <=( a16944a  and  a16935a );
 a4588a <=( a16926a  and  a16917a );
 a4589a <=( a16908a  and  a16899a );
 a4590a <=( a16890a  and  a16881a );
 a4591a <=( a16872a  and  a16863a );
 a4592a <=( a16854a  and  a16845a );
 a4593a <=( a16836a  and  a16827a );
 a4594a <=( a16818a  and  a16809a );
 a4595a <=( a16800a  and  a16791a );
 a4596a <=( a16782a  and  a16773a );
 a4597a <=( a16764a  and  a16755a );
 a4598a <=( a16746a  and  a16737a );
 a4599a <=( a16728a  and  a16719a );
 a4600a <=( a16710a  and  a16701a );
 a4601a <=( a16692a  and  a16683a );
 a4602a <=( a16674a  and  a16665a );
 a4603a <=( a16656a  and  a16647a );
 a4604a <=( a16638a  and  a16629a );
 a4605a <=( a16620a  and  a16611a );
 a4606a <=( a16602a  and  a16593a );
 a4607a <=( a16584a  and  a16575a );
 a4608a <=( a16566a  and  a16557a );
 a4609a <=( a16548a  and  a16539a );
 a4610a <=( a16530a  and  a16521a );
 a4611a <=( a16512a  and  a16503a );
 a4612a <=( a16494a  and  a16485a );
 a4613a <=( a16476a  and  a16467a );
 a4614a <=( a16458a  and  a16449a );
 a4615a <=( a16440a  and  a16431a );
 a4616a <=( a16422a  and  a16413a );
 a4617a <=( a16404a  and  a16395a );
 a4618a <=( a16386a  and  a16377a );
 a4619a <=( a16368a  and  a16359a );
 a4620a <=( a16350a  and  a16341a );
 a4621a <=( a16332a  and  a16323a );
 a4622a <=( a16314a  and  a16305a );
 a4623a <=( a16296a  and  a16287a );
 a4624a <=( a16278a  and  a16269a );
 a4625a <=( a16260a  and  a16251a );
 a4626a <=( a16242a  and  a16233a );
 a4627a <=( a16224a  and  a16215a );
 a4628a <=( a16206a  and  a16197a );
 a4629a <=( a16188a  and  a16179a );
 a4630a <=( a16170a  and  a16161a );
 a4631a <=( a16152a  and  a16143a );
 a4632a <=( a16134a  and  a16125a );
 a4633a <=( a16116a  and  a16107a );
 a4634a <=( a16098a  and  a16089a );
 a4635a <=( a16080a  and  a16071a );
 a4636a <=( a16062a  and  a16053a );
 a4637a <=( a16044a  and  a16035a );
 a4638a <=( a16026a  and  a16017a );
 a4639a <=( a16008a  and  a15999a );
 a4640a <=( a15990a  and  a15981a );
 a4641a <=( a15972a  and  a15963a );
 a4642a <=( a15954a  and  a15945a );
 a4643a <=( a15936a  and  a15927a );
 a4644a <=( a15918a  and  a15909a );
 a4645a <=( a15900a  and  a15891a );
 a4646a <=( a15882a  and  a15873a );
 a4647a <=( a15864a  and  a15855a );
 a4648a <=( a15846a  and  a15837a );
 a4649a <=( a15828a  and  a15819a );
 a4650a <=( a15810a  and  a15801a );
 a4651a <=( a15792a  and  a15783a );
 a4652a <=( a15774a  and  a15765a );
 a4653a <=( a15756a  and  a15747a );
 a4654a <=( a15738a  and  a15729a );
 a4655a <=( a15720a  and  a15711a );
 a4656a <=( a15702a  and  a15693a );
 a4657a <=( a15684a  and  a15675a );
 a4658a <=( a15666a  and  a15657a );
 a4659a <=( a15648a  and  a15639a );
 a4660a <=( a15630a  and  a15621a );
 a4661a <=( a15612a  and  a15603a );
 a4662a <=( a15594a  and  a15585a );
 a4663a <=( a15576a  and  a15567a );
 a4664a <=( a15558a  and  a15549a );
 a4665a <=( a15540a  and  a15531a );
 a4666a <=( a15522a  and  a15513a );
 a4667a <=( a15504a  and  a15495a );
 a4668a <=( a15486a  and  a15477a );
 a4669a <=( a15468a  and  a15459a );
 a4670a <=( a15450a  and  a15441a );
 a4671a <=( a15432a  and  a15423a );
 a4672a <=( a15414a  and  a15405a );
 a4673a <=( a15396a  and  a15387a );
 a4674a <=( a15380a  and  a15371a );
 a4675a <=( a15364a  and  a15355a );
 a4676a <=( a15348a  and  a15339a );
 a4677a <=( a15332a  and  a15323a );
 a4678a <=( a15316a  and  a15307a );
 a4679a <=( a15300a  and  a15291a );
 a4680a <=( a15284a  and  a15275a );
 a4681a <=( a15268a  and  a15259a );
 a4682a <=( a15252a  and  a15243a );
 a4683a <=( a15236a  and  a15227a );
 a4684a <=( a15220a  and  a15211a );
 a4685a <=( a15204a  and  a15195a );
 a4686a <=( a15188a  and  a15179a );
 a4687a <=( a15172a  and  a15163a );
 a4688a <=( a15156a  and  a15147a );
 a4689a <=( a15140a  and  a15131a );
 a4690a <=( a15124a  and  a15115a );
 a4691a <=( a15108a  and  a15099a );
 a4692a <=( a15092a  and  a15083a );
 a4693a <=( a15076a  and  a15067a );
 a4694a <=( a15060a  and  a15051a );
 a4695a <=( a15044a  and  a15035a );
 a4696a <=( a15028a  and  a15019a );
 a4697a <=( a15012a  and  a15003a );
 a4698a <=( a14996a  and  a14987a );
 a4699a <=( a14980a  and  a14971a );
 a4700a <=( a14964a  and  a14955a );
 a4701a <=( a14948a  and  a14939a );
 a4702a <=( a14932a  and  a14923a );
 a4703a <=( a14916a  and  a14907a );
 a4704a <=( a14900a  and  a14891a );
 a4705a <=( a14884a  and  a14877a );
 a4706a <=( a14870a  and  a14863a );
 a4707a <=( a14856a  and  a14849a );
 a4708a <=( a14842a  and  a14835a );
 a4709a <=( a14828a  and  a14821a );
 a4710a <=( a14814a  and  a14807a );
 a4711a <=( a14800a  and  a14793a );
 a4712a <=( a14786a  and  a14779a );
 a4713a <=( a14772a  and  a14765a );
 a4714a <=( a14758a  and  a14751a );
 a4715a <=( a14744a  and  a14737a );
 a4716a <=( a14730a  and  a14723a );
 a4717a <=( a14716a  and  a14709a );
 a4718a <=( a14702a  and  a14695a );
 a4719a <=( a14688a  and  a14681a );
 a4720a <=( a14674a  and  a14667a );
 a4721a <=( a14660a  and  a14653a );
 a4722a <=( a14646a  and  a14639a );
 a4723a <=( a14632a  and  a14625a );
 a4724a <=( a14618a  and  a14611a );
 a4725a <=( a14604a  and  a14597a );
 a4726a <=( a14590a  and  a14583a );
 a4727a <=( a14576a  and  a14569a );
 a4728a <=( a14562a  and  a14555a );
 a4729a <=( a14548a  and  a14543a );
 a4730a <=( a14538a  and  a14533a );
 a4731a <=( a14528a  and  a14523a );
 a4732a <=( a14518a  and  a14513a );
 a4733a <=( a14508a  and  a14503a );
 a4734a <=( a14498a  and  a14493a );
 a4735a <=( a14488a  and  a14483a );
 a4736a <=( a14478a  and  a14473a );
 a4737a <=( a14468a  and  a14463a );
 a4738a <=( a14458a  and  a14453a );
 a4739a <=( a14448a  and  a14443a );
 a4740a <=( a14438a  and  a14433a );
 a4741a <=( a14428a  and  a14423a );
 a4742a <=( a14418a  and  a14413a );
 a4743a <=( a14408a  and  a14403a );
 a4744a <=( a14398a  and  a14393a );
 a4745a <=( a14388a  and  a14383a );
 a4746a <=( a14378a  and  a14373a );
 a4747a <=( a14368a  and  a14363a );
 a4748a <=( a14358a  and  a14353a );
 a4749a <=( a14348a  and  a14343a );
 a4750a <=( a14338a  and  a14333a );
 a4751a <=( a14328a  and  a14323a );
 a4752a <=( a14318a  and  a14313a );
 a4753a <=( a14308a  and  a14305a );
 a4754a <=( a14302a  and  a14299a );
 a4755a <=( a14296a  and  a14293a );
 a4756a <=( a14290a  and  a14287a );
 a4757a <=( a14284a  and  a14281a );
 a4758a <=( a14278a  and  a14275a );
 a4761a <=( a4757a ) or ( a4758a );
 a4764a <=( a4755a ) or ( a4756a );
 a4765a <=( a4764a ) or ( a4761a );
 a4768a <=( a4753a ) or ( a4754a );
 a4772a <=( a4750a ) or ( a4751a );
 a4773a <=( a4752a ) or ( a4772a );
 a4774a <=( a4773a ) or ( a4768a );
 a4775a <=( a4774a ) or ( a4765a );
 a4778a <=( a4748a ) or ( a4749a );
 a4781a <=( a4746a ) or ( a4747a );
 a4782a <=( a4781a ) or ( a4778a );
 a4785a <=( a4744a ) or ( a4745a );
 a4789a <=( a4741a ) or ( a4742a );
 a4790a <=( a4743a ) or ( a4789a );
 a4791a <=( a4790a ) or ( a4785a );
 a4792a <=( a4791a ) or ( a4782a );
 a4793a <=( a4792a ) or ( a4775a );
 a4796a <=( a4739a ) or ( a4740a );
 a4799a <=( a4737a ) or ( a4738a );
 a4800a <=( a4799a ) or ( a4796a );
 a4803a <=( a4735a ) or ( a4736a );
 a4807a <=( a4732a ) or ( a4733a );
 a4808a <=( a4734a ) or ( a4807a );
 a4809a <=( a4808a ) or ( a4803a );
 a4810a <=( a4809a ) or ( a4800a );
 a4813a <=( a4730a ) or ( a4731a );
 a4817a <=( a4727a ) or ( a4728a );
 a4818a <=( a4729a ) or ( a4817a );
 a4819a <=( a4818a ) or ( a4813a );
 a4822a <=( a4725a ) or ( a4726a );
 a4826a <=( a4722a ) or ( a4723a );
 a4827a <=( a4724a ) or ( a4826a );
 a4828a <=( a4827a ) or ( a4822a );
 a4829a <=( a4828a ) or ( a4819a );
 a4830a <=( a4829a ) or ( a4810a );
 a4831a <=( a4830a ) or ( a4793a );
 a4834a <=( a4720a ) or ( a4721a );
 a4837a <=( a4718a ) or ( a4719a );
 a4838a <=( a4837a ) or ( a4834a );
 a4841a <=( a4716a ) or ( a4717a );
 a4845a <=( a4713a ) or ( a4714a );
 a4846a <=( a4715a ) or ( a4845a );
 a4847a <=( a4846a ) or ( a4841a );
 a4848a <=( a4847a ) or ( a4838a );
 a4851a <=( a4711a ) or ( a4712a );
 a4854a <=( a4709a ) or ( a4710a );
 a4855a <=( a4854a ) or ( a4851a );
 a4858a <=( a4707a ) or ( a4708a );
 a4862a <=( a4704a ) or ( a4705a );
 a4863a <=( a4706a ) or ( a4862a );
 a4864a <=( a4863a ) or ( a4858a );
 a4865a <=( a4864a ) or ( a4855a );
 a4866a <=( a4865a ) or ( a4848a );
 a4869a <=( a4702a ) or ( a4703a );
 a4872a <=( a4700a ) or ( a4701a );
 a4873a <=( a4872a ) or ( a4869a );
 a4876a <=( a4698a ) or ( a4699a );
 a4880a <=( a4695a ) or ( a4696a );
 a4881a <=( a4697a ) or ( a4880a );
 a4882a <=( a4881a ) or ( a4876a );
 a4883a <=( a4882a ) or ( a4873a );
 a4886a <=( a4693a ) or ( a4694a );
 a4890a <=( a4690a ) or ( a4691a );
 a4891a <=( a4692a ) or ( a4890a );
 a4892a <=( a4891a ) or ( a4886a );
 a4895a <=( a4688a ) or ( a4689a );
 a4899a <=( a4685a ) or ( a4686a );
 a4900a <=( a4687a ) or ( a4899a );
 a4901a <=( a4900a ) or ( a4895a );
 a4902a <=( a4901a ) or ( a4892a );
 a4903a <=( a4902a ) or ( a4883a );
 a4904a <=( a4903a ) or ( a4866a );
 a4905a <=( a4904a ) or ( a4831a );
 a4908a <=( a4683a ) or ( a4684a );
 a4911a <=( a4681a ) or ( a4682a );
 a4912a <=( a4911a ) or ( a4908a );
 a4915a <=( a4679a ) or ( a4680a );
 a4919a <=( a4676a ) or ( a4677a );
 a4920a <=( a4678a ) or ( a4919a );
 a4921a <=( a4920a ) or ( a4915a );
 a4922a <=( a4921a ) or ( a4912a );
 a4925a <=( a4674a ) or ( a4675a );
 a4928a <=( a4672a ) or ( a4673a );
 a4929a <=( a4928a ) or ( a4925a );
 a4932a <=( a4670a ) or ( a4671a );
 a4936a <=( a4667a ) or ( a4668a );
 a4937a <=( a4669a ) or ( a4936a );
 a4938a <=( a4937a ) or ( a4932a );
 a4939a <=( a4938a ) or ( a4929a );
 a4940a <=( a4939a ) or ( a4922a );
 a4943a <=( a4665a ) or ( a4666a );
 a4946a <=( a4663a ) or ( a4664a );
 a4947a <=( a4946a ) or ( a4943a );
 a4950a <=( a4661a ) or ( a4662a );
 a4954a <=( a4658a ) or ( a4659a );
 a4955a <=( a4660a ) or ( a4954a );
 a4956a <=( a4955a ) or ( a4950a );
 a4957a <=( a4956a ) or ( a4947a );
 a4960a <=( a4656a ) or ( a4657a );
 a4964a <=( a4653a ) or ( a4654a );
 a4965a <=( a4655a ) or ( a4964a );
 a4966a <=( a4965a ) or ( a4960a );
 a4969a <=( a4651a ) or ( a4652a );
 a4973a <=( a4648a ) or ( a4649a );
 a4974a <=( a4650a ) or ( a4973a );
 a4975a <=( a4974a ) or ( a4969a );
 a4976a <=( a4975a ) or ( a4966a );
 a4977a <=( a4976a ) or ( a4957a );
 a4978a <=( a4977a ) or ( a4940a );
 a4981a <=( a4646a ) or ( a4647a );
 a4984a <=( a4644a ) or ( a4645a );
 a4985a <=( a4984a ) or ( a4981a );
 a4988a <=( a4642a ) or ( a4643a );
 a4992a <=( a4639a ) or ( a4640a );
 a4993a <=( a4641a ) or ( a4992a );
 a4994a <=( a4993a ) or ( a4988a );
 a4995a <=( a4994a ) or ( a4985a );
 a4998a <=( a4637a ) or ( a4638a );
 a5001a <=( a4635a ) or ( a4636a );
 a5002a <=( a5001a ) or ( a4998a );
 a5005a <=( a4633a ) or ( a4634a );
 a5009a <=( a4630a ) or ( a4631a );
 a5010a <=( a4632a ) or ( a5009a );
 a5011a <=( a5010a ) or ( a5005a );
 a5012a <=( a5011a ) or ( a5002a );
 a5013a <=( a5012a ) or ( a4995a );
 a5016a <=( a4628a ) or ( a4629a );
 a5019a <=( a4626a ) or ( a4627a );
 a5020a <=( a5019a ) or ( a5016a );
 a5023a <=( a4624a ) or ( a4625a );
 a5027a <=( a4621a ) or ( a4622a );
 a5028a <=( a4623a ) or ( a5027a );
 a5029a <=( a5028a ) or ( a5023a );
 a5030a <=( a5029a ) or ( a5020a );
 a5033a <=( a4619a ) or ( a4620a );
 a5037a <=( a4616a ) or ( a4617a );
 a5038a <=( a4618a ) or ( a5037a );
 a5039a <=( a5038a ) or ( a5033a );
 a5042a <=( a4614a ) or ( a4615a );
 a5046a <=( a4611a ) or ( a4612a );
 a5047a <=( a4613a ) or ( a5046a );
 a5048a <=( a5047a ) or ( a5042a );
 a5049a <=( a5048a ) or ( a5039a );
 a5050a <=( a5049a ) or ( a5030a );
 a5051a <=( a5050a ) or ( a5013a );
 a5052a <=( a5051a ) or ( a4978a );
 a5053a <=( a5052a ) or ( a4905a );
 a5056a <=( a4609a ) or ( a4610a );
 a5059a <=( a4607a ) or ( a4608a );
 a5060a <=( a5059a ) or ( a5056a );
 a5063a <=( a4605a ) or ( a4606a );
 a5067a <=( a4602a ) or ( a4603a );
 a5068a <=( a4604a ) or ( a5067a );
 a5069a <=( a5068a ) or ( a5063a );
 a5070a <=( a5069a ) or ( a5060a );
 a5073a <=( a4600a ) or ( a4601a );
 a5076a <=( a4598a ) or ( a4599a );
 a5077a <=( a5076a ) or ( a5073a );
 a5080a <=( a4596a ) or ( a4597a );
 a5084a <=( a4593a ) or ( a4594a );
 a5085a <=( a4595a ) or ( a5084a );
 a5086a <=( a5085a ) or ( a5080a );
 a5087a <=( a5086a ) or ( a5077a );
 a5088a <=( a5087a ) or ( a5070a );
 a5091a <=( a4591a ) or ( a4592a );
 a5094a <=( a4589a ) or ( a4590a );
 a5095a <=( a5094a ) or ( a5091a );
 a5098a <=( a4587a ) or ( a4588a );
 a5102a <=( a4584a ) or ( a4585a );
 a5103a <=( a4586a ) or ( a5102a );
 a5104a <=( a5103a ) or ( a5098a );
 a5105a <=( a5104a ) or ( a5095a );
 a5108a <=( a4582a ) or ( a4583a );
 a5112a <=( a4579a ) or ( a4580a );
 a5113a <=( a4581a ) or ( a5112a );
 a5114a <=( a5113a ) or ( a5108a );
 a5117a <=( a4577a ) or ( a4578a );
 a5121a <=( a4574a ) or ( a4575a );
 a5122a <=( a4576a ) or ( a5121a );
 a5123a <=( a5122a ) or ( a5117a );
 a5124a <=( a5123a ) or ( a5114a );
 a5125a <=( a5124a ) or ( a5105a );
 a5126a <=( a5125a ) or ( a5088a );
 a5129a <=( a4572a ) or ( a4573a );
 a5132a <=( a4570a ) or ( a4571a );
 a5133a <=( a5132a ) or ( a5129a );
 a5136a <=( a4568a ) or ( a4569a );
 a5140a <=( a4565a ) or ( a4566a );
 a5141a <=( a4567a ) or ( a5140a );
 a5142a <=( a5141a ) or ( a5136a );
 a5143a <=( a5142a ) or ( a5133a );
 a5146a <=( a4563a ) or ( a4564a );
 a5149a <=( a4561a ) or ( a4562a );
 a5150a <=( a5149a ) or ( a5146a );
 a5153a <=( a4559a ) or ( a4560a );
 a5157a <=( a4556a ) or ( a4557a );
 a5158a <=( a4558a ) or ( a5157a );
 a5159a <=( a5158a ) or ( a5153a );
 a5160a <=( a5159a ) or ( a5150a );
 a5161a <=( a5160a ) or ( a5143a );
 a5164a <=( a4554a ) or ( a4555a );
 a5167a <=( a4552a ) or ( a4553a );
 a5168a <=( a5167a ) or ( a5164a );
 a5171a <=( a4550a ) or ( a4551a );
 a5175a <=( a4547a ) or ( a4548a );
 a5176a <=( a4549a ) or ( a5175a );
 a5177a <=( a5176a ) or ( a5171a );
 a5178a <=( a5177a ) or ( a5168a );
 a5181a <=( a4545a ) or ( a4546a );
 a5185a <=( a4542a ) or ( a4543a );
 a5186a <=( a4544a ) or ( a5185a );
 a5187a <=( a5186a ) or ( a5181a );
 a5190a <=( a4540a ) or ( a4541a );
 a5194a <=( a4537a ) or ( a4538a );
 a5195a <=( a4539a ) or ( a5194a );
 a5196a <=( a5195a ) or ( a5190a );
 a5197a <=( a5196a ) or ( a5187a );
 a5198a <=( a5197a ) or ( a5178a );
 a5199a <=( a5198a ) or ( a5161a );
 a5200a <=( a5199a ) or ( a5126a );
 a5203a <=( a4535a ) or ( a4536a );
 a5206a <=( a4533a ) or ( a4534a );
 a5207a <=( a5206a ) or ( a5203a );
 a5210a <=( a4531a ) or ( a4532a );
 a5214a <=( a4528a ) or ( a4529a );
 a5215a <=( a4530a ) or ( a5214a );
 a5216a <=( a5215a ) or ( a5210a );
 a5217a <=( a5216a ) or ( a5207a );
 a5220a <=( a4526a ) or ( a4527a );
 a5223a <=( a4524a ) or ( a4525a );
 a5224a <=( a5223a ) or ( a5220a );
 a5227a <=( a4522a ) or ( a4523a );
 a5231a <=( a4519a ) or ( a4520a );
 a5232a <=( a4521a ) or ( a5231a );
 a5233a <=( a5232a ) or ( a5227a );
 a5234a <=( a5233a ) or ( a5224a );
 a5235a <=( a5234a ) or ( a5217a );
 a5238a <=( a4517a ) or ( a4518a );
 a5241a <=( a4515a ) or ( a4516a );
 a5242a <=( a5241a ) or ( a5238a );
 a5245a <=( a4513a ) or ( a4514a );
 a5249a <=( a4510a ) or ( a4511a );
 a5250a <=( a4512a ) or ( a5249a );
 a5251a <=( a5250a ) or ( a5245a );
 a5252a <=( a5251a ) or ( a5242a );
 a5255a <=( a4508a ) or ( a4509a );
 a5259a <=( a4505a ) or ( a4506a );
 a5260a <=( a4507a ) or ( a5259a );
 a5261a <=( a5260a ) or ( a5255a );
 a5264a <=( a4503a ) or ( a4504a );
 a5268a <=( a4500a ) or ( a4501a );
 a5269a <=( a4502a ) or ( a5268a );
 a5270a <=( a5269a ) or ( a5264a );
 a5271a <=( a5270a ) or ( a5261a );
 a5272a <=( a5271a ) or ( a5252a );
 a5273a <=( a5272a ) or ( a5235a );
 a5276a <=( a4498a ) or ( a4499a );
 a5279a <=( a4496a ) or ( a4497a );
 a5280a <=( a5279a ) or ( a5276a );
 a5283a <=( a4494a ) or ( a4495a );
 a5287a <=( a4491a ) or ( a4492a );
 a5288a <=( a4493a ) or ( a5287a );
 a5289a <=( a5288a ) or ( a5283a );
 a5290a <=( a5289a ) or ( a5280a );
 a5293a <=( a4489a ) or ( a4490a );
 a5297a <=( a4486a ) or ( a4487a );
 a5298a <=( a4488a ) or ( a5297a );
 a5299a <=( a5298a ) or ( a5293a );
 a5302a <=( a4484a ) or ( a4485a );
 a5306a <=( a4481a ) or ( a4482a );
 a5307a <=( a4483a ) or ( a5306a );
 a5308a <=( a5307a ) or ( a5302a );
 a5309a <=( a5308a ) or ( a5299a );
 a5310a <=( a5309a ) or ( a5290a );
 a5313a <=( a4479a ) or ( a4480a );
 a5316a <=( a4477a ) or ( a4478a );
 a5317a <=( a5316a ) or ( a5313a );
 a5320a <=( a4475a ) or ( a4476a );
 a5324a <=( a4472a ) or ( a4473a );
 a5325a <=( a4474a ) or ( a5324a );
 a5326a <=( a5325a ) or ( a5320a );
 a5327a <=( a5326a ) or ( a5317a );
 a5330a <=( a4470a ) or ( a4471a );
 a5334a <=( a4467a ) or ( a4468a );
 a5335a <=( a4469a ) or ( a5334a );
 a5336a <=( a5335a ) or ( a5330a );
 a5339a <=( a4465a ) or ( a4466a );
 a5343a <=( a4462a ) or ( a4463a );
 a5344a <=( a4464a ) or ( a5343a );
 a5345a <=( a5344a ) or ( a5339a );
 a5346a <=( a5345a ) or ( a5336a );
 a5347a <=( a5346a ) or ( a5327a );
 a5348a <=( a5347a ) or ( a5310a );
 a5349a <=( a5348a ) or ( a5273a );
 a5350a <=( a5349a ) or ( a5200a );
 a5351a <=( a5350a ) or ( a5053a );
 a5354a <=( a4460a ) or ( a4461a );
 a5357a <=( a4458a ) or ( a4459a );
 a5358a <=( a5357a ) or ( a5354a );
 a5361a <=( a4456a ) or ( a4457a );
 a5365a <=( a4453a ) or ( a4454a );
 a5366a <=( a4455a ) or ( a5365a );
 a5367a <=( a5366a ) or ( a5361a );
 a5368a <=( a5367a ) or ( a5358a );
 a5371a <=( a4451a ) or ( a4452a );
 a5374a <=( a4449a ) or ( a4450a );
 a5375a <=( a5374a ) or ( a5371a );
 a5378a <=( a4447a ) or ( a4448a );
 a5382a <=( a4444a ) or ( a4445a );
 a5383a <=( a4446a ) or ( a5382a );
 a5384a <=( a5383a ) or ( a5378a );
 a5385a <=( a5384a ) or ( a5375a );
 a5386a <=( a5385a ) or ( a5368a );
 a5389a <=( a4442a ) or ( a4443a );
 a5392a <=( a4440a ) or ( a4441a );
 a5393a <=( a5392a ) or ( a5389a );
 a5396a <=( a4438a ) or ( a4439a );
 a5400a <=( a4435a ) or ( a4436a );
 a5401a <=( a4437a ) or ( a5400a );
 a5402a <=( a5401a ) or ( a5396a );
 a5403a <=( a5402a ) or ( a5393a );
 a5406a <=( a4433a ) or ( a4434a );
 a5410a <=( a4430a ) or ( a4431a );
 a5411a <=( a4432a ) or ( a5410a );
 a5412a <=( a5411a ) or ( a5406a );
 a5415a <=( a4428a ) or ( a4429a );
 a5419a <=( a4425a ) or ( a4426a );
 a5420a <=( a4427a ) or ( a5419a );
 a5421a <=( a5420a ) or ( a5415a );
 a5422a <=( a5421a ) or ( a5412a );
 a5423a <=( a5422a ) or ( a5403a );
 a5424a <=( a5423a ) or ( a5386a );
 a5427a <=( a4423a ) or ( a4424a );
 a5430a <=( a4421a ) or ( a4422a );
 a5431a <=( a5430a ) or ( a5427a );
 a5434a <=( a4419a ) or ( a4420a );
 a5438a <=( a4416a ) or ( a4417a );
 a5439a <=( a4418a ) or ( a5438a );
 a5440a <=( a5439a ) or ( a5434a );
 a5441a <=( a5440a ) or ( a5431a );
 a5444a <=( a4414a ) or ( a4415a );
 a5447a <=( a4412a ) or ( a4413a );
 a5448a <=( a5447a ) or ( a5444a );
 a5451a <=( a4410a ) or ( a4411a );
 a5455a <=( a4407a ) or ( a4408a );
 a5456a <=( a4409a ) or ( a5455a );
 a5457a <=( a5456a ) or ( a5451a );
 a5458a <=( a5457a ) or ( a5448a );
 a5459a <=( a5458a ) or ( a5441a );
 a5462a <=( a4405a ) or ( a4406a );
 a5465a <=( a4403a ) or ( a4404a );
 a5466a <=( a5465a ) or ( a5462a );
 a5469a <=( a4401a ) or ( a4402a );
 a5473a <=( a4398a ) or ( a4399a );
 a5474a <=( a4400a ) or ( a5473a );
 a5475a <=( a5474a ) or ( a5469a );
 a5476a <=( a5475a ) or ( a5466a );
 a5479a <=( a4396a ) or ( a4397a );
 a5483a <=( a4393a ) or ( a4394a );
 a5484a <=( a4395a ) or ( a5483a );
 a5485a <=( a5484a ) or ( a5479a );
 a5488a <=( a4391a ) or ( a4392a );
 a5492a <=( a4388a ) or ( a4389a );
 a5493a <=( a4390a ) or ( a5492a );
 a5494a <=( a5493a ) or ( a5488a );
 a5495a <=( a5494a ) or ( a5485a );
 a5496a <=( a5495a ) or ( a5476a );
 a5497a <=( a5496a ) or ( a5459a );
 a5498a <=( a5497a ) or ( a5424a );
 a5501a <=( a4386a ) or ( a4387a );
 a5504a <=( a4384a ) or ( a4385a );
 a5505a <=( a5504a ) or ( a5501a );
 a5508a <=( a4382a ) or ( a4383a );
 a5512a <=( a4379a ) or ( a4380a );
 a5513a <=( a4381a ) or ( a5512a );
 a5514a <=( a5513a ) or ( a5508a );
 a5515a <=( a5514a ) or ( a5505a );
 a5518a <=( a4377a ) or ( a4378a );
 a5521a <=( a4375a ) or ( a4376a );
 a5522a <=( a5521a ) or ( a5518a );
 a5525a <=( a4373a ) or ( a4374a );
 a5529a <=( a4370a ) or ( a4371a );
 a5530a <=( a4372a ) or ( a5529a );
 a5531a <=( a5530a ) or ( a5525a );
 a5532a <=( a5531a ) or ( a5522a );
 a5533a <=( a5532a ) or ( a5515a );
 a5536a <=( a4368a ) or ( a4369a );
 a5539a <=( a4366a ) or ( a4367a );
 a5540a <=( a5539a ) or ( a5536a );
 a5543a <=( a4364a ) or ( a4365a );
 a5547a <=( a4361a ) or ( a4362a );
 a5548a <=( a4363a ) or ( a5547a );
 a5549a <=( a5548a ) or ( a5543a );
 a5550a <=( a5549a ) or ( a5540a );
 a5553a <=( a4359a ) or ( a4360a );
 a5557a <=( a4356a ) or ( a4357a );
 a5558a <=( a4358a ) or ( a5557a );
 a5559a <=( a5558a ) or ( a5553a );
 a5562a <=( a4354a ) or ( a4355a );
 a5566a <=( a4351a ) or ( a4352a );
 a5567a <=( a4353a ) or ( a5566a );
 a5568a <=( a5567a ) or ( a5562a );
 a5569a <=( a5568a ) or ( a5559a );
 a5570a <=( a5569a ) or ( a5550a );
 a5571a <=( a5570a ) or ( a5533a );
 a5574a <=( a4349a ) or ( a4350a );
 a5577a <=( a4347a ) or ( a4348a );
 a5578a <=( a5577a ) or ( a5574a );
 a5581a <=( a4345a ) or ( a4346a );
 a5585a <=( a4342a ) or ( a4343a );
 a5586a <=( a4344a ) or ( a5585a );
 a5587a <=( a5586a ) or ( a5581a );
 a5588a <=( a5587a ) or ( a5578a );
 a5591a <=( a4340a ) or ( a4341a );
 a5594a <=( a4338a ) or ( a4339a );
 a5595a <=( a5594a ) or ( a5591a );
 a5598a <=( a4336a ) or ( a4337a );
 a5602a <=( a4333a ) or ( a4334a );
 a5603a <=( a4335a ) or ( a5602a );
 a5604a <=( a5603a ) or ( a5598a );
 a5605a <=( a5604a ) or ( a5595a );
 a5606a <=( a5605a ) or ( a5588a );
 a5609a <=( a4331a ) or ( a4332a );
 a5612a <=( a4329a ) or ( a4330a );
 a5613a <=( a5612a ) or ( a5609a );
 a5616a <=( a4327a ) or ( a4328a );
 a5620a <=( a4324a ) or ( a4325a );
 a5621a <=( a4326a ) or ( a5620a );
 a5622a <=( a5621a ) or ( a5616a );
 a5623a <=( a5622a ) or ( a5613a );
 a5626a <=( a4322a ) or ( a4323a );
 a5630a <=( a4319a ) or ( a4320a );
 a5631a <=( a4321a ) or ( a5630a );
 a5632a <=( a5631a ) or ( a5626a );
 a5635a <=( a4317a ) or ( a4318a );
 a5639a <=( a4314a ) or ( a4315a );
 a5640a <=( a4316a ) or ( a5639a );
 a5641a <=( a5640a ) or ( a5635a );
 a5642a <=( a5641a ) or ( a5632a );
 a5643a <=( a5642a ) or ( a5623a );
 a5644a <=( a5643a ) or ( a5606a );
 a5645a <=( a5644a ) or ( a5571a );
 a5646a <=( a5645a ) or ( a5498a );
 a5649a <=( a4312a ) or ( a4313a );
 a5652a <=( a4310a ) or ( a4311a );
 a5653a <=( a5652a ) or ( a5649a );
 a5656a <=( a4308a ) or ( a4309a );
 a5660a <=( a4305a ) or ( a4306a );
 a5661a <=( a4307a ) or ( a5660a );
 a5662a <=( a5661a ) or ( a5656a );
 a5663a <=( a5662a ) or ( a5653a );
 a5666a <=( a4303a ) or ( a4304a );
 a5669a <=( a4301a ) or ( a4302a );
 a5670a <=( a5669a ) or ( a5666a );
 a5673a <=( a4299a ) or ( a4300a );
 a5677a <=( a4296a ) or ( a4297a );
 a5678a <=( a4298a ) or ( a5677a );
 a5679a <=( a5678a ) or ( a5673a );
 a5680a <=( a5679a ) or ( a5670a );
 a5681a <=( a5680a ) or ( a5663a );
 a5684a <=( a4294a ) or ( a4295a );
 a5687a <=( a4292a ) or ( a4293a );
 a5688a <=( a5687a ) or ( a5684a );
 a5691a <=( a4290a ) or ( a4291a );
 a5695a <=( a4287a ) or ( a4288a );
 a5696a <=( a4289a ) or ( a5695a );
 a5697a <=( a5696a ) or ( a5691a );
 a5698a <=( a5697a ) or ( a5688a );
 a5701a <=( a4285a ) or ( a4286a );
 a5705a <=( a4282a ) or ( a4283a );
 a5706a <=( a4284a ) or ( a5705a );
 a5707a <=( a5706a ) or ( a5701a );
 a5710a <=( a4280a ) or ( a4281a );
 a5714a <=( a4277a ) or ( a4278a );
 a5715a <=( a4279a ) or ( a5714a );
 a5716a <=( a5715a ) or ( a5710a );
 a5717a <=( a5716a ) or ( a5707a );
 a5718a <=( a5717a ) or ( a5698a );
 a5719a <=( a5718a ) or ( a5681a );
 a5722a <=( a4275a ) or ( a4276a );
 a5725a <=( a4273a ) or ( a4274a );
 a5726a <=( a5725a ) or ( a5722a );
 a5729a <=( a4271a ) or ( a4272a );
 a5733a <=( a4268a ) or ( a4269a );
 a5734a <=( a4270a ) or ( a5733a );
 a5735a <=( a5734a ) or ( a5729a );
 a5736a <=( a5735a ) or ( a5726a );
 a5739a <=( a4266a ) or ( a4267a );
 a5742a <=( a4264a ) or ( a4265a );
 a5743a <=( a5742a ) or ( a5739a );
 a5746a <=( a4262a ) or ( a4263a );
 a5750a <=( a4259a ) or ( a4260a );
 a5751a <=( a4261a ) or ( a5750a );
 a5752a <=( a5751a ) or ( a5746a );
 a5753a <=( a5752a ) or ( a5743a );
 a5754a <=( a5753a ) or ( a5736a );
 a5757a <=( a4257a ) or ( a4258a );
 a5760a <=( a4255a ) or ( a4256a );
 a5761a <=( a5760a ) or ( a5757a );
 a5764a <=( a4253a ) or ( a4254a );
 a5768a <=( a4250a ) or ( a4251a );
 a5769a <=( a4252a ) or ( a5768a );
 a5770a <=( a5769a ) or ( a5764a );
 a5771a <=( a5770a ) or ( a5761a );
 a5774a <=( a4248a ) or ( a4249a );
 a5778a <=( a4245a ) or ( a4246a );
 a5779a <=( a4247a ) or ( a5778a );
 a5780a <=( a5779a ) or ( a5774a );
 a5783a <=( a4243a ) or ( a4244a );
 a5787a <=( a4240a ) or ( a4241a );
 a5788a <=( a4242a ) or ( a5787a );
 a5789a <=( a5788a ) or ( a5783a );
 a5790a <=( a5789a ) or ( a5780a );
 a5791a <=( a5790a ) or ( a5771a );
 a5792a <=( a5791a ) or ( a5754a );
 a5793a <=( a5792a ) or ( a5719a );
 a5796a <=( a4238a ) or ( a4239a );
 a5799a <=( a4236a ) or ( a4237a );
 a5800a <=( a5799a ) or ( a5796a );
 a5803a <=( a4234a ) or ( a4235a );
 a5807a <=( a4231a ) or ( a4232a );
 a5808a <=( a4233a ) or ( a5807a );
 a5809a <=( a5808a ) or ( a5803a );
 a5810a <=( a5809a ) or ( a5800a );
 a5813a <=( a4229a ) or ( a4230a );
 a5816a <=( a4227a ) or ( a4228a );
 a5817a <=( a5816a ) or ( a5813a );
 a5820a <=( a4225a ) or ( a4226a );
 a5824a <=( a4222a ) or ( a4223a );
 a5825a <=( a4224a ) or ( a5824a );
 a5826a <=( a5825a ) or ( a5820a );
 a5827a <=( a5826a ) or ( a5817a );
 a5828a <=( a5827a ) or ( a5810a );
 a5831a <=( a4220a ) or ( a4221a );
 a5834a <=( a4218a ) or ( a4219a );
 a5835a <=( a5834a ) or ( a5831a );
 a5838a <=( a4216a ) or ( a4217a );
 a5842a <=( a4213a ) or ( a4214a );
 a5843a <=( a4215a ) or ( a5842a );
 a5844a <=( a5843a ) or ( a5838a );
 a5845a <=( a5844a ) or ( a5835a );
 a5848a <=( a4211a ) or ( a4212a );
 a5852a <=( a4208a ) or ( a4209a );
 a5853a <=( a4210a ) or ( a5852a );
 a5854a <=( a5853a ) or ( a5848a );
 a5857a <=( a4206a ) or ( a4207a );
 a5861a <=( a4203a ) or ( a4204a );
 a5862a <=( a4205a ) or ( a5861a );
 a5863a <=( a5862a ) or ( a5857a );
 a5864a <=( a5863a ) or ( a5854a );
 a5865a <=( a5864a ) or ( a5845a );
 a5866a <=( a5865a ) or ( a5828a );
 a5869a <=( a4201a ) or ( a4202a );
 a5872a <=( a4199a ) or ( a4200a );
 a5873a <=( a5872a ) or ( a5869a );
 a5876a <=( a4197a ) or ( a4198a );
 a5880a <=( a4194a ) or ( a4195a );
 a5881a <=( a4196a ) or ( a5880a );
 a5882a <=( a5881a ) or ( a5876a );
 a5883a <=( a5882a ) or ( a5873a );
 a5886a <=( a4192a ) or ( a4193a );
 a5890a <=( a4189a ) or ( a4190a );
 a5891a <=( a4191a ) or ( a5890a );
 a5892a <=( a5891a ) or ( a5886a );
 a5895a <=( a4187a ) or ( a4188a );
 a5899a <=( a4184a ) or ( a4185a );
 a5900a <=( a4186a ) or ( a5899a );
 a5901a <=( a5900a ) or ( a5895a );
 a5902a <=( a5901a ) or ( a5892a );
 a5903a <=( a5902a ) or ( a5883a );
 a5906a <=( a4182a ) or ( a4183a );
 a5909a <=( a4180a ) or ( a4181a );
 a5910a <=( a5909a ) or ( a5906a );
 a5913a <=( a4178a ) or ( a4179a );
 a5917a <=( a4175a ) or ( a4176a );
 a5918a <=( a4177a ) or ( a5917a );
 a5919a <=( a5918a ) or ( a5913a );
 a5920a <=( a5919a ) or ( a5910a );
 a5923a <=( a4173a ) or ( a4174a );
 a5927a <=( a4170a ) or ( a4171a );
 a5928a <=( a4172a ) or ( a5927a );
 a5929a <=( a5928a ) or ( a5923a );
 a5932a <=( a4168a ) or ( a4169a );
 a5936a <=( a4165a ) or ( a4166a );
 a5937a <=( a4167a ) or ( a5936a );
 a5938a <=( a5937a ) or ( a5932a );
 a5939a <=( a5938a ) or ( a5929a );
 a5940a <=( a5939a ) or ( a5920a );
 a5941a <=( a5940a ) or ( a5903a );
 a5942a <=( a5941a ) or ( a5866a );
 a5943a <=( a5942a ) or ( a5793a );
 a5944a <=( a5943a ) or ( a5646a );
 a5945a <=( a5944a ) or ( a5351a );
 a5948a <=( a4163a ) or ( a4164a );
 a5951a <=( a4161a ) or ( a4162a );
 a5952a <=( a5951a ) or ( a5948a );
 a5955a <=( a4159a ) or ( a4160a );
 a5959a <=( a4156a ) or ( a4157a );
 a5960a <=( a4158a ) or ( a5959a );
 a5961a <=( a5960a ) or ( a5955a );
 a5962a <=( a5961a ) or ( a5952a );
 a5965a <=( a4154a ) or ( a4155a );
 a5968a <=( a4152a ) or ( a4153a );
 a5969a <=( a5968a ) or ( a5965a );
 a5972a <=( a4150a ) or ( a4151a );
 a5976a <=( a4147a ) or ( a4148a );
 a5977a <=( a4149a ) or ( a5976a );
 a5978a <=( a5977a ) or ( a5972a );
 a5979a <=( a5978a ) or ( a5969a );
 a5980a <=( a5979a ) or ( a5962a );
 a5983a <=( a4145a ) or ( a4146a );
 a5986a <=( a4143a ) or ( a4144a );
 a5987a <=( a5986a ) or ( a5983a );
 a5990a <=( a4141a ) or ( a4142a );
 a5994a <=( a4138a ) or ( a4139a );
 a5995a <=( a4140a ) or ( a5994a );
 a5996a <=( a5995a ) or ( a5990a );
 a5997a <=( a5996a ) or ( a5987a );
 a6000a <=( a4136a ) or ( a4137a );
 a6004a <=( a4133a ) or ( a4134a );
 a6005a <=( a4135a ) or ( a6004a );
 a6006a <=( a6005a ) or ( a6000a );
 a6009a <=( a4131a ) or ( a4132a );
 a6013a <=( a4128a ) or ( a4129a );
 a6014a <=( a4130a ) or ( a6013a );
 a6015a <=( a6014a ) or ( a6009a );
 a6016a <=( a6015a ) or ( a6006a );
 a6017a <=( a6016a ) or ( a5997a );
 a6018a <=( a6017a ) or ( a5980a );
 a6021a <=( a4126a ) or ( a4127a );
 a6024a <=( a4124a ) or ( a4125a );
 a6025a <=( a6024a ) or ( a6021a );
 a6028a <=( a4122a ) or ( a4123a );
 a6032a <=( a4119a ) or ( a4120a );
 a6033a <=( a4121a ) or ( a6032a );
 a6034a <=( a6033a ) or ( a6028a );
 a6035a <=( a6034a ) or ( a6025a );
 a6038a <=( a4117a ) or ( a4118a );
 a6041a <=( a4115a ) or ( a4116a );
 a6042a <=( a6041a ) or ( a6038a );
 a6045a <=( a4113a ) or ( a4114a );
 a6049a <=( a4110a ) or ( a4111a );
 a6050a <=( a4112a ) or ( a6049a );
 a6051a <=( a6050a ) or ( a6045a );
 a6052a <=( a6051a ) or ( a6042a );
 a6053a <=( a6052a ) or ( a6035a );
 a6056a <=( a4108a ) or ( a4109a );
 a6059a <=( a4106a ) or ( a4107a );
 a6060a <=( a6059a ) or ( a6056a );
 a6063a <=( a4104a ) or ( a4105a );
 a6067a <=( a4101a ) or ( a4102a );
 a6068a <=( a4103a ) or ( a6067a );
 a6069a <=( a6068a ) or ( a6063a );
 a6070a <=( a6069a ) or ( a6060a );
 a6073a <=( a4099a ) or ( a4100a );
 a6077a <=( a4096a ) or ( a4097a );
 a6078a <=( a4098a ) or ( a6077a );
 a6079a <=( a6078a ) or ( a6073a );
 a6082a <=( a4094a ) or ( a4095a );
 a6086a <=( a4091a ) or ( a4092a );
 a6087a <=( a4093a ) or ( a6086a );
 a6088a <=( a6087a ) or ( a6082a );
 a6089a <=( a6088a ) or ( a6079a );
 a6090a <=( a6089a ) or ( a6070a );
 a6091a <=( a6090a ) or ( a6053a );
 a6092a <=( a6091a ) or ( a6018a );
 a6095a <=( a4089a ) or ( a4090a );
 a6098a <=( a4087a ) or ( a4088a );
 a6099a <=( a6098a ) or ( a6095a );
 a6102a <=( a4085a ) or ( a4086a );
 a6106a <=( a4082a ) or ( a4083a );
 a6107a <=( a4084a ) or ( a6106a );
 a6108a <=( a6107a ) or ( a6102a );
 a6109a <=( a6108a ) or ( a6099a );
 a6112a <=( a4080a ) or ( a4081a );
 a6115a <=( a4078a ) or ( a4079a );
 a6116a <=( a6115a ) or ( a6112a );
 a6119a <=( a4076a ) or ( a4077a );
 a6123a <=( a4073a ) or ( a4074a );
 a6124a <=( a4075a ) or ( a6123a );
 a6125a <=( a6124a ) or ( a6119a );
 a6126a <=( a6125a ) or ( a6116a );
 a6127a <=( a6126a ) or ( a6109a );
 a6130a <=( a4071a ) or ( a4072a );
 a6133a <=( a4069a ) or ( a4070a );
 a6134a <=( a6133a ) or ( a6130a );
 a6137a <=( a4067a ) or ( a4068a );
 a6141a <=( a4064a ) or ( a4065a );
 a6142a <=( a4066a ) or ( a6141a );
 a6143a <=( a6142a ) or ( a6137a );
 a6144a <=( a6143a ) or ( a6134a );
 a6147a <=( a4062a ) or ( a4063a );
 a6151a <=( a4059a ) or ( a4060a );
 a6152a <=( a4061a ) or ( a6151a );
 a6153a <=( a6152a ) or ( a6147a );
 a6156a <=( a4057a ) or ( a4058a );
 a6160a <=( a4054a ) or ( a4055a );
 a6161a <=( a4056a ) or ( a6160a );
 a6162a <=( a6161a ) or ( a6156a );
 a6163a <=( a6162a ) or ( a6153a );
 a6164a <=( a6163a ) or ( a6144a );
 a6165a <=( a6164a ) or ( a6127a );
 a6168a <=( a4052a ) or ( a4053a );
 a6171a <=( a4050a ) or ( a4051a );
 a6172a <=( a6171a ) or ( a6168a );
 a6175a <=( a4048a ) or ( a4049a );
 a6179a <=( a4045a ) or ( a4046a );
 a6180a <=( a4047a ) or ( a6179a );
 a6181a <=( a6180a ) or ( a6175a );
 a6182a <=( a6181a ) or ( a6172a );
 a6185a <=( a4043a ) or ( a4044a );
 a6188a <=( a4041a ) or ( a4042a );
 a6189a <=( a6188a ) or ( a6185a );
 a6192a <=( a4039a ) or ( a4040a );
 a6196a <=( a4036a ) or ( a4037a );
 a6197a <=( a4038a ) or ( a6196a );
 a6198a <=( a6197a ) or ( a6192a );
 a6199a <=( a6198a ) or ( a6189a );
 a6200a <=( a6199a ) or ( a6182a );
 a6203a <=( a4034a ) or ( a4035a );
 a6206a <=( a4032a ) or ( a4033a );
 a6207a <=( a6206a ) or ( a6203a );
 a6210a <=( a4030a ) or ( a4031a );
 a6214a <=( a4027a ) or ( a4028a );
 a6215a <=( a4029a ) or ( a6214a );
 a6216a <=( a6215a ) or ( a6210a );
 a6217a <=( a6216a ) or ( a6207a );
 a6220a <=( a4025a ) or ( a4026a );
 a6224a <=( a4022a ) or ( a4023a );
 a6225a <=( a4024a ) or ( a6224a );
 a6226a <=( a6225a ) or ( a6220a );
 a6229a <=( a4020a ) or ( a4021a );
 a6233a <=( a4017a ) or ( a4018a );
 a6234a <=( a4019a ) or ( a6233a );
 a6235a <=( a6234a ) or ( a6229a );
 a6236a <=( a6235a ) or ( a6226a );
 a6237a <=( a6236a ) or ( a6217a );
 a6238a <=( a6237a ) or ( a6200a );
 a6239a <=( a6238a ) or ( a6165a );
 a6240a <=( a6239a ) or ( a6092a );
 a6243a <=( a4015a ) or ( a4016a );
 a6246a <=( a4013a ) or ( a4014a );
 a6247a <=( a6246a ) or ( a6243a );
 a6250a <=( a4011a ) or ( a4012a );
 a6254a <=( a4008a ) or ( a4009a );
 a6255a <=( a4010a ) or ( a6254a );
 a6256a <=( a6255a ) or ( a6250a );
 a6257a <=( a6256a ) or ( a6247a );
 a6260a <=( a4006a ) or ( a4007a );
 a6263a <=( a4004a ) or ( a4005a );
 a6264a <=( a6263a ) or ( a6260a );
 a6267a <=( a4002a ) or ( a4003a );
 a6271a <=( a3999a ) or ( a4000a );
 a6272a <=( a4001a ) or ( a6271a );
 a6273a <=( a6272a ) or ( a6267a );
 a6274a <=( a6273a ) or ( a6264a );
 a6275a <=( a6274a ) or ( a6257a );
 a6278a <=( a3997a ) or ( a3998a );
 a6281a <=( a3995a ) or ( a3996a );
 a6282a <=( a6281a ) or ( a6278a );
 a6285a <=( a3993a ) or ( a3994a );
 a6289a <=( a3990a ) or ( a3991a );
 a6290a <=( a3992a ) or ( a6289a );
 a6291a <=( a6290a ) or ( a6285a );
 a6292a <=( a6291a ) or ( a6282a );
 a6295a <=( a3988a ) or ( a3989a );
 a6299a <=( a3985a ) or ( a3986a );
 a6300a <=( a3987a ) or ( a6299a );
 a6301a <=( a6300a ) or ( a6295a );
 a6304a <=( a3983a ) or ( a3984a );
 a6308a <=( a3980a ) or ( a3981a );
 a6309a <=( a3982a ) or ( a6308a );
 a6310a <=( a6309a ) or ( a6304a );
 a6311a <=( a6310a ) or ( a6301a );
 a6312a <=( a6311a ) or ( a6292a );
 a6313a <=( a6312a ) or ( a6275a );
 a6316a <=( a3978a ) or ( a3979a );
 a6319a <=( a3976a ) or ( a3977a );
 a6320a <=( a6319a ) or ( a6316a );
 a6323a <=( a3974a ) or ( a3975a );
 a6327a <=( a3971a ) or ( a3972a );
 a6328a <=( a3973a ) or ( a6327a );
 a6329a <=( a6328a ) or ( a6323a );
 a6330a <=( a6329a ) or ( a6320a );
 a6333a <=( a3969a ) or ( a3970a );
 a6336a <=( a3967a ) or ( a3968a );
 a6337a <=( a6336a ) or ( a6333a );
 a6340a <=( a3965a ) or ( a3966a );
 a6344a <=( a3962a ) or ( a3963a );
 a6345a <=( a3964a ) or ( a6344a );
 a6346a <=( a6345a ) or ( a6340a );
 a6347a <=( a6346a ) or ( a6337a );
 a6348a <=( a6347a ) or ( a6330a );
 a6351a <=( a3960a ) or ( a3961a );
 a6354a <=( a3958a ) or ( a3959a );
 a6355a <=( a6354a ) or ( a6351a );
 a6358a <=( a3956a ) or ( a3957a );
 a6362a <=( a3953a ) or ( a3954a );
 a6363a <=( a3955a ) or ( a6362a );
 a6364a <=( a6363a ) or ( a6358a );
 a6365a <=( a6364a ) or ( a6355a );
 a6368a <=( a3951a ) or ( a3952a );
 a6372a <=( a3948a ) or ( a3949a );
 a6373a <=( a3950a ) or ( a6372a );
 a6374a <=( a6373a ) or ( a6368a );
 a6377a <=( a3946a ) or ( a3947a );
 a6381a <=( a3943a ) or ( a3944a );
 a6382a <=( a3945a ) or ( a6381a );
 a6383a <=( a6382a ) or ( a6377a );
 a6384a <=( a6383a ) or ( a6374a );
 a6385a <=( a6384a ) or ( a6365a );
 a6386a <=( a6385a ) or ( a6348a );
 a6387a <=( a6386a ) or ( a6313a );
 a6390a <=( a3941a ) or ( a3942a );
 a6393a <=( a3939a ) or ( a3940a );
 a6394a <=( a6393a ) or ( a6390a );
 a6397a <=( a3937a ) or ( a3938a );
 a6401a <=( a3934a ) or ( a3935a );
 a6402a <=( a3936a ) or ( a6401a );
 a6403a <=( a6402a ) or ( a6397a );
 a6404a <=( a6403a ) or ( a6394a );
 a6407a <=( a3932a ) or ( a3933a );
 a6410a <=( a3930a ) or ( a3931a );
 a6411a <=( a6410a ) or ( a6407a );
 a6414a <=( a3928a ) or ( a3929a );
 a6418a <=( a3925a ) or ( a3926a );
 a6419a <=( a3927a ) or ( a6418a );
 a6420a <=( a6419a ) or ( a6414a );
 a6421a <=( a6420a ) or ( a6411a );
 a6422a <=( a6421a ) or ( a6404a );
 a6425a <=( a3923a ) or ( a3924a );
 a6428a <=( a3921a ) or ( a3922a );
 a6429a <=( a6428a ) or ( a6425a );
 a6432a <=( a3919a ) or ( a3920a );
 a6436a <=( a3916a ) or ( a3917a );
 a6437a <=( a3918a ) or ( a6436a );
 a6438a <=( a6437a ) or ( a6432a );
 a6439a <=( a6438a ) or ( a6429a );
 a6442a <=( a3914a ) or ( a3915a );
 a6446a <=( a3911a ) or ( a3912a );
 a6447a <=( a3913a ) or ( a6446a );
 a6448a <=( a6447a ) or ( a6442a );
 a6451a <=( a3909a ) or ( a3910a );
 a6455a <=( a3906a ) or ( a3907a );
 a6456a <=( a3908a ) or ( a6455a );
 a6457a <=( a6456a ) or ( a6451a );
 a6458a <=( a6457a ) or ( a6448a );
 a6459a <=( a6458a ) or ( a6439a );
 a6460a <=( a6459a ) or ( a6422a );
 a6463a <=( a3904a ) or ( a3905a );
 a6466a <=( a3902a ) or ( a3903a );
 a6467a <=( a6466a ) or ( a6463a );
 a6470a <=( a3900a ) or ( a3901a );
 a6474a <=( a3897a ) or ( a3898a );
 a6475a <=( a3899a ) or ( a6474a );
 a6476a <=( a6475a ) or ( a6470a );
 a6477a <=( a6476a ) or ( a6467a );
 a6480a <=( a3895a ) or ( a3896a );
 a6484a <=( a3892a ) or ( a3893a );
 a6485a <=( a3894a ) or ( a6484a );
 a6486a <=( a6485a ) or ( a6480a );
 a6489a <=( a3890a ) or ( a3891a );
 a6493a <=( a3887a ) or ( a3888a );
 a6494a <=( a3889a ) or ( a6493a );
 a6495a <=( a6494a ) or ( a6489a );
 a6496a <=( a6495a ) or ( a6486a );
 a6497a <=( a6496a ) or ( a6477a );
 a6500a <=( a3885a ) or ( a3886a );
 a6503a <=( a3883a ) or ( a3884a );
 a6504a <=( a6503a ) or ( a6500a );
 a6507a <=( a3881a ) or ( a3882a );
 a6511a <=( a3878a ) or ( a3879a );
 a6512a <=( a3880a ) or ( a6511a );
 a6513a <=( a6512a ) or ( a6507a );
 a6514a <=( a6513a ) or ( a6504a );
 a6517a <=( a3876a ) or ( a3877a );
 a6521a <=( a3873a ) or ( a3874a );
 a6522a <=( a3875a ) or ( a6521a );
 a6523a <=( a6522a ) or ( a6517a );
 a6526a <=( a3871a ) or ( a3872a );
 a6530a <=( a3868a ) or ( a3869a );
 a6531a <=( a3870a ) or ( a6530a );
 a6532a <=( a6531a ) or ( a6526a );
 a6533a <=( a6532a ) or ( a6523a );
 a6534a <=( a6533a ) or ( a6514a );
 a6535a <=( a6534a ) or ( a6497a );
 a6536a <=( a6535a ) or ( a6460a );
 a6537a <=( a6536a ) or ( a6387a );
 a6538a <=( a6537a ) or ( a6240a );
 a6541a <=( a3866a ) or ( a3867a );
 a6544a <=( a3864a ) or ( a3865a );
 a6545a <=( a6544a ) or ( a6541a );
 a6548a <=( a3862a ) or ( a3863a );
 a6552a <=( a3859a ) or ( a3860a );
 a6553a <=( a3861a ) or ( a6552a );
 a6554a <=( a6553a ) or ( a6548a );
 a6555a <=( a6554a ) or ( a6545a );
 a6558a <=( a3857a ) or ( a3858a );
 a6561a <=( a3855a ) or ( a3856a );
 a6562a <=( a6561a ) or ( a6558a );
 a6565a <=( a3853a ) or ( a3854a );
 a6569a <=( a3850a ) or ( a3851a );
 a6570a <=( a3852a ) or ( a6569a );
 a6571a <=( a6570a ) or ( a6565a );
 a6572a <=( a6571a ) or ( a6562a );
 a6573a <=( a6572a ) or ( a6555a );
 a6576a <=( a3848a ) or ( a3849a );
 a6579a <=( a3846a ) or ( a3847a );
 a6580a <=( a6579a ) or ( a6576a );
 a6583a <=( a3844a ) or ( a3845a );
 a6587a <=( a3841a ) or ( a3842a );
 a6588a <=( a3843a ) or ( a6587a );
 a6589a <=( a6588a ) or ( a6583a );
 a6590a <=( a6589a ) or ( a6580a );
 a6593a <=( a3839a ) or ( a3840a );
 a6597a <=( a3836a ) or ( a3837a );
 a6598a <=( a3838a ) or ( a6597a );
 a6599a <=( a6598a ) or ( a6593a );
 a6602a <=( a3834a ) or ( a3835a );
 a6606a <=( a3831a ) or ( a3832a );
 a6607a <=( a3833a ) or ( a6606a );
 a6608a <=( a6607a ) or ( a6602a );
 a6609a <=( a6608a ) or ( a6599a );
 a6610a <=( a6609a ) or ( a6590a );
 a6611a <=( a6610a ) or ( a6573a );
 a6614a <=( a3829a ) or ( a3830a );
 a6617a <=( a3827a ) or ( a3828a );
 a6618a <=( a6617a ) or ( a6614a );
 a6621a <=( a3825a ) or ( a3826a );
 a6625a <=( a3822a ) or ( a3823a );
 a6626a <=( a3824a ) or ( a6625a );
 a6627a <=( a6626a ) or ( a6621a );
 a6628a <=( a6627a ) or ( a6618a );
 a6631a <=( a3820a ) or ( a3821a );
 a6634a <=( a3818a ) or ( a3819a );
 a6635a <=( a6634a ) or ( a6631a );
 a6638a <=( a3816a ) or ( a3817a );
 a6642a <=( a3813a ) or ( a3814a );
 a6643a <=( a3815a ) or ( a6642a );
 a6644a <=( a6643a ) or ( a6638a );
 a6645a <=( a6644a ) or ( a6635a );
 a6646a <=( a6645a ) or ( a6628a );
 a6649a <=( a3811a ) or ( a3812a );
 a6652a <=( a3809a ) or ( a3810a );
 a6653a <=( a6652a ) or ( a6649a );
 a6656a <=( a3807a ) or ( a3808a );
 a6660a <=( a3804a ) or ( a3805a );
 a6661a <=( a3806a ) or ( a6660a );
 a6662a <=( a6661a ) or ( a6656a );
 a6663a <=( a6662a ) or ( a6653a );
 a6666a <=( a3802a ) or ( a3803a );
 a6670a <=( a3799a ) or ( a3800a );
 a6671a <=( a3801a ) or ( a6670a );
 a6672a <=( a6671a ) or ( a6666a );
 a6675a <=( a3797a ) or ( a3798a );
 a6679a <=( a3794a ) or ( a3795a );
 a6680a <=( a3796a ) or ( a6679a );
 a6681a <=( a6680a ) or ( a6675a );
 a6682a <=( a6681a ) or ( a6672a );
 a6683a <=( a6682a ) or ( a6663a );
 a6684a <=( a6683a ) or ( a6646a );
 a6685a <=( a6684a ) or ( a6611a );
 a6688a <=( a3792a ) or ( a3793a );
 a6691a <=( a3790a ) or ( a3791a );
 a6692a <=( a6691a ) or ( a6688a );
 a6695a <=( a3788a ) or ( a3789a );
 a6699a <=( a3785a ) or ( a3786a );
 a6700a <=( a3787a ) or ( a6699a );
 a6701a <=( a6700a ) or ( a6695a );
 a6702a <=( a6701a ) or ( a6692a );
 a6705a <=( a3783a ) or ( a3784a );
 a6708a <=( a3781a ) or ( a3782a );
 a6709a <=( a6708a ) or ( a6705a );
 a6712a <=( a3779a ) or ( a3780a );
 a6716a <=( a3776a ) or ( a3777a );
 a6717a <=( a3778a ) or ( a6716a );
 a6718a <=( a6717a ) or ( a6712a );
 a6719a <=( a6718a ) or ( a6709a );
 a6720a <=( a6719a ) or ( a6702a );
 a6723a <=( a3774a ) or ( a3775a );
 a6726a <=( a3772a ) or ( a3773a );
 a6727a <=( a6726a ) or ( a6723a );
 a6730a <=( a3770a ) or ( a3771a );
 a6734a <=( a3767a ) or ( a3768a );
 a6735a <=( a3769a ) or ( a6734a );
 a6736a <=( a6735a ) or ( a6730a );
 a6737a <=( a6736a ) or ( a6727a );
 a6740a <=( a3765a ) or ( a3766a );
 a6744a <=( a3762a ) or ( a3763a );
 a6745a <=( a3764a ) or ( a6744a );
 a6746a <=( a6745a ) or ( a6740a );
 a6749a <=( a3760a ) or ( a3761a );
 a6753a <=( a3757a ) or ( a3758a );
 a6754a <=( a3759a ) or ( a6753a );
 a6755a <=( a6754a ) or ( a6749a );
 a6756a <=( a6755a ) or ( a6746a );
 a6757a <=( a6756a ) or ( a6737a );
 a6758a <=( a6757a ) or ( a6720a );
 a6761a <=( a3755a ) or ( a3756a );
 a6764a <=( a3753a ) or ( a3754a );
 a6765a <=( a6764a ) or ( a6761a );
 a6768a <=( a3751a ) or ( a3752a );
 a6772a <=( a3748a ) or ( a3749a );
 a6773a <=( a3750a ) or ( a6772a );
 a6774a <=( a6773a ) or ( a6768a );
 a6775a <=( a6774a ) or ( a6765a );
 a6778a <=( a3746a ) or ( a3747a );
 a6782a <=( a3743a ) or ( a3744a );
 a6783a <=( a3745a ) or ( a6782a );
 a6784a <=( a6783a ) or ( a6778a );
 a6787a <=( a3741a ) or ( a3742a );
 a6791a <=( a3738a ) or ( a3739a );
 a6792a <=( a3740a ) or ( a6791a );
 a6793a <=( a6792a ) or ( a6787a );
 a6794a <=( a6793a ) or ( a6784a );
 a6795a <=( a6794a ) or ( a6775a );
 a6798a <=( a3736a ) or ( a3737a );
 a6801a <=( a3734a ) or ( a3735a );
 a6802a <=( a6801a ) or ( a6798a );
 a6805a <=( a3732a ) or ( a3733a );
 a6809a <=( a3729a ) or ( a3730a );
 a6810a <=( a3731a ) or ( a6809a );
 a6811a <=( a6810a ) or ( a6805a );
 a6812a <=( a6811a ) or ( a6802a );
 a6815a <=( a3727a ) or ( a3728a );
 a6819a <=( a3724a ) or ( a3725a );
 a6820a <=( a3726a ) or ( a6819a );
 a6821a <=( a6820a ) or ( a6815a );
 a6824a <=( a3722a ) or ( a3723a );
 a6828a <=( a3719a ) or ( a3720a );
 a6829a <=( a3721a ) or ( a6828a );
 a6830a <=( a6829a ) or ( a6824a );
 a6831a <=( a6830a ) or ( a6821a );
 a6832a <=( a6831a ) or ( a6812a );
 a6833a <=( a6832a ) or ( a6795a );
 a6834a <=( a6833a ) or ( a6758a );
 a6835a <=( a6834a ) or ( a6685a );
 a6838a <=( a3717a ) or ( a3718a );
 a6841a <=( a3715a ) or ( a3716a );
 a6842a <=( a6841a ) or ( a6838a );
 a6845a <=( a3713a ) or ( a3714a );
 a6849a <=( a3710a ) or ( a3711a );
 a6850a <=( a3712a ) or ( a6849a );
 a6851a <=( a6850a ) or ( a6845a );
 a6852a <=( a6851a ) or ( a6842a );
 a6855a <=( a3708a ) or ( a3709a );
 a6858a <=( a3706a ) or ( a3707a );
 a6859a <=( a6858a ) or ( a6855a );
 a6862a <=( a3704a ) or ( a3705a );
 a6866a <=( a3701a ) or ( a3702a );
 a6867a <=( a3703a ) or ( a6866a );
 a6868a <=( a6867a ) or ( a6862a );
 a6869a <=( a6868a ) or ( a6859a );
 a6870a <=( a6869a ) or ( a6852a );
 a6873a <=( a3699a ) or ( a3700a );
 a6876a <=( a3697a ) or ( a3698a );
 a6877a <=( a6876a ) or ( a6873a );
 a6880a <=( a3695a ) or ( a3696a );
 a6884a <=( a3692a ) or ( a3693a );
 a6885a <=( a3694a ) or ( a6884a );
 a6886a <=( a6885a ) or ( a6880a );
 a6887a <=( a6886a ) or ( a6877a );
 a6890a <=( a3690a ) or ( a3691a );
 a6894a <=( a3687a ) or ( a3688a );
 a6895a <=( a3689a ) or ( a6894a );
 a6896a <=( a6895a ) or ( a6890a );
 a6899a <=( a3685a ) or ( a3686a );
 a6903a <=( a3682a ) or ( a3683a );
 a6904a <=( a3684a ) or ( a6903a );
 a6905a <=( a6904a ) or ( a6899a );
 a6906a <=( a6905a ) or ( a6896a );
 a6907a <=( a6906a ) or ( a6887a );
 a6908a <=( a6907a ) or ( a6870a );
 a6911a <=( a3680a ) or ( a3681a );
 a6914a <=( a3678a ) or ( a3679a );
 a6915a <=( a6914a ) or ( a6911a );
 a6918a <=( a3676a ) or ( a3677a );
 a6922a <=( a3673a ) or ( a3674a );
 a6923a <=( a3675a ) or ( a6922a );
 a6924a <=( a6923a ) or ( a6918a );
 a6925a <=( a6924a ) or ( a6915a );
 a6928a <=( a3671a ) or ( a3672a );
 a6931a <=( a3669a ) or ( a3670a );
 a6932a <=( a6931a ) or ( a6928a );
 a6935a <=( a3667a ) or ( a3668a );
 a6939a <=( a3664a ) or ( a3665a );
 a6940a <=( a3666a ) or ( a6939a );
 a6941a <=( a6940a ) or ( a6935a );
 a6942a <=( a6941a ) or ( a6932a );
 a6943a <=( a6942a ) or ( a6925a );
 a6946a <=( a3662a ) or ( a3663a );
 a6949a <=( a3660a ) or ( a3661a );
 a6950a <=( a6949a ) or ( a6946a );
 a6953a <=( a3658a ) or ( a3659a );
 a6957a <=( a3655a ) or ( a3656a );
 a6958a <=( a3657a ) or ( a6957a );
 a6959a <=( a6958a ) or ( a6953a );
 a6960a <=( a6959a ) or ( a6950a );
 a6963a <=( a3653a ) or ( a3654a );
 a6967a <=( a3650a ) or ( a3651a );
 a6968a <=( a3652a ) or ( a6967a );
 a6969a <=( a6968a ) or ( a6963a );
 a6972a <=( a3648a ) or ( a3649a );
 a6976a <=( a3645a ) or ( a3646a );
 a6977a <=( a3647a ) or ( a6976a );
 a6978a <=( a6977a ) or ( a6972a );
 a6979a <=( a6978a ) or ( a6969a );
 a6980a <=( a6979a ) or ( a6960a );
 a6981a <=( a6980a ) or ( a6943a );
 a6982a <=( a6981a ) or ( a6908a );
 a6985a <=( a3643a ) or ( a3644a );
 a6988a <=( a3641a ) or ( a3642a );
 a6989a <=( a6988a ) or ( a6985a );
 a6992a <=( a3639a ) or ( a3640a );
 a6996a <=( a3636a ) or ( a3637a );
 a6997a <=( a3638a ) or ( a6996a );
 a6998a <=( a6997a ) or ( a6992a );
 a6999a <=( a6998a ) or ( a6989a );
 a7002a <=( a3634a ) or ( a3635a );
 a7005a <=( a3632a ) or ( a3633a );
 a7006a <=( a7005a ) or ( a7002a );
 a7009a <=( a3630a ) or ( a3631a );
 a7013a <=( a3627a ) or ( a3628a );
 a7014a <=( a3629a ) or ( a7013a );
 a7015a <=( a7014a ) or ( a7009a );
 a7016a <=( a7015a ) or ( a7006a );
 a7017a <=( a7016a ) or ( a6999a );
 a7020a <=( a3625a ) or ( a3626a );
 a7023a <=( a3623a ) or ( a3624a );
 a7024a <=( a7023a ) or ( a7020a );
 a7027a <=( a3621a ) or ( a3622a );
 a7031a <=( a3618a ) or ( a3619a );
 a7032a <=( a3620a ) or ( a7031a );
 a7033a <=( a7032a ) or ( a7027a );
 a7034a <=( a7033a ) or ( a7024a );
 a7037a <=( a3616a ) or ( a3617a );
 a7041a <=( a3613a ) or ( a3614a );
 a7042a <=( a3615a ) or ( a7041a );
 a7043a <=( a7042a ) or ( a7037a );
 a7046a <=( a3611a ) or ( a3612a );
 a7050a <=( a3608a ) or ( a3609a );
 a7051a <=( a3610a ) or ( a7050a );
 a7052a <=( a7051a ) or ( a7046a );
 a7053a <=( a7052a ) or ( a7043a );
 a7054a <=( a7053a ) or ( a7034a );
 a7055a <=( a7054a ) or ( a7017a );
 a7058a <=( a3606a ) or ( a3607a );
 a7061a <=( a3604a ) or ( a3605a );
 a7062a <=( a7061a ) or ( a7058a );
 a7065a <=( a3602a ) or ( a3603a );
 a7069a <=( a3599a ) or ( a3600a );
 a7070a <=( a3601a ) or ( a7069a );
 a7071a <=( a7070a ) or ( a7065a );
 a7072a <=( a7071a ) or ( a7062a );
 a7075a <=( a3597a ) or ( a3598a );
 a7079a <=( a3594a ) or ( a3595a );
 a7080a <=( a3596a ) or ( a7079a );
 a7081a <=( a7080a ) or ( a7075a );
 a7084a <=( a3592a ) or ( a3593a );
 a7088a <=( a3589a ) or ( a3590a );
 a7089a <=( a3591a ) or ( a7088a );
 a7090a <=( a7089a ) or ( a7084a );
 a7091a <=( a7090a ) or ( a7081a );
 a7092a <=( a7091a ) or ( a7072a );
 a7095a <=( a3587a ) or ( a3588a );
 a7098a <=( a3585a ) or ( a3586a );
 a7099a <=( a7098a ) or ( a7095a );
 a7102a <=( a3583a ) or ( a3584a );
 a7106a <=( a3580a ) or ( a3581a );
 a7107a <=( a3582a ) or ( a7106a );
 a7108a <=( a7107a ) or ( a7102a );
 a7109a <=( a7108a ) or ( a7099a );
 a7112a <=( a3578a ) or ( a3579a );
 a7116a <=( a3575a ) or ( a3576a );
 a7117a <=( a3577a ) or ( a7116a );
 a7118a <=( a7117a ) or ( a7112a );
 a7121a <=( a3573a ) or ( a3574a );
 a7125a <=( a3570a ) or ( a3571a );
 a7126a <=( a3572a ) or ( a7125a );
 a7127a <=( a7126a ) or ( a7121a );
 a7128a <=( a7127a ) or ( a7118a );
 a7129a <=( a7128a ) or ( a7109a );
 a7130a <=( a7129a ) or ( a7092a );
 a7131a <=( a7130a ) or ( a7055a );
 a7132a <=( a7131a ) or ( a6982a );
 a7133a <=( a7132a ) or ( a6835a );
 a7134a <=( a7133a ) or ( a6538a );
 a7135a <=( a7134a ) or ( a5945a );
 a7138a <=( a3568a ) or ( a3569a );
 a7141a <=( a3566a ) or ( a3567a );
 a7142a <=( a7141a ) or ( a7138a );
 a7145a <=( a3564a ) or ( a3565a );
 a7149a <=( a3561a ) or ( a3562a );
 a7150a <=( a3563a ) or ( a7149a );
 a7151a <=( a7150a ) or ( a7145a );
 a7152a <=( a7151a ) or ( a7142a );
 a7155a <=( a3559a ) or ( a3560a );
 a7158a <=( a3557a ) or ( a3558a );
 a7159a <=( a7158a ) or ( a7155a );
 a7162a <=( a3555a ) or ( a3556a );
 a7166a <=( a3552a ) or ( a3553a );
 a7167a <=( a3554a ) or ( a7166a );
 a7168a <=( a7167a ) or ( a7162a );
 a7169a <=( a7168a ) or ( a7159a );
 a7170a <=( a7169a ) or ( a7152a );
 a7173a <=( a3550a ) or ( a3551a );
 a7176a <=( a3548a ) or ( a3549a );
 a7177a <=( a7176a ) or ( a7173a );
 a7180a <=( a3546a ) or ( a3547a );
 a7184a <=( a3543a ) or ( a3544a );
 a7185a <=( a3545a ) or ( a7184a );
 a7186a <=( a7185a ) or ( a7180a );
 a7187a <=( a7186a ) or ( a7177a );
 a7190a <=( a3541a ) or ( a3542a );
 a7194a <=( a3538a ) or ( a3539a );
 a7195a <=( a3540a ) or ( a7194a );
 a7196a <=( a7195a ) or ( a7190a );
 a7199a <=( a3536a ) or ( a3537a );
 a7203a <=( a3533a ) or ( a3534a );
 a7204a <=( a3535a ) or ( a7203a );
 a7205a <=( a7204a ) or ( a7199a );
 a7206a <=( a7205a ) or ( a7196a );
 a7207a <=( a7206a ) or ( a7187a );
 a7208a <=( a7207a ) or ( a7170a );
 a7211a <=( a3531a ) or ( a3532a );
 a7214a <=( a3529a ) or ( a3530a );
 a7215a <=( a7214a ) or ( a7211a );
 a7218a <=( a3527a ) or ( a3528a );
 a7222a <=( a3524a ) or ( a3525a );
 a7223a <=( a3526a ) or ( a7222a );
 a7224a <=( a7223a ) or ( a7218a );
 a7225a <=( a7224a ) or ( a7215a );
 a7228a <=( a3522a ) or ( a3523a );
 a7231a <=( a3520a ) or ( a3521a );
 a7232a <=( a7231a ) or ( a7228a );
 a7235a <=( a3518a ) or ( a3519a );
 a7239a <=( a3515a ) or ( a3516a );
 a7240a <=( a3517a ) or ( a7239a );
 a7241a <=( a7240a ) or ( a7235a );
 a7242a <=( a7241a ) or ( a7232a );
 a7243a <=( a7242a ) or ( a7225a );
 a7246a <=( a3513a ) or ( a3514a );
 a7249a <=( a3511a ) or ( a3512a );
 a7250a <=( a7249a ) or ( a7246a );
 a7253a <=( a3509a ) or ( a3510a );
 a7257a <=( a3506a ) or ( a3507a );
 a7258a <=( a3508a ) or ( a7257a );
 a7259a <=( a7258a ) or ( a7253a );
 a7260a <=( a7259a ) or ( a7250a );
 a7263a <=( a3504a ) or ( a3505a );
 a7267a <=( a3501a ) or ( a3502a );
 a7268a <=( a3503a ) or ( a7267a );
 a7269a <=( a7268a ) or ( a7263a );
 a7272a <=( a3499a ) or ( a3500a );
 a7276a <=( a3496a ) or ( a3497a );
 a7277a <=( a3498a ) or ( a7276a );
 a7278a <=( a7277a ) or ( a7272a );
 a7279a <=( a7278a ) or ( a7269a );
 a7280a <=( a7279a ) or ( a7260a );
 a7281a <=( a7280a ) or ( a7243a );
 a7282a <=( a7281a ) or ( a7208a );
 a7285a <=( a3494a ) or ( a3495a );
 a7288a <=( a3492a ) or ( a3493a );
 a7289a <=( a7288a ) or ( a7285a );
 a7292a <=( a3490a ) or ( a3491a );
 a7296a <=( a3487a ) or ( a3488a );
 a7297a <=( a3489a ) or ( a7296a );
 a7298a <=( a7297a ) or ( a7292a );
 a7299a <=( a7298a ) or ( a7289a );
 a7302a <=( a3485a ) or ( a3486a );
 a7305a <=( a3483a ) or ( a3484a );
 a7306a <=( a7305a ) or ( a7302a );
 a7309a <=( a3481a ) or ( a3482a );
 a7313a <=( a3478a ) or ( a3479a );
 a7314a <=( a3480a ) or ( a7313a );
 a7315a <=( a7314a ) or ( a7309a );
 a7316a <=( a7315a ) or ( a7306a );
 a7317a <=( a7316a ) or ( a7299a );
 a7320a <=( a3476a ) or ( a3477a );
 a7323a <=( a3474a ) or ( a3475a );
 a7324a <=( a7323a ) or ( a7320a );
 a7327a <=( a3472a ) or ( a3473a );
 a7331a <=( a3469a ) or ( a3470a );
 a7332a <=( a3471a ) or ( a7331a );
 a7333a <=( a7332a ) or ( a7327a );
 a7334a <=( a7333a ) or ( a7324a );
 a7337a <=( a3467a ) or ( a3468a );
 a7341a <=( a3464a ) or ( a3465a );
 a7342a <=( a3466a ) or ( a7341a );
 a7343a <=( a7342a ) or ( a7337a );
 a7346a <=( a3462a ) or ( a3463a );
 a7350a <=( a3459a ) or ( a3460a );
 a7351a <=( a3461a ) or ( a7350a );
 a7352a <=( a7351a ) or ( a7346a );
 a7353a <=( a7352a ) or ( a7343a );
 a7354a <=( a7353a ) or ( a7334a );
 a7355a <=( a7354a ) or ( a7317a );
 a7358a <=( a3457a ) or ( a3458a );
 a7361a <=( a3455a ) or ( a3456a );
 a7362a <=( a7361a ) or ( a7358a );
 a7365a <=( a3453a ) or ( a3454a );
 a7369a <=( a3450a ) or ( a3451a );
 a7370a <=( a3452a ) or ( a7369a );
 a7371a <=( a7370a ) or ( a7365a );
 a7372a <=( a7371a ) or ( a7362a );
 a7375a <=( a3448a ) or ( a3449a );
 a7378a <=( a3446a ) or ( a3447a );
 a7379a <=( a7378a ) or ( a7375a );
 a7382a <=( a3444a ) or ( a3445a );
 a7386a <=( a3441a ) or ( a3442a );
 a7387a <=( a3443a ) or ( a7386a );
 a7388a <=( a7387a ) or ( a7382a );
 a7389a <=( a7388a ) or ( a7379a );
 a7390a <=( a7389a ) or ( a7372a );
 a7393a <=( a3439a ) or ( a3440a );
 a7396a <=( a3437a ) or ( a3438a );
 a7397a <=( a7396a ) or ( a7393a );
 a7400a <=( a3435a ) or ( a3436a );
 a7404a <=( a3432a ) or ( a3433a );
 a7405a <=( a3434a ) or ( a7404a );
 a7406a <=( a7405a ) or ( a7400a );
 a7407a <=( a7406a ) or ( a7397a );
 a7410a <=( a3430a ) or ( a3431a );
 a7414a <=( a3427a ) or ( a3428a );
 a7415a <=( a3429a ) or ( a7414a );
 a7416a <=( a7415a ) or ( a7410a );
 a7419a <=( a3425a ) or ( a3426a );
 a7423a <=( a3422a ) or ( a3423a );
 a7424a <=( a3424a ) or ( a7423a );
 a7425a <=( a7424a ) or ( a7419a );
 a7426a <=( a7425a ) or ( a7416a );
 a7427a <=( a7426a ) or ( a7407a );
 a7428a <=( a7427a ) or ( a7390a );
 a7429a <=( a7428a ) or ( a7355a );
 a7430a <=( a7429a ) or ( a7282a );
 a7433a <=( a3420a ) or ( a3421a );
 a7436a <=( a3418a ) or ( a3419a );
 a7437a <=( a7436a ) or ( a7433a );
 a7440a <=( a3416a ) or ( a3417a );
 a7444a <=( a3413a ) or ( a3414a );
 a7445a <=( a3415a ) or ( a7444a );
 a7446a <=( a7445a ) or ( a7440a );
 a7447a <=( a7446a ) or ( a7437a );
 a7450a <=( a3411a ) or ( a3412a );
 a7453a <=( a3409a ) or ( a3410a );
 a7454a <=( a7453a ) or ( a7450a );
 a7457a <=( a3407a ) or ( a3408a );
 a7461a <=( a3404a ) or ( a3405a );
 a7462a <=( a3406a ) or ( a7461a );
 a7463a <=( a7462a ) or ( a7457a );
 a7464a <=( a7463a ) or ( a7454a );
 a7465a <=( a7464a ) or ( a7447a );
 a7468a <=( a3402a ) or ( a3403a );
 a7471a <=( a3400a ) or ( a3401a );
 a7472a <=( a7471a ) or ( a7468a );
 a7475a <=( a3398a ) or ( a3399a );
 a7479a <=( a3395a ) or ( a3396a );
 a7480a <=( a3397a ) or ( a7479a );
 a7481a <=( a7480a ) or ( a7475a );
 a7482a <=( a7481a ) or ( a7472a );
 a7485a <=( a3393a ) or ( a3394a );
 a7489a <=( a3390a ) or ( a3391a );
 a7490a <=( a3392a ) or ( a7489a );
 a7491a <=( a7490a ) or ( a7485a );
 a7494a <=( a3388a ) or ( a3389a );
 a7498a <=( a3385a ) or ( a3386a );
 a7499a <=( a3387a ) or ( a7498a );
 a7500a <=( a7499a ) or ( a7494a );
 a7501a <=( a7500a ) or ( a7491a );
 a7502a <=( a7501a ) or ( a7482a );
 a7503a <=( a7502a ) or ( a7465a );
 a7506a <=( a3383a ) or ( a3384a );
 a7509a <=( a3381a ) or ( a3382a );
 a7510a <=( a7509a ) or ( a7506a );
 a7513a <=( a3379a ) or ( a3380a );
 a7517a <=( a3376a ) or ( a3377a );
 a7518a <=( a3378a ) or ( a7517a );
 a7519a <=( a7518a ) or ( a7513a );
 a7520a <=( a7519a ) or ( a7510a );
 a7523a <=( a3374a ) or ( a3375a );
 a7526a <=( a3372a ) or ( a3373a );
 a7527a <=( a7526a ) or ( a7523a );
 a7530a <=( a3370a ) or ( a3371a );
 a7534a <=( a3367a ) or ( a3368a );
 a7535a <=( a3369a ) or ( a7534a );
 a7536a <=( a7535a ) or ( a7530a );
 a7537a <=( a7536a ) or ( a7527a );
 a7538a <=( a7537a ) or ( a7520a );
 a7541a <=( a3365a ) or ( a3366a );
 a7544a <=( a3363a ) or ( a3364a );
 a7545a <=( a7544a ) or ( a7541a );
 a7548a <=( a3361a ) or ( a3362a );
 a7552a <=( a3358a ) or ( a3359a );
 a7553a <=( a3360a ) or ( a7552a );
 a7554a <=( a7553a ) or ( a7548a );
 a7555a <=( a7554a ) or ( a7545a );
 a7558a <=( a3356a ) or ( a3357a );
 a7562a <=( a3353a ) or ( a3354a );
 a7563a <=( a3355a ) or ( a7562a );
 a7564a <=( a7563a ) or ( a7558a );
 a7567a <=( a3351a ) or ( a3352a );
 a7571a <=( a3348a ) or ( a3349a );
 a7572a <=( a3350a ) or ( a7571a );
 a7573a <=( a7572a ) or ( a7567a );
 a7574a <=( a7573a ) or ( a7564a );
 a7575a <=( a7574a ) or ( a7555a );
 a7576a <=( a7575a ) or ( a7538a );
 a7577a <=( a7576a ) or ( a7503a );
 a7580a <=( a3346a ) or ( a3347a );
 a7583a <=( a3344a ) or ( a3345a );
 a7584a <=( a7583a ) or ( a7580a );
 a7587a <=( a3342a ) or ( a3343a );
 a7591a <=( a3339a ) or ( a3340a );
 a7592a <=( a3341a ) or ( a7591a );
 a7593a <=( a7592a ) or ( a7587a );
 a7594a <=( a7593a ) or ( a7584a );
 a7597a <=( a3337a ) or ( a3338a );
 a7600a <=( a3335a ) or ( a3336a );
 a7601a <=( a7600a ) or ( a7597a );
 a7604a <=( a3333a ) or ( a3334a );
 a7608a <=( a3330a ) or ( a3331a );
 a7609a <=( a3332a ) or ( a7608a );
 a7610a <=( a7609a ) or ( a7604a );
 a7611a <=( a7610a ) or ( a7601a );
 a7612a <=( a7611a ) or ( a7594a );
 a7615a <=( a3328a ) or ( a3329a );
 a7618a <=( a3326a ) or ( a3327a );
 a7619a <=( a7618a ) or ( a7615a );
 a7622a <=( a3324a ) or ( a3325a );
 a7626a <=( a3321a ) or ( a3322a );
 a7627a <=( a3323a ) or ( a7626a );
 a7628a <=( a7627a ) or ( a7622a );
 a7629a <=( a7628a ) or ( a7619a );
 a7632a <=( a3319a ) or ( a3320a );
 a7636a <=( a3316a ) or ( a3317a );
 a7637a <=( a3318a ) or ( a7636a );
 a7638a <=( a7637a ) or ( a7632a );
 a7641a <=( a3314a ) or ( a3315a );
 a7645a <=( a3311a ) or ( a3312a );
 a7646a <=( a3313a ) or ( a7645a );
 a7647a <=( a7646a ) or ( a7641a );
 a7648a <=( a7647a ) or ( a7638a );
 a7649a <=( a7648a ) or ( a7629a );
 a7650a <=( a7649a ) or ( a7612a );
 a7653a <=( a3309a ) or ( a3310a );
 a7656a <=( a3307a ) or ( a3308a );
 a7657a <=( a7656a ) or ( a7653a );
 a7660a <=( a3305a ) or ( a3306a );
 a7664a <=( a3302a ) or ( a3303a );
 a7665a <=( a3304a ) or ( a7664a );
 a7666a <=( a7665a ) or ( a7660a );
 a7667a <=( a7666a ) or ( a7657a );
 a7670a <=( a3300a ) or ( a3301a );
 a7674a <=( a3297a ) or ( a3298a );
 a7675a <=( a3299a ) or ( a7674a );
 a7676a <=( a7675a ) or ( a7670a );
 a7679a <=( a3295a ) or ( a3296a );
 a7683a <=( a3292a ) or ( a3293a );
 a7684a <=( a3294a ) or ( a7683a );
 a7685a <=( a7684a ) or ( a7679a );
 a7686a <=( a7685a ) or ( a7676a );
 a7687a <=( a7686a ) or ( a7667a );
 a7690a <=( a3290a ) or ( a3291a );
 a7693a <=( a3288a ) or ( a3289a );
 a7694a <=( a7693a ) or ( a7690a );
 a7697a <=( a3286a ) or ( a3287a );
 a7701a <=( a3283a ) or ( a3284a );
 a7702a <=( a3285a ) or ( a7701a );
 a7703a <=( a7702a ) or ( a7697a );
 a7704a <=( a7703a ) or ( a7694a );
 a7707a <=( a3281a ) or ( a3282a );
 a7711a <=( a3278a ) or ( a3279a );
 a7712a <=( a3280a ) or ( a7711a );
 a7713a <=( a7712a ) or ( a7707a );
 a7716a <=( a3276a ) or ( a3277a );
 a7720a <=( a3273a ) or ( a3274a );
 a7721a <=( a3275a ) or ( a7720a );
 a7722a <=( a7721a ) or ( a7716a );
 a7723a <=( a7722a ) or ( a7713a );
 a7724a <=( a7723a ) or ( a7704a );
 a7725a <=( a7724a ) or ( a7687a );
 a7726a <=( a7725a ) or ( a7650a );
 a7727a <=( a7726a ) or ( a7577a );
 a7728a <=( a7727a ) or ( a7430a );
 a7731a <=( a3271a ) or ( a3272a );
 a7734a <=( a3269a ) or ( a3270a );
 a7735a <=( a7734a ) or ( a7731a );
 a7738a <=( a3267a ) or ( a3268a );
 a7742a <=( a3264a ) or ( a3265a );
 a7743a <=( a3266a ) or ( a7742a );
 a7744a <=( a7743a ) or ( a7738a );
 a7745a <=( a7744a ) or ( a7735a );
 a7748a <=( a3262a ) or ( a3263a );
 a7751a <=( a3260a ) or ( a3261a );
 a7752a <=( a7751a ) or ( a7748a );
 a7755a <=( a3258a ) or ( a3259a );
 a7759a <=( a3255a ) or ( a3256a );
 a7760a <=( a3257a ) or ( a7759a );
 a7761a <=( a7760a ) or ( a7755a );
 a7762a <=( a7761a ) or ( a7752a );
 a7763a <=( a7762a ) or ( a7745a );
 a7766a <=( a3253a ) or ( a3254a );
 a7769a <=( a3251a ) or ( a3252a );
 a7770a <=( a7769a ) or ( a7766a );
 a7773a <=( a3249a ) or ( a3250a );
 a7777a <=( a3246a ) or ( a3247a );
 a7778a <=( a3248a ) or ( a7777a );
 a7779a <=( a7778a ) or ( a7773a );
 a7780a <=( a7779a ) or ( a7770a );
 a7783a <=( a3244a ) or ( a3245a );
 a7787a <=( a3241a ) or ( a3242a );
 a7788a <=( a3243a ) or ( a7787a );
 a7789a <=( a7788a ) or ( a7783a );
 a7792a <=( a3239a ) or ( a3240a );
 a7796a <=( a3236a ) or ( a3237a );
 a7797a <=( a3238a ) or ( a7796a );
 a7798a <=( a7797a ) or ( a7792a );
 a7799a <=( a7798a ) or ( a7789a );
 a7800a <=( a7799a ) or ( a7780a );
 a7801a <=( a7800a ) or ( a7763a );
 a7804a <=( a3234a ) or ( a3235a );
 a7807a <=( a3232a ) or ( a3233a );
 a7808a <=( a7807a ) or ( a7804a );
 a7811a <=( a3230a ) or ( a3231a );
 a7815a <=( a3227a ) or ( a3228a );
 a7816a <=( a3229a ) or ( a7815a );
 a7817a <=( a7816a ) or ( a7811a );
 a7818a <=( a7817a ) or ( a7808a );
 a7821a <=( a3225a ) or ( a3226a );
 a7824a <=( a3223a ) or ( a3224a );
 a7825a <=( a7824a ) or ( a7821a );
 a7828a <=( a3221a ) or ( a3222a );
 a7832a <=( a3218a ) or ( a3219a );
 a7833a <=( a3220a ) or ( a7832a );
 a7834a <=( a7833a ) or ( a7828a );
 a7835a <=( a7834a ) or ( a7825a );
 a7836a <=( a7835a ) or ( a7818a );
 a7839a <=( a3216a ) or ( a3217a );
 a7842a <=( a3214a ) or ( a3215a );
 a7843a <=( a7842a ) or ( a7839a );
 a7846a <=( a3212a ) or ( a3213a );
 a7850a <=( a3209a ) or ( a3210a );
 a7851a <=( a3211a ) or ( a7850a );
 a7852a <=( a7851a ) or ( a7846a );
 a7853a <=( a7852a ) or ( a7843a );
 a7856a <=( a3207a ) or ( a3208a );
 a7860a <=( a3204a ) or ( a3205a );
 a7861a <=( a3206a ) or ( a7860a );
 a7862a <=( a7861a ) or ( a7856a );
 a7865a <=( a3202a ) or ( a3203a );
 a7869a <=( a3199a ) or ( a3200a );
 a7870a <=( a3201a ) or ( a7869a );
 a7871a <=( a7870a ) or ( a7865a );
 a7872a <=( a7871a ) or ( a7862a );
 a7873a <=( a7872a ) or ( a7853a );
 a7874a <=( a7873a ) or ( a7836a );
 a7875a <=( a7874a ) or ( a7801a );
 a7878a <=( a3197a ) or ( a3198a );
 a7881a <=( a3195a ) or ( a3196a );
 a7882a <=( a7881a ) or ( a7878a );
 a7885a <=( a3193a ) or ( a3194a );
 a7889a <=( a3190a ) or ( a3191a );
 a7890a <=( a3192a ) or ( a7889a );
 a7891a <=( a7890a ) or ( a7885a );
 a7892a <=( a7891a ) or ( a7882a );
 a7895a <=( a3188a ) or ( a3189a );
 a7898a <=( a3186a ) or ( a3187a );
 a7899a <=( a7898a ) or ( a7895a );
 a7902a <=( a3184a ) or ( a3185a );
 a7906a <=( a3181a ) or ( a3182a );
 a7907a <=( a3183a ) or ( a7906a );
 a7908a <=( a7907a ) or ( a7902a );
 a7909a <=( a7908a ) or ( a7899a );
 a7910a <=( a7909a ) or ( a7892a );
 a7913a <=( a3179a ) or ( a3180a );
 a7916a <=( a3177a ) or ( a3178a );
 a7917a <=( a7916a ) or ( a7913a );
 a7920a <=( a3175a ) or ( a3176a );
 a7924a <=( a3172a ) or ( a3173a );
 a7925a <=( a3174a ) or ( a7924a );
 a7926a <=( a7925a ) or ( a7920a );
 a7927a <=( a7926a ) or ( a7917a );
 a7930a <=( a3170a ) or ( a3171a );
 a7934a <=( a3167a ) or ( a3168a );
 a7935a <=( a3169a ) or ( a7934a );
 a7936a <=( a7935a ) or ( a7930a );
 a7939a <=( a3165a ) or ( a3166a );
 a7943a <=( a3162a ) or ( a3163a );
 a7944a <=( a3164a ) or ( a7943a );
 a7945a <=( a7944a ) or ( a7939a );
 a7946a <=( a7945a ) or ( a7936a );
 a7947a <=( a7946a ) or ( a7927a );
 a7948a <=( a7947a ) or ( a7910a );
 a7951a <=( a3160a ) or ( a3161a );
 a7954a <=( a3158a ) or ( a3159a );
 a7955a <=( a7954a ) or ( a7951a );
 a7958a <=( a3156a ) or ( a3157a );
 a7962a <=( a3153a ) or ( a3154a );
 a7963a <=( a3155a ) or ( a7962a );
 a7964a <=( a7963a ) or ( a7958a );
 a7965a <=( a7964a ) or ( a7955a );
 a7968a <=( a3151a ) or ( a3152a );
 a7972a <=( a3148a ) or ( a3149a );
 a7973a <=( a3150a ) or ( a7972a );
 a7974a <=( a7973a ) or ( a7968a );
 a7977a <=( a3146a ) or ( a3147a );
 a7981a <=( a3143a ) or ( a3144a );
 a7982a <=( a3145a ) or ( a7981a );
 a7983a <=( a7982a ) or ( a7977a );
 a7984a <=( a7983a ) or ( a7974a );
 a7985a <=( a7984a ) or ( a7965a );
 a7988a <=( a3141a ) or ( a3142a );
 a7991a <=( a3139a ) or ( a3140a );
 a7992a <=( a7991a ) or ( a7988a );
 a7995a <=( a3137a ) or ( a3138a );
 a7999a <=( a3134a ) or ( a3135a );
 a8000a <=( a3136a ) or ( a7999a );
 a8001a <=( a8000a ) or ( a7995a );
 a8002a <=( a8001a ) or ( a7992a );
 a8005a <=( a3132a ) or ( a3133a );
 a8009a <=( a3129a ) or ( a3130a );
 a8010a <=( a3131a ) or ( a8009a );
 a8011a <=( a8010a ) or ( a8005a );
 a8014a <=( a3127a ) or ( a3128a );
 a8018a <=( a3124a ) or ( a3125a );
 a8019a <=( a3126a ) or ( a8018a );
 a8020a <=( a8019a ) or ( a8014a );
 a8021a <=( a8020a ) or ( a8011a );
 a8022a <=( a8021a ) or ( a8002a );
 a8023a <=( a8022a ) or ( a7985a );
 a8024a <=( a8023a ) or ( a7948a );
 a8025a <=( a8024a ) or ( a7875a );
 a8028a <=( a3122a ) or ( a3123a );
 a8031a <=( a3120a ) or ( a3121a );
 a8032a <=( a8031a ) or ( a8028a );
 a8035a <=( a3118a ) or ( a3119a );
 a8039a <=( a3115a ) or ( a3116a );
 a8040a <=( a3117a ) or ( a8039a );
 a8041a <=( a8040a ) or ( a8035a );
 a8042a <=( a8041a ) or ( a8032a );
 a8045a <=( a3113a ) or ( a3114a );
 a8048a <=( a3111a ) or ( a3112a );
 a8049a <=( a8048a ) or ( a8045a );
 a8052a <=( a3109a ) or ( a3110a );
 a8056a <=( a3106a ) or ( a3107a );
 a8057a <=( a3108a ) or ( a8056a );
 a8058a <=( a8057a ) or ( a8052a );
 a8059a <=( a8058a ) or ( a8049a );
 a8060a <=( a8059a ) or ( a8042a );
 a8063a <=( a3104a ) or ( a3105a );
 a8066a <=( a3102a ) or ( a3103a );
 a8067a <=( a8066a ) or ( a8063a );
 a8070a <=( a3100a ) or ( a3101a );
 a8074a <=( a3097a ) or ( a3098a );
 a8075a <=( a3099a ) or ( a8074a );
 a8076a <=( a8075a ) or ( a8070a );
 a8077a <=( a8076a ) or ( a8067a );
 a8080a <=( a3095a ) or ( a3096a );
 a8084a <=( a3092a ) or ( a3093a );
 a8085a <=( a3094a ) or ( a8084a );
 a8086a <=( a8085a ) or ( a8080a );
 a8089a <=( a3090a ) or ( a3091a );
 a8093a <=( a3087a ) or ( a3088a );
 a8094a <=( a3089a ) or ( a8093a );
 a8095a <=( a8094a ) or ( a8089a );
 a8096a <=( a8095a ) or ( a8086a );
 a8097a <=( a8096a ) or ( a8077a );
 a8098a <=( a8097a ) or ( a8060a );
 a8101a <=( a3085a ) or ( a3086a );
 a8104a <=( a3083a ) or ( a3084a );
 a8105a <=( a8104a ) or ( a8101a );
 a8108a <=( a3081a ) or ( a3082a );
 a8112a <=( a3078a ) or ( a3079a );
 a8113a <=( a3080a ) or ( a8112a );
 a8114a <=( a8113a ) or ( a8108a );
 a8115a <=( a8114a ) or ( a8105a );
 a8118a <=( a3076a ) or ( a3077a );
 a8121a <=( a3074a ) or ( a3075a );
 a8122a <=( a8121a ) or ( a8118a );
 a8125a <=( a3072a ) or ( a3073a );
 a8129a <=( a3069a ) or ( a3070a );
 a8130a <=( a3071a ) or ( a8129a );
 a8131a <=( a8130a ) or ( a8125a );
 a8132a <=( a8131a ) or ( a8122a );
 a8133a <=( a8132a ) or ( a8115a );
 a8136a <=( a3067a ) or ( a3068a );
 a8139a <=( a3065a ) or ( a3066a );
 a8140a <=( a8139a ) or ( a8136a );
 a8143a <=( a3063a ) or ( a3064a );
 a8147a <=( a3060a ) or ( a3061a );
 a8148a <=( a3062a ) or ( a8147a );
 a8149a <=( a8148a ) or ( a8143a );
 a8150a <=( a8149a ) or ( a8140a );
 a8153a <=( a3058a ) or ( a3059a );
 a8157a <=( a3055a ) or ( a3056a );
 a8158a <=( a3057a ) or ( a8157a );
 a8159a <=( a8158a ) or ( a8153a );
 a8162a <=( a3053a ) or ( a3054a );
 a8166a <=( a3050a ) or ( a3051a );
 a8167a <=( a3052a ) or ( a8166a );
 a8168a <=( a8167a ) or ( a8162a );
 a8169a <=( a8168a ) or ( a8159a );
 a8170a <=( a8169a ) or ( a8150a );
 a8171a <=( a8170a ) or ( a8133a );
 a8172a <=( a8171a ) or ( a8098a );
 a8175a <=( a3048a ) or ( a3049a );
 a8178a <=( a3046a ) or ( a3047a );
 a8179a <=( a8178a ) or ( a8175a );
 a8182a <=( a3044a ) or ( a3045a );
 a8186a <=( a3041a ) or ( a3042a );
 a8187a <=( a3043a ) or ( a8186a );
 a8188a <=( a8187a ) or ( a8182a );
 a8189a <=( a8188a ) or ( a8179a );
 a8192a <=( a3039a ) or ( a3040a );
 a8195a <=( a3037a ) or ( a3038a );
 a8196a <=( a8195a ) or ( a8192a );
 a8199a <=( a3035a ) or ( a3036a );
 a8203a <=( a3032a ) or ( a3033a );
 a8204a <=( a3034a ) or ( a8203a );
 a8205a <=( a8204a ) or ( a8199a );
 a8206a <=( a8205a ) or ( a8196a );
 a8207a <=( a8206a ) or ( a8189a );
 a8210a <=( a3030a ) or ( a3031a );
 a8213a <=( a3028a ) or ( a3029a );
 a8214a <=( a8213a ) or ( a8210a );
 a8217a <=( a3026a ) or ( a3027a );
 a8221a <=( a3023a ) or ( a3024a );
 a8222a <=( a3025a ) or ( a8221a );
 a8223a <=( a8222a ) or ( a8217a );
 a8224a <=( a8223a ) or ( a8214a );
 a8227a <=( a3021a ) or ( a3022a );
 a8231a <=( a3018a ) or ( a3019a );
 a8232a <=( a3020a ) or ( a8231a );
 a8233a <=( a8232a ) or ( a8227a );
 a8236a <=( a3016a ) or ( a3017a );
 a8240a <=( a3013a ) or ( a3014a );
 a8241a <=( a3015a ) or ( a8240a );
 a8242a <=( a8241a ) or ( a8236a );
 a8243a <=( a8242a ) or ( a8233a );
 a8244a <=( a8243a ) or ( a8224a );
 a8245a <=( a8244a ) or ( a8207a );
 a8248a <=( a3011a ) or ( a3012a );
 a8251a <=( a3009a ) or ( a3010a );
 a8252a <=( a8251a ) or ( a8248a );
 a8255a <=( a3007a ) or ( a3008a );
 a8259a <=( a3004a ) or ( a3005a );
 a8260a <=( a3006a ) or ( a8259a );
 a8261a <=( a8260a ) or ( a8255a );
 a8262a <=( a8261a ) or ( a8252a );
 a8265a <=( a3002a ) or ( a3003a );
 a8269a <=( a2999a ) or ( a3000a );
 a8270a <=( a3001a ) or ( a8269a );
 a8271a <=( a8270a ) or ( a8265a );
 a8274a <=( a2997a ) or ( a2998a );
 a8278a <=( a2994a ) or ( a2995a );
 a8279a <=( a2996a ) or ( a8278a );
 a8280a <=( a8279a ) or ( a8274a );
 a8281a <=( a8280a ) or ( a8271a );
 a8282a <=( a8281a ) or ( a8262a );
 a8285a <=( a2992a ) or ( a2993a );
 a8288a <=( a2990a ) or ( a2991a );
 a8289a <=( a8288a ) or ( a8285a );
 a8292a <=( a2988a ) or ( a2989a );
 a8296a <=( a2985a ) or ( a2986a );
 a8297a <=( a2987a ) or ( a8296a );
 a8298a <=( a8297a ) or ( a8292a );
 a8299a <=( a8298a ) or ( a8289a );
 a8302a <=( a2983a ) or ( a2984a );
 a8306a <=( a2980a ) or ( a2981a );
 a8307a <=( a2982a ) or ( a8306a );
 a8308a <=( a8307a ) or ( a8302a );
 a8311a <=( a2978a ) or ( a2979a );
 a8315a <=( a2975a ) or ( a2976a );
 a8316a <=( a2977a ) or ( a8315a );
 a8317a <=( a8316a ) or ( a8311a );
 a8318a <=( a8317a ) or ( a8308a );
 a8319a <=( a8318a ) or ( a8299a );
 a8320a <=( a8319a ) or ( a8282a );
 a8321a <=( a8320a ) or ( a8245a );
 a8322a <=( a8321a ) or ( a8172a );
 a8323a <=( a8322a ) or ( a8025a );
 a8324a <=( a8323a ) or ( a7728a );
 a8327a <=( a2973a ) or ( a2974a );
 a8330a <=( a2971a ) or ( a2972a );
 a8331a <=( a8330a ) or ( a8327a );
 a8334a <=( a2969a ) or ( a2970a );
 a8338a <=( a2966a ) or ( a2967a );
 a8339a <=( a2968a ) or ( a8338a );
 a8340a <=( a8339a ) or ( a8334a );
 a8341a <=( a8340a ) or ( a8331a );
 a8344a <=( a2964a ) or ( a2965a );
 a8347a <=( a2962a ) or ( a2963a );
 a8348a <=( a8347a ) or ( a8344a );
 a8351a <=( a2960a ) or ( a2961a );
 a8355a <=( a2957a ) or ( a2958a );
 a8356a <=( a2959a ) or ( a8355a );
 a8357a <=( a8356a ) or ( a8351a );
 a8358a <=( a8357a ) or ( a8348a );
 a8359a <=( a8358a ) or ( a8341a );
 a8362a <=( a2955a ) or ( a2956a );
 a8365a <=( a2953a ) or ( a2954a );
 a8366a <=( a8365a ) or ( a8362a );
 a8369a <=( a2951a ) or ( a2952a );
 a8373a <=( a2948a ) or ( a2949a );
 a8374a <=( a2950a ) or ( a8373a );
 a8375a <=( a8374a ) or ( a8369a );
 a8376a <=( a8375a ) or ( a8366a );
 a8379a <=( a2946a ) or ( a2947a );
 a8383a <=( a2943a ) or ( a2944a );
 a8384a <=( a2945a ) or ( a8383a );
 a8385a <=( a8384a ) or ( a8379a );
 a8388a <=( a2941a ) or ( a2942a );
 a8392a <=( a2938a ) or ( a2939a );
 a8393a <=( a2940a ) or ( a8392a );
 a8394a <=( a8393a ) or ( a8388a );
 a8395a <=( a8394a ) or ( a8385a );
 a8396a <=( a8395a ) or ( a8376a );
 a8397a <=( a8396a ) or ( a8359a );
 a8400a <=( a2936a ) or ( a2937a );
 a8403a <=( a2934a ) or ( a2935a );
 a8404a <=( a8403a ) or ( a8400a );
 a8407a <=( a2932a ) or ( a2933a );
 a8411a <=( a2929a ) or ( a2930a );
 a8412a <=( a2931a ) or ( a8411a );
 a8413a <=( a8412a ) or ( a8407a );
 a8414a <=( a8413a ) or ( a8404a );
 a8417a <=( a2927a ) or ( a2928a );
 a8420a <=( a2925a ) or ( a2926a );
 a8421a <=( a8420a ) or ( a8417a );
 a8424a <=( a2923a ) or ( a2924a );
 a8428a <=( a2920a ) or ( a2921a );
 a8429a <=( a2922a ) or ( a8428a );
 a8430a <=( a8429a ) or ( a8424a );
 a8431a <=( a8430a ) or ( a8421a );
 a8432a <=( a8431a ) or ( a8414a );
 a8435a <=( a2918a ) or ( a2919a );
 a8438a <=( a2916a ) or ( a2917a );
 a8439a <=( a8438a ) or ( a8435a );
 a8442a <=( a2914a ) or ( a2915a );
 a8446a <=( a2911a ) or ( a2912a );
 a8447a <=( a2913a ) or ( a8446a );
 a8448a <=( a8447a ) or ( a8442a );
 a8449a <=( a8448a ) or ( a8439a );
 a8452a <=( a2909a ) or ( a2910a );
 a8456a <=( a2906a ) or ( a2907a );
 a8457a <=( a2908a ) or ( a8456a );
 a8458a <=( a8457a ) or ( a8452a );
 a8461a <=( a2904a ) or ( a2905a );
 a8465a <=( a2901a ) or ( a2902a );
 a8466a <=( a2903a ) or ( a8465a );
 a8467a <=( a8466a ) or ( a8461a );
 a8468a <=( a8467a ) or ( a8458a );
 a8469a <=( a8468a ) or ( a8449a );
 a8470a <=( a8469a ) or ( a8432a );
 a8471a <=( a8470a ) or ( a8397a );
 a8474a <=( a2899a ) or ( a2900a );
 a8477a <=( a2897a ) or ( a2898a );
 a8478a <=( a8477a ) or ( a8474a );
 a8481a <=( a2895a ) or ( a2896a );
 a8485a <=( a2892a ) or ( a2893a );
 a8486a <=( a2894a ) or ( a8485a );
 a8487a <=( a8486a ) or ( a8481a );
 a8488a <=( a8487a ) or ( a8478a );
 a8491a <=( a2890a ) or ( a2891a );
 a8494a <=( a2888a ) or ( a2889a );
 a8495a <=( a8494a ) or ( a8491a );
 a8498a <=( a2886a ) or ( a2887a );
 a8502a <=( a2883a ) or ( a2884a );
 a8503a <=( a2885a ) or ( a8502a );
 a8504a <=( a8503a ) or ( a8498a );
 a8505a <=( a8504a ) or ( a8495a );
 a8506a <=( a8505a ) or ( a8488a );
 a8509a <=( a2881a ) or ( a2882a );
 a8512a <=( a2879a ) or ( a2880a );
 a8513a <=( a8512a ) or ( a8509a );
 a8516a <=( a2877a ) or ( a2878a );
 a8520a <=( a2874a ) or ( a2875a );
 a8521a <=( a2876a ) or ( a8520a );
 a8522a <=( a8521a ) or ( a8516a );
 a8523a <=( a8522a ) or ( a8513a );
 a8526a <=( a2872a ) or ( a2873a );
 a8530a <=( a2869a ) or ( a2870a );
 a8531a <=( a2871a ) or ( a8530a );
 a8532a <=( a8531a ) or ( a8526a );
 a8535a <=( a2867a ) or ( a2868a );
 a8539a <=( a2864a ) or ( a2865a );
 a8540a <=( a2866a ) or ( a8539a );
 a8541a <=( a8540a ) or ( a8535a );
 a8542a <=( a8541a ) or ( a8532a );
 a8543a <=( a8542a ) or ( a8523a );
 a8544a <=( a8543a ) or ( a8506a );
 a8547a <=( a2862a ) or ( a2863a );
 a8550a <=( a2860a ) or ( a2861a );
 a8551a <=( a8550a ) or ( a8547a );
 a8554a <=( a2858a ) or ( a2859a );
 a8558a <=( a2855a ) or ( a2856a );
 a8559a <=( a2857a ) or ( a8558a );
 a8560a <=( a8559a ) or ( a8554a );
 a8561a <=( a8560a ) or ( a8551a );
 a8564a <=( a2853a ) or ( a2854a );
 a8567a <=( a2851a ) or ( a2852a );
 a8568a <=( a8567a ) or ( a8564a );
 a8571a <=( a2849a ) or ( a2850a );
 a8575a <=( a2846a ) or ( a2847a );
 a8576a <=( a2848a ) or ( a8575a );
 a8577a <=( a8576a ) or ( a8571a );
 a8578a <=( a8577a ) or ( a8568a );
 a8579a <=( a8578a ) or ( a8561a );
 a8582a <=( a2844a ) or ( a2845a );
 a8585a <=( a2842a ) or ( a2843a );
 a8586a <=( a8585a ) or ( a8582a );
 a8589a <=( a2840a ) or ( a2841a );
 a8593a <=( a2837a ) or ( a2838a );
 a8594a <=( a2839a ) or ( a8593a );
 a8595a <=( a8594a ) or ( a8589a );
 a8596a <=( a8595a ) or ( a8586a );
 a8599a <=( a2835a ) or ( a2836a );
 a8603a <=( a2832a ) or ( a2833a );
 a8604a <=( a2834a ) or ( a8603a );
 a8605a <=( a8604a ) or ( a8599a );
 a8608a <=( a2830a ) or ( a2831a );
 a8612a <=( a2827a ) or ( a2828a );
 a8613a <=( a2829a ) or ( a8612a );
 a8614a <=( a8613a ) or ( a8608a );
 a8615a <=( a8614a ) or ( a8605a );
 a8616a <=( a8615a ) or ( a8596a );
 a8617a <=( a8616a ) or ( a8579a );
 a8618a <=( a8617a ) or ( a8544a );
 a8619a <=( a8618a ) or ( a8471a );
 a8622a <=( a2825a ) or ( a2826a );
 a8625a <=( a2823a ) or ( a2824a );
 a8626a <=( a8625a ) or ( a8622a );
 a8629a <=( a2821a ) or ( a2822a );
 a8633a <=( a2818a ) or ( a2819a );
 a8634a <=( a2820a ) or ( a8633a );
 a8635a <=( a8634a ) or ( a8629a );
 a8636a <=( a8635a ) or ( a8626a );
 a8639a <=( a2816a ) or ( a2817a );
 a8642a <=( a2814a ) or ( a2815a );
 a8643a <=( a8642a ) or ( a8639a );
 a8646a <=( a2812a ) or ( a2813a );
 a8650a <=( a2809a ) or ( a2810a );
 a8651a <=( a2811a ) or ( a8650a );
 a8652a <=( a8651a ) or ( a8646a );
 a8653a <=( a8652a ) or ( a8643a );
 a8654a <=( a8653a ) or ( a8636a );
 a8657a <=( a2807a ) or ( a2808a );
 a8660a <=( a2805a ) or ( a2806a );
 a8661a <=( a8660a ) or ( a8657a );
 a8664a <=( a2803a ) or ( a2804a );
 a8668a <=( a2800a ) or ( a2801a );
 a8669a <=( a2802a ) or ( a8668a );
 a8670a <=( a8669a ) or ( a8664a );
 a8671a <=( a8670a ) or ( a8661a );
 a8674a <=( a2798a ) or ( a2799a );
 a8678a <=( a2795a ) or ( a2796a );
 a8679a <=( a2797a ) or ( a8678a );
 a8680a <=( a8679a ) or ( a8674a );
 a8683a <=( a2793a ) or ( a2794a );
 a8687a <=( a2790a ) or ( a2791a );
 a8688a <=( a2792a ) or ( a8687a );
 a8689a <=( a8688a ) or ( a8683a );
 a8690a <=( a8689a ) or ( a8680a );
 a8691a <=( a8690a ) or ( a8671a );
 a8692a <=( a8691a ) or ( a8654a );
 a8695a <=( a2788a ) or ( a2789a );
 a8698a <=( a2786a ) or ( a2787a );
 a8699a <=( a8698a ) or ( a8695a );
 a8702a <=( a2784a ) or ( a2785a );
 a8706a <=( a2781a ) or ( a2782a );
 a8707a <=( a2783a ) or ( a8706a );
 a8708a <=( a8707a ) or ( a8702a );
 a8709a <=( a8708a ) or ( a8699a );
 a8712a <=( a2779a ) or ( a2780a );
 a8715a <=( a2777a ) or ( a2778a );
 a8716a <=( a8715a ) or ( a8712a );
 a8719a <=( a2775a ) or ( a2776a );
 a8723a <=( a2772a ) or ( a2773a );
 a8724a <=( a2774a ) or ( a8723a );
 a8725a <=( a8724a ) or ( a8719a );
 a8726a <=( a8725a ) or ( a8716a );
 a8727a <=( a8726a ) or ( a8709a );
 a8730a <=( a2770a ) or ( a2771a );
 a8733a <=( a2768a ) or ( a2769a );
 a8734a <=( a8733a ) or ( a8730a );
 a8737a <=( a2766a ) or ( a2767a );
 a8741a <=( a2763a ) or ( a2764a );
 a8742a <=( a2765a ) or ( a8741a );
 a8743a <=( a8742a ) or ( a8737a );
 a8744a <=( a8743a ) or ( a8734a );
 a8747a <=( a2761a ) or ( a2762a );
 a8751a <=( a2758a ) or ( a2759a );
 a8752a <=( a2760a ) or ( a8751a );
 a8753a <=( a8752a ) or ( a8747a );
 a8756a <=( a2756a ) or ( a2757a );
 a8760a <=( a2753a ) or ( a2754a );
 a8761a <=( a2755a ) or ( a8760a );
 a8762a <=( a8761a ) or ( a8756a );
 a8763a <=( a8762a ) or ( a8753a );
 a8764a <=( a8763a ) or ( a8744a );
 a8765a <=( a8764a ) or ( a8727a );
 a8766a <=( a8765a ) or ( a8692a );
 a8769a <=( a2751a ) or ( a2752a );
 a8772a <=( a2749a ) or ( a2750a );
 a8773a <=( a8772a ) or ( a8769a );
 a8776a <=( a2747a ) or ( a2748a );
 a8780a <=( a2744a ) or ( a2745a );
 a8781a <=( a2746a ) or ( a8780a );
 a8782a <=( a8781a ) or ( a8776a );
 a8783a <=( a8782a ) or ( a8773a );
 a8786a <=( a2742a ) or ( a2743a );
 a8789a <=( a2740a ) or ( a2741a );
 a8790a <=( a8789a ) or ( a8786a );
 a8793a <=( a2738a ) or ( a2739a );
 a8797a <=( a2735a ) or ( a2736a );
 a8798a <=( a2737a ) or ( a8797a );
 a8799a <=( a8798a ) or ( a8793a );
 a8800a <=( a8799a ) or ( a8790a );
 a8801a <=( a8800a ) or ( a8783a );
 a8804a <=( a2733a ) or ( a2734a );
 a8807a <=( a2731a ) or ( a2732a );
 a8808a <=( a8807a ) or ( a8804a );
 a8811a <=( a2729a ) or ( a2730a );
 a8815a <=( a2726a ) or ( a2727a );
 a8816a <=( a2728a ) or ( a8815a );
 a8817a <=( a8816a ) or ( a8811a );
 a8818a <=( a8817a ) or ( a8808a );
 a8821a <=( a2724a ) or ( a2725a );
 a8825a <=( a2721a ) or ( a2722a );
 a8826a <=( a2723a ) or ( a8825a );
 a8827a <=( a8826a ) or ( a8821a );
 a8830a <=( a2719a ) or ( a2720a );
 a8834a <=( a2716a ) or ( a2717a );
 a8835a <=( a2718a ) or ( a8834a );
 a8836a <=( a8835a ) or ( a8830a );
 a8837a <=( a8836a ) or ( a8827a );
 a8838a <=( a8837a ) or ( a8818a );
 a8839a <=( a8838a ) or ( a8801a );
 a8842a <=( a2714a ) or ( a2715a );
 a8845a <=( a2712a ) or ( a2713a );
 a8846a <=( a8845a ) or ( a8842a );
 a8849a <=( a2710a ) or ( a2711a );
 a8853a <=( a2707a ) or ( a2708a );
 a8854a <=( a2709a ) or ( a8853a );
 a8855a <=( a8854a ) or ( a8849a );
 a8856a <=( a8855a ) or ( a8846a );
 a8859a <=( a2705a ) or ( a2706a );
 a8863a <=( a2702a ) or ( a2703a );
 a8864a <=( a2704a ) or ( a8863a );
 a8865a <=( a8864a ) or ( a8859a );
 a8868a <=( a2700a ) or ( a2701a );
 a8872a <=( a2697a ) or ( a2698a );
 a8873a <=( a2699a ) or ( a8872a );
 a8874a <=( a8873a ) or ( a8868a );
 a8875a <=( a8874a ) or ( a8865a );
 a8876a <=( a8875a ) or ( a8856a );
 a8879a <=( a2695a ) or ( a2696a );
 a8882a <=( a2693a ) or ( a2694a );
 a8883a <=( a8882a ) or ( a8879a );
 a8886a <=( a2691a ) or ( a2692a );
 a8890a <=( a2688a ) or ( a2689a );
 a8891a <=( a2690a ) or ( a8890a );
 a8892a <=( a8891a ) or ( a8886a );
 a8893a <=( a8892a ) or ( a8883a );
 a8896a <=( a2686a ) or ( a2687a );
 a8900a <=( a2683a ) or ( a2684a );
 a8901a <=( a2685a ) or ( a8900a );
 a8902a <=( a8901a ) or ( a8896a );
 a8905a <=( a2681a ) or ( a2682a );
 a8909a <=( a2678a ) or ( a2679a );
 a8910a <=( a2680a ) or ( a8909a );
 a8911a <=( a8910a ) or ( a8905a );
 a8912a <=( a8911a ) or ( a8902a );
 a8913a <=( a8912a ) or ( a8893a );
 a8914a <=( a8913a ) or ( a8876a );
 a8915a <=( a8914a ) or ( a8839a );
 a8916a <=( a8915a ) or ( a8766a );
 a8917a <=( a8916a ) or ( a8619a );
 a8920a <=( a2676a ) or ( a2677a );
 a8923a <=( a2674a ) or ( a2675a );
 a8924a <=( a8923a ) or ( a8920a );
 a8927a <=( a2672a ) or ( a2673a );
 a8931a <=( a2669a ) or ( a2670a );
 a8932a <=( a2671a ) or ( a8931a );
 a8933a <=( a8932a ) or ( a8927a );
 a8934a <=( a8933a ) or ( a8924a );
 a8937a <=( a2667a ) or ( a2668a );
 a8940a <=( a2665a ) or ( a2666a );
 a8941a <=( a8940a ) or ( a8937a );
 a8944a <=( a2663a ) or ( a2664a );
 a8948a <=( a2660a ) or ( a2661a );
 a8949a <=( a2662a ) or ( a8948a );
 a8950a <=( a8949a ) or ( a8944a );
 a8951a <=( a8950a ) or ( a8941a );
 a8952a <=( a8951a ) or ( a8934a );
 a8955a <=( a2658a ) or ( a2659a );
 a8958a <=( a2656a ) or ( a2657a );
 a8959a <=( a8958a ) or ( a8955a );
 a8962a <=( a2654a ) or ( a2655a );
 a8966a <=( a2651a ) or ( a2652a );
 a8967a <=( a2653a ) or ( a8966a );
 a8968a <=( a8967a ) or ( a8962a );
 a8969a <=( a8968a ) or ( a8959a );
 a8972a <=( a2649a ) or ( a2650a );
 a8976a <=( a2646a ) or ( a2647a );
 a8977a <=( a2648a ) or ( a8976a );
 a8978a <=( a8977a ) or ( a8972a );
 a8981a <=( a2644a ) or ( a2645a );
 a8985a <=( a2641a ) or ( a2642a );
 a8986a <=( a2643a ) or ( a8985a );
 a8987a <=( a8986a ) or ( a8981a );
 a8988a <=( a8987a ) or ( a8978a );
 a8989a <=( a8988a ) or ( a8969a );
 a8990a <=( a8989a ) or ( a8952a );
 a8993a <=( a2639a ) or ( a2640a );
 a8996a <=( a2637a ) or ( a2638a );
 a8997a <=( a8996a ) or ( a8993a );
 a9000a <=( a2635a ) or ( a2636a );
 a9004a <=( a2632a ) or ( a2633a );
 a9005a <=( a2634a ) or ( a9004a );
 a9006a <=( a9005a ) or ( a9000a );
 a9007a <=( a9006a ) or ( a8997a );
 a9010a <=( a2630a ) or ( a2631a );
 a9013a <=( a2628a ) or ( a2629a );
 a9014a <=( a9013a ) or ( a9010a );
 a9017a <=( a2626a ) or ( a2627a );
 a9021a <=( a2623a ) or ( a2624a );
 a9022a <=( a2625a ) or ( a9021a );
 a9023a <=( a9022a ) or ( a9017a );
 a9024a <=( a9023a ) or ( a9014a );
 a9025a <=( a9024a ) or ( a9007a );
 a9028a <=( a2621a ) or ( a2622a );
 a9031a <=( a2619a ) or ( a2620a );
 a9032a <=( a9031a ) or ( a9028a );
 a9035a <=( a2617a ) or ( a2618a );
 a9039a <=( a2614a ) or ( a2615a );
 a9040a <=( a2616a ) or ( a9039a );
 a9041a <=( a9040a ) or ( a9035a );
 a9042a <=( a9041a ) or ( a9032a );
 a9045a <=( a2612a ) or ( a2613a );
 a9049a <=( a2609a ) or ( a2610a );
 a9050a <=( a2611a ) or ( a9049a );
 a9051a <=( a9050a ) or ( a9045a );
 a9054a <=( a2607a ) or ( a2608a );
 a9058a <=( a2604a ) or ( a2605a );
 a9059a <=( a2606a ) or ( a9058a );
 a9060a <=( a9059a ) or ( a9054a );
 a9061a <=( a9060a ) or ( a9051a );
 a9062a <=( a9061a ) or ( a9042a );
 a9063a <=( a9062a ) or ( a9025a );
 a9064a <=( a9063a ) or ( a8990a );
 a9067a <=( a2602a ) or ( a2603a );
 a9070a <=( a2600a ) or ( a2601a );
 a9071a <=( a9070a ) or ( a9067a );
 a9074a <=( a2598a ) or ( a2599a );
 a9078a <=( a2595a ) or ( a2596a );
 a9079a <=( a2597a ) or ( a9078a );
 a9080a <=( a9079a ) or ( a9074a );
 a9081a <=( a9080a ) or ( a9071a );
 a9084a <=( a2593a ) or ( a2594a );
 a9087a <=( a2591a ) or ( a2592a );
 a9088a <=( a9087a ) or ( a9084a );
 a9091a <=( a2589a ) or ( a2590a );
 a9095a <=( a2586a ) or ( a2587a );
 a9096a <=( a2588a ) or ( a9095a );
 a9097a <=( a9096a ) or ( a9091a );
 a9098a <=( a9097a ) or ( a9088a );
 a9099a <=( a9098a ) or ( a9081a );
 a9102a <=( a2584a ) or ( a2585a );
 a9105a <=( a2582a ) or ( a2583a );
 a9106a <=( a9105a ) or ( a9102a );
 a9109a <=( a2580a ) or ( a2581a );
 a9113a <=( a2577a ) or ( a2578a );
 a9114a <=( a2579a ) or ( a9113a );
 a9115a <=( a9114a ) or ( a9109a );
 a9116a <=( a9115a ) or ( a9106a );
 a9119a <=( a2575a ) or ( a2576a );
 a9123a <=( a2572a ) or ( a2573a );
 a9124a <=( a2574a ) or ( a9123a );
 a9125a <=( a9124a ) or ( a9119a );
 a9128a <=( a2570a ) or ( a2571a );
 a9132a <=( a2567a ) or ( a2568a );
 a9133a <=( a2569a ) or ( a9132a );
 a9134a <=( a9133a ) or ( a9128a );
 a9135a <=( a9134a ) or ( a9125a );
 a9136a <=( a9135a ) or ( a9116a );
 a9137a <=( a9136a ) or ( a9099a );
 a9140a <=( a2565a ) or ( a2566a );
 a9143a <=( a2563a ) or ( a2564a );
 a9144a <=( a9143a ) or ( a9140a );
 a9147a <=( a2561a ) or ( a2562a );
 a9151a <=( a2558a ) or ( a2559a );
 a9152a <=( a2560a ) or ( a9151a );
 a9153a <=( a9152a ) or ( a9147a );
 a9154a <=( a9153a ) or ( a9144a );
 a9157a <=( a2556a ) or ( a2557a );
 a9161a <=( a2553a ) or ( a2554a );
 a9162a <=( a2555a ) or ( a9161a );
 a9163a <=( a9162a ) or ( a9157a );
 a9166a <=( a2551a ) or ( a2552a );
 a9170a <=( a2548a ) or ( a2549a );
 a9171a <=( a2550a ) or ( a9170a );
 a9172a <=( a9171a ) or ( a9166a );
 a9173a <=( a9172a ) or ( a9163a );
 a9174a <=( a9173a ) or ( a9154a );
 a9177a <=( a2546a ) or ( a2547a );
 a9180a <=( a2544a ) or ( a2545a );
 a9181a <=( a9180a ) or ( a9177a );
 a9184a <=( a2542a ) or ( a2543a );
 a9188a <=( a2539a ) or ( a2540a );
 a9189a <=( a2541a ) or ( a9188a );
 a9190a <=( a9189a ) or ( a9184a );
 a9191a <=( a9190a ) or ( a9181a );
 a9194a <=( a2537a ) or ( a2538a );
 a9198a <=( a2534a ) or ( a2535a );
 a9199a <=( a2536a ) or ( a9198a );
 a9200a <=( a9199a ) or ( a9194a );
 a9203a <=( a2532a ) or ( a2533a );
 a9207a <=( a2529a ) or ( a2530a );
 a9208a <=( a2531a ) or ( a9207a );
 a9209a <=( a9208a ) or ( a9203a );
 a9210a <=( a9209a ) or ( a9200a );
 a9211a <=( a9210a ) or ( a9191a );
 a9212a <=( a9211a ) or ( a9174a );
 a9213a <=( a9212a ) or ( a9137a );
 a9214a <=( a9213a ) or ( a9064a );
 a9217a <=( a2527a ) or ( a2528a );
 a9220a <=( a2525a ) or ( a2526a );
 a9221a <=( a9220a ) or ( a9217a );
 a9224a <=( a2523a ) or ( a2524a );
 a9228a <=( a2520a ) or ( a2521a );
 a9229a <=( a2522a ) or ( a9228a );
 a9230a <=( a9229a ) or ( a9224a );
 a9231a <=( a9230a ) or ( a9221a );
 a9234a <=( a2518a ) or ( a2519a );
 a9237a <=( a2516a ) or ( a2517a );
 a9238a <=( a9237a ) or ( a9234a );
 a9241a <=( a2514a ) or ( a2515a );
 a9245a <=( a2511a ) or ( a2512a );
 a9246a <=( a2513a ) or ( a9245a );
 a9247a <=( a9246a ) or ( a9241a );
 a9248a <=( a9247a ) or ( a9238a );
 a9249a <=( a9248a ) or ( a9231a );
 a9252a <=( a2509a ) or ( a2510a );
 a9255a <=( a2507a ) or ( a2508a );
 a9256a <=( a9255a ) or ( a9252a );
 a9259a <=( a2505a ) or ( a2506a );
 a9263a <=( a2502a ) or ( a2503a );
 a9264a <=( a2504a ) or ( a9263a );
 a9265a <=( a9264a ) or ( a9259a );
 a9266a <=( a9265a ) or ( a9256a );
 a9269a <=( a2500a ) or ( a2501a );
 a9273a <=( a2497a ) or ( a2498a );
 a9274a <=( a2499a ) or ( a9273a );
 a9275a <=( a9274a ) or ( a9269a );
 a9278a <=( a2495a ) or ( a2496a );
 a9282a <=( a2492a ) or ( a2493a );
 a9283a <=( a2494a ) or ( a9282a );
 a9284a <=( a9283a ) or ( a9278a );
 a9285a <=( a9284a ) or ( a9275a );
 a9286a <=( a9285a ) or ( a9266a );
 a9287a <=( a9286a ) or ( a9249a );
 a9290a <=( a2490a ) or ( a2491a );
 a9293a <=( a2488a ) or ( a2489a );
 a9294a <=( a9293a ) or ( a9290a );
 a9297a <=( a2486a ) or ( a2487a );
 a9301a <=( a2483a ) or ( a2484a );
 a9302a <=( a2485a ) or ( a9301a );
 a9303a <=( a9302a ) or ( a9297a );
 a9304a <=( a9303a ) or ( a9294a );
 a9307a <=( a2481a ) or ( a2482a );
 a9310a <=( a2479a ) or ( a2480a );
 a9311a <=( a9310a ) or ( a9307a );
 a9314a <=( a2477a ) or ( a2478a );
 a9318a <=( a2474a ) or ( a2475a );
 a9319a <=( a2476a ) or ( a9318a );
 a9320a <=( a9319a ) or ( a9314a );
 a9321a <=( a9320a ) or ( a9311a );
 a9322a <=( a9321a ) or ( a9304a );
 a9325a <=( a2472a ) or ( a2473a );
 a9328a <=( a2470a ) or ( a2471a );
 a9329a <=( a9328a ) or ( a9325a );
 a9332a <=( a2468a ) or ( a2469a );
 a9336a <=( a2465a ) or ( a2466a );
 a9337a <=( a2467a ) or ( a9336a );
 a9338a <=( a9337a ) or ( a9332a );
 a9339a <=( a9338a ) or ( a9329a );
 a9342a <=( a2463a ) or ( a2464a );
 a9346a <=( a2460a ) or ( a2461a );
 a9347a <=( a2462a ) or ( a9346a );
 a9348a <=( a9347a ) or ( a9342a );
 a9351a <=( a2458a ) or ( a2459a );
 a9355a <=( a2455a ) or ( a2456a );
 a9356a <=( a2457a ) or ( a9355a );
 a9357a <=( a9356a ) or ( a9351a );
 a9358a <=( a9357a ) or ( a9348a );
 a9359a <=( a9358a ) or ( a9339a );
 a9360a <=( a9359a ) or ( a9322a );
 a9361a <=( a9360a ) or ( a9287a );
 a9364a <=( a2453a ) or ( a2454a );
 a9367a <=( a2451a ) or ( a2452a );
 a9368a <=( a9367a ) or ( a9364a );
 a9371a <=( a2449a ) or ( a2450a );
 a9375a <=( a2446a ) or ( a2447a );
 a9376a <=( a2448a ) or ( a9375a );
 a9377a <=( a9376a ) or ( a9371a );
 a9378a <=( a9377a ) or ( a9368a );
 a9381a <=( a2444a ) or ( a2445a );
 a9384a <=( a2442a ) or ( a2443a );
 a9385a <=( a9384a ) or ( a9381a );
 a9388a <=( a2440a ) or ( a2441a );
 a9392a <=( a2437a ) or ( a2438a );
 a9393a <=( a2439a ) or ( a9392a );
 a9394a <=( a9393a ) or ( a9388a );
 a9395a <=( a9394a ) or ( a9385a );
 a9396a <=( a9395a ) or ( a9378a );
 a9399a <=( a2435a ) or ( a2436a );
 a9402a <=( a2433a ) or ( a2434a );
 a9403a <=( a9402a ) or ( a9399a );
 a9406a <=( a2431a ) or ( a2432a );
 a9410a <=( a2428a ) or ( a2429a );
 a9411a <=( a2430a ) or ( a9410a );
 a9412a <=( a9411a ) or ( a9406a );
 a9413a <=( a9412a ) or ( a9403a );
 a9416a <=( a2426a ) or ( a2427a );
 a9420a <=( a2423a ) or ( a2424a );
 a9421a <=( a2425a ) or ( a9420a );
 a9422a <=( a9421a ) or ( a9416a );
 a9425a <=( a2421a ) or ( a2422a );
 a9429a <=( a2418a ) or ( a2419a );
 a9430a <=( a2420a ) or ( a9429a );
 a9431a <=( a9430a ) or ( a9425a );
 a9432a <=( a9431a ) or ( a9422a );
 a9433a <=( a9432a ) or ( a9413a );
 a9434a <=( a9433a ) or ( a9396a );
 a9437a <=( a2416a ) or ( a2417a );
 a9440a <=( a2414a ) or ( a2415a );
 a9441a <=( a9440a ) or ( a9437a );
 a9444a <=( a2412a ) or ( a2413a );
 a9448a <=( a2409a ) or ( a2410a );
 a9449a <=( a2411a ) or ( a9448a );
 a9450a <=( a9449a ) or ( a9444a );
 a9451a <=( a9450a ) or ( a9441a );
 a9454a <=( a2407a ) or ( a2408a );
 a9458a <=( a2404a ) or ( a2405a );
 a9459a <=( a2406a ) or ( a9458a );
 a9460a <=( a9459a ) or ( a9454a );
 a9463a <=( a2402a ) or ( a2403a );
 a9467a <=( a2399a ) or ( a2400a );
 a9468a <=( a2401a ) or ( a9467a );
 a9469a <=( a9468a ) or ( a9463a );
 a9470a <=( a9469a ) or ( a9460a );
 a9471a <=( a9470a ) or ( a9451a );
 a9474a <=( a2397a ) or ( a2398a );
 a9477a <=( a2395a ) or ( a2396a );
 a9478a <=( a9477a ) or ( a9474a );
 a9481a <=( a2393a ) or ( a2394a );
 a9485a <=( a2390a ) or ( a2391a );
 a9486a <=( a2392a ) or ( a9485a );
 a9487a <=( a9486a ) or ( a9481a );
 a9488a <=( a9487a ) or ( a9478a );
 a9491a <=( a2388a ) or ( a2389a );
 a9495a <=( a2385a ) or ( a2386a );
 a9496a <=( a2387a ) or ( a9495a );
 a9497a <=( a9496a ) or ( a9491a );
 a9500a <=( a2383a ) or ( a2384a );
 a9504a <=( a2380a ) or ( a2381a );
 a9505a <=( a2382a ) or ( a9504a );
 a9506a <=( a9505a ) or ( a9500a );
 a9507a <=( a9506a ) or ( a9497a );
 a9508a <=( a9507a ) or ( a9488a );
 a9509a <=( a9508a ) or ( a9471a );
 a9510a <=( a9509a ) or ( a9434a );
 a9511a <=( a9510a ) or ( a9361a );
 a9512a <=( a9511a ) or ( a9214a );
 a9513a <=( a9512a ) or ( a8917a );
 a9514a <=( a9513a ) or ( a8324a );
 a9515a <=( a9514a ) or ( a7135a );
 a9518a <=( a2378a ) or ( a2379a );
 a9521a <=( a2376a ) or ( a2377a );
 a9522a <=( a9521a ) or ( a9518a );
 a9525a <=( a2374a ) or ( a2375a );
 a9529a <=( a2371a ) or ( a2372a );
 a9530a <=( a2373a ) or ( a9529a );
 a9531a <=( a9530a ) or ( a9525a );
 a9532a <=( a9531a ) or ( a9522a );
 a9535a <=( a2369a ) or ( a2370a );
 a9538a <=( a2367a ) or ( a2368a );
 a9539a <=( a9538a ) or ( a9535a );
 a9542a <=( a2365a ) or ( a2366a );
 a9546a <=( a2362a ) or ( a2363a );
 a9547a <=( a2364a ) or ( a9546a );
 a9548a <=( a9547a ) or ( a9542a );
 a9549a <=( a9548a ) or ( a9539a );
 a9550a <=( a9549a ) or ( a9532a );
 a9553a <=( a2360a ) or ( a2361a );
 a9556a <=( a2358a ) or ( a2359a );
 a9557a <=( a9556a ) or ( a9553a );
 a9560a <=( a2356a ) or ( a2357a );
 a9564a <=( a2353a ) or ( a2354a );
 a9565a <=( a2355a ) or ( a9564a );
 a9566a <=( a9565a ) or ( a9560a );
 a9567a <=( a9566a ) or ( a9557a );
 a9570a <=( a2351a ) or ( a2352a );
 a9574a <=( a2348a ) or ( a2349a );
 a9575a <=( a2350a ) or ( a9574a );
 a9576a <=( a9575a ) or ( a9570a );
 a9579a <=( a2346a ) or ( a2347a );
 a9583a <=( a2343a ) or ( a2344a );
 a9584a <=( a2345a ) or ( a9583a );
 a9585a <=( a9584a ) or ( a9579a );
 a9586a <=( a9585a ) or ( a9576a );
 a9587a <=( a9586a ) or ( a9567a );
 a9588a <=( a9587a ) or ( a9550a );
 a9591a <=( a2341a ) or ( a2342a );
 a9594a <=( a2339a ) or ( a2340a );
 a9595a <=( a9594a ) or ( a9591a );
 a9598a <=( a2337a ) or ( a2338a );
 a9602a <=( a2334a ) or ( a2335a );
 a9603a <=( a2336a ) or ( a9602a );
 a9604a <=( a9603a ) or ( a9598a );
 a9605a <=( a9604a ) or ( a9595a );
 a9608a <=( a2332a ) or ( a2333a );
 a9611a <=( a2330a ) or ( a2331a );
 a9612a <=( a9611a ) or ( a9608a );
 a9615a <=( a2328a ) or ( a2329a );
 a9619a <=( a2325a ) or ( a2326a );
 a9620a <=( a2327a ) or ( a9619a );
 a9621a <=( a9620a ) or ( a9615a );
 a9622a <=( a9621a ) or ( a9612a );
 a9623a <=( a9622a ) or ( a9605a );
 a9626a <=( a2323a ) or ( a2324a );
 a9629a <=( a2321a ) or ( a2322a );
 a9630a <=( a9629a ) or ( a9626a );
 a9633a <=( a2319a ) or ( a2320a );
 a9637a <=( a2316a ) or ( a2317a );
 a9638a <=( a2318a ) or ( a9637a );
 a9639a <=( a9638a ) or ( a9633a );
 a9640a <=( a9639a ) or ( a9630a );
 a9643a <=( a2314a ) or ( a2315a );
 a9647a <=( a2311a ) or ( a2312a );
 a9648a <=( a2313a ) or ( a9647a );
 a9649a <=( a9648a ) or ( a9643a );
 a9652a <=( a2309a ) or ( a2310a );
 a9656a <=( a2306a ) or ( a2307a );
 a9657a <=( a2308a ) or ( a9656a );
 a9658a <=( a9657a ) or ( a9652a );
 a9659a <=( a9658a ) or ( a9649a );
 a9660a <=( a9659a ) or ( a9640a );
 a9661a <=( a9660a ) or ( a9623a );
 a9662a <=( a9661a ) or ( a9588a );
 a9665a <=( a2304a ) or ( a2305a );
 a9668a <=( a2302a ) or ( a2303a );
 a9669a <=( a9668a ) or ( a9665a );
 a9672a <=( a2300a ) or ( a2301a );
 a9676a <=( a2297a ) or ( a2298a );
 a9677a <=( a2299a ) or ( a9676a );
 a9678a <=( a9677a ) or ( a9672a );
 a9679a <=( a9678a ) or ( a9669a );
 a9682a <=( a2295a ) or ( a2296a );
 a9685a <=( a2293a ) or ( a2294a );
 a9686a <=( a9685a ) or ( a9682a );
 a9689a <=( a2291a ) or ( a2292a );
 a9693a <=( a2288a ) or ( a2289a );
 a9694a <=( a2290a ) or ( a9693a );
 a9695a <=( a9694a ) or ( a9689a );
 a9696a <=( a9695a ) or ( a9686a );
 a9697a <=( a9696a ) or ( a9679a );
 a9700a <=( a2286a ) or ( a2287a );
 a9703a <=( a2284a ) or ( a2285a );
 a9704a <=( a9703a ) or ( a9700a );
 a9707a <=( a2282a ) or ( a2283a );
 a9711a <=( a2279a ) or ( a2280a );
 a9712a <=( a2281a ) or ( a9711a );
 a9713a <=( a9712a ) or ( a9707a );
 a9714a <=( a9713a ) or ( a9704a );
 a9717a <=( a2277a ) or ( a2278a );
 a9721a <=( a2274a ) or ( a2275a );
 a9722a <=( a2276a ) or ( a9721a );
 a9723a <=( a9722a ) or ( a9717a );
 a9726a <=( a2272a ) or ( a2273a );
 a9730a <=( a2269a ) or ( a2270a );
 a9731a <=( a2271a ) or ( a9730a );
 a9732a <=( a9731a ) or ( a9726a );
 a9733a <=( a9732a ) or ( a9723a );
 a9734a <=( a9733a ) or ( a9714a );
 a9735a <=( a9734a ) or ( a9697a );
 a9738a <=( a2267a ) or ( a2268a );
 a9741a <=( a2265a ) or ( a2266a );
 a9742a <=( a9741a ) or ( a9738a );
 a9745a <=( a2263a ) or ( a2264a );
 a9749a <=( a2260a ) or ( a2261a );
 a9750a <=( a2262a ) or ( a9749a );
 a9751a <=( a9750a ) or ( a9745a );
 a9752a <=( a9751a ) or ( a9742a );
 a9755a <=( a2258a ) or ( a2259a );
 a9758a <=( a2256a ) or ( a2257a );
 a9759a <=( a9758a ) or ( a9755a );
 a9762a <=( a2254a ) or ( a2255a );
 a9766a <=( a2251a ) or ( a2252a );
 a9767a <=( a2253a ) or ( a9766a );
 a9768a <=( a9767a ) or ( a9762a );
 a9769a <=( a9768a ) or ( a9759a );
 a9770a <=( a9769a ) or ( a9752a );
 a9773a <=( a2249a ) or ( a2250a );
 a9776a <=( a2247a ) or ( a2248a );
 a9777a <=( a9776a ) or ( a9773a );
 a9780a <=( a2245a ) or ( a2246a );
 a9784a <=( a2242a ) or ( a2243a );
 a9785a <=( a2244a ) or ( a9784a );
 a9786a <=( a9785a ) or ( a9780a );
 a9787a <=( a9786a ) or ( a9777a );
 a9790a <=( a2240a ) or ( a2241a );
 a9794a <=( a2237a ) or ( a2238a );
 a9795a <=( a2239a ) or ( a9794a );
 a9796a <=( a9795a ) or ( a9790a );
 a9799a <=( a2235a ) or ( a2236a );
 a9803a <=( a2232a ) or ( a2233a );
 a9804a <=( a2234a ) or ( a9803a );
 a9805a <=( a9804a ) or ( a9799a );
 a9806a <=( a9805a ) or ( a9796a );
 a9807a <=( a9806a ) or ( a9787a );
 a9808a <=( a9807a ) or ( a9770a );
 a9809a <=( a9808a ) or ( a9735a );
 a9810a <=( a9809a ) or ( a9662a );
 a9813a <=( a2230a ) or ( a2231a );
 a9816a <=( a2228a ) or ( a2229a );
 a9817a <=( a9816a ) or ( a9813a );
 a9820a <=( a2226a ) or ( a2227a );
 a9824a <=( a2223a ) or ( a2224a );
 a9825a <=( a2225a ) or ( a9824a );
 a9826a <=( a9825a ) or ( a9820a );
 a9827a <=( a9826a ) or ( a9817a );
 a9830a <=( a2221a ) or ( a2222a );
 a9833a <=( a2219a ) or ( a2220a );
 a9834a <=( a9833a ) or ( a9830a );
 a9837a <=( a2217a ) or ( a2218a );
 a9841a <=( a2214a ) or ( a2215a );
 a9842a <=( a2216a ) or ( a9841a );
 a9843a <=( a9842a ) or ( a9837a );
 a9844a <=( a9843a ) or ( a9834a );
 a9845a <=( a9844a ) or ( a9827a );
 a9848a <=( a2212a ) or ( a2213a );
 a9851a <=( a2210a ) or ( a2211a );
 a9852a <=( a9851a ) or ( a9848a );
 a9855a <=( a2208a ) or ( a2209a );
 a9859a <=( a2205a ) or ( a2206a );
 a9860a <=( a2207a ) or ( a9859a );
 a9861a <=( a9860a ) or ( a9855a );
 a9862a <=( a9861a ) or ( a9852a );
 a9865a <=( a2203a ) or ( a2204a );
 a9869a <=( a2200a ) or ( a2201a );
 a9870a <=( a2202a ) or ( a9869a );
 a9871a <=( a9870a ) or ( a9865a );
 a9874a <=( a2198a ) or ( a2199a );
 a9878a <=( a2195a ) or ( a2196a );
 a9879a <=( a2197a ) or ( a9878a );
 a9880a <=( a9879a ) or ( a9874a );
 a9881a <=( a9880a ) or ( a9871a );
 a9882a <=( a9881a ) or ( a9862a );
 a9883a <=( a9882a ) or ( a9845a );
 a9886a <=( a2193a ) or ( a2194a );
 a9889a <=( a2191a ) or ( a2192a );
 a9890a <=( a9889a ) or ( a9886a );
 a9893a <=( a2189a ) or ( a2190a );
 a9897a <=( a2186a ) or ( a2187a );
 a9898a <=( a2188a ) or ( a9897a );
 a9899a <=( a9898a ) or ( a9893a );
 a9900a <=( a9899a ) or ( a9890a );
 a9903a <=( a2184a ) or ( a2185a );
 a9906a <=( a2182a ) or ( a2183a );
 a9907a <=( a9906a ) or ( a9903a );
 a9910a <=( a2180a ) or ( a2181a );
 a9914a <=( a2177a ) or ( a2178a );
 a9915a <=( a2179a ) or ( a9914a );
 a9916a <=( a9915a ) or ( a9910a );
 a9917a <=( a9916a ) or ( a9907a );
 a9918a <=( a9917a ) or ( a9900a );
 a9921a <=( a2175a ) or ( a2176a );
 a9924a <=( a2173a ) or ( a2174a );
 a9925a <=( a9924a ) or ( a9921a );
 a9928a <=( a2171a ) or ( a2172a );
 a9932a <=( a2168a ) or ( a2169a );
 a9933a <=( a2170a ) or ( a9932a );
 a9934a <=( a9933a ) or ( a9928a );
 a9935a <=( a9934a ) or ( a9925a );
 a9938a <=( a2166a ) or ( a2167a );
 a9942a <=( a2163a ) or ( a2164a );
 a9943a <=( a2165a ) or ( a9942a );
 a9944a <=( a9943a ) or ( a9938a );
 a9947a <=( a2161a ) or ( a2162a );
 a9951a <=( a2158a ) or ( a2159a );
 a9952a <=( a2160a ) or ( a9951a );
 a9953a <=( a9952a ) or ( a9947a );
 a9954a <=( a9953a ) or ( a9944a );
 a9955a <=( a9954a ) or ( a9935a );
 a9956a <=( a9955a ) or ( a9918a );
 a9957a <=( a9956a ) or ( a9883a );
 a9960a <=( a2156a ) or ( a2157a );
 a9963a <=( a2154a ) or ( a2155a );
 a9964a <=( a9963a ) or ( a9960a );
 a9967a <=( a2152a ) or ( a2153a );
 a9971a <=( a2149a ) or ( a2150a );
 a9972a <=( a2151a ) or ( a9971a );
 a9973a <=( a9972a ) or ( a9967a );
 a9974a <=( a9973a ) or ( a9964a );
 a9977a <=( a2147a ) or ( a2148a );
 a9980a <=( a2145a ) or ( a2146a );
 a9981a <=( a9980a ) or ( a9977a );
 a9984a <=( a2143a ) or ( a2144a );
 a9988a <=( a2140a ) or ( a2141a );
 a9989a <=( a2142a ) or ( a9988a );
 a9990a <=( a9989a ) or ( a9984a );
 a9991a <=( a9990a ) or ( a9981a );
 a9992a <=( a9991a ) or ( a9974a );
 a9995a <=( a2138a ) or ( a2139a );
 a9998a <=( a2136a ) or ( a2137a );
 a9999a <=( a9998a ) or ( a9995a );
 a10002a <=( a2134a ) or ( a2135a );
 a10006a <=( a2131a ) or ( a2132a );
 a10007a <=( a2133a ) or ( a10006a );
 a10008a <=( a10007a ) or ( a10002a );
 a10009a <=( a10008a ) or ( a9999a );
 a10012a <=( a2129a ) or ( a2130a );
 a10016a <=( a2126a ) or ( a2127a );
 a10017a <=( a2128a ) or ( a10016a );
 a10018a <=( a10017a ) or ( a10012a );
 a10021a <=( a2124a ) or ( a2125a );
 a10025a <=( a2121a ) or ( a2122a );
 a10026a <=( a2123a ) or ( a10025a );
 a10027a <=( a10026a ) or ( a10021a );
 a10028a <=( a10027a ) or ( a10018a );
 a10029a <=( a10028a ) or ( a10009a );
 a10030a <=( a10029a ) or ( a9992a );
 a10033a <=( a2119a ) or ( a2120a );
 a10036a <=( a2117a ) or ( a2118a );
 a10037a <=( a10036a ) or ( a10033a );
 a10040a <=( a2115a ) or ( a2116a );
 a10044a <=( a2112a ) or ( a2113a );
 a10045a <=( a2114a ) or ( a10044a );
 a10046a <=( a10045a ) or ( a10040a );
 a10047a <=( a10046a ) or ( a10037a );
 a10050a <=( a2110a ) or ( a2111a );
 a10054a <=( a2107a ) or ( a2108a );
 a10055a <=( a2109a ) or ( a10054a );
 a10056a <=( a10055a ) or ( a10050a );
 a10059a <=( a2105a ) or ( a2106a );
 a10063a <=( a2102a ) or ( a2103a );
 a10064a <=( a2104a ) or ( a10063a );
 a10065a <=( a10064a ) or ( a10059a );
 a10066a <=( a10065a ) or ( a10056a );
 a10067a <=( a10066a ) or ( a10047a );
 a10070a <=( a2100a ) or ( a2101a );
 a10073a <=( a2098a ) or ( a2099a );
 a10074a <=( a10073a ) or ( a10070a );
 a10077a <=( a2096a ) or ( a2097a );
 a10081a <=( a2093a ) or ( a2094a );
 a10082a <=( a2095a ) or ( a10081a );
 a10083a <=( a10082a ) or ( a10077a );
 a10084a <=( a10083a ) or ( a10074a );
 a10087a <=( a2091a ) or ( a2092a );
 a10091a <=( a2088a ) or ( a2089a );
 a10092a <=( a2090a ) or ( a10091a );
 a10093a <=( a10092a ) or ( a10087a );
 a10096a <=( a2086a ) or ( a2087a );
 a10100a <=( a2083a ) or ( a2084a );
 a10101a <=( a2085a ) or ( a10100a );
 a10102a <=( a10101a ) or ( a10096a );
 a10103a <=( a10102a ) or ( a10093a );
 a10104a <=( a10103a ) or ( a10084a );
 a10105a <=( a10104a ) or ( a10067a );
 a10106a <=( a10105a ) or ( a10030a );
 a10107a <=( a10106a ) or ( a9957a );
 a10108a <=( a10107a ) or ( a9810a );
 a10111a <=( a2081a ) or ( a2082a );
 a10114a <=( a2079a ) or ( a2080a );
 a10115a <=( a10114a ) or ( a10111a );
 a10118a <=( a2077a ) or ( a2078a );
 a10122a <=( a2074a ) or ( a2075a );
 a10123a <=( a2076a ) or ( a10122a );
 a10124a <=( a10123a ) or ( a10118a );
 a10125a <=( a10124a ) or ( a10115a );
 a10128a <=( a2072a ) or ( a2073a );
 a10131a <=( a2070a ) or ( a2071a );
 a10132a <=( a10131a ) or ( a10128a );
 a10135a <=( a2068a ) or ( a2069a );
 a10139a <=( a2065a ) or ( a2066a );
 a10140a <=( a2067a ) or ( a10139a );
 a10141a <=( a10140a ) or ( a10135a );
 a10142a <=( a10141a ) or ( a10132a );
 a10143a <=( a10142a ) or ( a10125a );
 a10146a <=( a2063a ) or ( a2064a );
 a10149a <=( a2061a ) or ( a2062a );
 a10150a <=( a10149a ) or ( a10146a );
 a10153a <=( a2059a ) or ( a2060a );
 a10157a <=( a2056a ) or ( a2057a );
 a10158a <=( a2058a ) or ( a10157a );
 a10159a <=( a10158a ) or ( a10153a );
 a10160a <=( a10159a ) or ( a10150a );
 a10163a <=( a2054a ) or ( a2055a );
 a10167a <=( a2051a ) or ( a2052a );
 a10168a <=( a2053a ) or ( a10167a );
 a10169a <=( a10168a ) or ( a10163a );
 a10172a <=( a2049a ) or ( a2050a );
 a10176a <=( a2046a ) or ( a2047a );
 a10177a <=( a2048a ) or ( a10176a );
 a10178a <=( a10177a ) or ( a10172a );
 a10179a <=( a10178a ) or ( a10169a );
 a10180a <=( a10179a ) or ( a10160a );
 a10181a <=( a10180a ) or ( a10143a );
 a10184a <=( a2044a ) or ( a2045a );
 a10187a <=( a2042a ) or ( a2043a );
 a10188a <=( a10187a ) or ( a10184a );
 a10191a <=( a2040a ) or ( a2041a );
 a10195a <=( a2037a ) or ( a2038a );
 a10196a <=( a2039a ) or ( a10195a );
 a10197a <=( a10196a ) or ( a10191a );
 a10198a <=( a10197a ) or ( a10188a );
 a10201a <=( a2035a ) or ( a2036a );
 a10204a <=( a2033a ) or ( a2034a );
 a10205a <=( a10204a ) or ( a10201a );
 a10208a <=( a2031a ) or ( a2032a );
 a10212a <=( a2028a ) or ( a2029a );
 a10213a <=( a2030a ) or ( a10212a );
 a10214a <=( a10213a ) or ( a10208a );
 a10215a <=( a10214a ) or ( a10205a );
 a10216a <=( a10215a ) or ( a10198a );
 a10219a <=( a2026a ) or ( a2027a );
 a10222a <=( a2024a ) or ( a2025a );
 a10223a <=( a10222a ) or ( a10219a );
 a10226a <=( a2022a ) or ( a2023a );
 a10230a <=( a2019a ) or ( a2020a );
 a10231a <=( a2021a ) or ( a10230a );
 a10232a <=( a10231a ) or ( a10226a );
 a10233a <=( a10232a ) or ( a10223a );
 a10236a <=( a2017a ) or ( a2018a );
 a10240a <=( a2014a ) or ( a2015a );
 a10241a <=( a2016a ) or ( a10240a );
 a10242a <=( a10241a ) or ( a10236a );
 a10245a <=( a2012a ) or ( a2013a );
 a10249a <=( a2009a ) or ( a2010a );
 a10250a <=( a2011a ) or ( a10249a );
 a10251a <=( a10250a ) or ( a10245a );
 a10252a <=( a10251a ) or ( a10242a );
 a10253a <=( a10252a ) or ( a10233a );
 a10254a <=( a10253a ) or ( a10216a );
 a10255a <=( a10254a ) or ( a10181a );
 a10258a <=( a2007a ) or ( a2008a );
 a10261a <=( a2005a ) or ( a2006a );
 a10262a <=( a10261a ) or ( a10258a );
 a10265a <=( a2003a ) or ( a2004a );
 a10269a <=( a2000a ) or ( a2001a );
 a10270a <=( a2002a ) or ( a10269a );
 a10271a <=( a10270a ) or ( a10265a );
 a10272a <=( a10271a ) or ( a10262a );
 a10275a <=( a1998a ) or ( a1999a );
 a10278a <=( a1996a ) or ( a1997a );
 a10279a <=( a10278a ) or ( a10275a );
 a10282a <=( a1994a ) or ( a1995a );
 a10286a <=( a1991a ) or ( a1992a );
 a10287a <=( a1993a ) or ( a10286a );
 a10288a <=( a10287a ) or ( a10282a );
 a10289a <=( a10288a ) or ( a10279a );
 a10290a <=( a10289a ) or ( a10272a );
 a10293a <=( a1989a ) or ( a1990a );
 a10296a <=( a1987a ) or ( a1988a );
 a10297a <=( a10296a ) or ( a10293a );
 a10300a <=( a1985a ) or ( a1986a );
 a10304a <=( a1982a ) or ( a1983a );
 a10305a <=( a1984a ) or ( a10304a );
 a10306a <=( a10305a ) or ( a10300a );
 a10307a <=( a10306a ) or ( a10297a );
 a10310a <=( a1980a ) or ( a1981a );
 a10314a <=( a1977a ) or ( a1978a );
 a10315a <=( a1979a ) or ( a10314a );
 a10316a <=( a10315a ) or ( a10310a );
 a10319a <=( a1975a ) or ( a1976a );
 a10323a <=( a1972a ) or ( a1973a );
 a10324a <=( a1974a ) or ( a10323a );
 a10325a <=( a10324a ) or ( a10319a );
 a10326a <=( a10325a ) or ( a10316a );
 a10327a <=( a10326a ) or ( a10307a );
 a10328a <=( a10327a ) or ( a10290a );
 a10331a <=( a1970a ) or ( a1971a );
 a10334a <=( a1968a ) or ( a1969a );
 a10335a <=( a10334a ) or ( a10331a );
 a10338a <=( a1966a ) or ( a1967a );
 a10342a <=( a1963a ) or ( a1964a );
 a10343a <=( a1965a ) or ( a10342a );
 a10344a <=( a10343a ) or ( a10338a );
 a10345a <=( a10344a ) or ( a10335a );
 a10348a <=( a1961a ) or ( a1962a );
 a10351a <=( a1959a ) or ( a1960a );
 a10352a <=( a10351a ) or ( a10348a );
 a10355a <=( a1957a ) or ( a1958a );
 a10359a <=( a1954a ) or ( a1955a );
 a10360a <=( a1956a ) or ( a10359a );
 a10361a <=( a10360a ) or ( a10355a );
 a10362a <=( a10361a ) or ( a10352a );
 a10363a <=( a10362a ) or ( a10345a );
 a10366a <=( a1952a ) or ( a1953a );
 a10369a <=( a1950a ) or ( a1951a );
 a10370a <=( a10369a ) or ( a10366a );
 a10373a <=( a1948a ) or ( a1949a );
 a10377a <=( a1945a ) or ( a1946a );
 a10378a <=( a1947a ) or ( a10377a );
 a10379a <=( a10378a ) or ( a10373a );
 a10380a <=( a10379a ) or ( a10370a );
 a10383a <=( a1943a ) or ( a1944a );
 a10387a <=( a1940a ) or ( a1941a );
 a10388a <=( a1942a ) or ( a10387a );
 a10389a <=( a10388a ) or ( a10383a );
 a10392a <=( a1938a ) or ( a1939a );
 a10396a <=( a1935a ) or ( a1936a );
 a10397a <=( a1937a ) or ( a10396a );
 a10398a <=( a10397a ) or ( a10392a );
 a10399a <=( a10398a ) or ( a10389a );
 a10400a <=( a10399a ) or ( a10380a );
 a10401a <=( a10400a ) or ( a10363a );
 a10402a <=( a10401a ) or ( a10328a );
 a10403a <=( a10402a ) or ( a10255a );
 a10406a <=( a1933a ) or ( a1934a );
 a10409a <=( a1931a ) or ( a1932a );
 a10410a <=( a10409a ) or ( a10406a );
 a10413a <=( a1929a ) or ( a1930a );
 a10417a <=( a1926a ) or ( a1927a );
 a10418a <=( a1928a ) or ( a10417a );
 a10419a <=( a10418a ) or ( a10413a );
 a10420a <=( a10419a ) or ( a10410a );
 a10423a <=( a1924a ) or ( a1925a );
 a10426a <=( a1922a ) or ( a1923a );
 a10427a <=( a10426a ) or ( a10423a );
 a10430a <=( a1920a ) or ( a1921a );
 a10434a <=( a1917a ) or ( a1918a );
 a10435a <=( a1919a ) or ( a10434a );
 a10436a <=( a10435a ) or ( a10430a );
 a10437a <=( a10436a ) or ( a10427a );
 a10438a <=( a10437a ) or ( a10420a );
 a10441a <=( a1915a ) or ( a1916a );
 a10444a <=( a1913a ) or ( a1914a );
 a10445a <=( a10444a ) or ( a10441a );
 a10448a <=( a1911a ) or ( a1912a );
 a10452a <=( a1908a ) or ( a1909a );
 a10453a <=( a1910a ) or ( a10452a );
 a10454a <=( a10453a ) or ( a10448a );
 a10455a <=( a10454a ) or ( a10445a );
 a10458a <=( a1906a ) or ( a1907a );
 a10462a <=( a1903a ) or ( a1904a );
 a10463a <=( a1905a ) or ( a10462a );
 a10464a <=( a10463a ) or ( a10458a );
 a10467a <=( a1901a ) or ( a1902a );
 a10471a <=( a1898a ) or ( a1899a );
 a10472a <=( a1900a ) or ( a10471a );
 a10473a <=( a10472a ) or ( a10467a );
 a10474a <=( a10473a ) or ( a10464a );
 a10475a <=( a10474a ) or ( a10455a );
 a10476a <=( a10475a ) or ( a10438a );
 a10479a <=( a1896a ) or ( a1897a );
 a10482a <=( a1894a ) or ( a1895a );
 a10483a <=( a10482a ) or ( a10479a );
 a10486a <=( a1892a ) or ( a1893a );
 a10490a <=( a1889a ) or ( a1890a );
 a10491a <=( a1891a ) or ( a10490a );
 a10492a <=( a10491a ) or ( a10486a );
 a10493a <=( a10492a ) or ( a10483a );
 a10496a <=( a1887a ) or ( a1888a );
 a10499a <=( a1885a ) or ( a1886a );
 a10500a <=( a10499a ) or ( a10496a );
 a10503a <=( a1883a ) or ( a1884a );
 a10507a <=( a1880a ) or ( a1881a );
 a10508a <=( a1882a ) or ( a10507a );
 a10509a <=( a10508a ) or ( a10503a );
 a10510a <=( a10509a ) or ( a10500a );
 a10511a <=( a10510a ) or ( a10493a );
 a10514a <=( a1878a ) or ( a1879a );
 a10517a <=( a1876a ) or ( a1877a );
 a10518a <=( a10517a ) or ( a10514a );
 a10521a <=( a1874a ) or ( a1875a );
 a10525a <=( a1871a ) or ( a1872a );
 a10526a <=( a1873a ) or ( a10525a );
 a10527a <=( a10526a ) or ( a10521a );
 a10528a <=( a10527a ) or ( a10518a );
 a10531a <=( a1869a ) or ( a1870a );
 a10535a <=( a1866a ) or ( a1867a );
 a10536a <=( a1868a ) or ( a10535a );
 a10537a <=( a10536a ) or ( a10531a );
 a10540a <=( a1864a ) or ( a1865a );
 a10544a <=( a1861a ) or ( a1862a );
 a10545a <=( a1863a ) or ( a10544a );
 a10546a <=( a10545a ) or ( a10540a );
 a10547a <=( a10546a ) or ( a10537a );
 a10548a <=( a10547a ) or ( a10528a );
 a10549a <=( a10548a ) or ( a10511a );
 a10550a <=( a10549a ) or ( a10476a );
 a10553a <=( a1859a ) or ( a1860a );
 a10556a <=( a1857a ) or ( a1858a );
 a10557a <=( a10556a ) or ( a10553a );
 a10560a <=( a1855a ) or ( a1856a );
 a10564a <=( a1852a ) or ( a1853a );
 a10565a <=( a1854a ) or ( a10564a );
 a10566a <=( a10565a ) or ( a10560a );
 a10567a <=( a10566a ) or ( a10557a );
 a10570a <=( a1850a ) or ( a1851a );
 a10573a <=( a1848a ) or ( a1849a );
 a10574a <=( a10573a ) or ( a10570a );
 a10577a <=( a1846a ) or ( a1847a );
 a10581a <=( a1843a ) or ( a1844a );
 a10582a <=( a1845a ) or ( a10581a );
 a10583a <=( a10582a ) or ( a10577a );
 a10584a <=( a10583a ) or ( a10574a );
 a10585a <=( a10584a ) or ( a10567a );
 a10588a <=( a1841a ) or ( a1842a );
 a10591a <=( a1839a ) or ( a1840a );
 a10592a <=( a10591a ) or ( a10588a );
 a10595a <=( a1837a ) or ( a1838a );
 a10599a <=( a1834a ) or ( a1835a );
 a10600a <=( a1836a ) or ( a10599a );
 a10601a <=( a10600a ) or ( a10595a );
 a10602a <=( a10601a ) or ( a10592a );
 a10605a <=( a1832a ) or ( a1833a );
 a10609a <=( a1829a ) or ( a1830a );
 a10610a <=( a1831a ) or ( a10609a );
 a10611a <=( a10610a ) or ( a10605a );
 a10614a <=( a1827a ) or ( a1828a );
 a10618a <=( a1824a ) or ( a1825a );
 a10619a <=( a1826a ) or ( a10618a );
 a10620a <=( a10619a ) or ( a10614a );
 a10621a <=( a10620a ) or ( a10611a );
 a10622a <=( a10621a ) or ( a10602a );
 a10623a <=( a10622a ) or ( a10585a );
 a10626a <=( a1822a ) or ( a1823a );
 a10629a <=( a1820a ) or ( a1821a );
 a10630a <=( a10629a ) or ( a10626a );
 a10633a <=( a1818a ) or ( a1819a );
 a10637a <=( a1815a ) or ( a1816a );
 a10638a <=( a1817a ) or ( a10637a );
 a10639a <=( a10638a ) or ( a10633a );
 a10640a <=( a10639a ) or ( a10630a );
 a10643a <=( a1813a ) or ( a1814a );
 a10647a <=( a1810a ) or ( a1811a );
 a10648a <=( a1812a ) or ( a10647a );
 a10649a <=( a10648a ) or ( a10643a );
 a10652a <=( a1808a ) or ( a1809a );
 a10656a <=( a1805a ) or ( a1806a );
 a10657a <=( a1807a ) or ( a10656a );
 a10658a <=( a10657a ) or ( a10652a );
 a10659a <=( a10658a ) or ( a10649a );
 a10660a <=( a10659a ) or ( a10640a );
 a10663a <=( a1803a ) or ( a1804a );
 a10666a <=( a1801a ) or ( a1802a );
 a10667a <=( a10666a ) or ( a10663a );
 a10670a <=( a1799a ) or ( a1800a );
 a10674a <=( a1796a ) or ( a1797a );
 a10675a <=( a1798a ) or ( a10674a );
 a10676a <=( a10675a ) or ( a10670a );
 a10677a <=( a10676a ) or ( a10667a );
 a10680a <=( a1794a ) or ( a1795a );
 a10684a <=( a1791a ) or ( a1792a );
 a10685a <=( a1793a ) or ( a10684a );
 a10686a <=( a10685a ) or ( a10680a );
 a10689a <=( a1789a ) or ( a1790a );
 a10693a <=( a1786a ) or ( a1787a );
 a10694a <=( a1788a ) or ( a10693a );
 a10695a <=( a10694a ) or ( a10689a );
 a10696a <=( a10695a ) or ( a10686a );
 a10697a <=( a10696a ) or ( a10677a );
 a10698a <=( a10697a ) or ( a10660a );
 a10699a <=( a10698a ) or ( a10623a );
 a10700a <=( a10699a ) or ( a10550a );
 a10701a <=( a10700a ) or ( a10403a );
 a10702a <=( a10701a ) or ( a10108a );
 a10705a <=( a1784a ) or ( a1785a );
 a10708a <=( a1782a ) or ( a1783a );
 a10709a <=( a10708a ) or ( a10705a );
 a10712a <=( a1780a ) or ( a1781a );
 a10716a <=( a1777a ) or ( a1778a );
 a10717a <=( a1779a ) or ( a10716a );
 a10718a <=( a10717a ) or ( a10712a );
 a10719a <=( a10718a ) or ( a10709a );
 a10722a <=( a1775a ) or ( a1776a );
 a10725a <=( a1773a ) or ( a1774a );
 a10726a <=( a10725a ) or ( a10722a );
 a10729a <=( a1771a ) or ( a1772a );
 a10733a <=( a1768a ) or ( a1769a );
 a10734a <=( a1770a ) or ( a10733a );
 a10735a <=( a10734a ) or ( a10729a );
 a10736a <=( a10735a ) or ( a10726a );
 a10737a <=( a10736a ) or ( a10719a );
 a10740a <=( a1766a ) or ( a1767a );
 a10743a <=( a1764a ) or ( a1765a );
 a10744a <=( a10743a ) or ( a10740a );
 a10747a <=( a1762a ) or ( a1763a );
 a10751a <=( a1759a ) or ( a1760a );
 a10752a <=( a1761a ) or ( a10751a );
 a10753a <=( a10752a ) or ( a10747a );
 a10754a <=( a10753a ) or ( a10744a );
 a10757a <=( a1757a ) or ( a1758a );
 a10761a <=( a1754a ) or ( a1755a );
 a10762a <=( a1756a ) or ( a10761a );
 a10763a <=( a10762a ) or ( a10757a );
 a10766a <=( a1752a ) or ( a1753a );
 a10770a <=( a1749a ) or ( a1750a );
 a10771a <=( a1751a ) or ( a10770a );
 a10772a <=( a10771a ) or ( a10766a );
 a10773a <=( a10772a ) or ( a10763a );
 a10774a <=( a10773a ) or ( a10754a );
 a10775a <=( a10774a ) or ( a10737a );
 a10778a <=( a1747a ) or ( a1748a );
 a10781a <=( a1745a ) or ( a1746a );
 a10782a <=( a10781a ) or ( a10778a );
 a10785a <=( a1743a ) or ( a1744a );
 a10789a <=( a1740a ) or ( a1741a );
 a10790a <=( a1742a ) or ( a10789a );
 a10791a <=( a10790a ) or ( a10785a );
 a10792a <=( a10791a ) or ( a10782a );
 a10795a <=( a1738a ) or ( a1739a );
 a10798a <=( a1736a ) or ( a1737a );
 a10799a <=( a10798a ) or ( a10795a );
 a10802a <=( a1734a ) or ( a1735a );
 a10806a <=( a1731a ) or ( a1732a );
 a10807a <=( a1733a ) or ( a10806a );
 a10808a <=( a10807a ) or ( a10802a );
 a10809a <=( a10808a ) or ( a10799a );
 a10810a <=( a10809a ) or ( a10792a );
 a10813a <=( a1729a ) or ( a1730a );
 a10816a <=( a1727a ) or ( a1728a );
 a10817a <=( a10816a ) or ( a10813a );
 a10820a <=( a1725a ) or ( a1726a );
 a10824a <=( a1722a ) or ( a1723a );
 a10825a <=( a1724a ) or ( a10824a );
 a10826a <=( a10825a ) or ( a10820a );
 a10827a <=( a10826a ) or ( a10817a );
 a10830a <=( a1720a ) or ( a1721a );
 a10834a <=( a1717a ) or ( a1718a );
 a10835a <=( a1719a ) or ( a10834a );
 a10836a <=( a10835a ) or ( a10830a );
 a10839a <=( a1715a ) or ( a1716a );
 a10843a <=( a1712a ) or ( a1713a );
 a10844a <=( a1714a ) or ( a10843a );
 a10845a <=( a10844a ) or ( a10839a );
 a10846a <=( a10845a ) or ( a10836a );
 a10847a <=( a10846a ) or ( a10827a );
 a10848a <=( a10847a ) or ( a10810a );
 a10849a <=( a10848a ) or ( a10775a );
 a10852a <=( a1710a ) or ( a1711a );
 a10855a <=( a1708a ) or ( a1709a );
 a10856a <=( a10855a ) or ( a10852a );
 a10859a <=( a1706a ) or ( a1707a );
 a10863a <=( a1703a ) or ( a1704a );
 a10864a <=( a1705a ) or ( a10863a );
 a10865a <=( a10864a ) or ( a10859a );
 a10866a <=( a10865a ) or ( a10856a );
 a10869a <=( a1701a ) or ( a1702a );
 a10872a <=( a1699a ) or ( a1700a );
 a10873a <=( a10872a ) or ( a10869a );
 a10876a <=( a1697a ) or ( a1698a );
 a10880a <=( a1694a ) or ( a1695a );
 a10881a <=( a1696a ) or ( a10880a );
 a10882a <=( a10881a ) or ( a10876a );
 a10883a <=( a10882a ) or ( a10873a );
 a10884a <=( a10883a ) or ( a10866a );
 a10887a <=( a1692a ) or ( a1693a );
 a10890a <=( a1690a ) or ( a1691a );
 a10891a <=( a10890a ) or ( a10887a );
 a10894a <=( a1688a ) or ( a1689a );
 a10898a <=( a1685a ) or ( a1686a );
 a10899a <=( a1687a ) or ( a10898a );
 a10900a <=( a10899a ) or ( a10894a );
 a10901a <=( a10900a ) or ( a10891a );
 a10904a <=( a1683a ) or ( a1684a );
 a10908a <=( a1680a ) or ( a1681a );
 a10909a <=( a1682a ) or ( a10908a );
 a10910a <=( a10909a ) or ( a10904a );
 a10913a <=( a1678a ) or ( a1679a );
 a10917a <=( a1675a ) or ( a1676a );
 a10918a <=( a1677a ) or ( a10917a );
 a10919a <=( a10918a ) or ( a10913a );
 a10920a <=( a10919a ) or ( a10910a );
 a10921a <=( a10920a ) or ( a10901a );
 a10922a <=( a10921a ) or ( a10884a );
 a10925a <=( a1673a ) or ( a1674a );
 a10928a <=( a1671a ) or ( a1672a );
 a10929a <=( a10928a ) or ( a10925a );
 a10932a <=( a1669a ) or ( a1670a );
 a10936a <=( a1666a ) or ( a1667a );
 a10937a <=( a1668a ) or ( a10936a );
 a10938a <=( a10937a ) or ( a10932a );
 a10939a <=( a10938a ) or ( a10929a );
 a10942a <=( a1664a ) or ( a1665a );
 a10945a <=( a1662a ) or ( a1663a );
 a10946a <=( a10945a ) or ( a10942a );
 a10949a <=( a1660a ) or ( a1661a );
 a10953a <=( a1657a ) or ( a1658a );
 a10954a <=( a1659a ) or ( a10953a );
 a10955a <=( a10954a ) or ( a10949a );
 a10956a <=( a10955a ) or ( a10946a );
 a10957a <=( a10956a ) or ( a10939a );
 a10960a <=( a1655a ) or ( a1656a );
 a10963a <=( a1653a ) or ( a1654a );
 a10964a <=( a10963a ) or ( a10960a );
 a10967a <=( a1651a ) or ( a1652a );
 a10971a <=( a1648a ) or ( a1649a );
 a10972a <=( a1650a ) or ( a10971a );
 a10973a <=( a10972a ) or ( a10967a );
 a10974a <=( a10973a ) or ( a10964a );
 a10977a <=( a1646a ) or ( a1647a );
 a10981a <=( a1643a ) or ( a1644a );
 a10982a <=( a1645a ) or ( a10981a );
 a10983a <=( a10982a ) or ( a10977a );
 a10986a <=( a1641a ) or ( a1642a );
 a10990a <=( a1638a ) or ( a1639a );
 a10991a <=( a1640a ) or ( a10990a );
 a10992a <=( a10991a ) or ( a10986a );
 a10993a <=( a10992a ) or ( a10983a );
 a10994a <=( a10993a ) or ( a10974a );
 a10995a <=( a10994a ) or ( a10957a );
 a10996a <=( a10995a ) or ( a10922a );
 a10997a <=( a10996a ) or ( a10849a );
 a11000a <=( a1636a ) or ( a1637a );
 a11003a <=( a1634a ) or ( a1635a );
 a11004a <=( a11003a ) or ( a11000a );
 a11007a <=( a1632a ) or ( a1633a );
 a11011a <=( a1629a ) or ( a1630a );
 a11012a <=( a1631a ) or ( a11011a );
 a11013a <=( a11012a ) or ( a11007a );
 a11014a <=( a11013a ) or ( a11004a );
 a11017a <=( a1627a ) or ( a1628a );
 a11020a <=( a1625a ) or ( a1626a );
 a11021a <=( a11020a ) or ( a11017a );
 a11024a <=( a1623a ) or ( a1624a );
 a11028a <=( a1620a ) or ( a1621a );
 a11029a <=( a1622a ) or ( a11028a );
 a11030a <=( a11029a ) or ( a11024a );
 a11031a <=( a11030a ) or ( a11021a );
 a11032a <=( a11031a ) or ( a11014a );
 a11035a <=( a1618a ) or ( a1619a );
 a11038a <=( a1616a ) or ( a1617a );
 a11039a <=( a11038a ) or ( a11035a );
 a11042a <=( a1614a ) or ( a1615a );
 a11046a <=( a1611a ) or ( a1612a );
 a11047a <=( a1613a ) or ( a11046a );
 a11048a <=( a11047a ) or ( a11042a );
 a11049a <=( a11048a ) or ( a11039a );
 a11052a <=( a1609a ) or ( a1610a );
 a11056a <=( a1606a ) or ( a1607a );
 a11057a <=( a1608a ) or ( a11056a );
 a11058a <=( a11057a ) or ( a11052a );
 a11061a <=( a1604a ) or ( a1605a );
 a11065a <=( a1601a ) or ( a1602a );
 a11066a <=( a1603a ) or ( a11065a );
 a11067a <=( a11066a ) or ( a11061a );
 a11068a <=( a11067a ) or ( a11058a );
 a11069a <=( a11068a ) or ( a11049a );
 a11070a <=( a11069a ) or ( a11032a );
 a11073a <=( a1599a ) or ( a1600a );
 a11076a <=( a1597a ) or ( a1598a );
 a11077a <=( a11076a ) or ( a11073a );
 a11080a <=( a1595a ) or ( a1596a );
 a11084a <=( a1592a ) or ( a1593a );
 a11085a <=( a1594a ) or ( a11084a );
 a11086a <=( a11085a ) or ( a11080a );
 a11087a <=( a11086a ) or ( a11077a );
 a11090a <=( a1590a ) or ( a1591a );
 a11093a <=( a1588a ) or ( a1589a );
 a11094a <=( a11093a ) or ( a11090a );
 a11097a <=( a1586a ) or ( a1587a );
 a11101a <=( a1583a ) or ( a1584a );
 a11102a <=( a1585a ) or ( a11101a );
 a11103a <=( a11102a ) or ( a11097a );
 a11104a <=( a11103a ) or ( a11094a );
 a11105a <=( a11104a ) or ( a11087a );
 a11108a <=( a1581a ) or ( a1582a );
 a11111a <=( a1579a ) or ( a1580a );
 a11112a <=( a11111a ) or ( a11108a );
 a11115a <=( a1577a ) or ( a1578a );
 a11119a <=( a1574a ) or ( a1575a );
 a11120a <=( a1576a ) or ( a11119a );
 a11121a <=( a11120a ) or ( a11115a );
 a11122a <=( a11121a ) or ( a11112a );
 a11125a <=( a1572a ) or ( a1573a );
 a11129a <=( a1569a ) or ( a1570a );
 a11130a <=( a1571a ) or ( a11129a );
 a11131a <=( a11130a ) or ( a11125a );
 a11134a <=( a1567a ) or ( a1568a );
 a11138a <=( a1564a ) or ( a1565a );
 a11139a <=( a1566a ) or ( a11138a );
 a11140a <=( a11139a ) or ( a11134a );
 a11141a <=( a11140a ) or ( a11131a );
 a11142a <=( a11141a ) or ( a11122a );
 a11143a <=( a11142a ) or ( a11105a );
 a11144a <=( a11143a ) or ( a11070a );
 a11147a <=( a1562a ) or ( a1563a );
 a11150a <=( a1560a ) or ( a1561a );
 a11151a <=( a11150a ) or ( a11147a );
 a11154a <=( a1558a ) or ( a1559a );
 a11158a <=( a1555a ) or ( a1556a );
 a11159a <=( a1557a ) or ( a11158a );
 a11160a <=( a11159a ) or ( a11154a );
 a11161a <=( a11160a ) or ( a11151a );
 a11164a <=( a1553a ) or ( a1554a );
 a11167a <=( a1551a ) or ( a1552a );
 a11168a <=( a11167a ) or ( a11164a );
 a11171a <=( a1549a ) or ( a1550a );
 a11175a <=( a1546a ) or ( a1547a );
 a11176a <=( a1548a ) or ( a11175a );
 a11177a <=( a11176a ) or ( a11171a );
 a11178a <=( a11177a ) or ( a11168a );
 a11179a <=( a11178a ) or ( a11161a );
 a11182a <=( a1544a ) or ( a1545a );
 a11185a <=( a1542a ) or ( a1543a );
 a11186a <=( a11185a ) or ( a11182a );
 a11189a <=( a1540a ) or ( a1541a );
 a11193a <=( a1537a ) or ( a1538a );
 a11194a <=( a1539a ) or ( a11193a );
 a11195a <=( a11194a ) or ( a11189a );
 a11196a <=( a11195a ) or ( a11186a );
 a11199a <=( a1535a ) or ( a1536a );
 a11203a <=( a1532a ) or ( a1533a );
 a11204a <=( a1534a ) or ( a11203a );
 a11205a <=( a11204a ) or ( a11199a );
 a11208a <=( a1530a ) or ( a1531a );
 a11212a <=( a1527a ) or ( a1528a );
 a11213a <=( a1529a ) or ( a11212a );
 a11214a <=( a11213a ) or ( a11208a );
 a11215a <=( a11214a ) or ( a11205a );
 a11216a <=( a11215a ) or ( a11196a );
 a11217a <=( a11216a ) or ( a11179a );
 a11220a <=( a1525a ) or ( a1526a );
 a11223a <=( a1523a ) or ( a1524a );
 a11224a <=( a11223a ) or ( a11220a );
 a11227a <=( a1521a ) or ( a1522a );
 a11231a <=( a1518a ) or ( a1519a );
 a11232a <=( a1520a ) or ( a11231a );
 a11233a <=( a11232a ) or ( a11227a );
 a11234a <=( a11233a ) or ( a11224a );
 a11237a <=( a1516a ) or ( a1517a );
 a11241a <=( a1513a ) or ( a1514a );
 a11242a <=( a1515a ) or ( a11241a );
 a11243a <=( a11242a ) or ( a11237a );
 a11246a <=( a1511a ) or ( a1512a );
 a11250a <=( a1508a ) or ( a1509a );
 a11251a <=( a1510a ) or ( a11250a );
 a11252a <=( a11251a ) or ( a11246a );
 a11253a <=( a11252a ) or ( a11243a );
 a11254a <=( a11253a ) or ( a11234a );
 a11257a <=( a1506a ) or ( a1507a );
 a11260a <=( a1504a ) or ( a1505a );
 a11261a <=( a11260a ) or ( a11257a );
 a11264a <=( a1502a ) or ( a1503a );
 a11268a <=( a1499a ) or ( a1500a );
 a11269a <=( a1501a ) or ( a11268a );
 a11270a <=( a11269a ) or ( a11264a );
 a11271a <=( a11270a ) or ( a11261a );
 a11274a <=( a1497a ) or ( a1498a );
 a11278a <=( a1494a ) or ( a1495a );
 a11279a <=( a1496a ) or ( a11278a );
 a11280a <=( a11279a ) or ( a11274a );
 a11283a <=( a1492a ) or ( a1493a );
 a11287a <=( a1489a ) or ( a1490a );
 a11288a <=( a1491a ) or ( a11287a );
 a11289a <=( a11288a ) or ( a11283a );
 a11290a <=( a11289a ) or ( a11280a );
 a11291a <=( a11290a ) or ( a11271a );
 a11292a <=( a11291a ) or ( a11254a );
 a11293a <=( a11292a ) or ( a11217a );
 a11294a <=( a11293a ) or ( a11144a );
 a11295a <=( a11294a ) or ( a10997a );
 a11298a <=( a1487a ) or ( a1488a );
 a11301a <=( a1485a ) or ( a1486a );
 a11302a <=( a11301a ) or ( a11298a );
 a11305a <=( a1483a ) or ( a1484a );
 a11309a <=( a1480a ) or ( a1481a );
 a11310a <=( a1482a ) or ( a11309a );
 a11311a <=( a11310a ) or ( a11305a );
 a11312a <=( a11311a ) or ( a11302a );
 a11315a <=( a1478a ) or ( a1479a );
 a11318a <=( a1476a ) or ( a1477a );
 a11319a <=( a11318a ) or ( a11315a );
 a11322a <=( a1474a ) or ( a1475a );
 a11326a <=( a1471a ) or ( a1472a );
 a11327a <=( a1473a ) or ( a11326a );
 a11328a <=( a11327a ) or ( a11322a );
 a11329a <=( a11328a ) or ( a11319a );
 a11330a <=( a11329a ) or ( a11312a );
 a11333a <=( a1469a ) or ( a1470a );
 a11336a <=( a1467a ) or ( a1468a );
 a11337a <=( a11336a ) or ( a11333a );
 a11340a <=( a1465a ) or ( a1466a );
 a11344a <=( a1462a ) or ( a1463a );
 a11345a <=( a1464a ) or ( a11344a );
 a11346a <=( a11345a ) or ( a11340a );
 a11347a <=( a11346a ) or ( a11337a );
 a11350a <=( a1460a ) or ( a1461a );
 a11354a <=( a1457a ) or ( a1458a );
 a11355a <=( a1459a ) or ( a11354a );
 a11356a <=( a11355a ) or ( a11350a );
 a11359a <=( a1455a ) or ( a1456a );
 a11363a <=( a1452a ) or ( a1453a );
 a11364a <=( a1454a ) or ( a11363a );
 a11365a <=( a11364a ) or ( a11359a );
 a11366a <=( a11365a ) or ( a11356a );
 a11367a <=( a11366a ) or ( a11347a );
 a11368a <=( a11367a ) or ( a11330a );
 a11371a <=( a1450a ) or ( a1451a );
 a11374a <=( a1448a ) or ( a1449a );
 a11375a <=( a11374a ) or ( a11371a );
 a11378a <=( a1446a ) or ( a1447a );
 a11382a <=( a1443a ) or ( a1444a );
 a11383a <=( a1445a ) or ( a11382a );
 a11384a <=( a11383a ) or ( a11378a );
 a11385a <=( a11384a ) or ( a11375a );
 a11388a <=( a1441a ) or ( a1442a );
 a11391a <=( a1439a ) or ( a1440a );
 a11392a <=( a11391a ) or ( a11388a );
 a11395a <=( a1437a ) or ( a1438a );
 a11399a <=( a1434a ) or ( a1435a );
 a11400a <=( a1436a ) or ( a11399a );
 a11401a <=( a11400a ) or ( a11395a );
 a11402a <=( a11401a ) or ( a11392a );
 a11403a <=( a11402a ) or ( a11385a );
 a11406a <=( a1432a ) or ( a1433a );
 a11409a <=( a1430a ) or ( a1431a );
 a11410a <=( a11409a ) or ( a11406a );
 a11413a <=( a1428a ) or ( a1429a );
 a11417a <=( a1425a ) or ( a1426a );
 a11418a <=( a1427a ) or ( a11417a );
 a11419a <=( a11418a ) or ( a11413a );
 a11420a <=( a11419a ) or ( a11410a );
 a11423a <=( a1423a ) or ( a1424a );
 a11427a <=( a1420a ) or ( a1421a );
 a11428a <=( a1422a ) or ( a11427a );
 a11429a <=( a11428a ) or ( a11423a );
 a11432a <=( a1418a ) or ( a1419a );
 a11436a <=( a1415a ) or ( a1416a );
 a11437a <=( a1417a ) or ( a11436a );
 a11438a <=( a11437a ) or ( a11432a );
 a11439a <=( a11438a ) or ( a11429a );
 a11440a <=( a11439a ) or ( a11420a );
 a11441a <=( a11440a ) or ( a11403a );
 a11442a <=( a11441a ) or ( a11368a );
 a11445a <=( a1413a ) or ( a1414a );
 a11448a <=( a1411a ) or ( a1412a );
 a11449a <=( a11448a ) or ( a11445a );
 a11452a <=( a1409a ) or ( a1410a );
 a11456a <=( a1406a ) or ( a1407a );
 a11457a <=( a1408a ) or ( a11456a );
 a11458a <=( a11457a ) or ( a11452a );
 a11459a <=( a11458a ) or ( a11449a );
 a11462a <=( a1404a ) or ( a1405a );
 a11465a <=( a1402a ) or ( a1403a );
 a11466a <=( a11465a ) or ( a11462a );
 a11469a <=( a1400a ) or ( a1401a );
 a11473a <=( a1397a ) or ( a1398a );
 a11474a <=( a1399a ) or ( a11473a );
 a11475a <=( a11474a ) or ( a11469a );
 a11476a <=( a11475a ) or ( a11466a );
 a11477a <=( a11476a ) or ( a11459a );
 a11480a <=( a1395a ) or ( a1396a );
 a11483a <=( a1393a ) or ( a1394a );
 a11484a <=( a11483a ) or ( a11480a );
 a11487a <=( a1391a ) or ( a1392a );
 a11491a <=( a1388a ) or ( a1389a );
 a11492a <=( a1390a ) or ( a11491a );
 a11493a <=( a11492a ) or ( a11487a );
 a11494a <=( a11493a ) or ( a11484a );
 a11497a <=( a1386a ) or ( a1387a );
 a11501a <=( a1383a ) or ( a1384a );
 a11502a <=( a1385a ) or ( a11501a );
 a11503a <=( a11502a ) or ( a11497a );
 a11506a <=( a1381a ) or ( a1382a );
 a11510a <=( a1378a ) or ( a1379a );
 a11511a <=( a1380a ) or ( a11510a );
 a11512a <=( a11511a ) or ( a11506a );
 a11513a <=( a11512a ) or ( a11503a );
 a11514a <=( a11513a ) or ( a11494a );
 a11515a <=( a11514a ) or ( a11477a );
 a11518a <=( a1376a ) or ( a1377a );
 a11521a <=( a1374a ) or ( a1375a );
 a11522a <=( a11521a ) or ( a11518a );
 a11525a <=( a1372a ) or ( a1373a );
 a11529a <=( a1369a ) or ( a1370a );
 a11530a <=( a1371a ) or ( a11529a );
 a11531a <=( a11530a ) or ( a11525a );
 a11532a <=( a11531a ) or ( a11522a );
 a11535a <=( a1367a ) or ( a1368a );
 a11539a <=( a1364a ) or ( a1365a );
 a11540a <=( a1366a ) or ( a11539a );
 a11541a <=( a11540a ) or ( a11535a );
 a11544a <=( a1362a ) or ( a1363a );
 a11548a <=( a1359a ) or ( a1360a );
 a11549a <=( a1361a ) or ( a11548a );
 a11550a <=( a11549a ) or ( a11544a );
 a11551a <=( a11550a ) or ( a11541a );
 a11552a <=( a11551a ) or ( a11532a );
 a11555a <=( a1357a ) or ( a1358a );
 a11558a <=( a1355a ) or ( a1356a );
 a11559a <=( a11558a ) or ( a11555a );
 a11562a <=( a1353a ) or ( a1354a );
 a11566a <=( a1350a ) or ( a1351a );
 a11567a <=( a1352a ) or ( a11566a );
 a11568a <=( a11567a ) or ( a11562a );
 a11569a <=( a11568a ) or ( a11559a );
 a11572a <=( a1348a ) or ( a1349a );
 a11576a <=( a1345a ) or ( a1346a );
 a11577a <=( a1347a ) or ( a11576a );
 a11578a <=( a11577a ) or ( a11572a );
 a11581a <=( a1343a ) or ( a1344a );
 a11585a <=( a1340a ) or ( a1341a );
 a11586a <=( a1342a ) or ( a11585a );
 a11587a <=( a11586a ) or ( a11581a );
 a11588a <=( a11587a ) or ( a11578a );
 a11589a <=( a11588a ) or ( a11569a );
 a11590a <=( a11589a ) or ( a11552a );
 a11591a <=( a11590a ) or ( a11515a );
 a11592a <=( a11591a ) or ( a11442a );
 a11595a <=( a1338a ) or ( a1339a );
 a11598a <=( a1336a ) or ( a1337a );
 a11599a <=( a11598a ) or ( a11595a );
 a11602a <=( a1334a ) or ( a1335a );
 a11606a <=( a1331a ) or ( a1332a );
 a11607a <=( a1333a ) or ( a11606a );
 a11608a <=( a11607a ) or ( a11602a );
 a11609a <=( a11608a ) or ( a11599a );
 a11612a <=( a1329a ) or ( a1330a );
 a11615a <=( a1327a ) or ( a1328a );
 a11616a <=( a11615a ) or ( a11612a );
 a11619a <=( a1325a ) or ( a1326a );
 a11623a <=( a1322a ) or ( a1323a );
 a11624a <=( a1324a ) or ( a11623a );
 a11625a <=( a11624a ) or ( a11619a );
 a11626a <=( a11625a ) or ( a11616a );
 a11627a <=( a11626a ) or ( a11609a );
 a11630a <=( a1320a ) or ( a1321a );
 a11633a <=( a1318a ) or ( a1319a );
 a11634a <=( a11633a ) or ( a11630a );
 a11637a <=( a1316a ) or ( a1317a );
 a11641a <=( a1313a ) or ( a1314a );
 a11642a <=( a1315a ) or ( a11641a );
 a11643a <=( a11642a ) or ( a11637a );
 a11644a <=( a11643a ) or ( a11634a );
 a11647a <=( a1311a ) or ( a1312a );
 a11651a <=( a1308a ) or ( a1309a );
 a11652a <=( a1310a ) or ( a11651a );
 a11653a <=( a11652a ) or ( a11647a );
 a11656a <=( a1306a ) or ( a1307a );
 a11660a <=( a1303a ) or ( a1304a );
 a11661a <=( a1305a ) or ( a11660a );
 a11662a <=( a11661a ) or ( a11656a );
 a11663a <=( a11662a ) or ( a11653a );
 a11664a <=( a11663a ) or ( a11644a );
 a11665a <=( a11664a ) or ( a11627a );
 a11668a <=( a1301a ) or ( a1302a );
 a11671a <=( a1299a ) or ( a1300a );
 a11672a <=( a11671a ) or ( a11668a );
 a11675a <=( a1297a ) or ( a1298a );
 a11679a <=( a1294a ) or ( a1295a );
 a11680a <=( a1296a ) or ( a11679a );
 a11681a <=( a11680a ) or ( a11675a );
 a11682a <=( a11681a ) or ( a11672a );
 a11685a <=( a1292a ) or ( a1293a );
 a11688a <=( a1290a ) or ( a1291a );
 a11689a <=( a11688a ) or ( a11685a );
 a11692a <=( a1288a ) or ( a1289a );
 a11696a <=( a1285a ) or ( a1286a );
 a11697a <=( a1287a ) or ( a11696a );
 a11698a <=( a11697a ) or ( a11692a );
 a11699a <=( a11698a ) or ( a11689a );
 a11700a <=( a11699a ) or ( a11682a );
 a11703a <=( a1283a ) or ( a1284a );
 a11706a <=( a1281a ) or ( a1282a );
 a11707a <=( a11706a ) or ( a11703a );
 a11710a <=( a1279a ) or ( a1280a );
 a11714a <=( a1276a ) or ( a1277a );
 a11715a <=( a1278a ) or ( a11714a );
 a11716a <=( a11715a ) or ( a11710a );
 a11717a <=( a11716a ) or ( a11707a );
 a11720a <=( a1274a ) or ( a1275a );
 a11724a <=( a1271a ) or ( a1272a );
 a11725a <=( a1273a ) or ( a11724a );
 a11726a <=( a11725a ) or ( a11720a );
 a11729a <=( a1269a ) or ( a1270a );
 a11733a <=( a1266a ) or ( a1267a );
 a11734a <=( a1268a ) or ( a11733a );
 a11735a <=( a11734a ) or ( a11729a );
 a11736a <=( a11735a ) or ( a11726a );
 a11737a <=( a11736a ) or ( a11717a );
 a11738a <=( a11737a ) or ( a11700a );
 a11739a <=( a11738a ) or ( a11665a );
 a11742a <=( a1264a ) or ( a1265a );
 a11745a <=( a1262a ) or ( a1263a );
 a11746a <=( a11745a ) or ( a11742a );
 a11749a <=( a1260a ) or ( a1261a );
 a11753a <=( a1257a ) or ( a1258a );
 a11754a <=( a1259a ) or ( a11753a );
 a11755a <=( a11754a ) or ( a11749a );
 a11756a <=( a11755a ) or ( a11746a );
 a11759a <=( a1255a ) or ( a1256a );
 a11762a <=( a1253a ) or ( a1254a );
 a11763a <=( a11762a ) or ( a11759a );
 a11766a <=( a1251a ) or ( a1252a );
 a11770a <=( a1248a ) or ( a1249a );
 a11771a <=( a1250a ) or ( a11770a );
 a11772a <=( a11771a ) or ( a11766a );
 a11773a <=( a11772a ) or ( a11763a );
 a11774a <=( a11773a ) or ( a11756a );
 a11777a <=( a1246a ) or ( a1247a );
 a11780a <=( a1244a ) or ( a1245a );
 a11781a <=( a11780a ) or ( a11777a );
 a11784a <=( a1242a ) or ( a1243a );
 a11788a <=( a1239a ) or ( a1240a );
 a11789a <=( a1241a ) or ( a11788a );
 a11790a <=( a11789a ) or ( a11784a );
 a11791a <=( a11790a ) or ( a11781a );
 a11794a <=( a1237a ) or ( a1238a );
 a11798a <=( a1234a ) or ( a1235a );
 a11799a <=( a1236a ) or ( a11798a );
 a11800a <=( a11799a ) or ( a11794a );
 a11803a <=( a1232a ) or ( a1233a );
 a11807a <=( a1229a ) or ( a1230a );
 a11808a <=( a1231a ) or ( a11807a );
 a11809a <=( a11808a ) or ( a11803a );
 a11810a <=( a11809a ) or ( a11800a );
 a11811a <=( a11810a ) or ( a11791a );
 a11812a <=( a11811a ) or ( a11774a );
 a11815a <=( a1227a ) or ( a1228a );
 a11818a <=( a1225a ) or ( a1226a );
 a11819a <=( a11818a ) or ( a11815a );
 a11822a <=( a1223a ) or ( a1224a );
 a11826a <=( a1220a ) or ( a1221a );
 a11827a <=( a1222a ) or ( a11826a );
 a11828a <=( a11827a ) or ( a11822a );
 a11829a <=( a11828a ) or ( a11819a );
 a11832a <=( a1218a ) or ( a1219a );
 a11836a <=( a1215a ) or ( a1216a );
 a11837a <=( a1217a ) or ( a11836a );
 a11838a <=( a11837a ) or ( a11832a );
 a11841a <=( a1213a ) or ( a1214a );
 a11845a <=( a1210a ) or ( a1211a );
 a11846a <=( a1212a ) or ( a11845a );
 a11847a <=( a11846a ) or ( a11841a );
 a11848a <=( a11847a ) or ( a11838a );
 a11849a <=( a11848a ) or ( a11829a );
 a11852a <=( a1208a ) or ( a1209a );
 a11855a <=( a1206a ) or ( a1207a );
 a11856a <=( a11855a ) or ( a11852a );
 a11859a <=( a1204a ) or ( a1205a );
 a11863a <=( a1201a ) or ( a1202a );
 a11864a <=( a1203a ) or ( a11863a );
 a11865a <=( a11864a ) or ( a11859a );
 a11866a <=( a11865a ) or ( a11856a );
 a11869a <=( a1199a ) or ( a1200a );
 a11873a <=( a1196a ) or ( a1197a );
 a11874a <=( a1198a ) or ( a11873a );
 a11875a <=( a11874a ) or ( a11869a );
 a11878a <=( a1194a ) or ( a1195a );
 a11882a <=( a1191a ) or ( a1192a );
 a11883a <=( a1193a ) or ( a11882a );
 a11884a <=( a11883a ) or ( a11878a );
 a11885a <=( a11884a ) or ( a11875a );
 a11886a <=( a11885a ) or ( a11866a );
 a11887a <=( a11886a ) or ( a11849a );
 a11888a <=( a11887a ) or ( a11812a );
 a11889a <=( a11888a ) or ( a11739a );
 a11890a <=( a11889a ) or ( a11592a );
 a11891a <=( a11890a ) or ( a11295a );
 a11892a <=( a11891a ) or ( a10702a );
 a11895a <=( a1189a ) or ( a1190a );
 a11898a <=( a1187a ) or ( a1188a );
 a11899a <=( a11898a ) or ( a11895a );
 a11902a <=( a1185a ) or ( a1186a );
 a11906a <=( a1182a ) or ( a1183a );
 a11907a <=( a1184a ) or ( a11906a );
 a11908a <=( a11907a ) or ( a11902a );
 a11909a <=( a11908a ) or ( a11899a );
 a11912a <=( a1180a ) or ( a1181a );
 a11915a <=( a1178a ) or ( a1179a );
 a11916a <=( a11915a ) or ( a11912a );
 a11919a <=( a1176a ) or ( a1177a );
 a11923a <=( a1173a ) or ( a1174a );
 a11924a <=( a1175a ) or ( a11923a );
 a11925a <=( a11924a ) or ( a11919a );
 a11926a <=( a11925a ) or ( a11916a );
 a11927a <=( a11926a ) or ( a11909a );
 a11930a <=( a1171a ) or ( a1172a );
 a11933a <=( a1169a ) or ( a1170a );
 a11934a <=( a11933a ) or ( a11930a );
 a11937a <=( a1167a ) or ( a1168a );
 a11941a <=( a1164a ) or ( a1165a );
 a11942a <=( a1166a ) or ( a11941a );
 a11943a <=( a11942a ) or ( a11937a );
 a11944a <=( a11943a ) or ( a11934a );
 a11947a <=( a1162a ) or ( a1163a );
 a11951a <=( a1159a ) or ( a1160a );
 a11952a <=( a1161a ) or ( a11951a );
 a11953a <=( a11952a ) or ( a11947a );
 a11956a <=( a1157a ) or ( a1158a );
 a11960a <=( a1154a ) or ( a1155a );
 a11961a <=( a1156a ) or ( a11960a );
 a11962a <=( a11961a ) or ( a11956a );
 a11963a <=( a11962a ) or ( a11953a );
 a11964a <=( a11963a ) or ( a11944a );
 a11965a <=( a11964a ) or ( a11927a );
 a11968a <=( a1152a ) or ( a1153a );
 a11971a <=( a1150a ) or ( a1151a );
 a11972a <=( a11971a ) or ( a11968a );
 a11975a <=( a1148a ) or ( a1149a );
 a11979a <=( a1145a ) or ( a1146a );
 a11980a <=( a1147a ) or ( a11979a );
 a11981a <=( a11980a ) or ( a11975a );
 a11982a <=( a11981a ) or ( a11972a );
 a11985a <=( a1143a ) or ( a1144a );
 a11988a <=( a1141a ) or ( a1142a );
 a11989a <=( a11988a ) or ( a11985a );
 a11992a <=( a1139a ) or ( a1140a );
 a11996a <=( a1136a ) or ( a1137a );
 a11997a <=( a1138a ) or ( a11996a );
 a11998a <=( a11997a ) or ( a11992a );
 a11999a <=( a11998a ) or ( a11989a );
 a12000a <=( a11999a ) or ( a11982a );
 a12003a <=( a1134a ) or ( a1135a );
 a12006a <=( a1132a ) or ( a1133a );
 a12007a <=( a12006a ) or ( a12003a );
 a12010a <=( a1130a ) or ( a1131a );
 a12014a <=( a1127a ) or ( a1128a );
 a12015a <=( a1129a ) or ( a12014a );
 a12016a <=( a12015a ) or ( a12010a );
 a12017a <=( a12016a ) or ( a12007a );
 a12020a <=( a1125a ) or ( a1126a );
 a12024a <=( a1122a ) or ( a1123a );
 a12025a <=( a1124a ) or ( a12024a );
 a12026a <=( a12025a ) or ( a12020a );
 a12029a <=( a1120a ) or ( a1121a );
 a12033a <=( a1117a ) or ( a1118a );
 a12034a <=( a1119a ) or ( a12033a );
 a12035a <=( a12034a ) or ( a12029a );
 a12036a <=( a12035a ) or ( a12026a );
 a12037a <=( a12036a ) or ( a12017a );
 a12038a <=( a12037a ) or ( a12000a );
 a12039a <=( a12038a ) or ( a11965a );
 a12042a <=( a1115a ) or ( a1116a );
 a12045a <=( a1113a ) or ( a1114a );
 a12046a <=( a12045a ) or ( a12042a );
 a12049a <=( a1111a ) or ( a1112a );
 a12053a <=( a1108a ) or ( a1109a );
 a12054a <=( a1110a ) or ( a12053a );
 a12055a <=( a12054a ) or ( a12049a );
 a12056a <=( a12055a ) or ( a12046a );
 a12059a <=( a1106a ) or ( a1107a );
 a12062a <=( a1104a ) or ( a1105a );
 a12063a <=( a12062a ) or ( a12059a );
 a12066a <=( a1102a ) or ( a1103a );
 a12070a <=( a1099a ) or ( a1100a );
 a12071a <=( a1101a ) or ( a12070a );
 a12072a <=( a12071a ) or ( a12066a );
 a12073a <=( a12072a ) or ( a12063a );
 a12074a <=( a12073a ) or ( a12056a );
 a12077a <=( a1097a ) or ( a1098a );
 a12080a <=( a1095a ) or ( a1096a );
 a12081a <=( a12080a ) or ( a12077a );
 a12084a <=( a1093a ) or ( a1094a );
 a12088a <=( a1090a ) or ( a1091a );
 a12089a <=( a1092a ) or ( a12088a );
 a12090a <=( a12089a ) or ( a12084a );
 a12091a <=( a12090a ) or ( a12081a );
 a12094a <=( a1088a ) or ( a1089a );
 a12098a <=( a1085a ) or ( a1086a );
 a12099a <=( a1087a ) or ( a12098a );
 a12100a <=( a12099a ) or ( a12094a );
 a12103a <=( a1083a ) or ( a1084a );
 a12107a <=( a1080a ) or ( a1081a );
 a12108a <=( a1082a ) or ( a12107a );
 a12109a <=( a12108a ) or ( a12103a );
 a12110a <=( a12109a ) or ( a12100a );
 a12111a <=( a12110a ) or ( a12091a );
 a12112a <=( a12111a ) or ( a12074a );
 a12115a <=( a1078a ) or ( a1079a );
 a12118a <=( a1076a ) or ( a1077a );
 a12119a <=( a12118a ) or ( a12115a );
 a12122a <=( a1074a ) or ( a1075a );
 a12126a <=( a1071a ) or ( a1072a );
 a12127a <=( a1073a ) or ( a12126a );
 a12128a <=( a12127a ) or ( a12122a );
 a12129a <=( a12128a ) or ( a12119a );
 a12132a <=( a1069a ) or ( a1070a );
 a12135a <=( a1067a ) or ( a1068a );
 a12136a <=( a12135a ) or ( a12132a );
 a12139a <=( a1065a ) or ( a1066a );
 a12143a <=( a1062a ) or ( a1063a );
 a12144a <=( a1064a ) or ( a12143a );
 a12145a <=( a12144a ) or ( a12139a );
 a12146a <=( a12145a ) or ( a12136a );
 a12147a <=( a12146a ) or ( a12129a );
 a12150a <=( a1060a ) or ( a1061a );
 a12153a <=( a1058a ) or ( a1059a );
 a12154a <=( a12153a ) or ( a12150a );
 a12157a <=( a1056a ) or ( a1057a );
 a12161a <=( a1053a ) or ( a1054a );
 a12162a <=( a1055a ) or ( a12161a );
 a12163a <=( a12162a ) or ( a12157a );
 a12164a <=( a12163a ) or ( a12154a );
 a12167a <=( a1051a ) or ( a1052a );
 a12171a <=( a1048a ) or ( a1049a );
 a12172a <=( a1050a ) or ( a12171a );
 a12173a <=( a12172a ) or ( a12167a );
 a12176a <=( a1046a ) or ( a1047a );
 a12180a <=( a1043a ) or ( a1044a );
 a12181a <=( a1045a ) or ( a12180a );
 a12182a <=( a12181a ) or ( a12176a );
 a12183a <=( a12182a ) or ( a12173a );
 a12184a <=( a12183a ) or ( a12164a );
 a12185a <=( a12184a ) or ( a12147a );
 a12186a <=( a12185a ) or ( a12112a );
 a12187a <=( a12186a ) or ( a12039a );
 a12190a <=( a1041a ) or ( a1042a );
 a12193a <=( a1039a ) or ( a1040a );
 a12194a <=( a12193a ) or ( a12190a );
 a12197a <=( a1037a ) or ( a1038a );
 a12201a <=( a1034a ) or ( a1035a );
 a12202a <=( a1036a ) or ( a12201a );
 a12203a <=( a12202a ) or ( a12197a );
 a12204a <=( a12203a ) or ( a12194a );
 a12207a <=( a1032a ) or ( a1033a );
 a12210a <=( a1030a ) or ( a1031a );
 a12211a <=( a12210a ) or ( a12207a );
 a12214a <=( a1028a ) or ( a1029a );
 a12218a <=( a1025a ) or ( a1026a );
 a12219a <=( a1027a ) or ( a12218a );
 a12220a <=( a12219a ) or ( a12214a );
 a12221a <=( a12220a ) or ( a12211a );
 a12222a <=( a12221a ) or ( a12204a );
 a12225a <=( a1023a ) or ( a1024a );
 a12228a <=( a1021a ) or ( a1022a );
 a12229a <=( a12228a ) or ( a12225a );
 a12232a <=( a1019a ) or ( a1020a );
 a12236a <=( a1016a ) or ( a1017a );
 a12237a <=( a1018a ) or ( a12236a );
 a12238a <=( a12237a ) or ( a12232a );
 a12239a <=( a12238a ) or ( a12229a );
 a12242a <=( a1014a ) or ( a1015a );
 a12246a <=( a1011a ) or ( a1012a );
 a12247a <=( a1013a ) or ( a12246a );
 a12248a <=( a12247a ) or ( a12242a );
 a12251a <=( a1009a ) or ( a1010a );
 a12255a <=( a1006a ) or ( a1007a );
 a12256a <=( a1008a ) or ( a12255a );
 a12257a <=( a12256a ) or ( a12251a );
 a12258a <=( a12257a ) or ( a12248a );
 a12259a <=( a12258a ) or ( a12239a );
 a12260a <=( a12259a ) or ( a12222a );
 a12263a <=( a1004a ) or ( a1005a );
 a12266a <=( a1002a ) or ( a1003a );
 a12267a <=( a12266a ) or ( a12263a );
 a12270a <=( a1000a ) or ( a1001a );
 a12274a <=( a997a ) or ( a998a );
 a12275a <=( a999a ) or ( a12274a );
 a12276a <=( a12275a ) or ( a12270a );
 a12277a <=( a12276a ) or ( a12267a );
 a12280a <=( a995a ) or ( a996a );
 a12283a <=( a993a ) or ( a994a );
 a12284a <=( a12283a ) or ( a12280a );
 a12287a <=( a991a ) or ( a992a );
 a12291a <=( a988a ) or ( a989a );
 a12292a <=( a990a ) or ( a12291a );
 a12293a <=( a12292a ) or ( a12287a );
 a12294a <=( a12293a ) or ( a12284a );
 a12295a <=( a12294a ) or ( a12277a );
 a12298a <=( a986a ) or ( a987a );
 a12301a <=( a984a ) or ( a985a );
 a12302a <=( a12301a ) or ( a12298a );
 a12305a <=( a982a ) or ( a983a );
 a12309a <=( a979a ) or ( a980a );
 a12310a <=( a981a ) or ( a12309a );
 a12311a <=( a12310a ) or ( a12305a );
 a12312a <=( a12311a ) or ( a12302a );
 a12315a <=( a977a ) or ( a978a );
 a12319a <=( a974a ) or ( a975a );
 a12320a <=( a976a ) or ( a12319a );
 a12321a <=( a12320a ) or ( a12315a );
 a12324a <=( a972a ) or ( a973a );
 a12328a <=( a969a ) or ( a970a );
 a12329a <=( a971a ) or ( a12328a );
 a12330a <=( a12329a ) or ( a12324a );
 a12331a <=( a12330a ) or ( a12321a );
 a12332a <=( a12331a ) or ( a12312a );
 a12333a <=( a12332a ) or ( a12295a );
 a12334a <=( a12333a ) or ( a12260a );
 a12337a <=( a967a ) or ( a968a );
 a12340a <=( a965a ) or ( a966a );
 a12341a <=( a12340a ) or ( a12337a );
 a12344a <=( a963a ) or ( a964a );
 a12348a <=( a960a ) or ( a961a );
 a12349a <=( a962a ) or ( a12348a );
 a12350a <=( a12349a ) or ( a12344a );
 a12351a <=( a12350a ) or ( a12341a );
 a12354a <=( a958a ) or ( a959a );
 a12357a <=( a956a ) or ( a957a );
 a12358a <=( a12357a ) or ( a12354a );
 a12361a <=( a954a ) or ( a955a );
 a12365a <=( a951a ) or ( a952a );
 a12366a <=( a953a ) or ( a12365a );
 a12367a <=( a12366a ) or ( a12361a );
 a12368a <=( a12367a ) or ( a12358a );
 a12369a <=( a12368a ) or ( a12351a );
 a12372a <=( a949a ) or ( a950a );
 a12375a <=( a947a ) or ( a948a );
 a12376a <=( a12375a ) or ( a12372a );
 a12379a <=( a945a ) or ( a946a );
 a12383a <=( a942a ) or ( a943a );
 a12384a <=( a944a ) or ( a12383a );
 a12385a <=( a12384a ) or ( a12379a );
 a12386a <=( a12385a ) or ( a12376a );
 a12389a <=( a940a ) or ( a941a );
 a12393a <=( a937a ) or ( a938a );
 a12394a <=( a939a ) or ( a12393a );
 a12395a <=( a12394a ) or ( a12389a );
 a12398a <=( a935a ) or ( a936a );
 a12402a <=( a932a ) or ( a933a );
 a12403a <=( a934a ) or ( a12402a );
 a12404a <=( a12403a ) or ( a12398a );
 a12405a <=( a12404a ) or ( a12395a );
 a12406a <=( a12405a ) or ( a12386a );
 a12407a <=( a12406a ) or ( a12369a );
 a12410a <=( a930a ) or ( a931a );
 a12413a <=( a928a ) or ( a929a );
 a12414a <=( a12413a ) or ( a12410a );
 a12417a <=( a926a ) or ( a927a );
 a12421a <=( a923a ) or ( a924a );
 a12422a <=( a925a ) or ( a12421a );
 a12423a <=( a12422a ) or ( a12417a );
 a12424a <=( a12423a ) or ( a12414a );
 a12427a <=( a921a ) or ( a922a );
 a12431a <=( a918a ) or ( a919a );
 a12432a <=( a920a ) or ( a12431a );
 a12433a <=( a12432a ) or ( a12427a );
 a12436a <=( a916a ) or ( a917a );
 a12440a <=( a913a ) or ( a914a );
 a12441a <=( a915a ) or ( a12440a );
 a12442a <=( a12441a ) or ( a12436a );
 a12443a <=( a12442a ) or ( a12433a );
 a12444a <=( a12443a ) or ( a12424a );
 a12447a <=( a911a ) or ( a912a );
 a12450a <=( a909a ) or ( a910a );
 a12451a <=( a12450a ) or ( a12447a );
 a12454a <=( a907a ) or ( a908a );
 a12458a <=( a904a ) or ( a905a );
 a12459a <=( a906a ) or ( a12458a );
 a12460a <=( a12459a ) or ( a12454a );
 a12461a <=( a12460a ) or ( a12451a );
 a12464a <=( a902a ) or ( a903a );
 a12468a <=( a899a ) or ( a900a );
 a12469a <=( a901a ) or ( a12468a );
 a12470a <=( a12469a ) or ( a12464a );
 a12473a <=( a897a ) or ( a898a );
 a12477a <=( a894a ) or ( a895a );
 a12478a <=( a896a ) or ( a12477a );
 a12479a <=( a12478a ) or ( a12473a );
 a12480a <=( a12479a ) or ( a12470a );
 a12481a <=( a12480a ) or ( a12461a );
 a12482a <=( a12481a ) or ( a12444a );
 a12483a <=( a12482a ) or ( a12407a );
 a12484a <=( a12483a ) or ( a12334a );
 a12485a <=( a12484a ) or ( a12187a );
 a12488a <=( a892a ) or ( a893a );
 a12491a <=( a890a ) or ( a891a );
 a12492a <=( a12491a ) or ( a12488a );
 a12495a <=( a888a ) or ( a889a );
 a12499a <=( a885a ) or ( a886a );
 a12500a <=( a887a ) or ( a12499a );
 a12501a <=( a12500a ) or ( a12495a );
 a12502a <=( a12501a ) or ( a12492a );
 a12505a <=( a883a ) or ( a884a );
 a12508a <=( a881a ) or ( a882a );
 a12509a <=( a12508a ) or ( a12505a );
 a12512a <=( a879a ) or ( a880a );
 a12516a <=( a876a ) or ( a877a );
 a12517a <=( a878a ) or ( a12516a );
 a12518a <=( a12517a ) or ( a12512a );
 a12519a <=( a12518a ) or ( a12509a );
 a12520a <=( a12519a ) or ( a12502a );
 a12523a <=( a874a ) or ( a875a );
 a12526a <=( a872a ) or ( a873a );
 a12527a <=( a12526a ) or ( a12523a );
 a12530a <=( a870a ) or ( a871a );
 a12534a <=( a867a ) or ( a868a );
 a12535a <=( a869a ) or ( a12534a );
 a12536a <=( a12535a ) or ( a12530a );
 a12537a <=( a12536a ) or ( a12527a );
 a12540a <=( a865a ) or ( a866a );
 a12544a <=( a862a ) or ( a863a );
 a12545a <=( a864a ) or ( a12544a );
 a12546a <=( a12545a ) or ( a12540a );
 a12549a <=( a860a ) or ( a861a );
 a12553a <=( a857a ) or ( a858a );
 a12554a <=( a859a ) or ( a12553a );
 a12555a <=( a12554a ) or ( a12549a );
 a12556a <=( a12555a ) or ( a12546a );
 a12557a <=( a12556a ) or ( a12537a );
 a12558a <=( a12557a ) or ( a12520a );
 a12561a <=( a855a ) or ( a856a );
 a12564a <=( a853a ) or ( a854a );
 a12565a <=( a12564a ) or ( a12561a );
 a12568a <=( a851a ) or ( a852a );
 a12572a <=( a848a ) or ( a849a );
 a12573a <=( a850a ) or ( a12572a );
 a12574a <=( a12573a ) or ( a12568a );
 a12575a <=( a12574a ) or ( a12565a );
 a12578a <=( a846a ) or ( a847a );
 a12581a <=( a844a ) or ( a845a );
 a12582a <=( a12581a ) or ( a12578a );
 a12585a <=( a842a ) or ( a843a );
 a12589a <=( a839a ) or ( a840a );
 a12590a <=( a841a ) or ( a12589a );
 a12591a <=( a12590a ) or ( a12585a );
 a12592a <=( a12591a ) or ( a12582a );
 a12593a <=( a12592a ) or ( a12575a );
 a12596a <=( a837a ) or ( a838a );
 a12599a <=( a835a ) or ( a836a );
 a12600a <=( a12599a ) or ( a12596a );
 a12603a <=( a833a ) or ( a834a );
 a12607a <=( a830a ) or ( a831a );
 a12608a <=( a832a ) or ( a12607a );
 a12609a <=( a12608a ) or ( a12603a );
 a12610a <=( a12609a ) or ( a12600a );
 a12613a <=( a828a ) or ( a829a );
 a12617a <=( a825a ) or ( a826a );
 a12618a <=( a827a ) or ( a12617a );
 a12619a <=( a12618a ) or ( a12613a );
 a12622a <=( a823a ) or ( a824a );
 a12626a <=( a820a ) or ( a821a );
 a12627a <=( a822a ) or ( a12626a );
 a12628a <=( a12627a ) or ( a12622a );
 a12629a <=( a12628a ) or ( a12619a );
 a12630a <=( a12629a ) or ( a12610a );
 a12631a <=( a12630a ) or ( a12593a );
 a12632a <=( a12631a ) or ( a12558a );
 a12635a <=( a818a ) or ( a819a );
 a12638a <=( a816a ) or ( a817a );
 a12639a <=( a12638a ) or ( a12635a );
 a12642a <=( a814a ) or ( a815a );
 a12646a <=( a811a ) or ( a812a );
 a12647a <=( a813a ) or ( a12646a );
 a12648a <=( a12647a ) or ( a12642a );
 a12649a <=( a12648a ) or ( a12639a );
 a12652a <=( a809a ) or ( a810a );
 a12655a <=( a807a ) or ( a808a );
 a12656a <=( a12655a ) or ( a12652a );
 a12659a <=( a805a ) or ( a806a );
 a12663a <=( a802a ) or ( a803a );
 a12664a <=( a804a ) or ( a12663a );
 a12665a <=( a12664a ) or ( a12659a );
 a12666a <=( a12665a ) or ( a12656a );
 a12667a <=( a12666a ) or ( a12649a );
 a12670a <=( a800a ) or ( a801a );
 a12673a <=( a798a ) or ( a799a );
 a12674a <=( a12673a ) or ( a12670a );
 a12677a <=( a796a ) or ( a797a );
 a12681a <=( a793a ) or ( a794a );
 a12682a <=( a795a ) or ( a12681a );
 a12683a <=( a12682a ) or ( a12677a );
 a12684a <=( a12683a ) or ( a12674a );
 a12687a <=( a791a ) or ( a792a );
 a12691a <=( a788a ) or ( a789a );
 a12692a <=( a790a ) or ( a12691a );
 a12693a <=( a12692a ) or ( a12687a );
 a12696a <=( a786a ) or ( a787a );
 a12700a <=( a783a ) or ( a784a );
 a12701a <=( a785a ) or ( a12700a );
 a12702a <=( a12701a ) or ( a12696a );
 a12703a <=( a12702a ) or ( a12693a );
 a12704a <=( a12703a ) or ( a12684a );
 a12705a <=( a12704a ) or ( a12667a );
 a12708a <=( a781a ) or ( a782a );
 a12711a <=( a779a ) or ( a780a );
 a12712a <=( a12711a ) or ( a12708a );
 a12715a <=( a777a ) or ( a778a );
 a12719a <=( a774a ) or ( a775a );
 a12720a <=( a776a ) or ( a12719a );
 a12721a <=( a12720a ) or ( a12715a );
 a12722a <=( a12721a ) or ( a12712a );
 a12725a <=( a772a ) or ( a773a );
 a12729a <=( a769a ) or ( a770a );
 a12730a <=( a771a ) or ( a12729a );
 a12731a <=( a12730a ) or ( a12725a );
 a12734a <=( a767a ) or ( a768a );
 a12738a <=( a764a ) or ( a765a );
 a12739a <=( a766a ) or ( a12738a );
 a12740a <=( a12739a ) or ( a12734a );
 a12741a <=( a12740a ) or ( a12731a );
 a12742a <=( a12741a ) or ( a12722a );
 a12745a <=( a762a ) or ( a763a );
 a12748a <=( a760a ) or ( a761a );
 a12749a <=( a12748a ) or ( a12745a );
 a12752a <=( a758a ) or ( a759a );
 a12756a <=( a755a ) or ( a756a );
 a12757a <=( a757a ) or ( a12756a );
 a12758a <=( a12757a ) or ( a12752a );
 a12759a <=( a12758a ) or ( a12749a );
 a12762a <=( a753a ) or ( a754a );
 a12766a <=( a750a ) or ( a751a );
 a12767a <=( a752a ) or ( a12766a );
 a12768a <=( a12767a ) or ( a12762a );
 a12771a <=( a748a ) or ( a749a );
 a12775a <=( a745a ) or ( a746a );
 a12776a <=( a747a ) or ( a12775a );
 a12777a <=( a12776a ) or ( a12771a );
 a12778a <=( a12777a ) or ( a12768a );
 a12779a <=( a12778a ) or ( a12759a );
 a12780a <=( a12779a ) or ( a12742a );
 a12781a <=( a12780a ) or ( a12705a );
 a12782a <=( a12781a ) or ( a12632a );
 a12785a <=( a743a ) or ( a744a );
 a12788a <=( a741a ) or ( a742a );
 a12789a <=( a12788a ) or ( a12785a );
 a12792a <=( a739a ) or ( a740a );
 a12796a <=( a736a ) or ( a737a );
 a12797a <=( a738a ) or ( a12796a );
 a12798a <=( a12797a ) or ( a12792a );
 a12799a <=( a12798a ) or ( a12789a );
 a12802a <=( a734a ) or ( a735a );
 a12805a <=( a732a ) or ( a733a );
 a12806a <=( a12805a ) or ( a12802a );
 a12809a <=( a730a ) or ( a731a );
 a12813a <=( a727a ) or ( a728a );
 a12814a <=( a729a ) or ( a12813a );
 a12815a <=( a12814a ) or ( a12809a );
 a12816a <=( a12815a ) or ( a12806a );
 a12817a <=( a12816a ) or ( a12799a );
 a12820a <=( a725a ) or ( a726a );
 a12823a <=( a723a ) or ( a724a );
 a12824a <=( a12823a ) or ( a12820a );
 a12827a <=( a721a ) or ( a722a );
 a12831a <=( a718a ) or ( a719a );
 a12832a <=( a720a ) or ( a12831a );
 a12833a <=( a12832a ) or ( a12827a );
 a12834a <=( a12833a ) or ( a12824a );
 a12837a <=( a716a ) or ( a717a );
 a12841a <=( a713a ) or ( a714a );
 a12842a <=( a715a ) or ( a12841a );
 a12843a <=( a12842a ) or ( a12837a );
 a12846a <=( a711a ) or ( a712a );
 a12850a <=( a708a ) or ( a709a );
 a12851a <=( a710a ) or ( a12850a );
 a12852a <=( a12851a ) or ( a12846a );
 a12853a <=( a12852a ) or ( a12843a );
 a12854a <=( a12853a ) or ( a12834a );
 a12855a <=( a12854a ) or ( a12817a );
 a12858a <=( a706a ) or ( a707a );
 a12861a <=( a704a ) or ( a705a );
 a12862a <=( a12861a ) or ( a12858a );
 a12865a <=( a702a ) or ( a703a );
 a12869a <=( a699a ) or ( a700a );
 a12870a <=( a701a ) or ( a12869a );
 a12871a <=( a12870a ) or ( a12865a );
 a12872a <=( a12871a ) or ( a12862a );
 a12875a <=( a697a ) or ( a698a );
 a12878a <=( a695a ) or ( a696a );
 a12879a <=( a12878a ) or ( a12875a );
 a12882a <=( a693a ) or ( a694a );
 a12886a <=( a690a ) or ( a691a );
 a12887a <=( a692a ) or ( a12886a );
 a12888a <=( a12887a ) or ( a12882a );
 a12889a <=( a12888a ) or ( a12879a );
 a12890a <=( a12889a ) or ( a12872a );
 a12893a <=( a688a ) or ( a689a );
 a12896a <=( a686a ) or ( a687a );
 a12897a <=( a12896a ) or ( a12893a );
 a12900a <=( a684a ) or ( a685a );
 a12904a <=( a681a ) or ( a682a );
 a12905a <=( a683a ) or ( a12904a );
 a12906a <=( a12905a ) or ( a12900a );
 a12907a <=( a12906a ) or ( a12897a );
 a12910a <=( a679a ) or ( a680a );
 a12914a <=( a676a ) or ( a677a );
 a12915a <=( a678a ) or ( a12914a );
 a12916a <=( a12915a ) or ( a12910a );
 a12919a <=( a674a ) or ( a675a );
 a12923a <=( a671a ) or ( a672a );
 a12924a <=( a673a ) or ( a12923a );
 a12925a <=( a12924a ) or ( a12919a );
 a12926a <=( a12925a ) or ( a12916a );
 a12927a <=( a12926a ) or ( a12907a );
 a12928a <=( a12927a ) or ( a12890a );
 a12929a <=( a12928a ) or ( a12855a );
 a12932a <=( a669a ) or ( a670a );
 a12935a <=( a667a ) or ( a668a );
 a12936a <=( a12935a ) or ( a12932a );
 a12939a <=( a665a ) or ( a666a );
 a12943a <=( a662a ) or ( a663a );
 a12944a <=( a664a ) or ( a12943a );
 a12945a <=( a12944a ) or ( a12939a );
 a12946a <=( a12945a ) or ( a12936a );
 a12949a <=( a660a ) or ( a661a );
 a12952a <=( a658a ) or ( a659a );
 a12953a <=( a12952a ) or ( a12949a );
 a12956a <=( a656a ) or ( a657a );
 a12960a <=( a653a ) or ( a654a );
 a12961a <=( a655a ) or ( a12960a );
 a12962a <=( a12961a ) or ( a12956a );
 a12963a <=( a12962a ) or ( a12953a );
 a12964a <=( a12963a ) or ( a12946a );
 a12967a <=( a651a ) or ( a652a );
 a12970a <=( a649a ) or ( a650a );
 a12971a <=( a12970a ) or ( a12967a );
 a12974a <=( a647a ) or ( a648a );
 a12978a <=( a644a ) or ( a645a );
 a12979a <=( a646a ) or ( a12978a );
 a12980a <=( a12979a ) or ( a12974a );
 a12981a <=( a12980a ) or ( a12971a );
 a12984a <=( a642a ) or ( a643a );
 a12988a <=( a639a ) or ( a640a );
 a12989a <=( a641a ) or ( a12988a );
 a12990a <=( a12989a ) or ( a12984a );
 a12993a <=( a637a ) or ( a638a );
 a12997a <=( a634a ) or ( a635a );
 a12998a <=( a636a ) or ( a12997a );
 a12999a <=( a12998a ) or ( a12993a );
 a13000a <=( a12999a ) or ( a12990a );
 a13001a <=( a13000a ) or ( a12981a );
 a13002a <=( a13001a ) or ( a12964a );
 a13005a <=( a632a ) or ( a633a );
 a13008a <=( a630a ) or ( a631a );
 a13009a <=( a13008a ) or ( a13005a );
 a13012a <=( a628a ) or ( a629a );
 a13016a <=( a625a ) or ( a626a );
 a13017a <=( a627a ) or ( a13016a );
 a13018a <=( a13017a ) or ( a13012a );
 a13019a <=( a13018a ) or ( a13009a );
 a13022a <=( a623a ) or ( a624a );
 a13026a <=( a620a ) or ( a621a );
 a13027a <=( a622a ) or ( a13026a );
 a13028a <=( a13027a ) or ( a13022a );
 a13031a <=( a618a ) or ( a619a );
 a13035a <=( a615a ) or ( a616a );
 a13036a <=( a617a ) or ( a13035a );
 a13037a <=( a13036a ) or ( a13031a );
 a13038a <=( a13037a ) or ( a13028a );
 a13039a <=( a13038a ) or ( a13019a );
 a13042a <=( a613a ) or ( a614a );
 a13045a <=( a611a ) or ( a612a );
 a13046a <=( a13045a ) or ( a13042a );
 a13049a <=( a609a ) or ( a610a );
 a13053a <=( a606a ) or ( a607a );
 a13054a <=( a608a ) or ( a13053a );
 a13055a <=( a13054a ) or ( a13049a );
 a13056a <=( a13055a ) or ( a13046a );
 a13059a <=( a604a ) or ( a605a );
 a13063a <=( a601a ) or ( a602a );
 a13064a <=( a603a ) or ( a13063a );
 a13065a <=( a13064a ) or ( a13059a );
 a13068a <=( a599a ) or ( a600a );
 a13072a <=( a596a ) or ( a597a );
 a13073a <=( a598a ) or ( a13072a );
 a13074a <=( a13073a ) or ( a13068a );
 a13075a <=( a13074a ) or ( a13065a );
 a13076a <=( a13075a ) or ( a13056a );
 a13077a <=( a13076a ) or ( a13039a );
 a13078a <=( a13077a ) or ( a13002a );
 a13079a <=( a13078a ) or ( a12929a );
 a13080a <=( a13079a ) or ( a12782a );
 a13081a <=( a13080a ) or ( a12485a );
 a13084a <=( a594a ) or ( a595a );
 a13087a <=( a592a ) or ( a593a );
 a13088a <=( a13087a ) or ( a13084a );
 a13091a <=( a590a ) or ( a591a );
 a13095a <=( a587a ) or ( a588a );
 a13096a <=( a589a ) or ( a13095a );
 a13097a <=( a13096a ) or ( a13091a );
 a13098a <=( a13097a ) or ( a13088a );
 a13101a <=( a585a ) or ( a586a );
 a13104a <=( a583a ) or ( a584a );
 a13105a <=( a13104a ) or ( a13101a );
 a13108a <=( a581a ) or ( a582a );
 a13112a <=( a578a ) or ( a579a );
 a13113a <=( a580a ) or ( a13112a );
 a13114a <=( a13113a ) or ( a13108a );
 a13115a <=( a13114a ) or ( a13105a );
 a13116a <=( a13115a ) or ( a13098a );
 a13119a <=( a576a ) or ( a577a );
 a13122a <=( a574a ) or ( a575a );
 a13123a <=( a13122a ) or ( a13119a );
 a13126a <=( a572a ) or ( a573a );
 a13130a <=( a569a ) or ( a570a );
 a13131a <=( a571a ) or ( a13130a );
 a13132a <=( a13131a ) or ( a13126a );
 a13133a <=( a13132a ) or ( a13123a );
 a13136a <=( a567a ) or ( a568a );
 a13140a <=( a564a ) or ( a565a );
 a13141a <=( a566a ) or ( a13140a );
 a13142a <=( a13141a ) or ( a13136a );
 a13145a <=( a562a ) or ( a563a );
 a13149a <=( a559a ) or ( a560a );
 a13150a <=( a561a ) or ( a13149a );
 a13151a <=( a13150a ) or ( a13145a );
 a13152a <=( a13151a ) or ( a13142a );
 a13153a <=( a13152a ) or ( a13133a );
 a13154a <=( a13153a ) or ( a13116a );
 a13157a <=( a557a ) or ( a558a );
 a13160a <=( a555a ) or ( a556a );
 a13161a <=( a13160a ) or ( a13157a );
 a13164a <=( a553a ) or ( a554a );
 a13168a <=( a550a ) or ( a551a );
 a13169a <=( a552a ) or ( a13168a );
 a13170a <=( a13169a ) or ( a13164a );
 a13171a <=( a13170a ) or ( a13161a );
 a13174a <=( a548a ) or ( a549a );
 a13177a <=( a546a ) or ( a547a );
 a13178a <=( a13177a ) or ( a13174a );
 a13181a <=( a544a ) or ( a545a );
 a13185a <=( a541a ) or ( a542a );
 a13186a <=( a543a ) or ( a13185a );
 a13187a <=( a13186a ) or ( a13181a );
 a13188a <=( a13187a ) or ( a13178a );
 a13189a <=( a13188a ) or ( a13171a );
 a13192a <=( a539a ) or ( a540a );
 a13195a <=( a537a ) or ( a538a );
 a13196a <=( a13195a ) or ( a13192a );
 a13199a <=( a535a ) or ( a536a );
 a13203a <=( a532a ) or ( a533a );
 a13204a <=( a534a ) or ( a13203a );
 a13205a <=( a13204a ) or ( a13199a );
 a13206a <=( a13205a ) or ( a13196a );
 a13209a <=( a530a ) or ( a531a );
 a13213a <=( a527a ) or ( a528a );
 a13214a <=( a529a ) or ( a13213a );
 a13215a <=( a13214a ) or ( a13209a );
 a13218a <=( a525a ) or ( a526a );
 a13222a <=( a522a ) or ( a523a );
 a13223a <=( a524a ) or ( a13222a );
 a13224a <=( a13223a ) or ( a13218a );
 a13225a <=( a13224a ) or ( a13215a );
 a13226a <=( a13225a ) or ( a13206a );
 a13227a <=( a13226a ) or ( a13189a );
 a13228a <=( a13227a ) or ( a13154a );
 a13231a <=( a520a ) or ( a521a );
 a13234a <=( a518a ) or ( a519a );
 a13235a <=( a13234a ) or ( a13231a );
 a13238a <=( a516a ) or ( a517a );
 a13242a <=( a513a ) or ( a514a );
 a13243a <=( a515a ) or ( a13242a );
 a13244a <=( a13243a ) or ( a13238a );
 a13245a <=( a13244a ) or ( a13235a );
 a13248a <=( a511a ) or ( a512a );
 a13251a <=( a509a ) or ( a510a );
 a13252a <=( a13251a ) or ( a13248a );
 a13255a <=( a507a ) or ( a508a );
 a13259a <=( a504a ) or ( a505a );
 a13260a <=( a506a ) or ( a13259a );
 a13261a <=( a13260a ) or ( a13255a );
 a13262a <=( a13261a ) or ( a13252a );
 a13263a <=( a13262a ) or ( a13245a );
 a13266a <=( a502a ) or ( a503a );
 a13269a <=( a500a ) or ( a501a );
 a13270a <=( a13269a ) or ( a13266a );
 a13273a <=( a498a ) or ( a499a );
 a13277a <=( a495a ) or ( a496a );
 a13278a <=( a497a ) or ( a13277a );
 a13279a <=( a13278a ) or ( a13273a );
 a13280a <=( a13279a ) or ( a13270a );
 a13283a <=( a493a ) or ( a494a );
 a13287a <=( a490a ) or ( a491a );
 a13288a <=( a492a ) or ( a13287a );
 a13289a <=( a13288a ) or ( a13283a );
 a13292a <=( a488a ) or ( a489a );
 a13296a <=( a485a ) or ( a486a );
 a13297a <=( a487a ) or ( a13296a );
 a13298a <=( a13297a ) or ( a13292a );
 a13299a <=( a13298a ) or ( a13289a );
 a13300a <=( a13299a ) or ( a13280a );
 a13301a <=( a13300a ) or ( a13263a );
 a13304a <=( a483a ) or ( a484a );
 a13307a <=( a481a ) or ( a482a );
 a13308a <=( a13307a ) or ( a13304a );
 a13311a <=( a479a ) or ( a480a );
 a13315a <=( a476a ) or ( a477a );
 a13316a <=( a478a ) or ( a13315a );
 a13317a <=( a13316a ) or ( a13311a );
 a13318a <=( a13317a ) or ( a13308a );
 a13321a <=( a474a ) or ( a475a );
 a13324a <=( a472a ) or ( a473a );
 a13325a <=( a13324a ) or ( a13321a );
 a13328a <=( a470a ) or ( a471a );
 a13332a <=( a467a ) or ( a468a );
 a13333a <=( a469a ) or ( a13332a );
 a13334a <=( a13333a ) or ( a13328a );
 a13335a <=( a13334a ) or ( a13325a );
 a13336a <=( a13335a ) or ( a13318a );
 a13339a <=( a465a ) or ( a466a );
 a13342a <=( a463a ) or ( a464a );
 a13343a <=( a13342a ) or ( a13339a );
 a13346a <=( a461a ) or ( a462a );
 a13350a <=( a458a ) or ( a459a );
 a13351a <=( a460a ) or ( a13350a );
 a13352a <=( a13351a ) or ( a13346a );
 a13353a <=( a13352a ) or ( a13343a );
 a13356a <=( a456a ) or ( a457a );
 a13360a <=( a453a ) or ( a454a );
 a13361a <=( a455a ) or ( a13360a );
 a13362a <=( a13361a ) or ( a13356a );
 a13365a <=( a451a ) or ( a452a );
 a13369a <=( a448a ) or ( a449a );
 a13370a <=( a450a ) or ( a13369a );
 a13371a <=( a13370a ) or ( a13365a );
 a13372a <=( a13371a ) or ( a13362a );
 a13373a <=( a13372a ) or ( a13353a );
 a13374a <=( a13373a ) or ( a13336a );
 a13375a <=( a13374a ) or ( a13301a );
 a13376a <=( a13375a ) or ( a13228a );
 a13379a <=( a446a ) or ( a447a );
 a13382a <=( a444a ) or ( a445a );
 a13383a <=( a13382a ) or ( a13379a );
 a13386a <=( a442a ) or ( a443a );
 a13390a <=( a439a ) or ( a440a );
 a13391a <=( a441a ) or ( a13390a );
 a13392a <=( a13391a ) or ( a13386a );
 a13393a <=( a13392a ) or ( a13383a );
 a13396a <=( a437a ) or ( a438a );
 a13399a <=( a435a ) or ( a436a );
 a13400a <=( a13399a ) or ( a13396a );
 a13403a <=( a433a ) or ( a434a );
 a13407a <=( a430a ) or ( a431a );
 a13408a <=( a432a ) or ( a13407a );
 a13409a <=( a13408a ) or ( a13403a );
 a13410a <=( a13409a ) or ( a13400a );
 a13411a <=( a13410a ) or ( a13393a );
 a13414a <=( a428a ) or ( a429a );
 a13417a <=( a426a ) or ( a427a );
 a13418a <=( a13417a ) or ( a13414a );
 a13421a <=( a424a ) or ( a425a );
 a13425a <=( a421a ) or ( a422a );
 a13426a <=( a423a ) or ( a13425a );
 a13427a <=( a13426a ) or ( a13421a );
 a13428a <=( a13427a ) or ( a13418a );
 a13431a <=( a419a ) or ( a420a );
 a13435a <=( a416a ) or ( a417a );
 a13436a <=( a418a ) or ( a13435a );
 a13437a <=( a13436a ) or ( a13431a );
 a13440a <=( a414a ) or ( a415a );
 a13444a <=( a411a ) or ( a412a );
 a13445a <=( a413a ) or ( a13444a );
 a13446a <=( a13445a ) or ( a13440a );
 a13447a <=( a13446a ) or ( a13437a );
 a13448a <=( a13447a ) or ( a13428a );
 a13449a <=( a13448a ) or ( a13411a );
 a13452a <=( a409a ) or ( a410a );
 a13455a <=( a407a ) or ( a408a );
 a13456a <=( a13455a ) or ( a13452a );
 a13459a <=( a405a ) or ( a406a );
 a13463a <=( a402a ) or ( a403a );
 a13464a <=( a404a ) or ( a13463a );
 a13465a <=( a13464a ) or ( a13459a );
 a13466a <=( a13465a ) or ( a13456a );
 a13469a <=( a400a ) or ( a401a );
 a13472a <=( a398a ) or ( a399a );
 a13473a <=( a13472a ) or ( a13469a );
 a13476a <=( a396a ) or ( a397a );
 a13480a <=( a393a ) or ( a394a );
 a13481a <=( a395a ) or ( a13480a );
 a13482a <=( a13481a ) or ( a13476a );
 a13483a <=( a13482a ) or ( a13473a );
 a13484a <=( a13483a ) or ( a13466a );
 a13487a <=( a391a ) or ( a392a );
 a13490a <=( a389a ) or ( a390a );
 a13491a <=( a13490a ) or ( a13487a );
 a13494a <=( a387a ) or ( a388a );
 a13498a <=( a384a ) or ( a385a );
 a13499a <=( a386a ) or ( a13498a );
 a13500a <=( a13499a ) or ( a13494a );
 a13501a <=( a13500a ) or ( a13491a );
 a13504a <=( a382a ) or ( a383a );
 a13508a <=( a379a ) or ( a380a );
 a13509a <=( a381a ) or ( a13508a );
 a13510a <=( a13509a ) or ( a13504a );
 a13513a <=( a377a ) or ( a378a );
 a13517a <=( a374a ) or ( a375a );
 a13518a <=( a376a ) or ( a13517a );
 a13519a <=( a13518a ) or ( a13513a );
 a13520a <=( a13519a ) or ( a13510a );
 a13521a <=( a13520a ) or ( a13501a );
 a13522a <=( a13521a ) or ( a13484a );
 a13523a <=( a13522a ) or ( a13449a );
 a13526a <=( a372a ) or ( a373a );
 a13529a <=( a370a ) or ( a371a );
 a13530a <=( a13529a ) or ( a13526a );
 a13533a <=( a368a ) or ( a369a );
 a13537a <=( a365a ) or ( a366a );
 a13538a <=( a367a ) or ( a13537a );
 a13539a <=( a13538a ) or ( a13533a );
 a13540a <=( a13539a ) or ( a13530a );
 a13543a <=( a363a ) or ( a364a );
 a13546a <=( a361a ) or ( a362a );
 a13547a <=( a13546a ) or ( a13543a );
 a13550a <=( a359a ) or ( a360a );
 a13554a <=( a356a ) or ( a357a );
 a13555a <=( a358a ) or ( a13554a );
 a13556a <=( a13555a ) or ( a13550a );
 a13557a <=( a13556a ) or ( a13547a );
 a13558a <=( a13557a ) or ( a13540a );
 a13561a <=( a354a ) or ( a355a );
 a13564a <=( a352a ) or ( a353a );
 a13565a <=( a13564a ) or ( a13561a );
 a13568a <=( a350a ) or ( a351a );
 a13572a <=( a347a ) or ( a348a );
 a13573a <=( a349a ) or ( a13572a );
 a13574a <=( a13573a ) or ( a13568a );
 a13575a <=( a13574a ) or ( a13565a );
 a13578a <=( a345a ) or ( a346a );
 a13582a <=( a342a ) or ( a343a );
 a13583a <=( a344a ) or ( a13582a );
 a13584a <=( a13583a ) or ( a13578a );
 a13587a <=( a340a ) or ( a341a );
 a13591a <=( a337a ) or ( a338a );
 a13592a <=( a339a ) or ( a13591a );
 a13593a <=( a13592a ) or ( a13587a );
 a13594a <=( a13593a ) or ( a13584a );
 a13595a <=( a13594a ) or ( a13575a );
 a13596a <=( a13595a ) or ( a13558a );
 a13599a <=( a335a ) or ( a336a );
 a13602a <=( a333a ) or ( a334a );
 a13603a <=( a13602a ) or ( a13599a );
 a13606a <=( a331a ) or ( a332a );
 a13610a <=( a328a ) or ( a329a );
 a13611a <=( a330a ) or ( a13610a );
 a13612a <=( a13611a ) or ( a13606a );
 a13613a <=( a13612a ) or ( a13603a );
 a13616a <=( a326a ) or ( a327a );
 a13620a <=( a323a ) or ( a324a );
 a13621a <=( a325a ) or ( a13620a );
 a13622a <=( a13621a ) or ( a13616a );
 a13625a <=( a321a ) or ( a322a );
 a13629a <=( a318a ) or ( a319a );
 a13630a <=( a320a ) or ( a13629a );
 a13631a <=( a13630a ) or ( a13625a );
 a13632a <=( a13631a ) or ( a13622a );
 a13633a <=( a13632a ) or ( a13613a );
 a13636a <=( a316a ) or ( a317a );
 a13639a <=( a314a ) or ( a315a );
 a13640a <=( a13639a ) or ( a13636a );
 a13643a <=( a312a ) or ( a313a );
 a13647a <=( a309a ) or ( a310a );
 a13648a <=( a311a ) or ( a13647a );
 a13649a <=( a13648a ) or ( a13643a );
 a13650a <=( a13649a ) or ( a13640a );
 a13653a <=( a307a ) or ( a308a );
 a13657a <=( a304a ) or ( a305a );
 a13658a <=( a306a ) or ( a13657a );
 a13659a <=( a13658a ) or ( a13653a );
 a13662a <=( a302a ) or ( a303a );
 a13666a <=( a299a ) or ( a300a );
 a13667a <=( a301a ) or ( a13666a );
 a13668a <=( a13667a ) or ( a13662a );
 a13669a <=( a13668a ) or ( a13659a );
 a13670a <=( a13669a ) or ( a13650a );
 a13671a <=( a13670a ) or ( a13633a );
 a13672a <=( a13671a ) or ( a13596a );
 a13673a <=( a13672a ) or ( a13523a );
 a13674a <=( a13673a ) or ( a13376a );
 a13677a <=( a297a ) or ( a298a );
 a13680a <=( a295a ) or ( a296a );
 a13681a <=( a13680a ) or ( a13677a );
 a13684a <=( a293a ) or ( a294a );
 a13688a <=( a290a ) or ( a291a );
 a13689a <=( a292a ) or ( a13688a );
 a13690a <=( a13689a ) or ( a13684a );
 a13691a <=( a13690a ) or ( a13681a );
 a13694a <=( a288a ) or ( a289a );
 a13697a <=( a286a ) or ( a287a );
 a13698a <=( a13697a ) or ( a13694a );
 a13701a <=( a284a ) or ( a285a );
 a13705a <=( a281a ) or ( a282a );
 a13706a <=( a283a ) or ( a13705a );
 a13707a <=( a13706a ) or ( a13701a );
 a13708a <=( a13707a ) or ( a13698a );
 a13709a <=( a13708a ) or ( a13691a );
 a13712a <=( a279a ) or ( a280a );
 a13715a <=( a277a ) or ( a278a );
 a13716a <=( a13715a ) or ( a13712a );
 a13719a <=( a275a ) or ( a276a );
 a13723a <=( a272a ) or ( a273a );
 a13724a <=( a274a ) or ( a13723a );
 a13725a <=( a13724a ) or ( a13719a );
 a13726a <=( a13725a ) or ( a13716a );
 a13729a <=( a270a ) or ( a271a );
 a13733a <=( a267a ) or ( a268a );
 a13734a <=( a269a ) or ( a13733a );
 a13735a <=( a13734a ) or ( a13729a );
 a13738a <=( a265a ) or ( a266a );
 a13742a <=( a262a ) or ( a263a );
 a13743a <=( a264a ) or ( a13742a );
 a13744a <=( a13743a ) or ( a13738a );
 a13745a <=( a13744a ) or ( a13735a );
 a13746a <=( a13745a ) or ( a13726a );
 a13747a <=( a13746a ) or ( a13709a );
 a13750a <=( a260a ) or ( a261a );
 a13753a <=( a258a ) or ( a259a );
 a13754a <=( a13753a ) or ( a13750a );
 a13757a <=( a256a ) or ( a257a );
 a13761a <=( a253a ) or ( a254a );
 a13762a <=( a255a ) or ( a13761a );
 a13763a <=( a13762a ) or ( a13757a );
 a13764a <=( a13763a ) or ( a13754a );
 a13767a <=( a251a ) or ( a252a );
 a13770a <=( a249a ) or ( a250a );
 a13771a <=( a13770a ) or ( a13767a );
 a13774a <=( a247a ) or ( a248a );
 a13778a <=( a244a ) or ( a245a );
 a13779a <=( a246a ) or ( a13778a );
 a13780a <=( a13779a ) or ( a13774a );
 a13781a <=( a13780a ) or ( a13771a );
 a13782a <=( a13781a ) or ( a13764a );
 a13785a <=( a242a ) or ( a243a );
 a13788a <=( a240a ) or ( a241a );
 a13789a <=( a13788a ) or ( a13785a );
 a13792a <=( a238a ) or ( a239a );
 a13796a <=( a235a ) or ( a236a );
 a13797a <=( a237a ) or ( a13796a );
 a13798a <=( a13797a ) or ( a13792a );
 a13799a <=( a13798a ) or ( a13789a );
 a13802a <=( a233a ) or ( a234a );
 a13806a <=( a230a ) or ( a231a );
 a13807a <=( a232a ) or ( a13806a );
 a13808a <=( a13807a ) or ( a13802a );
 a13811a <=( a228a ) or ( a229a );
 a13815a <=( a225a ) or ( a226a );
 a13816a <=( a227a ) or ( a13815a );
 a13817a <=( a13816a ) or ( a13811a );
 a13818a <=( a13817a ) or ( a13808a );
 a13819a <=( a13818a ) or ( a13799a );
 a13820a <=( a13819a ) or ( a13782a );
 a13821a <=( a13820a ) or ( a13747a );
 a13824a <=( a223a ) or ( a224a );
 a13827a <=( a221a ) or ( a222a );
 a13828a <=( a13827a ) or ( a13824a );
 a13831a <=( a219a ) or ( a220a );
 a13835a <=( a216a ) or ( a217a );
 a13836a <=( a218a ) or ( a13835a );
 a13837a <=( a13836a ) or ( a13831a );
 a13838a <=( a13837a ) or ( a13828a );
 a13841a <=( a214a ) or ( a215a );
 a13844a <=( a212a ) or ( a213a );
 a13845a <=( a13844a ) or ( a13841a );
 a13848a <=( a210a ) or ( a211a );
 a13852a <=( a207a ) or ( a208a );
 a13853a <=( a209a ) or ( a13852a );
 a13854a <=( a13853a ) or ( a13848a );
 a13855a <=( a13854a ) or ( a13845a );
 a13856a <=( a13855a ) or ( a13838a );
 a13859a <=( a205a ) or ( a206a );
 a13862a <=( a203a ) or ( a204a );
 a13863a <=( a13862a ) or ( a13859a );
 a13866a <=( a201a ) or ( a202a );
 a13870a <=( a198a ) or ( a199a );
 a13871a <=( a200a ) or ( a13870a );
 a13872a <=( a13871a ) or ( a13866a );
 a13873a <=( a13872a ) or ( a13863a );
 a13876a <=( a196a ) or ( a197a );
 a13880a <=( a193a ) or ( a194a );
 a13881a <=( a195a ) or ( a13880a );
 a13882a <=( a13881a ) or ( a13876a );
 a13885a <=( a191a ) or ( a192a );
 a13889a <=( a188a ) or ( a189a );
 a13890a <=( a190a ) or ( a13889a );
 a13891a <=( a13890a ) or ( a13885a );
 a13892a <=( a13891a ) or ( a13882a );
 a13893a <=( a13892a ) or ( a13873a );
 a13894a <=( a13893a ) or ( a13856a );
 a13897a <=( a186a ) or ( a187a );
 a13900a <=( a184a ) or ( a185a );
 a13901a <=( a13900a ) or ( a13897a );
 a13904a <=( a182a ) or ( a183a );
 a13908a <=( a179a ) or ( a180a );
 a13909a <=( a181a ) or ( a13908a );
 a13910a <=( a13909a ) or ( a13904a );
 a13911a <=( a13910a ) or ( a13901a );
 a13914a <=( a177a ) or ( a178a );
 a13918a <=( a174a ) or ( a175a );
 a13919a <=( a176a ) or ( a13918a );
 a13920a <=( a13919a ) or ( a13914a );
 a13923a <=( a172a ) or ( a173a );
 a13927a <=( a169a ) or ( a170a );
 a13928a <=( a171a ) or ( a13927a );
 a13929a <=( a13928a ) or ( a13923a );
 a13930a <=( a13929a ) or ( a13920a );
 a13931a <=( a13930a ) or ( a13911a );
 a13934a <=( a167a ) or ( a168a );
 a13937a <=( a165a ) or ( a166a );
 a13938a <=( a13937a ) or ( a13934a );
 a13941a <=( a163a ) or ( a164a );
 a13945a <=( a160a ) or ( a161a );
 a13946a <=( a162a ) or ( a13945a );
 a13947a <=( a13946a ) or ( a13941a );
 a13948a <=( a13947a ) or ( a13938a );
 a13951a <=( a158a ) or ( a159a );
 a13955a <=( a155a ) or ( a156a );
 a13956a <=( a157a ) or ( a13955a );
 a13957a <=( a13956a ) or ( a13951a );
 a13960a <=( a153a ) or ( a154a );
 a13964a <=( a150a ) or ( a151a );
 a13965a <=( a152a ) or ( a13964a );
 a13966a <=( a13965a ) or ( a13960a );
 a13967a <=( a13966a ) or ( a13957a );
 a13968a <=( a13967a ) or ( a13948a );
 a13969a <=( a13968a ) or ( a13931a );
 a13970a <=( a13969a ) or ( a13894a );
 a13971a <=( a13970a ) or ( a13821a );
 a13974a <=( a148a ) or ( a149a );
 a13977a <=( a146a ) or ( a147a );
 a13978a <=( a13977a ) or ( a13974a );
 a13981a <=( a144a ) or ( a145a );
 a13985a <=( a141a ) or ( a142a );
 a13986a <=( a143a ) or ( a13985a );
 a13987a <=( a13986a ) or ( a13981a );
 a13988a <=( a13987a ) or ( a13978a );
 a13991a <=( a139a ) or ( a140a );
 a13994a <=( a137a ) or ( a138a );
 a13995a <=( a13994a ) or ( a13991a );
 a13998a <=( a135a ) or ( a136a );
 a14002a <=( a132a ) or ( a133a );
 a14003a <=( a134a ) or ( a14002a );
 a14004a <=( a14003a ) or ( a13998a );
 a14005a <=( a14004a ) or ( a13995a );
 a14006a <=( a14005a ) or ( a13988a );
 a14009a <=( a130a ) or ( a131a );
 a14012a <=( a128a ) or ( a129a );
 a14013a <=( a14012a ) or ( a14009a );
 a14016a <=( a126a ) or ( a127a );
 a14020a <=( a123a ) or ( a124a );
 a14021a <=( a125a ) or ( a14020a );
 a14022a <=( a14021a ) or ( a14016a );
 a14023a <=( a14022a ) or ( a14013a );
 a14026a <=( a121a ) or ( a122a );
 a14030a <=( a118a ) or ( a119a );
 a14031a <=( a120a ) or ( a14030a );
 a14032a <=( a14031a ) or ( a14026a );
 a14035a <=( a116a ) or ( a117a );
 a14039a <=( a113a ) or ( a114a );
 a14040a <=( a115a ) or ( a14039a );
 a14041a <=( a14040a ) or ( a14035a );
 a14042a <=( a14041a ) or ( a14032a );
 a14043a <=( a14042a ) or ( a14023a );
 a14044a <=( a14043a ) or ( a14006a );
 a14047a <=( a111a ) or ( a112a );
 a14050a <=( a109a ) or ( a110a );
 a14051a <=( a14050a ) or ( a14047a );
 a14054a <=( a107a ) or ( a108a );
 a14058a <=( a104a ) or ( a105a );
 a14059a <=( a106a ) or ( a14058a );
 a14060a <=( a14059a ) or ( a14054a );
 a14061a <=( a14060a ) or ( a14051a );
 a14064a <=( a102a ) or ( a103a );
 a14067a <=( a100a ) or ( a101a );
 a14068a <=( a14067a ) or ( a14064a );
 a14071a <=( a98a ) or ( a99a );
 a14075a <=( a95a ) or ( a96a );
 a14076a <=( a97a ) or ( a14075a );
 a14077a <=( a14076a ) or ( a14071a );
 a14078a <=( a14077a ) or ( a14068a );
 a14079a <=( a14078a ) or ( a14061a );
 a14082a <=( a93a ) or ( a94a );
 a14085a <=( a91a ) or ( a92a );
 a14086a <=( a14085a ) or ( a14082a );
 a14089a <=( a89a ) or ( a90a );
 a14093a <=( a86a ) or ( a87a );
 a14094a <=( a88a ) or ( a14093a );
 a14095a <=( a14094a ) or ( a14089a );
 a14096a <=( a14095a ) or ( a14086a );
 a14099a <=( a84a ) or ( a85a );
 a14103a <=( a81a ) or ( a82a );
 a14104a <=( a83a ) or ( a14103a );
 a14105a <=( a14104a ) or ( a14099a );
 a14108a <=( a79a ) or ( a80a );
 a14112a <=( a76a ) or ( a77a );
 a14113a <=( a78a ) or ( a14112a );
 a14114a <=( a14113a ) or ( a14108a );
 a14115a <=( a14114a ) or ( a14105a );
 a14116a <=( a14115a ) or ( a14096a );
 a14117a <=( a14116a ) or ( a14079a );
 a14118a <=( a14117a ) or ( a14044a );
 a14121a <=( a74a ) or ( a75a );
 a14124a <=( a72a ) or ( a73a );
 a14125a <=( a14124a ) or ( a14121a );
 a14128a <=( a70a ) or ( a71a );
 a14132a <=( a67a ) or ( a68a );
 a14133a <=( a69a ) or ( a14132a );
 a14134a <=( a14133a ) or ( a14128a );
 a14135a <=( a14134a ) or ( a14125a );
 a14138a <=( a65a ) or ( a66a );
 a14141a <=( a63a ) or ( a64a );
 a14142a <=( a14141a ) or ( a14138a );
 a14145a <=( a61a ) or ( a62a );
 a14149a <=( a58a ) or ( a59a );
 a14150a <=( a60a ) or ( a14149a );
 a14151a <=( a14150a ) or ( a14145a );
 a14152a <=( a14151a ) or ( a14142a );
 a14153a <=( a14152a ) or ( a14135a );
 a14156a <=( a56a ) or ( a57a );
 a14159a <=( a54a ) or ( a55a );
 a14160a <=( a14159a ) or ( a14156a );
 a14163a <=( a52a ) or ( a53a );
 a14167a <=( a49a ) or ( a50a );
 a14168a <=( a51a ) or ( a14167a );
 a14169a <=( a14168a ) or ( a14163a );
 a14170a <=( a14169a ) or ( a14160a );
 a14173a <=( a47a ) or ( a48a );
 a14177a <=( a44a ) or ( a45a );
 a14178a <=( a46a ) or ( a14177a );
 a14179a <=( a14178a ) or ( a14173a );
 a14182a <=( a42a ) or ( a43a );
 a14186a <=( a39a ) or ( a40a );
 a14187a <=( a41a ) or ( a14186a );
 a14188a <=( a14187a ) or ( a14182a );
 a14189a <=( a14188a ) or ( a14179a );
 a14190a <=( a14189a ) or ( a14170a );
 a14191a <=( a14190a ) or ( a14153a );
 a14194a <=( a37a ) or ( a38a );
 a14197a <=( a35a ) or ( a36a );
 a14198a <=( a14197a ) or ( a14194a );
 a14201a <=( a33a ) or ( a34a );
 a14205a <=( a30a ) or ( a31a );
 a14206a <=( a32a ) or ( a14205a );
 a14207a <=( a14206a ) or ( a14201a );
 a14208a <=( a14207a ) or ( a14198a );
 a14211a <=( a28a ) or ( a29a );
 a14215a <=( a25a ) or ( a26a );
 a14216a <=( a27a ) or ( a14215a );
 a14217a <=( a14216a ) or ( a14211a );
 a14220a <=( a23a ) or ( a24a );
 a14224a <=( a20a ) or ( a21a );
 a14225a <=( a22a ) or ( a14224a );
 a14226a <=( a14225a ) or ( a14220a );
 a14227a <=( a14226a ) or ( a14217a );
 a14228a <=( a14227a ) or ( a14208a );
 a14231a <=( a18a ) or ( a19a );
 a14234a <=( a16a ) or ( a17a );
 a14235a <=( a14234a ) or ( a14231a );
 a14238a <=( a14a ) or ( a15a );
 a14242a <=( a11a ) or ( a12a );
 a14243a <=( a13a ) or ( a14242a );
 a14244a <=( a14243a ) or ( a14238a );
 a14245a <=( a14244a ) or ( a14235a );
 a14248a <=( a9a ) or ( a10a );
 a14252a <=( a6a ) or ( a7a );
 a14253a <=( a8a ) or ( a14252a );
 a14254a <=( a14253a ) or ( a14248a );
 a14257a <=( a4a ) or ( a5a );
 a14261a <=( a1a ) or ( a2a );
 a14262a <=( a3a ) or ( a14261a );
 a14263a <=( a14262a ) or ( a14257a );
 a14264a <=( a14263a ) or ( a14254a );
 a14265a <=( a14264a ) or ( a14245a );
 a14266a <=( a14265a ) or ( a14228a );
 a14267a <=( a14266a ) or ( a14191a );
 a14268a <=( a14267a ) or ( a14118a );
 a14269a <=( a14268a ) or ( a13971a );
 a14270a <=( a14269a ) or ( a13674a );
 a14271a <=( a14270a ) or ( a13081a );
 a14272a <=( a14271a ) or ( a11892a );
 a14275a <=( A201  and  A199 );
 a14278a <=( A234  and  A232 );
 a14281a <=( A201  and  A199 );
 a14284a <=( A234  and  A233 );
 a14287a <=( A201  and  A200 );
 a14290a <=( A234  and  A232 );
 a14293a <=( A201  and  A200 );
 a14296a <=( A234  and  A233 );
 a14299a <=( (not A166)  and  A167 );
 a14302a <=( A234  and  A232 );
 a14305a <=( (not A166)  and  A167 );
 a14308a <=( A234  and  A233 );
 a14312a <=( A232  and  A201 );
 a14313a <=( A199  and  a14312a );
 a14317a <=( (not A236)  and  A235 );
 a14318a <=( A233  and  a14317a );
 a14322a <=( (not A232)  and  A201 );
 a14323a <=( A199  and  a14322a );
 a14327a <=( A236  and  (not A235) );
 a14328a <=( A233  and  a14327a );
 a14332a <=( A232  and  A201 );
 a14333a <=( A199  and  a14332a );
 a14337a <=( A236  and  (not A235) );
 a14338a <=( (not A233)  and  a14337a );
 a14342a <=( (not A232)  and  A201 );
 a14343a <=( A199  and  a14342a );
 a14347a <=( (not A236)  and  A235 );
 a14348a <=( (not A233)  and  a14347a );
 a14352a <=( A232  and  A201 );
 a14353a <=( A200  and  a14352a );
 a14357a <=( (not A236)  and  A235 );
 a14358a <=( A233  and  a14357a );
 a14362a <=( (not A232)  and  A201 );
 a14363a <=( A200  and  a14362a );
 a14367a <=( A236  and  (not A235) );
 a14368a <=( A233  and  a14367a );
 a14372a <=( A232  and  A201 );
 a14373a <=( A200  and  a14372a );
 a14377a <=( A236  and  (not A235) );
 a14378a <=( (not A233)  and  a14377a );
 a14382a <=( (not A232)  and  A201 );
 a14383a <=( A200  and  a14382a );
 a14387a <=( (not A236)  and  A235 );
 a14388a <=( (not A233)  and  a14387a );
 a14392a <=( A202  and  A200 );
 a14393a <=( A199  and  a14392a );
 a14397a <=( A234  and  A232 );
 a14398a <=( (not A203)  and  a14397a );
 a14402a <=( A202  and  A200 );
 a14403a <=( A199  and  a14402a );
 a14407a <=( A234  and  A233 );
 a14408a <=( (not A203)  and  a14407a );
 a14412a <=( (not A202)  and  A200 );
 a14413a <=( (not A199)  and  a14412a );
 a14417a <=( A234  and  A232 );
 a14418a <=( A203  and  a14417a );
 a14422a <=( (not A202)  and  A200 );
 a14423a <=( (not A199)  and  a14422a );
 a14427a <=( A234  and  A233 );
 a14428a <=( A203  and  a14427a );
 a14432a <=( (not A202)  and  (not A200) );
 a14433a <=( A199  and  a14432a );
 a14437a <=( A234  and  A232 );
 a14438a <=( A203  and  a14437a );
 a14442a <=( (not A202)  and  (not A200) );
 a14443a <=( A199  and  a14442a );
 a14447a <=( A234  and  A233 );
 a14448a <=( A203  and  a14447a );
 a14452a <=( A202  and  (not A200) );
 a14453a <=( (not A199)  and  a14452a );
 a14457a <=( A234  and  A232 );
 a14458a <=( (not A203)  and  a14457a );
 a14462a <=( A202  and  (not A200) );
 a14463a <=( (not A199)  and  a14462a );
 a14467a <=( A234  and  A233 );
 a14468a <=( (not A203)  and  a14467a );
 a14472a <=( A232  and  (not A166) );
 a14473a <=( A167  and  a14472a );
 a14477a <=( (not A236)  and  A235 );
 a14478a <=( A233  and  a14477a );
 a14482a <=( (not A232)  and  (not A166) );
 a14483a <=( A167  and  a14482a );
 a14487a <=( A236  and  (not A235) );
 a14488a <=( A233  and  a14487a );
 a14492a <=( A232  and  (not A166) );
 a14493a <=( A167  and  a14492a );
 a14497a <=( A236  and  (not A235) );
 a14498a <=( (not A233)  and  a14497a );
 a14502a <=( (not A232)  and  (not A166) );
 a14503a <=( A167  and  a14502a );
 a14507a <=( (not A236)  and  A235 );
 a14508a <=( (not A233)  and  a14507a );
 a14512a <=( (not A167)  and  A168 );
 a14513a <=( A170  and  a14512a );
 a14517a <=( A234  and  A232 );
 a14518a <=( A166  and  a14517a );
 a14522a <=( (not A167)  and  A168 );
 a14523a <=( A170  and  a14522a );
 a14527a <=( A234  and  A233 );
 a14528a <=( A166  and  a14527a );
 a14532a <=( (not A167)  and  A168 );
 a14533a <=( A169  and  a14532a );
 a14537a <=( A234  and  A232 );
 a14538a <=( A166  and  a14537a );
 a14542a <=( (not A167)  and  A168 );
 a14543a <=( A169  and  a14542a );
 a14547a <=( A234  and  A233 );
 a14548a <=( A166  and  a14547a );
 a14551a <=( A200  and  A199 );
 a14554a <=( (not A203)  and  A202 );
 a14555a <=( a14554a  and  a14551a );
 a14558a <=( A233  and  A232 );
 a14561a <=( (not A236)  and  A235 );
 a14562a <=( a14561a  and  a14558a );
 a14565a <=( A200  and  A199 );
 a14568a <=( (not A203)  and  A202 );
 a14569a <=( a14568a  and  a14565a );
 a14572a <=( A233  and  (not A232) );
 a14575a <=( A236  and  (not A235) );
 a14576a <=( a14575a  and  a14572a );
 a14579a <=( A200  and  A199 );
 a14582a <=( (not A203)  and  A202 );
 a14583a <=( a14582a  and  a14579a );
 a14586a <=( (not A233)  and  A232 );
 a14589a <=( A236  and  (not A235) );
 a14590a <=( a14589a  and  a14586a );
 a14593a <=( A200  and  A199 );
 a14596a <=( (not A203)  and  A202 );
 a14597a <=( a14596a  and  a14593a );
 a14600a <=( (not A233)  and  (not A232) );
 a14603a <=( (not A236)  and  A235 );
 a14604a <=( a14603a  and  a14600a );
 a14607a <=( A200  and  (not A199) );
 a14610a <=( A203  and  (not A202) );
 a14611a <=( a14610a  and  a14607a );
 a14614a <=( A233  and  A232 );
 a14617a <=( (not A236)  and  A235 );
 a14618a <=( a14617a  and  a14614a );
 a14621a <=( A200  and  (not A199) );
 a14624a <=( A203  and  (not A202) );
 a14625a <=( a14624a  and  a14621a );
 a14628a <=( A233  and  (not A232) );
 a14631a <=( A236  and  (not A235) );
 a14632a <=( a14631a  and  a14628a );
 a14635a <=( A200  and  (not A199) );
 a14638a <=( A203  and  (not A202) );
 a14639a <=( a14638a  and  a14635a );
 a14642a <=( (not A233)  and  A232 );
 a14645a <=( A236  and  (not A235) );
 a14646a <=( a14645a  and  a14642a );
 a14649a <=( A200  and  (not A199) );
 a14652a <=( A203  and  (not A202) );
 a14653a <=( a14652a  and  a14649a );
 a14656a <=( (not A233)  and  (not A232) );
 a14659a <=( (not A236)  and  A235 );
 a14660a <=( a14659a  and  a14656a );
 a14663a <=( (not A200)  and  A199 );
 a14666a <=( A203  and  (not A202) );
 a14667a <=( a14666a  and  a14663a );
 a14670a <=( A233  and  A232 );
 a14673a <=( (not A236)  and  A235 );
 a14674a <=( a14673a  and  a14670a );
 a14677a <=( (not A200)  and  A199 );
 a14680a <=( A203  and  (not A202) );
 a14681a <=( a14680a  and  a14677a );
 a14684a <=( A233  and  (not A232) );
 a14687a <=( A236  and  (not A235) );
 a14688a <=( a14687a  and  a14684a );
 a14691a <=( (not A200)  and  A199 );
 a14694a <=( A203  and  (not A202) );
 a14695a <=( a14694a  and  a14691a );
 a14698a <=( (not A233)  and  A232 );
 a14701a <=( A236  and  (not A235) );
 a14702a <=( a14701a  and  a14698a );
 a14705a <=( (not A200)  and  A199 );
 a14708a <=( A203  and  (not A202) );
 a14709a <=( a14708a  and  a14705a );
 a14712a <=( (not A233)  and  (not A232) );
 a14715a <=( (not A236)  and  A235 );
 a14716a <=( a14715a  and  a14712a );
 a14719a <=( (not A200)  and  (not A199) );
 a14722a <=( (not A203)  and  A202 );
 a14723a <=( a14722a  and  a14719a );
 a14726a <=( A233  and  A232 );
 a14729a <=( (not A236)  and  A235 );
 a14730a <=( a14729a  and  a14726a );
 a14733a <=( (not A200)  and  (not A199) );
 a14736a <=( (not A203)  and  A202 );
 a14737a <=( a14736a  and  a14733a );
 a14740a <=( A233  and  (not A232) );
 a14743a <=( A236  and  (not A235) );
 a14744a <=( a14743a  and  a14740a );
 a14747a <=( (not A200)  and  (not A199) );
 a14750a <=( (not A203)  and  A202 );
 a14751a <=( a14750a  and  a14747a );
 a14754a <=( (not A233)  and  A232 );
 a14757a <=( A236  and  (not A235) );
 a14758a <=( a14757a  and  a14754a );
 a14761a <=( (not A200)  and  (not A199) );
 a14764a <=( (not A203)  and  A202 );
 a14765a <=( a14764a  and  a14761a );
 a14768a <=( (not A233)  and  (not A232) );
 a14771a <=( (not A236)  and  A235 );
 a14772a <=( a14771a  and  a14768a );
 a14775a <=( A168  and  A170 );
 a14778a <=( A166  and  (not A167) );
 a14779a <=( a14778a  and  a14775a );
 a14782a <=( A233  and  A232 );
 a14785a <=( (not A236)  and  A235 );
 a14786a <=( a14785a  and  a14782a );
 a14789a <=( A168  and  A170 );
 a14792a <=( A166  and  (not A167) );
 a14793a <=( a14792a  and  a14789a );
 a14796a <=( A233  and  (not A232) );
 a14799a <=( A236  and  (not A235) );
 a14800a <=( a14799a  and  a14796a );
 a14803a <=( A168  and  A170 );
 a14806a <=( A166  and  (not A167) );
 a14807a <=( a14806a  and  a14803a );
 a14810a <=( (not A233)  and  A232 );
 a14813a <=( A236  and  (not A235) );
 a14814a <=( a14813a  and  a14810a );
 a14817a <=( A168  and  A170 );
 a14820a <=( A166  and  (not A167) );
 a14821a <=( a14820a  and  a14817a );
 a14824a <=( (not A233)  and  (not A232) );
 a14827a <=( (not A236)  and  A235 );
 a14828a <=( a14827a  and  a14824a );
 a14831a <=( A168  and  A169 );
 a14834a <=( A166  and  (not A167) );
 a14835a <=( a14834a  and  a14831a );
 a14838a <=( A233  and  A232 );
 a14841a <=( (not A236)  and  A235 );
 a14842a <=( a14841a  and  a14838a );
 a14845a <=( A168  and  A169 );
 a14848a <=( A166  and  (not A167) );
 a14849a <=( a14848a  and  a14845a );
 a14852a <=( A233  and  (not A232) );
 a14855a <=( A236  and  (not A235) );
 a14856a <=( a14855a  and  a14852a );
 a14859a <=( A168  and  A169 );
 a14862a <=( A166  and  (not A167) );
 a14863a <=( a14862a  and  a14859a );
 a14866a <=( (not A233)  and  A232 );
 a14869a <=( A236  and  (not A235) );
 a14870a <=( a14869a  and  a14866a );
 a14873a <=( A168  and  A169 );
 a14876a <=( A166  and  (not A167) );
 a14877a <=( a14876a  and  a14873a );
 a14880a <=( (not A233)  and  (not A232) );
 a14883a <=( (not A236)  and  A235 );
 a14884a <=( a14883a  and  a14880a );
 a14887a <=( A166  and  A167 );
 a14890a <=( A201  and  A199 );
 a14891a <=( a14890a  and  a14887a );
 a14894a <=( (not A266)  and  (not A265) );
 a14898a <=( A300  and  A299 );
 a14899a <=( (not A268)  and  a14898a );
 a14900a <=( a14899a  and  a14894a );
 a14903a <=( A166  and  A167 );
 a14906a <=( A201  and  A199 );
 a14907a <=( a14906a  and  a14903a );
 a14910a <=( (not A266)  and  (not A265) );
 a14914a <=( A300  and  A298 );
 a14915a <=( (not A268)  and  a14914a );
 a14916a <=( a14915a  and  a14910a );
 a14919a <=( A166  and  A167 );
 a14922a <=( A201  and  A199 );
 a14923a <=( a14922a  and  a14919a );
 a14926a <=( (not A266)  and  (not A265) );
 a14930a <=( A300  and  A299 );
 a14931a <=( A269  and  a14930a );
 a14932a <=( a14931a  and  a14926a );
 a14935a <=( A166  and  A167 );
 a14938a <=( A201  and  A199 );
 a14939a <=( a14938a  and  a14935a );
 a14942a <=( (not A266)  and  (not A265) );
 a14946a <=( A300  and  A298 );
 a14947a <=( A269  and  a14946a );
 a14948a <=( a14947a  and  a14942a );
 a14951a <=( A166  and  A167 );
 a14954a <=( A201  and  A200 );
 a14955a <=( a14954a  and  a14951a );
 a14958a <=( (not A266)  and  (not A265) );
 a14962a <=( A300  and  A299 );
 a14963a <=( (not A268)  and  a14962a );
 a14964a <=( a14963a  and  a14958a );
 a14967a <=( A166  and  A167 );
 a14970a <=( A201  and  A200 );
 a14971a <=( a14970a  and  a14967a );
 a14974a <=( (not A266)  and  (not A265) );
 a14978a <=( A300  and  A298 );
 a14979a <=( (not A268)  and  a14978a );
 a14980a <=( a14979a  and  a14974a );
 a14983a <=( A166  and  A167 );
 a14986a <=( A201  and  A200 );
 a14987a <=( a14986a  and  a14983a );
 a14990a <=( (not A266)  and  (not A265) );
 a14994a <=( A300  and  A299 );
 a14995a <=( A269  and  a14994a );
 a14996a <=( a14995a  and  a14990a );
 a14999a <=( A166  and  A167 );
 a15002a <=( A201  and  A200 );
 a15003a <=( a15002a  and  a14999a );
 a15006a <=( (not A266)  and  (not A265) );
 a15010a <=( A300  and  A298 );
 a15011a <=( A269  and  a15010a );
 a15012a <=( a15011a  and  a15006a );
 a15015a <=( (not A166)  and  A167 );
 a15018a <=( A201  and  A199 );
 a15019a <=( a15018a  and  a15015a );
 a15022a <=( A267  and  A265 );
 a15026a <=( (not A301)  and  (not A299) );
 a15027a <=( (not A298)  and  a15026a );
 a15028a <=( a15027a  and  a15022a );
 a15031a <=( (not A166)  and  A167 );
 a15034a <=( A201  and  A199 );
 a15035a <=( a15034a  and  a15031a );
 a15038a <=( A267  and  A265 );
 a15042a <=( A302  and  (not A299) );
 a15043a <=( (not A298)  and  a15042a );
 a15044a <=( a15043a  and  a15038a );
 a15047a <=( (not A166)  and  A167 );
 a15050a <=( A201  and  A199 );
 a15051a <=( a15050a  and  a15047a );
 a15054a <=( A267  and  A266 );
 a15058a <=( (not A301)  and  (not A299) );
 a15059a <=( (not A298)  and  a15058a );
 a15060a <=( a15059a  and  a15054a );
 a15063a <=( (not A166)  and  A167 );
 a15066a <=( A201  and  A199 );
 a15067a <=( a15066a  and  a15063a );
 a15070a <=( A267  and  A266 );
 a15074a <=( A302  and  (not A299) );
 a15075a <=( (not A298)  and  a15074a );
 a15076a <=( a15075a  and  a15070a );
 a15079a <=( (not A166)  and  A167 );
 a15082a <=( A201  and  A200 );
 a15083a <=( a15082a  and  a15079a );
 a15086a <=( A267  and  A265 );
 a15090a <=( (not A301)  and  (not A299) );
 a15091a <=( (not A298)  and  a15090a );
 a15092a <=( a15091a  and  a15086a );
 a15095a <=( (not A166)  and  A167 );
 a15098a <=( A201  and  A200 );
 a15099a <=( a15098a  and  a15095a );
 a15102a <=( A267  and  A265 );
 a15106a <=( A302  and  (not A299) );
 a15107a <=( (not A298)  and  a15106a );
 a15108a <=( a15107a  and  a15102a );
 a15111a <=( (not A166)  and  A167 );
 a15114a <=( A201  and  A200 );
 a15115a <=( a15114a  and  a15111a );
 a15118a <=( A267  and  A266 );
 a15122a <=( (not A301)  and  (not A299) );
 a15123a <=( (not A298)  and  a15122a );
 a15124a <=( a15123a  and  a15118a );
 a15127a <=( (not A166)  and  A167 );
 a15130a <=( A201  and  A200 );
 a15131a <=( a15130a  and  a15127a );
 a15134a <=( A267  and  A266 );
 a15138a <=( A302  and  (not A299) );
 a15139a <=( (not A298)  and  a15138a );
 a15140a <=( a15139a  and  a15134a );
 a15143a <=( (not A166)  and  (not A167) );
 a15146a <=( A201  and  A199 );
 a15147a <=( a15146a  and  a15143a );
 a15150a <=( (not A266)  and  (not A265) );
 a15154a <=( A300  and  A299 );
 a15155a <=( (not A268)  and  a15154a );
 a15156a <=( a15155a  and  a15150a );
 a15159a <=( (not A166)  and  (not A167) );
 a15162a <=( A201  and  A199 );
 a15163a <=( a15162a  and  a15159a );
 a15166a <=( (not A266)  and  (not A265) );
 a15170a <=( A300  and  A298 );
 a15171a <=( (not A268)  and  a15170a );
 a15172a <=( a15171a  and  a15166a );
 a15175a <=( (not A166)  and  (not A167) );
 a15178a <=( A201  and  A199 );
 a15179a <=( a15178a  and  a15175a );
 a15182a <=( (not A266)  and  (not A265) );
 a15186a <=( A300  and  A299 );
 a15187a <=( A269  and  a15186a );
 a15188a <=( a15187a  and  a15182a );
 a15191a <=( (not A166)  and  (not A167) );
 a15194a <=( A201  and  A199 );
 a15195a <=( a15194a  and  a15191a );
 a15198a <=( (not A266)  and  (not A265) );
 a15202a <=( A300  and  A298 );
 a15203a <=( A269  and  a15202a );
 a15204a <=( a15203a  and  a15198a );
 a15207a <=( (not A166)  and  (not A167) );
 a15210a <=( A201  and  A200 );
 a15211a <=( a15210a  and  a15207a );
 a15214a <=( (not A266)  and  (not A265) );
 a15218a <=( A300  and  A299 );
 a15219a <=( (not A268)  and  a15218a );
 a15220a <=( a15219a  and  a15214a );
 a15223a <=( (not A166)  and  (not A167) );
 a15226a <=( A201  and  A200 );
 a15227a <=( a15226a  and  a15223a );
 a15230a <=( (not A266)  and  (not A265) );
 a15234a <=( A300  and  A298 );
 a15235a <=( (not A268)  and  a15234a );
 a15236a <=( a15235a  and  a15230a );
 a15239a <=( (not A166)  and  (not A167) );
 a15242a <=( A201  and  A200 );
 a15243a <=( a15242a  and  a15239a );
 a15246a <=( (not A266)  and  (not A265) );
 a15250a <=( A300  and  A299 );
 a15251a <=( A269  and  a15250a );
 a15252a <=( a15251a  and  a15246a );
 a15255a <=( (not A166)  and  (not A167) );
 a15258a <=( A201  and  A200 );
 a15259a <=( a15258a  and  a15255a );
 a15262a <=( (not A266)  and  (not A265) );
 a15266a <=( A300  and  A298 );
 a15267a <=( A269  and  a15266a );
 a15268a <=( a15267a  and  a15262a );
 a15271a <=( (not A167)  and  (not A168) );
 a15274a <=( A201  and  A199 );
 a15275a <=( a15274a  and  a15271a );
 a15278a <=( (not A266)  and  (not A265) );
 a15282a <=( A300  and  A299 );
 a15283a <=( (not A268)  and  a15282a );
 a15284a <=( a15283a  and  a15278a );
 a15287a <=( (not A167)  and  (not A168) );
 a15290a <=( A201  and  A199 );
 a15291a <=( a15290a  and  a15287a );
 a15294a <=( (not A266)  and  (not A265) );
 a15298a <=( A300  and  A298 );
 a15299a <=( (not A268)  and  a15298a );
 a15300a <=( a15299a  and  a15294a );
 a15303a <=( (not A167)  and  (not A168) );
 a15306a <=( A201  and  A199 );
 a15307a <=( a15306a  and  a15303a );
 a15310a <=( (not A266)  and  (not A265) );
 a15314a <=( A300  and  A299 );
 a15315a <=( A269  and  a15314a );
 a15316a <=( a15315a  and  a15310a );
 a15319a <=( (not A167)  and  (not A168) );
 a15322a <=( A201  and  A199 );
 a15323a <=( a15322a  and  a15319a );
 a15326a <=( (not A266)  and  (not A265) );
 a15330a <=( A300  and  A298 );
 a15331a <=( A269  and  a15330a );
 a15332a <=( a15331a  and  a15326a );
 a15335a <=( (not A167)  and  (not A168) );
 a15338a <=( A201  and  A200 );
 a15339a <=( a15338a  and  a15335a );
 a15342a <=( (not A266)  and  (not A265) );
 a15346a <=( A300  and  A299 );
 a15347a <=( (not A268)  and  a15346a );
 a15348a <=( a15347a  and  a15342a );
 a15351a <=( (not A167)  and  (not A168) );
 a15354a <=( A201  and  A200 );
 a15355a <=( a15354a  and  a15351a );
 a15358a <=( (not A266)  and  (not A265) );
 a15362a <=( A300  and  A298 );
 a15363a <=( (not A268)  and  a15362a );
 a15364a <=( a15363a  and  a15358a );
 a15367a <=( (not A167)  and  (not A168) );
 a15370a <=( A201  and  A200 );
 a15371a <=( a15370a  and  a15367a );
 a15374a <=( (not A266)  and  (not A265) );
 a15378a <=( A300  and  A299 );
 a15379a <=( A269  and  a15378a );
 a15380a <=( a15379a  and  a15374a );
 a15383a <=( (not A167)  and  (not A168) );
 a15386a <=( A201  and  A200 );
 a15387a <=( a15386a  and  a15383a );
 a15390a <=( (not A266)  and  (not A265) );
 a15394a <=( A300  and  A298 );
 a15395a <=( A269  and  a15394a );
 a15396a <=( a15395a  and  a15390a );
 a15399a <=( A166  and  A167 );
 a15403a <=( A265  and  A201 );
 a15404a <=( A199  and  a15403a );
 a15405a <=( a15404a  and  a15399a );
 a15408a <=( (not A267)  and  A266 );
 a15412a <=( A300  and  A299 );
 a15413a <=( (not A268)  and  a15412a );
 a15414a <=( a15413a  and  a15408a );
 a15417a <=( A166  and  A167 );
 a15421a <=( A265  and  A201 );
 a15422a <=( A199  and  a15421a );
 a15423a <=( a15422a  and  a15417a );
 a15426a <=( (not A267)  and  A266 );
 a15430a <=( A300  and  A298 );
 a15431a <=( (not A268)  and  a15430a );
 a15432a <=( a15431a  and  a15426a );
 a15435a <=( A166  and  A167 );
 a15439a <=( A265  and  A201 );
 a15440a <=( A199  and  a15439a );
 a15441a <=( a15440a  and  a15435a );
 a15444a <=( (not A267)  and  A266 );
 a15448a <=( A300  and  A299 );
 a15449a <=( A269  and  a15448a );
 a15450a <=( a15449a  and  a15444a );
 a15453a <=( A166  and  A167 );
 a15457a <=( A265  and  A201 );
 a15458a <=( A199  and  a15457a );
 a15459a <=( a15458a  and  a15453a );
 a15462a <=( (not A267)  and  A266 );
 a15466a <=( A300  and  A298 );
 a15467a <=( A269  and  a15466a );
 a15468a <=( a15467a  and  a15462a );
 a15471a <=( A166  and  A167 );
 a15475a <=( (not A265)  and  A201 );
 a15476a <=( A199  and  a15475a );
 a15477a <=( a15476a  and  a15471a );
 a15480a <=( (not A267)  and  A266 );
 a15484a <=( A300  and  A299 );
 a15485a <=( A268  and  a15484a );
 a15486a <=( a15485a  and  a15480a );
 a15489a <=( A166  and  A167 );
 a15493a <=( (not A265)  and  A201 );
 a15494a <=( A199  and  a15493a );
 a15495a <=( a15494a  and  a15489a );
 a15498a <=( (not A267)  and  A266 );
 a15502a <=( A300  and  A298 );
 a15503a <=( A268  and  a15502a );
 a15504a <=( a15503a  and  a15498a );
 a15507a <=( A166  and  A167 );
 a15511a <=( (not A265)  and  A201 );
 a15512a <=( A199  and  a15511a );
 a15513a <=( a15512a  and  a15507a );
 a15516a <=( (not A267)  and  A266 );
 a15520a <=( A300  and  A299 );
 a15521a <=( (not A269)  and  a15520a );
 a15522a <=( a15521a  and  a15516a );
 a15525a <=( A166  and  A167 );
 a15529a <=( (not A265)  and  A201 );
 a15530a <=( A199  and  a15529a );
 a15531a <=( a15530a  and  a15525a );
 a15534a <=( (not A267)  and  A266 );
 a15538a <=( A300  and  A298 );
 a15539a <=( (not A269)  and  a15538a );
 a15540a <=( a15539a  and  a15534a );
 a15543a <=( A166  and  A167 );
 a15547a <=( A265  and  A201 );
 a15548a <=( A199  and  a15547a );
 a15549a <=( a15548a  and  a15543a );
 a15552a <=( (not A267)  and  (not A266) );
 a15556a <=( A300  and  A299 );
 a15557a <=( A268  and  a15556a );
 a15558a <=( a15557a  and  a15552a );
 a15561a <=( A166  and  A167 );
 a15565a <=( A265  and  A201 );
 a15566a <=( A199  and  a15565a );
 a15567a <=( a15566a  and  a15561a );
 a15570a <=( (not A267)  and  (not A266) );
 a15574a <=( A300  and  A298 );
 a15575a <=( A268  and  a15574a );
 a15576a <=( a15575a  and  a15570a );
 a15579a <=( A166  and  A167 );
 a15583a <=( A265  and  A201 );
 a15584a <=( A199  and  a15583a );
 a15585a <=( a15584a  and  a15579a );
 a15588a <=( (not A267)  and  (not A266) );
 a15592a <=( A300  and  A299 );
 a15593a <=( (not A269)  and  a15592a );
 a15594a <=( a15593a  and  a15588a );
 a15597a <=( A166  and  A167 );
 a15601a <=( A265  and  A201 );
 a15602a <=( A199  and  a15601a );
 a15603a <=( a15602a  and  a15597a );
 a15606a <=( (not A267)  and  (not A266) );
 a15610a <=( A300  and  A298 );
 a15611a <=( (not A269)  and  a15610a );
 a15612a <=( a15611a  and  a15606a );
 a15615a <=( A166  and  A167 );
 a15619a <=( A265  and  A201 );
 a15620a <=( A200  and  a15619a );
 a15621a <=( a15620a  and  a15615a );
 a15624a <=( (not A267)  and  A266 );
 a15628a <=( A300  and  A299 );
 a15629a <=( (not A268)  and  a15628a );
 a15630a <=( a15629a  and  a15624a );
 a15633a <=( A166  and  A167 );
 a15637a <=( A265  and  A201 );
 a15638a <=( A200  and  a15637a );
 a15639a <=( a15638a  and  a15633a );
 a15642a <=( (not A267)  and  A266 );
 a15646a <=( A300  and  A298 );
 a15647a <=( (not A268)  and  a15646a );
 a15648a <=( a15647a  and  a15642a );
 a15651a <=( A166  and  A167 );
 a15655a <=( A265  and  A201 );
 a15656a <=( A200  and  a15655a );
 a15657a <=( a15656a  and  a15651a );
 a15660a <=( (not A267)  and  A266 );
 a15664a <=( A300  and  A299 );
 a15665a <=( A269  and  a15664a );
 a15666a <=( a15665a  and  a15660a );
 a15669a <=( A166  and  A167 );
 a15673a <=( A265  and  A201 );
 a15674a <=( A200  and  a15673a );
 a15675a <=( a15674a  and  a15669a );
 a15678a <=( (not A267)  and  A266 );
 a15682a <=( A300  and  A298 );
 a15683a <=( A269  and  a15682a );
 a15684a <=( a15683a  and  a15678a );
 a15687a <=( A166  and  A167 );
 a15691a <=( (not A265)  and  A201 );
 a15692a <=( A200  and  a15691a );
 a15693a <=( a15692a  and  a15687a );
 a15696a <=( (not A267)  and  A266 );
 a15700a <=( A300  and  A299 );
 a15701a <=( A268  and  a15700a );
 a15702a <=( a15701a  and  a15696a );
 a15705a <=( A166  and  A167 );
 a15709a <=( (not A265)  and  A201 );
 a15710a <=( A200  and  a15709a );
 a15711a <=( a15710a  and  a15705a );
 a15714a <=( (not A267)  and  A266 );
 a15718a <=( A300  and  A298 );
 a15719a <=( A268  and  a15718a );
 a15720a <=( a15719a  and  a15714a );
 a15723a <=( A166  and  A167 );
 a15727a <=( (not A265)  and  A201 );
 a15728a <=( A200  and  a15727a );
 a15729a <=( a15728a  and  a15723a );
 a15732a <=( (not A267)  and  A266 );
 a15736a <=( A300  and  A299 );
 a15737a <=( (not A269)  and  a15736a );
 a15738a <=( a15737a  and  a15732a );
 a15741a <=( A166  and  A167 );
 a15745a <=( (not A265)  and  A201 );
 a15746a <=( A200  and  a15745a );
 a15747a <=( a15746a  and  a15741a );
 a15750a <=( (not A267)  and  A266 );
 a15754a <=( A300  and  A298 );
 a15755a <=( (not A269)  and  a15754a );
 a15756a <=( a15755a  and  a15750a );
 a15759a <=( A166  and  A167 );
 a15763a <=( A265  and  A201 );
 a15764a <=( A200  and  a15763a );
 a15765a <=( a15764a  and  a15759a );
 a15768a <=( (not A267)  and  (not A266) );
 a15772a <=( A300  and  A299 );
 a15773a <=( A268  and  a15772a );
 a15774a <=( a15773a  and  a15768a );
 a15777a <=( A166  and  A167 );
 a15781a <=( A265  and  A201 );
 a15782a <=( A200  and  a15781a );
 a15783a <=( a15782a  and  a15777a );
 a15786a <=( (not A267)  and  (not A266) );
 a15790a <=( A300  and  A298 );
 a15791a <=( A268  and  a15790a );
 a15792a <=( a15791a  and  a15786a );
 a15795a <=( A166  and  A167 );
 a15799a <=( A265  and  A201 );
 a15800a <=( A200  and  a15799a );
 a15801a <=( a15800a  and  a15795a );
 a15804a <=( (not A267)  and  (not A266) );
 a15808a <=( A300  and  A299 );
 a15809a <=( (not A269)  and  a15808a );
 a15810a <=( a15809a  and  a15804a );
 a15813a <=( A166  and  A167 );
 a15817a <=( A265  and  A201 );
 a15818a <=( A200  and  a15817a );
 a15819a <=( a15818a  and  a15813a );
 a15822a <=( (not A267)  and  (not A266) );
 a15826a <=( A300  and  A298 );
 a15827a <=( (not A269)  and  a15826a );
 a15828a <=( a15827a  and  a15822a );
 a15831a <=( A166  and  A167 );
 a15835a <=( (not A202)  and  (not A200) );
 a15836a <=( (not A199)  and  a15835a );
 a15837a <=( a15836a  and  a15831a );
 a15840a <=( A267  and  A265 );
 a15844a <=( (not A301)  and  (not A299) );
 a15845a <=( (not A298)  and  a15844a );
 a15846a <=( a15845a  and  a15840a );
 a15849a <=( A166  and  A167 );
 a15853a <=( (not A202)  and  (not A200) );
 a15854a <=( (not A199)  and  a15853a );
 a15855a <=( a15854a  and  a15849a );
 a15858a <=( A267  and  A265 );
 a15862a <=( A302  and  (not A299) );
 a15863a <=( (not A298)  and  a15862a );
 a15864a <=( a15863a  and  a15858a );
 a15867a <=( A166  and  A167 );
 a15871a <=( (not A202)  and  (not A200) );
 a15872a <=( (not A199)  and  a15871a );
 a15873a <=( a15872a  and  a15867a );
 a15876a <=( A267  and  A266 );
 a15880a <=( (not A301)  and  (not A299) );
 a15881a <=( (not A298)  and  a15880a );
 a15882a <=( a15881a  and  a15876a );
 a15885a <=( A166  and  A167 );
 a15889a <=( (not A202)  and  (not A200) );
 a15890a <=( (not A199)  and  a15889a );
 a15891a <=( a15890a  and  a15885a );
 a15894a <=( A267  and  A266 );
 a15898a <=( A302  and  (not A299) );
 a15899a <=( (not A298)  and  a15898a );
 a15900a <=( a15899a  and  a15894a );
 a15903a <=( A166  and  A167 );
 a15907a <=( A203  and  (not A200) );
 a15908a <=( (not A199)  and  a15907a );
 a15909a <=( a15908a  and  a15903a );
 a15912a <=( A267  and  A265 );
 a15916a <=( (not A301)  and  (not A299) );
 a15917a <=( (not A298)  and  a15916a );
 a15918a <=( a15917a  and  a15912a );
 a15921a <=( A166  and  A167 );
 a15925a <=( A203  and  (not A200) );
 a15926a <=( (not A199)  and  a15925a );
 a15927a <=( a15926a  and  a15921a );
 a15930a <=( A267  and  A265 );
 a15934a <=( A302  and  (not A299) );
 a15935a <=( (not A298)  and  a15934a );
 a15936a <=( a15935a  and  a15930a );
 a15939a <=( A166  and  A167 );
 a15943a <=( A203  and  (not A200) );
 a15944a <=( (not A199)  and  a15943a );
 a15945a <=( a15944a  and  a15939a );
 a15948a <=( A267  and  A266 );
 a15952a <=( (not A301)  and  (not A299) );
 a15953a <=( (not A298)  and  a15952a );
 a15954a <=( a15953a  and  a15948a );
 a15957a <=( A166  and  A167 );
 a15961a <=( A203  and  (not A200) );
 a15962a <=( (not A199)  and  a15961a );
 a15963a <=( a15962a  and  a15957a );
 a15966a <=( A267  and  A266 );
 a15970a <=( A302  and  (not A299) );
 a15971a <=( (not A298)  and  a15970a );
 a15972a <=( a15971a  and  a15966a );
 a15975a <=( (not A166)  and  A167 );
 a15979a <=( A265  and  A201 );
 a15980a <=( A199  and  a15979a );
 a15981a <=( a15980a  and  a15975a );
 a15984a <=( A298  and  A267 );
 a15988a <=( (not A301)  and  (not A300) );
 a15989a <=( A299  and  a15988a );
 a15990a <=( a15989a  and  a15984a );
 a15993a <=( (not A166)  and  A167 );
 a15997a <=( A265  and  A201 );
 a15998a <=( A199  and  a15997a );
 a15999a <=( a15998a  and  a15993a );
 a16002a <=( A298  and  A267 );
 a16006a <=( A302  and  (not A300) );
 a16007a <=( A299  and  a16006a );
 a16008a <=( a16007a  and  a16002a );
 a16011a <=( (not A166)  and  A167 );
 a16015a <=( A265  and  A201 );
 a16016a <=( A199  and  a16015a );
 a16017a <=( a16016a  and  a16011a );
 a16020a <=( A298  and  A267 );
 a16024a <=( A301  and  (not A300) );
 a16025a <=( (not A299)  and  a16024a );
 a16026a <=( a16025a  and  a16020a );
 a16029a <=( (not A166)  and  A167 );
 a16033a <=( A265  and  A201 );
 a16034a <=( A199  and  a16033a );
 a16035a <=( a16034a  and  a16029a );
 a16038a <=( A298  and  A267 );
 a16042a <=( (not A302)  and  (not A300) );
 a16043a <=( (not A299)  and  a16042a );
 a16044a <=( a16043a  and  a16038a );
 a16047a <=( (not A166)  and  A167 );
 a16051a <=( A265  and  A201 );
 a16052a <=( A199  and  a16051a );
 a16053a <=( a16052a  and  a16047a );
 a16056a <=( (not A298)  and  A267 );
 a16060a <=( A301  and  (not A300) );
 a16061a <=( A299  and  a16060a );
 a16062a <=( a16061a  and  a16056a );
 a16065a <=( (not A166)  and  A167 );
 a16069a <=( A265  and  A201 );
 a16070a <=( A199  and  a16069a );
 a16071a <=( a16070a  and  a16065a );
 a16074a <=( (not A298)  and  A267 );
 a16078a <=( (not A302)  and  (not A300) );
 a16079a <=( A299  and  a16078a );
 a16080a <=( a16079a  and  a16074a );
 a16083a <=( (not A166)  and  A167 );
 a16087a <=( A266  and  A201 );
 a16088a <=( A199  and  a16087a );
 a16089a <=( a16088a  and  a16083a );
 a16092a <=( A298  and  A267 );
 a16096a <=( (not A301)  and  (not A300) );
 a16097a <=( A299  and  a16096a );
 a16098a <=( a16097a  and  a16092a );
 a16101a <=( (not A166)  and  A167 );
 a16105a <=( A266  and  A201 );
 a16106a <=( A199  and  a16105a );
 a16107a <=( a16106a  and  a16101a );
 a16110a <=( A298  and  A267 );
 a16114a <=( A302  and  (not A300) );
 a16115a <=( A299  and  a16114a );
 a16116a <=( a16115a  and  a16110a );
 a16119a <=( (not A166)  and  A167 );
 a16123a <=( A266  and  A201 );
 a16124a <=( A199  and  a16123a );
 a16125a <=( a16124a  and  a16119a );
 a16128a <=( A298  and  A267 );
 a16132a <=( A301  and  (not A300) );
 a16133a <=( (not A299)  and  a16132a );
 a16134a <=( a16133a  and  a16128a );
 a16137a <=( (not A166)  and  A167 );
 a16141a <=( A266  and  A201 );
 a16142a <=( A199  and  a16141a );
 a16143a <=( a16142a  and  a16137a );
 a16146a <=( A298  and  A267 );
 a16150a <=( (not A302)  and  (not A300) );
 a16151a <=( (not A299)  and  a16150a );
 a16152a <=( a16151a  and  a16146a );
 a16155a <=( (not A166)  and  A167 );
 a16159a <=( A266  and  A201 );
 a16160a <=( A199  and  a16159a );
 a16161a <=( a16160a  and  a16155a );
 a16164a <=( (not A298)  and  A267 );
 a16168a <=( A301  and  (not A300) );
 a16169a <=( A299  and  a16168a );
 a16170a <=( a16169a  and  a16164a );
 a16173a <=( (not A166)  and  A167 );
 a16177a <=( A266  and  A201 );
 a16178a <=( A199  and  a16177a );
 a16179a <=( a16178a  and  a16173a );
 a16182a <=( (not A298)  and  A267 );
 a16186a <=( (not A302)  and  (not A300) );
 a16187a <=( A299  and  a16186a );
 a16188a <=( a16187a  and  a16182a );
 a16191a <=( (not A166)  and  A167 );
 a16195a <=( A265  and  A201 );
 a16196a <=( A200  and  a16195a );
 a16197a <=( a16196a  and  a16191a );
 a16200a <=( A298  and  A267 );
 a16204a <=( (not A301)  and  (not A300) );
 a16205a <=( A299  and  a16204a );
 a16206a <=( a16205a  and  a16200a );
 a16209a <=( (not A166)  and  A167 );
 a16213a <=( A265  and  A201 );
 a16214a <=( A200  and  a16213a );
 a16215a <=( a16214a  and  a16209a );
 a16218a <=( A298  and  A267 );
 a16222a <=( A302  and  (not A300) );
 a16223a <=( A299  and  a16222a );
 a16224a <=( a16223a  and  a16218a );
 a16227a <=( (not A166)  and  A167 );
 a16231a <=( A265  and  A201 );
 a16232a <=( A200  and  a16231a );
 a16233a <=( a16232a  and  a16227a );
 a16236a <=( A298  and  A267 );
 a16240a <=( A301  and  (not A300) );
 a16241a <=( (not A299)  and  a16240a );
 a16242a <=( a16241a  and  a16236a );
 a16245a <=( (not A166)  and  A167 );
 a16249a <=( A265  and  A201 );
 a16250a <=( A200  and  a16249a );
 a16251a <=( a16250a  and  a16245a );
 a16254a <=( A298  and  A267 );
 a16258a <=( (not A302)  and  (not A300) );
 a16259a <=( (not A299)  and  a16258a );
 a16260a <=( a16259a  and  a16254a );
 a16263a <=( (not A166)  and  A167 );
 a16267a <=( A265  and  A201 );
 a16268a <=( A200  and  a16267a );
 a16269a <=( a16268a  and  a16263a );
 a16272a <=( (not A298)  and  A267 );
 a16276a <=( A301  and  (not A300) );
 a16277a <=( A299  and  a16276a );
 a16278a <=( a16277a  and  a16272a );
 a16281a <=( (not A166)  and  A167 );
 a16285a <=( A265  and  A201 );
 a16286a <=( A200  and  a16285a );
 a16287a <=( a16286a  and  a16281a );
 a16290a <=( (not A298)  and  A267 );
 a16294a <=( (not A302)  and  (not A300) );
 a16295a <=( A299  and  a16294a );
 a16296a <=( a16295a  and  a16290a );
 a16299a <=( (not A166)  and  A167 );
 a16303a <=( A266  and  A201 );
 a16304a <=( A200  and  a16303a );
 a16305a <=( a16304a  and  a16299a );
 a16308a <=( A298  and  A267 );
 a16312a <=( (not A301)  and  (not A300) );
 a16313a <=( A299  and  a16312a );
 a16314a <=( a16313a  and  a16308a );
 a16317a <=( (not A166)  and  A167 );
 a16321a <=( A266  and  A201 );
 a16322a <=( A200  and  a16321a );
 a16323a <=( a16322a  and  a16317a );
 a16326a <=( A298  and  A267 );
 a16330a <=( A302  and  (not A300) );
 a16331a <=( A299  and  a16330a );
 a16332a <=( a16331a  and  a16326a );
 a16335a <=( (not A166)  and  A167 );
 a16339a <=( A266  and  A201 );
 a16340a <=( A200  and  a16339a );
 a16341a <=( a16340a  and  a16335a );
 a16344a <=( A298  and  A267 );
 a16348a <=( A301  and  (not A300) );
 a16349a <=( (not A299)  and  a16348a );
 a16350a <=( a16349a  and  a16344a );
 a16353a <=( (not A166)  and  A167 );
 a16357a <=( A266  and  A201 );
 a16358a <=( A200  and  a16357a );
 a16359a <=( a16358a  and  a16353a );
 a16362a <=( A298  and  A267 );
 a16366a <=( (not A302)  and  (not A300) );
 a16367a <=( (not A299)  and  a16366a );
 a16368a <=( a16367a  and  a16362a );
 a16371a <=( (not A166)  and  A167 );
 a16375a <=( A266  and  A201 );
 a16376a <=( A200  and  a16375a );
 a16377a <=( a16376a  and  a16371a );
 a16380a <=( (not A298)  and  A267 );
 a16384a <=( A301  and  (not A300) );
 a16385a <=( A299  and  a16384a );
 a16386a <=( a16385a  and  a16380a );
 a16389a <=( (not A166)  and  A167 );
 a16393a <=( A266  and  A201 );
 a16394a <=( A200  and  a16393a );
 a16395a <=( a16394a  and  a16389a );
 a16398a <=( (not A298)  and  A267 );
 a16402a <=( (not A302)  and  (not A300) );
 a16403a <=( A299  and  a16402a );
 a16404a <=( a16403a  and  a16398a );
 a16407a <=( (not A166)  and  A167 );
 a16411a <=( (not A202)  and  (not A200) );
 a16412a <=( (not A199)  and  a16411a );
 a16413a <=( a16412a  and  a16407a );
 a16416a <=( (not A266)  and  (not A265) );
 a16420a <=( A300  and  A299 );
 a16421a <=( (not A268)  and  a16420a );
 a16422a <=( a16421a  and  a16416a );
 a16425a <=( (not A166)  and  A167 );
 a16429a <=( (not A202)  and  (not A200) );
 a16430a <=( (not A199)  and  a16429a );
 a16431a <=( a16430a  and  a16425a );
 a16434a <=( (not A266)  and  (not A265) );
 a16438a <=( A300  and  A298 );
 a16439a <=( (not A268)  and  a16438a );
 a16440a <=( a16439a  and  a16434a );
 a16443a <=( (not A166)  and  A167 );
 a16447a <=( (not A202)  and  (not A200) );
 a16448a <=( (not A199)  and  a16447a );
 a16449a <=( a16448a  and  a16443a );
 a16452a <=( (not A266)  and  (not A265) );
 a16456a <=( A300  and  A299 );
 a16457a <=( A269  and  a16456a );
 a16458a <=( a16457a  and  a16452a );
 a16461a <=( (not A166)  and  A167 );
 a16465a <=( (not A202)  and  (not A200) );
 a16466a <=( (not A199)  and  a16465a );
 a16467a <=( a16466a  and  a16461a );
 a16470a <=( (not A266)  and  (not A265) );
 a16474a <=( A300  and  A298 );
 a16475a <=( A269  and  a16474a );
 a16476a <=( a16475a  and  a16470a );
 a16479a <=( (not A166)  and  A167 );
 a16483a <=( A203  and  (not A200) );
 a16484a <=( (not A199)  and  a16483a );
 a16485a <=( a16484a  and  a16479a );
 a16488a <=( (not A266)  and  (not A265) );
 a16492a <=( A300  and  A299 );
 a16493a <=( (not A268)  and  a16492a );
 a16494a <=( a16493a  and  a16488a );
 a16497a <=( (not A166)  and  A167 );
 a16501a <=( A203  and  (not A200) );
 a16502a <=( (not A199)  and  a16501a );
 a16503a <=( a16502a  and  a16497a );
 a16506a <=( (not A266)  and  (not A265) );
 a16510a <=( A300  and  A298 );
 a16511a <=( (not A268)  and  a16510a );
 a16512a <=( a16511a  and  a16506a );
 a16515a <=( (not A166)  and  A167 );
 a16519a <=( A203  and  (not A200) );
 a16520a <=( (not A199)  and  a16519a );
 a16521a <=( a16520a  and  a16515a );
 a16524a <=( (not A266)  and  (not A265) );
 a16528a <=( A300  and  A299 );
 a16529a <=( A269  and  a16528a );
 a16530a <=( a16529a  and  a16524a );
 a16533a <=( (not A166)  and  A167 );
 a16537a <=( A203  and  (not A200) );
 a16538a <=( (not A199)  and  a16537a );
 a16539a <=( a16538a  and  a16533a );
 a16542a <=( (not A266)  and  (not A265) );
 a16546a <=( A300  and  A298 );
 a16547a <=( A269  and  a16546a );
 a16548a <=( a16547a  and  a16542a );
 a16551a <=( (not A166)  and  (not A167) );
 a16555a <=( A265  and  A201 );
 a16556a <=( A199  and  a16555a );
 a16557a <=( a16556a  and  a16551a );
 a16560a <=( (not A267)  and  A266 );
 a16564a <=( A300  and  A299 );
 a16565a <=( (not A268)  and  a16564a );
 a16566a <=( a16565a  and  a16560a );
 a16569a <=( (not A166)  and  (not A167) );
 a16573a <=( A265  and  A201 );
 a16574a <=( A199  and  a16573a );
 a16575a <=( a16574a  and  a16569a );
 a16578a <=( (not A267)  and  A266 );
 a16582a <=( A300  and  A298 );
 a16583a <=( (not A268)  and  a16582a );
 a16584a <=( a16583a  and  a16578a );
 a16587a <=( (not A166)  and  (not A167) );
 a16591a <=( A265  and  A201 );
 a16592a <=( A199  and  a16591a );
 a16593a <=( a16592a  and  a16587a );
 a16596a <=( (not A267)  and  A266 );
 a16600a <=( A300  and  A299 );
 a16601a <=( A269  and  a16600a );
 a16602a <=( a16601a  and  a16596a );
 a16605a <=( (not A166)  and  (not A167) );
 a16609a <=( A265  and  A201 );
 a16610a <=( A199  and  a16609a );
 a16611a <=( a16610a  and  a16605a );
 a16614a <=( (not A267)  and  A266 );
 a16618a <=( A300  and  A298 );
 a16619a <=( A269  and  a16618a );
 a16620a <=( a16619a  and  a16614a );
 a16623a <=( (not A166)  and  (not A167) );
 a16627a <=( (not A265)  and  A201 );
 a16628a <=( A199  and  a16627a );
 a16629a <=( a16628a  and  a16623a );
 a16632a <=( (not A267)  and  A266 );
 a16636a <=( A300  and  A299 );
 a16637a <=( A268  and  a16636a );
 a16638a <=( a16637a  and  a16632a );
 a16641a <=( (not A166)  and  (not A167) );
 a16645a <=( (not A265)  and  A201 );
 a16646a <=( A199  and  a16645a );
 a16647a <=( a16646a  and  a16641a );
 a16650a <=( (not A267)  and  A266 );
 a16654a <=( A300  and  A298 );
 a16655a <=( A268  and  a16654a );
 a16656a <=( a16655a  and  a16650a );
 a16659a <=( (not A166)  and  (not A167) );
 a16663a <=( (not A265)  and  A201 );
 a16664a <=( A199  and  a16663a );
 a16665a <=( a16664a  and  a16659a );
 a16668a <=( (not A267)  and  A266 );
 a16672a <=( A300  and  A299 );
 a16673a <=( (not A269)  and  a16672a );
 a16674a <=( a16673a  and  a16668a );
 a16677a <=( (not A166)  and  (not A167) );
 a16681a <=( (not A265)  and  A201 );
 a16682a <=( A199  and  a16681a );
 a16683a <=( a16682a  and  a16677a );
 a16686a <=( (not A267)  and  A266 );
 a16690a <=( A300  and  A298 );
 a16691a <=( (not A269)  and  a16690a );
 a16692a <=( a16691a  and  a16686a );
 a16695a <=( (not A166)  and  (not A167) );
 a16699a <=( A265  and  A201 );
 a16700a <=( A199  and  a16699a );
 a16701a <=( a16700a  and  a16695a );
 a16704a <=( (not A267)  and  (not A266) );
 a16708a <=( A300  and  A299 );
 a16709a <=( A268  and  a16708a );
 a16710a <=( a16709a  and  a16704a );
 a16713a <=( (not A166)  and  (not A167) );
 a16717a <=( A265  and  A201 );
 a16718a <=( A199  and  a16717a );
 a16719a <=( a16718a  and  a16713a );
 a16722a <=( (not A267)  and  (not A266) );
 a16726a <=( A300  and  A298 );
 a16727a <=( A268  and  a16726a );
 a16728a <=( a16727a  and  a16722a );
 a16731a <=( (not A166)  and  (not A167) );
 a16735a <=( A265  and  A201 );
 a16736a <=( A199  and  a16735a );
 a16737a <=( a16736a  and  a16731a );
 a16740a <=( (not A267)  and  (not A266) );
 a16744a <=( A300  and  A299 );
 a16745a <=( (not A269)  and  a16744a );
 a16746a <=( a16745a  and  a16740a );
 a16749a <=( (not A166)  and  (not A167) );
 a16753a <=( A265  and  A201 );
 a16754a <=( A199  and  a16753a );
 a16755a <=( a16754a  and  a16749a );
 a16758a <=( (not A267)  and  (not A266) );
 a16762a <=( A300  and  A298 );
 a16763a <=( (not A269)  and  a16762a );
 a16764a <=( a16763a  and  a16758a );
 a16767a <=( (not A166)  and  (not A167) );
 a16771a <=( A265  and  A201 );
 a16772a <=( A200  and  a16771a );
 a16773a <=( a16772a  and  a16767a );
 a16776a <=( (not A267)  and  A266 );
 a16780a <=( A300  and  A299 );
 a16781a <=( (not A268)  and  a16780a );
 a16782a <=( a16781a  and  a16776a );
 a16785a <=( (not A166)  and  (not A167) );
 a16789a <=( A265  and  A201 );
 a16790a <=( A200  and  a16789a );
 a16791a <=( a16790a  and  a16785a );
 a16794a <=( (not A267)  and  A266 );
 a16798a <=( A300  and  A298 );
 a16799a <=( (not A268)  and  a16798a );
 a16800a <=( a16799a  and  a16794a );
 a16803a <=( (not A166)  and  (not A167) );
 a16807a <=( A265  and  A201 );
 a16808a <=( A200  and  a16807a );
 a16809a <=( a16808a  and  a16803a );
 a16812a <=( (not A267)  and  A266 );
 a16816a <=( A300  and  A299 );
 a16817a <=( A269  and  a16816a );
 a16818a <=( a16817a  and  a16812a );
 a16821a <=( (not A166)  and  (not A167) );
 a16825a <=( A265  and  A201 );
 a16826a <=( A200  and  a16825a );
 a16827a <=( a16826a  and  a16821a );
 a16830a <=( (not A267)  and  A266 );
 a16834a <=( A300  and  A298 );
 a16835a <=( A269  and  a16834a );
 a16836a <=( a16835a  and  a16830a );
 a16839a <=( (not A166)  and  (not A167) );
 a16843a <=( (not A265)  and  A201 );
 a16844a <=( A200  and  a16843a );
 a16845a <=( a16844a  and  a16839a );
 a16848a <=( (not A267)  and  A266 );
 a16852a <=( A300  and  A299 );
 a16853a <=( A268  and  a16852a );
 a16854a <=( a16853a  and  a16848a );
 a16857a <=( (not A166)  and  (not A167) );
 a16861a <=( (not A265)  and  A201 );
 a16862a <=( A200  and  a16861a );
 a16863a <=( a16862a  and  a16857a );
 a16866a <=( (not A267)  and  A266 );
 a16870a <=( A300  and  A298 );
 a16871a <=( A268  and  a16870a );
 a16872a <=( a16871a  and  a16866a );
 a16875a <=( (not A166)  and  (not A167) );
 a16879a <=( (not A265)  and  A201 );
 a16880a <=( A200  and  a16879a );
 a16881a <=( a16880a  and  a16875a );
 a16884a <=( (not A267)  and  A266 );
 a16888a <=( A300  and  A299 );
 a16889a <=( (not A269)  and  a16888a );
 a16890a <=( a16889a  and  a16884a );
 a16893a <=( (not A166)  and  (not A167) );
 a16897a <=( (not A265)  and  A201 );
 a16898a <=( A200  and  a16897a );
 a16899a <=( a16898a  and  a16893a );
 a16902a <=( (not A267)  and  A266 );
 a16906a <=( A300  and  A298 );
 a16907a <=( (not A269)  and  a16906a );
 a16908a <=( a16907a  and  a16902a );
 a16911a <=( (not A166)  and  (not A167) );
 a16915a <=( A265  and  A201 );
 a16916a <=( A200  and  a16915a );
 a16917a <=( a16916a  and  a16911a );
 a16920a <=( (not A267)  and  (not A266) );
 a16924a <=( A300  and  A299 );
 a16925a <=( A268  and  a16924a );
 a16926a <=( a16925a  and  a16920a );
 a16929a <=( (not A166)  and  (not A167) );
 a16933a <=( A265  and  A201 );
 a16934a <=( A200  and  a16933a );
 a16935a <=( a16934a  and  a16929a );
 a16938a <=( (not A267)  and  (not A266) );
 a16942a <=( A300  and  A298 );
 a16943a <=( A268  and  a16942a );
 a16944a <=( a16943a  and  a16938a );
 a16947a <=( (not A166)  and  (not A167) );
 a16951a <=( A265  and  A201 );
 a16952a <=( A200  and  a16951a );
 a16953a <=( a16952a  and  a16947a );
 a16956a <=( (not A267)  and  (not A266) );
 a16960a <=( A300  and  A299 );
 a16961a <=( (not A269)  and  a16960a );
 a16962a <=( a16961a  and  a16956a );
 a16965a <=( (not A166)  and  (not A167) );
 a16969a <=( A265  and  A201 );
 a16970a <=( A200  and  a16969a );
 a16971a <=( a16970a  and  a16965a );
 a16974a <=( (not A267)  and  (not A266) );
 a16978a <=( A300  and  A298 );
 a16979a <=( (not A269)  and  a16978a );
 a16980a <=( a16979a  and  a16974a );
 a16983a <=( (not A166)  and  (not A167) );
 a16987a <=( (not A202)  and  (not A200) );
 a16988a <=( (not A199)  and  a16987a );
 a16989a <=( a16988a  and  a16983a );
 a16992a <=( A267  and  A265 );
 a16996a <=( (not A301)  and  (not A299) );
 a16997a <=( (not A298)  and  a16996a );
 a16998a <=( a16997a  and  a16992a );
 a17001a <=( (not A166)  and  (not A167) );
 a17005a <=( (not A202)  and  (not A200) );
 a17006a <=( (not A199)  and  a17005a );
 a17007a <=( a17006a  and  a17001a );
 a17010a <=( A267  and  A265 );
 a17014a <=( A302  and  (not A299) );
 a17015a <=( (not A298)  and  a17014a );
 a17016a <=( a17015a  and  a17010a );
 a17019a <=( (not A166)  and  (not A167) );
 a17023a <=( (not A202)  and  (not A200) );
 a17024a <=( (not A199)  and  a17023a );
 a17025a <=( a17024a  and  a17019a );
 a17028a <=( A267  and  A266 );
 a17032a <=( (not A301)  and  (not A299) );
 a17033a <=( (not A298)  and  a17032a );
 a17034a <=( a17033a  and  a17028a );
 a17037a <=( (not A166)  and  (not A167) );
 a17041a <=( (not A202)  and  (not A200) );
 a17042a <=( (not A199)  and  a17041a );
 a17043a <=( a17042a  and  a17037a );
 a17046a <=( A267  and  A266 );
 a17050a <=( A302  and  (not A299) );
 a17051a <=( (not A298)  and  a17050a );
 a17052a <=( a17051a  and  a17046a );
 a17055a <=( (not A166)  and  (not A167) );
 a17059a <=( A203  and  (not A200) );
 a17060a <=( (not A199)  and  a17059a );
 a17061a <=( a17060a  and  a17055a );
 a17064a <=( A267  and  A265 );
 a17068a <=( (not A301)  and  (not A299) );
 a17069a <=( (not A298)  and  a17068a );
 a17070a <=( a17069a  and  a17064a );
 a17073a <=( (not A166)  and  (not A167) );
 a17077a <=( A203  and  (not A200) );
 a17078a <=( (not A199)  and  a17077a );
 a17079a <=( a17078a  and  a17073a );
 a17082a <=( A267  and  A265 );
 a17086a <=( A302  and  (not A299) );
 a17087a <=( (not A298)  and  a17086a );
 a17088a <=( a17087a  and  a17082a );
 a17091a <=( (not A166)  and  (not A167) );
 a17095a <=( A203  and  (not A200) );
 a17096a <=( (not A199)  and  a17095a );
 a17097a <=( a17096a  and  a17091a );
 a17100a <=( A267  and  A266 );
 a17104a <=( (not A301)  and  (not A299) );
 a17105a <=( (not A298)  and  a17104a );
 a17106a <=( a17105a  and  a17100a );
 a17109a <=( (not A166)  and  (not A167) );
 a17113a <=( A203  and  (not A200) );
 a17114a <=( (not A199)  and  a17113a );
 a17115a <=( a17114a  and  a17109a );
 a17118a <=( A267  and  A266 );
 a17122a <=( A302  and  (not A299) );
 a17123a <=( (not A298)  and  a17122a );
 a17124a <=( a17123a  and  a17118a );
 a17127a <=( (not A167)  and  (not A168) );
 a17131a <=( A265  and  A201 );
 a17132a <=( A199  and  a17131a );
 a17133a <=( a17132a  and  a17127a );
 a17136a <=( (not A267)  and  A266 );
 a17140a <=( A300  and  A299 );
 a17141a <=( (not A268)  and  a17140a );
 a17142a <=( a17141a  and  a17136a );
 a17145a <=( (not A167)  and  (not A168) );
 a17149a <=( A265  and  A201 );
 a17150a <=( A199  and  a17149a );
 a17151a <=( a17150a  and  a17145a );
 a17154a <=( (not A267)  and  A266 );
 a17158a <=( A300  and  A298 );
 a17159a <=( (not A268)  and  a17158a );
 a17160a <=( a17159a  and  a17154a );
 a17163a <=( (not A167)  and  (not A168) );
 a17167a <=( A265  and  A201 );
 a17168a <=( A199  and  a17167a );
 a17169a <=( a17168a  and  a17163a );
 a17172a <=( (not A267)  and  A266 );
 a17176a <=( A300  and  A299 );
 a17177a <=( A269  and  a17176a );
 a17178a <=( a17177a  and  a17172a );
 a17181a <=( (not A167)  and  (not A168) );
 a17185a <=( A265  and  A201 );
 a17186a <=( A199  and  a17185a );
 a17187a <=( a17186a  and  a17181a );
 a17190a <=( (not A267)  and  A266 );
 a17194a <=( A300  and  A298 );
 a17195a <=( A269  and  a17194a );
 a17196a <=( a17195a  and  a17190a );
 a17199a <=( (not A167)  and  (not A168) );
 a17203a <=( (not A265)  and  A201 );
 a17204a <=( A199  and  a17203a );
 a17205a <=( a17204a  and  a17199a );
 a17208a <=( (not A267)  and  A266 );
 a17212a <=( A300  and  A299 );
 a17213a <=( A268  and  a17212a );
 a17214a <=( a17213a  and  a17208a );
 a17217a <=( (not A167)  and  (not A168) );
 a17221a <=( (not A265)  and  A201 );
 a17222a <=( A199  and  a17221a );
 a17223a <=( a17222a  and  a17217a );
 a17226a <=( (not A267)  and  A266 );
 a17230a <=( A300  and  A298 );
 a17231a <=( A268  and  a17230a );
 a17232a <=( a17231a  and  a17226a );
 a17235a <=( (not A167)  and  (not A168) );
 a17239a <=( (not A265)  and  A201 );
 a17240a <=( A199  and  a17239a );
 a17241a <=( a17240a  and  a17235a );
 a17244a <=( (not A267)  and  A266 );
 a17248a <=( A300  and  A299 );
 a17249a <=( (not A269)  and  a17248a );
 a17250a <=( a17249a  and  a17244a );
 a17253a <=( (not A167)  and  (not A168) );
 a17257a <=( (not A265)  and  A201 );
 a17258a <=( A199  and  a17257a );
 a17259a <=( a17258a  and  a17253a );
 a17262a <=( (not A267)  and  A266 );
 a17266a <=( A300  and  A298 );
 a17267a <=( (not A269)  and  a17266a );
 a17268a <=( a17267a  and  a17262a );
 a17271a <=( (not A167)  and  (not A168) );
 a17275a <=( A265  and  A201 );
 a17276a <=( A199  and  a17275a );
 a17277a <=( a17276a  and  a17271a );
 a17280a <=( (not A267)  and  (not A266) );
 a17284a <=( A300  and  A299 );
 a17285a <=( A268  and  a17284a );
 a17286a <=( a17285a  and  a17280a );
 a17289a <=( (not A167)  and  (not A168) );
 a17293a <=( A265  and  A201 );
 a17294a <=( A199  and  a17293a );
 a17295a <=( a17294a  and  a17289a );
 a17298a <=( (not A267)  and  (not A266) );
 a17302a <=( A300  and  A298 );
 a17303a <=( A268  and  a17302a );
 a17304a <=( a17303a  and  a17298a );
 a17307a <=( (not A167)  and  (not A168) );
 a17311a <=( A265  and  A201 );
 a17312a <=( A199  and  a17311a );
 a17313a <=( a17312a  and  a17307a );
 a17316a <=( (not A267)  and  (not A266) );
 a17320a <=( A300  and  A299 );
 a17321a <=( (not A269)  and  a17320a );
 a17322a <=( a17321a  and  a17316a );
 a17325a <=( (not A167)  and  (not A168) );
 a17329a <=( A265  and  A201 );
 a17330a <=( A199  and  a17329a );
 a17331a <=( a17330a  and  a17325a );
 a17334a <=( (not A267)  and  (not A266) );
 a17338a <=( A300  and  A298 );
 a17339a <=( (not A269)  and  a17338a );
 a17340a <=( a17339a  and  a17334a );
 a17343a <=( (not A167)  and  (not A168) );
 a17347a <=( A265  and  A201 );
 a17348a <=( A200  and  a17347a );
 a17349a <=( a17348a  and  a17343a );
 a17352a <=( (not A267)  and  A266 );
 a17356a <=( A300  and  A299 );
 a17357a <=( (not A268)  and  a17356a );
 a17358a <=( a17357a  and  a17352a );
 a17361a <=( (not A167)  and  (not A168) );
 a17365a <=( A265  and  A201 );
 a17366a <=( A200  and  a17365a );
 a17367a <=( a17366a  and  a17361a );
 a17370a <=( (not A267)  and  A266 );
 a17374a <=( A300  and  A298 );
 a17375a <=( (not A268)  and  a17374a );
 a17376a <=( a17375a  and  a17370a );
 a17379a <=( (not A167)  and  (not A168) );
 a17383a <=( A265  and  A201 );
 a17384a <=( A200  and  a17383a );
 a17385a <=( a17384a  and  a17379a );
 a17388a <=( (not A267)  and  A266 );
 a17392a <=( A300  and  A299 );
 a17393a <=( A269  and  a17392a );
 a17394a <=( a17393a  and  a17388a );
 a17397a <=( (not A167)  and  (not A168) );
 a17401a <=( A265  and  A201 );
 a17402a <=( A200  and  a17401a );
 a17403a <=( a17402a  and  a17397a );
 a17406a <=( (not A267)  and  A266 );
 a17410a <=( A300  and  A298 );
 a17411a <=( A269  and  a17410a );
 a17412a <=( a17411a  and  a17406a );
 a17415a <=( (not A167)  and  (not A168) );
 a17419a <=( (not A265)  and  A201 );
 a17420a <=( A200  and  a17419a );
 a17421a <=( a17420a  and  a17415a );
 a17424a <=( (not A267)  and  A266 );
 a17428a <=( A300  and  A299 );
 a17429a <=( A268  and  a17428a );
 a17430a <=( a17429a  and  a17424a );
 a17433a <=( (not A167)  and  (not A168) );
 a17437a <=( (not A265)  and  A201 );
 a17438a <=( A200  and  a17437a );
 a17439a <=( a17438a  and  a17433a );
 a17442a <=( (not A267)  and  A266 );
 a17446a <=( A300  and  A298 );
 a17447a <=( A268  and  a17446a );
 a17448a <=( a17447a  and  a17442a );
 a17451a <=( (not A167)  and  (not A168) );
 a17455a <=( (not A265)  and  A201 );
 a17456a <=( A200  and  a17455a );
 a17457a <=( a17456a  and  a17451a );
 a17460a <=( (not A267)  and  A266 );
 a17464a <=( A300  and  A299 );
 a17465a <=( (not A269)  and  a17464a );
 a17466a <=( a17465a  and  a17460a );
 a17469a <=( (not A167)  and  (not A168) );
 a17473a <=( (not A265)  and  A201 );
 a17474a <=( A200  and  a17473a );
 a17475a <=( a17474a  and  a17469a );
 a17478a <=( (not A267)  and  A266 );
 a17482a <=( A300  and  A298 );
 a17483a <=( (not A269)  and  a17482a );
 a17484a <=( a17483a  and  a17478a );
 a17487a <=( (not A167)  and  (not A168) );
 a17491a <=( A265  and  A201 );
 a17492a <=( A200  and  a17491a );
 a17493a <=( a17492a  and  a17487a );
 a17496a <=( (not A267)  and  (not A266) );
 a17500a <=( A300  and  A299 );
 a17501a <=( A268  and  a17500a );
 a17502a <=( a17501a  and  a17496a );
 a17505a <=( (not A167)  and  (not A168) );
 a17509a <=( A265  and  A201 );
 a17510a <=( A200  and  a17509a );
 a17511a <=( a17510a  and  a17505a );
 a17514a <=( (not A267)  and  (not A266) );
 a17518a <=( A300  and  A298 );
 a17519a <=( A268  and  a17518a );
 a17520a <=( a17519a  and  a17514a );
 a17523a <=( (not A167)  and  (not A168) );
 a17527a <=( A265  and  A201 );
 a17528a <=( A200  and  a17527a );
 a17529a <=( a17528a  and  a17523a );
 a17532a <=( (not A267)  and  (not A266) );
 a17536a <=( A300  and  A299 );
 a17537a <=( (not A269)  and  a17536a );
 a17538a <=( a17537a  and  a17532a );
 a17541a <=( (not A167)  and  (not A168) );
 a17545a <=( A265  and  A201 );
 a17546a <=( A200  and  a17545a );
 a17547a <=( a17546a  and  a17541a );
 a17550a <=( (not A267)  and  (not A266) );
 a17554a <=( A300  and  A298 );
 a17555a <=( (not A269)  and  a17554a );
 a17556a <=( a17555a  and  a17550a );
 a17559a <=( (not A167)  and  (not A168) );
 a17563a <=( (not A202)  and  (not A200) );
 a17564a <=( (not A199)  and  a17563a );
 a17565a <=( a17564a  and  a17559a );
 a17568a <=( A267  and  A265 );
 a17572a <=( (not A301)  and  (not A299) );
 a17573a <=( (not A298)  and  a17572a );
 a17574a <=( a17573a  and  a17568a );
 a17577a <=( (not A167)  and  (not A168) );
 a17581a <=( (not A202)  and  (not A200) );
 a17582a <=( (not A199)  and  a17581a );
 a17583a <=( a17582a  and  a17577a );
 a17586a <=( A267  and  A265 );
 a17590a <=( A302  and  (not A299) );
 a17591a <=( (not A298)  and  a17590a );
 a17592a <=( a17591a  and  a17586a );
 a17595a <=( (not A167)  and  (not A168) );
 a17599a <=( (not A202)  and  (not A200) );
 a17600a <=( (not A199)  and  a17599a );
 a17601a <=( a17600a  and  a17595a );
 a17604a <=( A267  and  A266 );
 a17608a <=( (not A301)  and  (not A299) );
 a17609a <=( (not A298)  and  a17608a );
 a17610a <=( a17609a  and  a17604a );
 a17613a <=( (not A167)  and  (not A168) );
 a17617a <=( (not A202)  and  (not A200) );
 a17618a <=( (not A199)  and  a17617a );
 a17619a <=( a17618a  and  a17613a );
 a17622a <=( A267  and  A266 );
 a17626a <=( A302  and  (not A299) );
 a17627a <=( (not A298)  and  a17626a );
 a17628a <=( a17627a  and  a17622a );
 a17631a <=( (not A167)  and  (not A168) );
 a17635a <=( A203  and  (not A200) );
 a17636a <=( (not A199)  and  a17635a );
 a17637a <=( a17636a  and  a17631a );
 a17640a <=( A267  and  A265 );
 a17644a <=( (not A301)  and  (not A299) );
 a17645a <=( (not A298)  and  a17644a );
 a17646a <=( a17645a  and  a17640a );
 a17649a <=( (not A167)  and  (not A168) );
 a17653a <=( A203  and  (not A200) );
 a17654a <=( (not A199)  and  a17653a );
 a17655a <=( a17654a  and  a17649a );
 a17658a <=( A267  and  A265 );
 a17662a <=( A302  and  (not A299) );
 a17663a <=( (not A298)  and  a17662a );
 a17664a <=( a17663a  and  a17658a );
 a17667a <=( (not A167)  and  (not A168) );
 a17671a <=( A203  and  (not A200) );
 a17672a <=( (not A199)  and  a17671a );
 a17673a <=( a17672a  and  a17667a );
 a17676a <=( A267  and  A266 );
 a17680a <=( (not A301)  and  (not A299) );
 a17681a <=( (not A298)  and  a17680a );
 a17682a <=( a17681a  and  a17676a );
 a17685a <=( (not A167)  and  (not A168) );
 a17689a <=( A203  and  (not A200) );
 a17690a <=( (not A199)  and  a17689a );
 a17691a <=( a17690a  and  a17685a );
 a17694a <=( A267  and  A266 );
 a17698a <=( A302  and  (not A299) );
 a17699a <=( (not A298)  and  a17698a );
 a17700a <=( a17699a  and  a17694a );
 a17703a <=( (not A169)  and  (not A170) );
 a17707a <=( A201  and  A199 );
 a17708a <=( (not A167)  and  a17707a );
 a17709a <=( a17708a  and  a17703a );
 a17712a <=( (not A266)  and  (not A265) );
 a17716a <=( A300  and  A299 );
 a17717a <=( (not A268)  and  a17716a );
 a17718a <=( a17717a  and  a17712a );
 a17721a <=( (not A169)  and  (not A170) );
 a17725a <=( A201  and  A199 );
 a17726a <=( (not A167)  and  a17725a );
 a17727a <=( a17726a  and  a17721a );
 a17730a <=( (not A266)  and  (not A265) );
 a17734a <=( A300  and  A298 );
 a17735a <=( (not A268)  and  a17734a );
 a17736a <=( a17735a  and  a17730a );
 a17739a <=( (not A169)  and  (not A170) );
 a17743a <=( A201  and  A199 );
 a17744a <=( (not A167)  and  a17743a );
 a17745a <=( a17744a  and  a17739a );
 a17748a <=( (not A266)  and  (not A265) );
 a17752a <=( A300  and  A299 );
 a17753a <=( A269  and  a17752a );
 a17754a <=( a17753a  and  a17748a );
 a17757a <=( (not A169)  and  (not A170) );
 a17761a <=( A201  and  A199 );
 a17762a <=( (not A167)  and  a17761a );
 a17763a <=( a17762a  and  a17757a );
 a17766a <=( (not A266)  and  (not A265) );
 a17770a <=( A300  and  A298 );
 a17771a <=( A269  and  a17770a );
 a17772a <=( a17771a  and  a17766a );
 a17775a <=( (not A169)  and  (not A170) );
 a17779a <=( A201  and  A200 );
 a17780a <=( (not A167)  and  a17779a );
 a17781a <=( a17780a  and  a17775a );
 a17784a <=( (not A266)  and  (not A265) );
 a17788a <=( A300  and  A299 );
 a17789a <=( (not A268)  and  a17788a );
 a17790a <=( a17789a  and  a17784a );
 a17793a <=( (not A169)  and  (not A170) );
 a17797a <=( A201  and  A200 );
 a17798a <=( (not A167)  and  a17797a );
 a17799a <=( a17798a  and  a17793a );
 a17802a <=( (not A266)  and  (not A265) );
 a17806a <=( A300  and  A298 );
 a17807a <=( (not A268)  and  a17806a );
 a17808a <=( a17807a  and  a17802a );
 a17811a <=( (not A169)  and  (not A170) );
 a17815a <=( A201  and  A200 );
 a17816a <=( (not A167)  and  a17815a );
 a17817a <=( a17816a  and  a17811a );
 a17820a <=( (not A266)  and  (not A265) );
 a17824a <=( A300  and  A299 );
 a17825a <=( A269  and  a17824a );
 a17826a <=( a17825a  and  a17820a );
 a17829a <=( (not A169)  and  (not A170) );
 a17833a <=( A201  and  A200 );
 a17834a <=( (not A167)  and  a17833a );
 a17835a <=( a17834a  and  a17829a );
 a17838a <=( (not A266)  and  (not A265) );
 a17842a <=( A300  and  A298 );
 a17843a <=( A269  and  a17842a );
 a17844a <=( a17843a  and  a17838a );
 a17847a <=( A166  and  A167 );
 a17851a <=( (not A265)  and  A201 );
 a17852a <=( A199  and  a17851a );
 a17853a <=( a17852a  and  a17847a );
 a17857a <=( A298  and  (not A268) );
 a17858a <=( (not A266)  and  a17857a );
 a17862a <=( (not A302)  and  A301 );
 a17863a <=( A299  and  a17862a );
 a17864a <=( a17863a  and  a17858a );
 a17867a <=( A166  and  A167 );
 a17871a <=( (not A265)  and  A201 );
 a17872a <=( A199  and  a17871a );
 a17873a <=( a17872a  and  a17867a );
 a17877a <=( A298  and  (not A268) );
 a17878a <=( (not A266)  and  a17877a );
 a17882a <=( A302  and  (not A301) );
 a17883a <=( (not A299)  and  a17882a );
 a17884a <=( a17883a  and  a17878a );
 a17887a <=( A166  and  A167 );
 a17891a <=( (not A265)  and  A201 );
 a17892a <=( A199  and  a17891a );
 a17893a <=( a17892a  and  a17887a );
 a17897a <=( (not A298)  and  (not A268) );
 a17898a <=( (not A266)  and  a17897a );
 a17902a <=( A302  and  (not A301) );
 a17903a <=( A299  and  a17902a );
 a17904a <=( a17903a  and  a17898a );
 a17907a <=( A166  and  A167 );
 a17911a <=( (not A265)  and  A201 );
 a17912a <=( A199  and  a17911a );
 a17913a <=( a17912a  and  a17907a );
 a17917a <=( (not A298)  and  (not A268) );
 a17918a <=( (not A266)  and  a17917a );
 a17922a <=( (not A302)  and  A301 );
 a17923a <=( (not A299)  and  a17922a );
 a17924a <=( a17923a  and  a17918a );
 a17927a <=( A166  and  A167 );
 a17931a <=( (not A265)  and  A201 );
 a17932a <=( A199  and  a17931a );
 a17933a <=( a17932a  and  a17927a );
 a17937a <=( A298  and  A269 );
 a17938a <=( (not A266)  and  a17937a );
 a17942a <=( (not A302)  and  A301 );
 a17943a <=( A299  and  a17942a );
 a17944a <=( a17943a  and  a17938a );
 a17947a <=( A166  and  A167 );
 a17951a <=( (not A265)  and  A201 );
 a17952a <=( A199  and  a17951a );
 a17953a <=( a17952a  and  a17947a );
 a17957a <=( A298  and  A269 );
 a17958a <=( (not A266)  and  a17957a );
 a17962a <=( A302  and  (not A301) );
 a17963a <=( (not A299)  and  a17962a );
 a17964a <=( a17963a  and  a17958a );
 a17967a <=( A166  and  A167 );
 a17971a <=( (not A265)  and  A201 );
 a17972a <=( A199  and  a17971a );
 a17973a <=( a17972a  and  a17967a );
 a17977a <=( (not A298)  and  A269 );
 a17978a <=( (not A266)  and  a17977a );
 a17982a <=( A302  and  (not A301) );
 a17983a <=( A299  and  a17982a );
 a17984a <=( a17983a  and  a17978a );
 a17987a <=( A166  and  A167 );
 a17991a <=( (not A265)  and  A201 );
 a17992a <=( A199  and  a17991a );
 a17993a <=( a17992a  and  a17987a );
 a17997a <=( (not A298)  and  A269 );
 a17998a <=( (not A266)  and  a17997a );
 a18002a <=( (not A302)  and  A301 );
 a18003a <=( (not A299)  and  a18002a );
 a18004a <=( a18003a  and  a17998a );
 a18007a <=( A166  and  A167 );
 a18011a <=( (not A265)  and  A201 );
 a18012a <=( A200  and  a18011a );
 a18013a <=( a18012a  and  a18007a );
 a18017a <=( A298  and  (not A268) );
 a18018a <=( (not A266)  and  a18017a );
 a18022a <=( (not A302)  and  A301 );
 a18023a <=( A299  and  a18022a );
 a18024a <=( a18023a  and  a18018a );
 a18027a <=( A166  and  A167 );
 a18031a <=( (not A265)  and  A201 );
 a18032a <=( A200  and  a18031a );
 a18033a <=( a18032a  and  a18027a );
 a18037a <=( A298  and  (not A268) );
 a18038a <=( (not A266)  and  a18037a );
 a18042a <=( A302  and  (not A301) );
 a18043a <=( (not A299)  and  a18042a );
 a18044a <=( a18043a  and  a18038a );
 a18047a <=( A166  and  A167 );
 a18051a <=( (not A265)  and  A201 );
 a18052a <=( A200  and  a18051a );
 a18053a <=( a18052a  and  a18047a );
 a18057a <=( (not A298)  and  (not A268) );
 a18058a <=( (not A266)  and  a18057a );
 a18062a <=( A302  and  (not A301) );
 a18063a <=( A299  and  a18062a );
 a18064a <=( a18063a  and  a18058a );
 a18067a <=( A166  and  A167 );
 a18071a <=( (not A265)  and  A201 );
 a18072a <=( A200  and  a18071a );
 a18073a <=( a18072a  and  a18067a );
 a18077a <=( (not A298)  and  (not A268) );
 a18078a <=( (not A266)  and  a18077a );
 a18082a <=( (not A302)  and  A301 );
 a18083a <=( (not A299)  and  a18082a );
 a18084a <=( a18083a  and  a18078a );
 a18087a <=( A166  and  A167 );
 a18091a <=( (not A265)  and  A201 );
 a18092a <=( A200  and  a18091a );
 a18093a <=( a18092a  and  a18087a );
 a18097a <=( A298  and  A269 );
 a18098a <=( (not A266)  and  a18097a );
 a18102a <=( (not A302)  and  A301 );
 a18103a <=( A299  and  a18102a );
 a18104a <=( a18103a  and  a18098a );
 a18107a <=( A166  and  A167 );
 a18111a <=( (not A265)  and  A201 );
 a18112a <=( A200  and  a18111a );
 a18113a <=( a18112a  and  a18107a );
 a18117a <=( A298  and  A269 );
 a18118a <=( (not A266)  and  a18117a );
 a18122a <=( A302  and  (not A301) );
 a18123a <=( (not A299)  and  a18122a );
 a18124a <=( a18123a  and  a18118a );
 a18127a <=( A166  and  A167 );
 a18131a <=( (not A265)  and  A201 );
 a18132a <=( A200  and  a18131a );
 a18133a <=( a18132a  and  a18127a );
 a18137a <=( (not A298)  and  A269 );
 a18138a <=( (not A266)  and  a18137a );
 a18142a <=( A302  and  (not A301) );
 a18143a <=( A299  and  a18142a );
 a18144a <=( a18143a  and  a18138a );
 a18147a <=( A166  and  A167 );
 a18151a <=( (not A265)  and  A201 );
 a18152a <=( A200  and  a18151a );
 a18153a <=( a18152a  and  a18147a );
 a18157a <=( (not A298)  and  A269 );
 a18158a <=( (not A266)  and  a18157a );
 a18162a <=( (not A302)  and  A301 );
 a18163a <=( (not A299)  and  a18162a );
 a18164a <=( a18163a  and  a18158a );
 a18167a <=( A166  and  A167 );
 a18171a <=( A202  and  A200 );
 a18172a <=( A199  and  a18171a );
 a18173a <=( a18172a  and  a18167a );
 a18177a <=( (not A266)  and  (not A265) );
 a18178a <=( (not A203)  and  a18177a );
 a18182a <=( A300  and  A299 );
 a18183a <=( (not A268)  and  a18182a );
 a18184a <=( a18183a  and  a18178a );
 a18187a <=( A166  and  A167 );
 a18191a <=( A202  and  A200 );
 a18192a <=( A199  and  a18191a );
 a18193a <=( a18192a  and  a18187a );
 a18197a <=( (not A266)  and  (not A265) );
 a18198a <=( (not A203)  and  a18197a );
 a18202a <=( A300  and  A298 );
 a18203a <=( (not A268)  and  a18202a );
 a18204a <=( a18203a  and  a18198a );
 a18207a <=( A166  and  A167 );
 a18211a <=( A202  and  A200 );
 a18212a <=( A199  and  a18211a );
 a18213a <=( a18212a  and  a18207a );
 a18217a <=( (not A266)  and  (not A265) );
 a18218a <=( (not A203)  and  a18217a );
 a18222a <=( A300  and  A299 );
 a18223a <=( A269  and  a18222a );
 a18224a <=( a18223a  and  a18218a );
 a18227a <=( A166  and  A167 );
 a18231a <=( A202  and  A200 );
 a18232a <=( A199  and  a18231a );
 a18233a <=( a18232a  and  a18227a );
 a18237a <=( (not A266)  and  (not A265) );
 a18238a <=( (not A203)  and  a18237a );
 a18242a <=( A300  and  A298 );
 a18243a <=( A269  and  a18242a );
 a18244a <=( a18243a  and  a18238a );
 a18247a <=( A166  and  A167 );
 a18251a <=( (not A201)  and  A200 );
 a18252a <=( A199  and  a18251a );
 a18253a <=( a18252a  and  a18247a );
 a18257a <=( A267  and  A265 );
 a18258a <=( (not A202)  and  a18257a );
 a18262a <=( (not A301)  and  (not A299) );
 a18263a <=( (not A298)  and  a18262a );
 a18264a <=( a18263a  and  a18258a );
 a18267a <=( A166  and  A167 );
 a18271a <=( (not A201)  and  A200 );
 a18272a <=( A199  and  a18271a );
 a18273a <=( a18272a  and  a18267a );
 a18277a <=( A267  and  A265 );
 a18278a <=( (not A202)  and  a18277a );
 a18282a <=( A302  and  (not A299) );
 a18283a <=( (not A298)  and  a18282a );
 a18284a <=( a18283a  and  a18278a );
 a18287a <=( A166  and  A167 );
 a18291a <=( (not A201)  and  A200 );
 a18292a <=( A199  and  a18291a );
 a18293a <=( a18292a  and  a18287a );
 a18297a <=( A267  and  A266 );
 a18298a <=( (not A202)  and  a18297a );
 a18302a <=( (not A301)  and  (not A299) );
 a18303a <=( (not A298)  and  a18302a );
 a18304a <=( a18303a  and  a18298a );
 a18307a <=( A166  and  A167 );
 a18311a <=( (not A201)  and  A200 );
 a18312a <=( A199  and  a18311a );
 a18313a <=( a18312a  and  a18307a );
 a18317a <=( A267  and  A266 );
 a18318a <=( (not A202)  and  a18317a );
 a18322a <=( A302  and  (not A299) );
 a18323a <=( (not A298)  and  a18322a );
 a18324a <=( a18323a  and  a18318a );
 a18327a <=( A166  and  A167 );
 a18331a <=( (not A201)  and  A200 );
 a18332a <=( A199  and  a18331a );
 a18333a <=( a18332a  and  a18327a );
 a18337a <=( A267  and  A265 );
 a18338a <=( A203  and  a18337a );
 a18342a <=( (not A301)  and  (not A299) );
 a18343a <=( (not A298)  and  a18342a );
 a18344a <=( a18343a  and  a18338a );
 a18347a <=( A166  and  A167 );
 a18351a <=( (not A201)  and  A200 );
 a18352a <=( A199  and  a18351a );
 a18353a <=( a18352a  and  a18347a );
 a18357a <=( A267  and  A265 );
 a18358a <=( A203  and  a18357a );
 a18362a <=( A302  and  (not A299) );
 a18363a <=( (not A298)  and  a18362a );
 a18364a <=( a18363a  and  a18358a );
 a18367a <=( A166  and  A167 );
 a18371a <=( (not A201)  and  A200 );
 a18372a <=( A199  and  a18371a );
 a18373a <=( a18372a  and  a18367a );
 a18377a <=( A267  and  A266 );
 a18378a <=( A203  and  a18377a );
 a18382a <=( (not A301)  and  (not A299) );
 a18383a <=( (not A298)  and  a18382a );
 a18384a <=( a18383a  and  a18378a );
 a18387a <=( A166  and  A167 );
 a18391a <=( (not A201)  and  A200 );
 a18392a <=( A199  and  a18391a );
 a18393a <=( a18392a  and  a18387a );
 a18397a <=( A267  and  A266 );
 a18398a <=( A203  and  a18397a );
 a18402a <=( A302  and  (not A299) );
 a18403a <=( (not A298)  and  a18402a );
 a18404a <=( a18403a  and  a18398a );
 a18407a <=( A166  and  A167 );
 a18411a <=( (not A202)  and  A200 );
 a18412a <=( (not A199)  and  a18411a );
 a18413a <=( a18412a  and  a18407a );
 a18417a <=( (not A266)  and  (not A265) );
 a18418a <=( A203  and  a18417a );
 a18422a <=( A300  and  A299 );
 a18423a <=( (not A268)  and  a18422a );
 a18424a <=( a18423a  and  a18418a );
 a18427a <=( A166  and  A167 );
 a18431a <=( (not A202)  and  A200 );
 a18432a <=( (not A199)  and  a18431a );
 a18433a <=( a18432a  and  a18427a );
 a18437a <=( (not A266)  and  (not A265) );
 a18438a <=( A203  and  a18437a );
 a18442a <=( A300  and  A298 );
 a18443a <=( (not A268)  and  a18442a );
 a18444a <=( a18443a  and  a18438a );
 a18447a <=( A166  and  A167 );
 a18451a <=( (not A202)  and  A200 );
 a18452a <=( (not A199)  and  a18451a );
 a18453a <=( a18452a  and  a18447a );
 a18457a <=( (not A266)  and  (not A265) );
 a18458a <=( A203  and  a18457a );
 a18462a <=( A300  and  A299 );
 a18463a <=( A269  and  a18462a );
 a18464a <=( a18463a  and  a18458a );
 a18467a <=( A166  and  A167 );
 a18471a <=( (not A202)  and  A200 );
 a18472a <=( (not A199)  and  a18471a );
 a18473a <=( a18472a  and  a18467a );
 a18477a <=( (not A266)  and  (not A265) );
 a18478a <=( A203  and  a18477a );
 a18482a <=( A300  and  A298 );
 a18483a <=( A269  and  a18482a );
 a18484a <=( a18483a  and  a18478a );
 a18487a <=( A166  and  A167 );
 a18491a <=( (not A201)  and  A200 );
 a18492a <=( (not A199)  and  a18491a );
 a18493a <=( a18492a  and  a18487a );
 a18497a <=( A267  and  A265 );
 a18498a <=( A202  and  a18497a );
 a18502a <=( (not A301)  and  (not A299) );
 a18503a <=( (not A298)  and  a18502a );
 a18504a <=( a18503a  and  a18498a );
 a18507a <=( A166  and  A167 );
 a18511a <=( (not A201)  and  A200 );
 a18512a <=( (not A199)  and  a18511a );
 a18513a <=( a18512a  and  a18507a );
 a18517a <=( A267  and  A265 );
 a18518a <=( A202  and  a18517a );
 a18522a <=( A302  and  (not A299) );
 a18523a <=( (not A298)  and  a18522a );
 a18524a <=( a18523a  and  a18518a );
 a18527a <=( A166  and  A167 );
 a18531a <=( (not A201)  and  A200 );
 a18532a <=( (not A199)  and  a18531a );
 a18533a <=( a18532a  and  a18527a );
 a18537a <=( A267  and  A266 );
 a18538a <=( A202  and  a18537a );
 a18542a <=( (not A301)  and  (not A299) );
 a18543a <=( (not A298)  and  a18542a );
 a18544a <=( a18543a  and  a18538a );
 a18547a <=( A166  and  A167 );
 a18551a <=( (not A201)  and  A200 );
 a18552a <=( (not A199)  and  a18551a );
 a18553a <=( a18552a  and  a18547a );
 a18557a <=( A267  and  A266 );
 a18558a <=( A202  and  a18557a );
 a18562a <=( A302  and  (not A299) );
 a18563a <=( (not A298)  and  a18562a );
 a18564a <=( a18563a  and  a18558a );
 a18567a <=( A166  and  A167 );
 a18571a <=( (not A201)  and  A200 );
 a18572a <=( (not A199)  and  a18571a );
 a18573a <=( a18572a  and  a18567a );
 a18577a <=( A267  and  A265 );
 a18578a <=( (not A203)  and  a18577a );
 a18582a <=( (not A301)  and  (not A299) );
 a18583a <=( (not A298)  and  a18582a );
 a18584a <=( a18583a  and  a18578a );
 a18587a <=( A166  and  A167 );
 a18591a <=( (not A201)  and  A200 );
 a18592a <=( (not A199)  and  a18591a );
 a18593a <=( a18592a  and  a18587a );
 a18597a <=( A267  and  A265 );
 a18598a <=( (not A203)  and  a18597a );
 a18602a <=( A302  and  (not A299) );
 a18603a <=( (not A298)  and  a18602a );
 a18604a <=( a18603a  and  a18598a );
 a18607a <=( A166  and  A167 );
 a18611a <=( (not A201)  and  A200 );
 a18612a <=( (not A199)  and  a18611a );
 a18613a <=( a18612a  and  a18607a );
 a18617a <=( A267  and  A266 );
 a18618a <=( (not A203)  and  a18617a );
 a18622a <=( (not A301)  and  (not A299) );
 a18623a <=( (not A298)  and  a18622a );
 a18624a <=( a18623a  and  a18618a );
 a18627a <=( A166  and  A167 );
 a18631a <=( (not A201)  and  A200 );
 a18632a <=( (not A199)  and  a18631a );
 a18633a <=( a18632a  and  a18627a );
 a18637a <=( A267  and  A266 );
 a18638a <=( (not A203)  and  a18637a );
 a18642a <=( A302  and  (not A299) );
 a18643a <=( (not A298)  and  a18642a );
 a18644a <=( a18643a  and  a18638a );
 a18647a <=( A166  and  A167 );
 a18651a <=( (not A202)  and  (not A200) );
 a18652a <=( A199  and  a18651a );
 a18653a <=( a18652a  and  a18647a );
 a18657a <=( (not A266)  and  (not A265) );
 a18658a <=( A203  and  a18657a );
 a18662a <=( A300  and  A299 );
 a18663a <=( (not A268)  and  a18662a );
 a18664a <=( a18663a  and  a18658a );
 a18667a <=( A166  and  A167 );
 a18671a <=( (not A202)  and  (not A200) );
 a18672a <=( A199  and  a18671a );
 a18673a <=( a18672a  and  a18667a );
 a18677a <=( (not A266)  and  (not A265) );
 a18678a <=( A203  and  a18677a );
 a18682a <=( A300  and  A298 );
 a18683a <=( (not A268)  and  a18682a );
 a18684a <=( a18683a  and  a18678a );
 a18687a <=( A166  and  A167 );
 a18691a <=( (not A202)  and  (not A200) );
 a18692a <=( A199  and  a18691a );
 a18693a <=( a18692a  and  a18687a );
 a18697a <=( (not A266)  and  (not A265) );
 a18698a <=( A203  and  a18697a );
 a18702a <=( A300  and  A299 );
 a18703a <=( A269  and  a18702a );
 a18704a <=( a18703a  and  a18698a );
 a18707a <=( A166  and  A167 );
 a18711a <=( (not A202)  and  (not A200) );
 a18712a <=( A199  and  a18711a );
 a18713a <=( a18712a  and  a18707a );
 a18717a <=( (not A266)  and  (not A265) );
 a18718a <=( A203  and  a18717a );
 a18722a <=( A300  and  A298 );
 a18723a <=( A269  and  a18722a );
 a18724a <=( a18723a  and  a18718a );
 a18727a <=( A166  and  A167 );
 a18731a <=( (not A201)  and  (not A200) );
 a18732a <=( A199  and  a18731a );
 a18733a <=( a18732a  and  a18727a );
 a18737a <=( A267  and  A265 );
 a18738a <=( A202  and  a18737a );
 a18742a <=( (not A301)  and  (not A299) );
 a18743a <=( (not A298)  and  a18742a );
 a18744a <=( a18743a  and  a18738a );
 a18747a <=( A166  and  A167 );
 a18751a <=( (not A201)  and  (not A200) );
 a18752a <=( A199  and  a18751a );
 a18753a <=( a18752a  and  a18747a );
 a18757a <=( A267  and  A265 );
 a18758a <=( A202  and  a18757a );
 a18762a <=( A302  and  (not A299) );
 a18763a <=( (not A298)  and  a18762a );
 a18764a <=( a18763a  and  a18758a );
 a18767a <=( A166  and  A167 );
 a18771a <=( (not A201)  and  (not A200) );
 a18772a <=( A199  and  a18771a );
 a18773a <=( a18772a  and  a18767a );
 a18777a <=( A267  and  A266 );
 a18778a <=( A202  and  a18777a );
 a18782a <=( (not A301)  and  (not A299) );
 a18783a <=( (not A298)  and  a18782a );
 a18784a <=( a18783a  and  a18778a );
 a18787a <=( A166  and  A167 );
 a18791a <=( (not A201)  and  (not A200) );
 a18792a <=( A199  and  a18791a );
 a18793a <=( a18792a  and  a18787a );
 a18797a <=( A267  and  A266 );
 a18798a <=( A202  and  a18797a );
 a18802a <=( A302  and  (not A299) );
 a18803a <=( (not A298)  and  a18802a );
 a18804a <=( a18803a  and  a18798a );
 a18807a <=( A166  and  A167 );
 a18811a <=( (not A201)  and  (not A200) );
 a18812a <=( A199  and  a18811a );
 a18813a <=( a18812a  and  a18807a );
 a18817a <=( A267  and  A265 );
 a18818a <=( (not A203)  and  a18817a );
 a18822a <=( (not A301)  and  (not A299) );
 a18823a <=( (not A298)  and  a18822a );
 a18824a <=( a18823a  and  a18818a );
 a18827a <=( A166  and  A167 );
 a18831a <=( (not A201)  and  (not A200) );
 a18832a <=( A199  and  a18831a );
 a18833a <=( a18832a  and  a18827a );
 a18837a <=( A267  and  A265 );
 a18838a <=( (not A203)  and  a18837a );
 a18842a <=( A302  and  (not A299) );
 a18843a <=( (not A298)  and  a18842a );
 a18844a <=( a18843a  and  a18838a );
 a18847a <=( A166  and  A167 );
 a18851a <=( (not A201)  and  (not A200) );
 a18852a <=( A199  and  a18851a );
 a18853a <=( a18852a  and  a18847a );
 a18857a <=( A267  and  A266 );
 a18858a <=( (not A203)  and  a18857a );
 a18862a <=( (not A301)  and  (not A299) );
 a18863a <=( (not A298)  and  a18862a );
 a18864a <=( a18863a  and  a18858a );
 a18867a <=( A166  and  A167 );
 a18871a <=( (not A201)  and  (not A200) );
 a18872a <=( A199  and  a18871a );
 a18873a <=( a18872a  and  a18867a );
 a18877a <=( A267  and  A266 );
 a18878a <=( (not A203)  and  a18877a );
 a18882a <=( A302  and  (not A299) );
 a18883a <=( (not A298)  and  a18882a );
 a18884a <=( a18883a  and  a18878a );
 a18887a <=( A166  and  A167 );
 a18891a <=( (not A202)  and  (not A200) );
 a18892a <=( (not A199)  and  a18891a );
 a18893a <=( a18892a  and  a18887a );
 a18897a <=( A298  and  A267 );
 a18898a <=( A265  and  a18897a );
 a18902a <=( (not A301)  and  (not A300) );
 a18903a <=( A299  and  a18902a );
 a18904a <=( a18903a  and  a18898a );
 a18907a <=( A166  and  A167 );
 a18911a <=( (not A202)  and  (not A200) );
 a18912a <=( (not A199)  and  a18911a );
 a18913a <=( a18912a  and  a18907a );
 a18917a <=( A298  and  A267 );
 a18918a <=( A265  and  a18917a );
 a18922a <=( A302  and  (not A300) );
 a18923a <=( A299  and  a18922a );
 a18924a <=( a18923a  and  a18918a );
 a18927a <=( A166  and  A167 );
 a18931a <=( (not A202)  and  (not A200) );
 a18932a <=( (not A199)  and  a18931a );
 a18933a <=( a18932a  and  a18927a );
 a18937a <=( A298  and  A267 );
 a18938a <=( A265  and  a18937a );
 a18942a <=( A301  and  (not A300) );
 a18943a <=( (not A299)  and  a18942a );
 a18944a <=( a18943a  and  a18938a );
 a18947a <=( A166  and  A167 );
 a18951a <=( (not A202)  and  (not A200) );
 a18952a <=( (not A199)  and  a18951a );
 a18953a <=( a18952a  and  a18947a );
 a18957a <=( A298  and  A267 );
 a18958a <=( A265  and  a18957a );
 a18962a <=( (not A302)  and  (not A300) );
 a18963a <=( (not A299)  and  a18962a );
 a18964a <=( a18963a  and  a18958a );
 a18967a <=( A166  and  A167 );
 a18971a <=( (not A202)  and  (not A200) );
 a18972a <=( (not A199)  and  a18971a );
 a18973a <=( a18972a  and  a18967a );
 a18977a <=( (not A298)  and  A267 );
 a18978a <=( A265  and  a18977a );
 a18982a <=( A301  and  (not A300) );
 a18983a <=( A299  and  a18982a );
 a18984a <=( a18983a  and  a18978a );
 a18987a <=( A166  and  A167 );
 a18991a <=( (not A202)  and  (not A200) );
 a18992a <=( (not A199)  and  a18991a );
 a18993a <=( a18992a  and  a18987a );
 a18997a <=( (not A298)  and  A267 );
 a18998a <=( A265  and  a18997a );
 a19002a <=( (not A302)  and  (not A300) );
 a19003a <=( A299  and  a19002a );
 a19004a <=( a19003a  and  a18998a );
 a19007a <=( A166  and  A167 );
 a19011a <=( (not A202)  and  (not A200) );
 a19012a <=( (not A199)  and  a19011a );
 a19013a <=( a19012a  and  a19007a );
 a19017a <=( A298  and  A267 );
 a19018a <=( A266  and  a19017a );
 a19022a <=( (not A301)  and  (not A300) );
 a19023a <=( A299  and  a19022a );
 a19024a <=( a19023a  and  a19018a );
 a19027a <=( A166  and  A167 );
 a19031a <=( (not A202)  and  (not A200) );
 a19032a <=( (not A199)  and  a19031a );
 a19033a <=( a19032a  and  a19027a );
 a19037a <=( A298  and  A267 );
 a19038a <=( A266  and  a19037a );
 a19042a <=( A302  and  (not A300) );
 a19043a <=( A299  and  a19042a );
 a19044a <=( a19043a  and  a19038a );
 a19047a <=( A166  and  A167 );
 a19051a <=( (not A202)  and  (not A200) );
 a19052a <=( (not A199)  and  a19051a );
 a19053a <=( a19052a  and  a19047a );
 a19057a <=( A298  and  A267 );
 a19058a <=( A266  and  a19057a );
 a19062a <=( A301  and  (not A300) );
 a19063a <=( (not A299)  and  a19062a );
 a19064a <=( a19063a  and  a19058a );
 a19067a <=( A166  and  A167 );
 a19071a <=( (not A202)  and  (not A200) );
 a19072a <=( (not A199)  and  a19071a );
 a19073a <=( a19072a  and  a19067a );
 a19077a <=( A298  and  A267 );
 a19078a <=( A266  and  a19077a );
 a19082a <=( (not A302)  and  (not A300) );
 a19083a <=( (not A299)  and  a19082a );
 a19084a <=( a19083a  and  a19078a );
 a19087a <=( A166  and  A167 );
 a19091a <=( (not A202)  and  (not A200) );
 a19092a <=( (not A199)  and  a19091a );
 a19093a <=( a19092a  and  a19087a );
 a19097a <=( (not A298)  and  A267 );
 a19098a <=( A266  and  a19097a );
 a19102a <=( A301  and  (not A300) );
 a19103a <=( A299  and  a19102a );
 a19104a <=( a19103a  and  a19098a );
 a19107a <=( A166  and  A167 );
 a19111a <=( (not A202)  and  (not A200) );
 a19112a <=( (not A199)  and  a19111a );
 a19113a <=( a19112a  and  a19107a );
 a19117a <=( (not A298)  and  A267 );
 a19118a <=( A266  and  a19117a );
 a19122a <=( (not A302)  and  (not A300) );
 a19123a <=( A299  and  a19122a );
 a19124a <=( a19123a  and  a19118a );
 a19127a <=( A166  and  A167 );
 a19131a <=( A203  and  (not A200) );
 a19132a <=( (not A199)  and  a19131a );
 a19133a <=( a19132a  and  a19127a );
 a19137a <=( A298  and  A267 );
 a19138a <=( A265  and  a19137a );
 a19142a <=( (not A301)  and  (not A300) );
 a19143a <=( A299  and  a19142a );
 a19144a <=( a19143a  and  a19138a );
 a19147a <=( A166  and  A167 );
 a19151a <=( A203  and  (not A200) );
 a19152a <=( (not A199)  and  a19151a );
 a19153a <=( a19152a  and  a19147a );
 a19157a <=( A298  and  A267 );
 a19158a <=( A265  and  a19157a );
 a19162a <=( A302  and  (not A300) );
 a19163a <=( A299  and  a19162a );
 a19164a <=( a19163a  and  a19158a );
 a19167a <=( A166  and  A167 );
 a19171a <=( A203  and  (not A200) );
 a19172a <=( (not A199)  and  a19171a );
 a19173a <=( a19172a  and  a19167a );
 a19177a <=( A298  and  A267 );
 a19178a <=( A265  and  a19177a );
 a19182a <=( A301  and  (not A300) );
 a19183a <=( (not A299)  and  a19182a );
 a19184a <=( a19183a  and  a19178a );
 a19187a <=( A166  and  A167 );
 a19191a <=( A203  and  (not A200) );
 a19192a <=( (not A199)  and  a19191a );
 a19193a <=( a19192a  and  a19187a );
 a19197a <=( A298  and  A267 );
 a19198a <=( A265  and  a19197a );
 a19202a <=( (not A302)  and  (not A300) );
 a19203a <=( (not A299)  and  a19202a );
 a19204a <=( a19203a  and  a19198a );
 a19207a <=( A166  and  A167 );
 a19211a <=( A203  and  (not A200) );
 a19212a <=( (not A199)  and  a19211a );
 a19213a <=( a19212a  and  a19207a );
 a19217a <=( (not A298)  and  A267 );
 a19218a <=( A265  and  a19217a );
 a19222a <=( A301  and  (not A300) );
 a19223a <=( A299  and  a19222a );
 a19224a <=( a19223a  and  a19218a );
 a19227a <=( A166  and  A167 );
 a19231a <=( A203  and  (not A200) );
 a19232a <=( (not A199)  and  a19231a );
 a19233a <=( a19232a  and  a19227a );
 a19237a <=( (not A298)  and  A267 );
 a19238a <=( A265  and  a19237a );
 a19242a <=( (not A302)  and  (not A300) );
 a19243a <=( A299  and  a19242a );
 a19244a <=( a19243a  and  a19238a );
 a19247a <=( A166  and  A167 );
 a19251a <=( A203  and  (not A200) );
 a19252a <=( (not A199)  and  a19251a );
 a19253a <=( a19252a  and  a19247a );
 a19257a <=( A298  and  A267 );
 a19258a <=( A266  and  a19257a );
 a19262a <=( (not A301)  and  (not A300) );
 a19263a <=( A299  and  a19262a );
 a19264a <=( a19263a  and  a19258a );
 a19267a <=( A166  and  A167 );
 a19271a <=( A203  and  (not A200) );
 a19272a <=( (not A199)  and  a19271a );
 a19273a <=( a19272a  and  a19267a );
 a19277a <=( A298  and  A267 );
 a19278a <=( A266  and  a19277a );
 a19282a <=( A302  and  (not A300) );
 a19283a <=( A299  and  a19282a );
 a19284a <=( a19283a  and  a19278a );
 a19287a <=( A166  and  A167 );
 a19291a <=( A203  and  (not A200) );
 a19292a <=( (not A199)  and  a19291a );
 a19293a <=( a19292a  and  a19287a );
 a19297a <=( A298  and  A267 );
 a19298a <=( A266  and  a19297a );
 a19302a <=( A301  and  (not A300) );
 a19303a <=( (not A299)  and  a19302a );
 a19304a <=( a19303a  and  a19298a );
 a19307a <=( A166  and  A167 );
 a19311a <=( A203  and  (not A200) );
 a19312a <=( (not A199)  and  a19311a );
 a19313a <=( a19312a  and  a19307a );
 a19317a <=( A298  and  A267 );
 a19318a <=( A266  and  a19317a );
 a19322a <=( (not A302)  and  (not A300) );
 a19323a <=( (not A299)  and  a19322a );
 a19324a <=( a19323a  and  a19318a );
 a19327a <=( A166  and  A167 );
 a19331a <=( A203  and  (not A200) );
 a19332a <=( (not A199)  and  a19331a );
 a19333a <=( a19332a  and  a19327a );
 a19337a <=( (not A298)  and  A267 );
 a19338a <=( A266  and  a19337a );
 a19342a <=( A301  and  (not A300) );
 a19343a <=( A299  and  a19342a );
 a19344a <=( a19343a  and  a19338a );
 a19347a <=( A166  and  A167 );
 a19351a <=( A203  and  (not A200) );
 a19352a <=( (not A199)  and  a19351a );
 a19353a <=( a19352a  and  a19347a );
 a19357a <=( (not A298)  and  A267 );
 a19358a <=( A266  and  a19357a );
 a19362a <=( (not A302)  and  (not A300) );
 a19363a <=( A299  and  a19362a );
 a19364a <=( a19363a  and  a19358a );
 a19367a <=( A166  and  A167 );
 a19371a <=( A202  and  (not A200) );
 a19372a <=( (not A199)  and  a19371a );
 a19373a <=( a19372a  and  a19367a );
 a19377a <=( (not A266)  and  (not A265) );
 a19378a <=( (not A203)  and  a19377a );
 a19382a <=( A300  and  A299 );
 a19383a <=( (not A268)  and  a19382a );
 a19384a <=( a19383a  and  a19378a );
 a19387a <=( A166  and  A167 );
 a19391a <=( A202  and  (not A200) );
 a19392a <=( (not A199)  and  a19391a );
 a19393a <=( a19392a  and  a19387a );
 a19397a <=( (not A266)  and  (not A265) );
 a19398a <=( (not A203)  and  a19397a );
 a19402a <=( A300  and  A298 );
 a19403a <=( (not A268)  and  a19402a );
 a19404a <=( a19403a  and  a19398a );
 a19407a <=( A166  and  A167 );
 a19411a <=( A202  and  (not A200) );
 a19412a <=( (not A199)  and  a19411a );
 a19413a <=( a19412a  and  a19407a );
 a19417a <=( (not A266)  and  (not A265) );
 a19418a <=( (not A203)  and  a19417a );
 a19422a <=( A300  and  A299 );
 a19423a <=( A269  and  a19422a );
 a19424a <=( a19423a  and  a19418a );
 a19427a <=( A166  and  A167 );
 a19431a <=( A202  and  (not A200) );
 a19432a <=( (not A199)  and  a19431a );
 a19433a <=( a19432a  and  a19427a );
 a19437a <=( (not A266)  and  (not A265) );
 a19438a <=( (not A203)  and  a19437a );
 a19442a <=( A300  and  A298 );
 a19443a <=( A269  and  a19442a );
 a19444a <=( a19443a  and  a19438a );
 a19447a <=( (not A166)  and  A167 );
 a19451a <=( A265  and  A201 );
 a19452a <=( A199  and  a19451a );
 a19453a <=( a19452a  and  a19447a );
 a19457a <=( (not A269)  and  A268 );
 a19458a <=( A266  and  a19457a );
 a19462a <=( (not A301)  and  (not A299) );
 a19463a <=( (not A298)  and  a19462a );
 a19464a <=( a19463a  and  a19458a );
 a19467a <=( (not A166)  and  A167 );
 a19471a <=( A265  and  A201 );
 a19472a <=( A199  and  a19471a );
 a19473a <=( a19472a  and  a19467a );
 a19477a <=( (not A269)  and  A268 );
 a19478a <=( A266  and  a19477a );
 a19482a <=( A302  and  (not A299) );
 a19483a <=( (not A298)  and  a19482a );
 a19484a <=( a19483a  and  a19478a );
 a19487a <=( (not A166)  and  A167 );
 a19491a <=( (not A265)  and  A201 );
 a19492a <=( A199  and  a19491a );
 a19493a <=( a19492a  and  a19487a );
 a19497a <=( A269  and  (not A268) );
 a19498a <=( A266  and  a19497a );
 a19502a <=( (not A301)  and  (not A299) );
 a19503a <=( (not A298)  and  a19502a );
 a19504a <=( a19503a  and  a19498a );
 a19507a <=( (not A166)  and  A167 );
 a19511a <=( (not A265)  and  A201 );
 a19512a <=( A199  and  a19511a );
 a19513a <=( a19512a  and  a19507a );
 a19517a <=( A269  and  (not A268) );
 a19518a <=( A266  and  a19517a );
 a19522a <=( A302  and  (not A299) );
 a19523a <=( (not A298)  and  a19522a );
 a19524a <=( a19523a  and  a19518a );
 a19527a <=( (not A166)  and  A167 );
 a19531a <=( A265  and  A201 );
 a19532a <=( A199  and  a19531a );
 a19533a <=( a19532a  and  a19527a );
 a19537a <=( A269  and  (not A268) );
 a19538a <=( (not A266)  and  a19537a );
 a19542a <=( (not A301)  and  (not A299) );
 a19543a <=( (not A298)  and  a19542a );
 a19544a <=( a19543a  and  a19538a );
 a19547a <=( (not A166)  and  A167 );
 a19551a <=( A265  and  A201 );
 a19552a <=( A199  and  a19551a );
 a19553a <=( a19552a  and  a19547a );
 a19557a <=( A269  and  (not A268) );
 a19558a <=( (not A266)  and  a19557a );
 a19562a <=( A302  and  (not A299) );
 a19563a <=( (not A298)  and  a19562a );
 a19564a <=( a19563a  and  a19558a );
 a19567a <=( (not A166)  and  A167 );
 a19571a <=( (not A265)  and  A201 );
 a19572a <=( A199  and  a19571a );
 a19573a <=( a19572a  and  a19567a );
 a19577a <=( (not A269)  and  A268 );
 a19578a <=( (not A266)  and  a19577a );
 a19582a <=( (not A301)  and  (not A299) );
 a19583a <=( (not A298)  and  a19582a );
 a19584a <=( a19583a  and  a19578a );
 a19587a <=( (not A166)  and  A167 );
 a19591a <=( (not A265)  and  A201 );
 a19592a <=( A199  and  a19591a );
 a19593a <=( a19592a  and  a19587a );
 a19597a <=( (not A269)  and  A268 );
 a19598a <=( (not A266)  and  a19597a );
 a19602a <=( A302  and  (not A299) );
 a19603a <=( (not A298)  and  a19602a );
 a19604a <=( a19603a  and  a19598a );
 a19607a <=( (not A166)  and  A167 );
 a19611a <=( A265  and  A201 );
 a19612a <=( A200  and  a19611a );
 a19613a <=( a19612a  and  a19607a );
 a19617a <=( (not A269)  and  A268 );
 a19618a <=( A266  and  a19617a );
 a19622a <=( (not A301)  and  (not A299) );
 a19623a <=( (not A298)  and  a19622a );
 a19624a <=( a19623a  and  a19618a );
 a19627a <=( (not A166)  and  A167 );
 a19631a <=( A265  and  A201 );
 a19632a <=( A200  and  a19631a );
 a19633a <=( a19632a  and  a19627a );
 a19637a <=( (not A269)  and  A268 );
 a19638a <=( A266  and  a19637a );
 a19642a <=( A302  and  (not A299) );
 a19643a <=( (not A298)  and  a19642a );
 a19644a <=( a19643a  and  a19638a );
 a19647a <=( (not A166)  and  A167 );
 a19651a <=( (not A265)  and  A201 );
 a19652a <=( A200  and  a19651a );
 a19653a <=( a19652a  and  a19647a );
 a19657a <=( A269  and  (not A268) );
 a19658a <=( A266  and  a19657a );
 a19662a <=( (not A301)  and  (not A299) );
 a19663a <=( (not A298)  and  a19662a );
 a19664a <=( a19663a  and  a19658a );
 a19667a <=( (not A166)  and  A167 );
 a19671a <=( (not A265)  and  A201 );
 a19672a <=( A200  and  a19671a );
 a19673a <=( a19672a  and  a19667a );
 a19677a <=( A269  and  (not A268) );
 a19678a <=( A266  and  a19677a );
 a19682a <=( A302  and  (not A299) );
 a19683a <=( (not A298)  and  a19682a );
 a19684a <=( a19683a  and  a19678a );
 a19687a <=( (not A166)  and  A167 );
 a19691a <=( A265  and  A201 );
 a19692a <=( A200  and  a19691a );
 a19693a <=( a19692a  and  a19687a );
 a19697a <=( A269  and  (not A268) );
 a19698a <=( (not A266)  and  a19697a );
 a19702a <=( (not A301)  and  (not A299) );
 a19703a <=( (not A298)  and  a19702a );
 a19704a <=( a19703a  and  a19698a );
 a19707a <=( (not A166)  and  A167 );
 a19711a <=( A265  and  A201 );
 a19712a <=( A200  and  a19711a );
 a19713a <=( a19712a  and  a19707a );
 a19717a <=( A269  and  (not A268) );
 a19718a <=( (not A266)  and  a19717a );
 a19722a <=( A302  and  (not A299) );
 a19723a <=( (not A298)  and  a19722a );
 a19724a <=( a19723a  and  a19718a );
 a19727a <=( (not A166)  and  A167 );
 a19731a <=( (not A265)  and  A201 );
 a19732a <=( A200  and  a19731a );
 a19733a <=( a19732a  and  a19727a );
 a19737a <=( (not A269)  and  A268 );
 a19738a <=( (not A266)  and  a19737a );
 a19742a <=( (not A301)  and  (not A299) );
 a19743a <=( (not A298)  and  a19742a );
 a19744a <=( a19743a  and  a19738a );
 a19747a <=( (not A166)  and  A167 );
 a19751a <=( (not A265)  and  A201 );
 a19752a <=( A200  and  a19751a );
 a19753a <=( a19752a  and  a19747a );
 a19757a <=( (not A269)  and  A268 );
 a19758a <=( (not A266)  and  a19757a );
 a19762a <=( A302  and  (not A299) );
 a19763a <=( (not A298)  and  a19762a );
 a19764a <=( a19763a  and  a19758a );
 a19767a <=( (not A166)  and  A167 );
 a19771a <=( A202  and  A200 );
 a19772a <=( A199  and  a19771a );
 a19773a <=( a19772a  and  a19767a );
 a19777a <=( A267  and  A265 );
 a19778a <=( (not A203)  and  a19777a );
 a19782a <=( (not A301)  and  (not A299) );
 a19783a <=( (not A298)  and  a19782a );
 a19784a <=( a19783a  and  a19778a );
 a19787a <=( (not A166)  and  A167 );
 a19791a <=( A202  and  A200 );
 a19792a <=( A199  and  a19791a );
 a19793a <=( a19792a  and  a19787a );
 a19797a <=( A267  and  A265 );
 a19798a <=( (not A203)  and  a19797a );
 a19802a <=( A302  and  (not A299) );
 a19803a <=( (not A298)  and  a19802a );
 a19804a <=( a19803a  and  a19798a );
 a19807a <=( (not A166)  and  A167 );
 a19811a <=( A202  and  A200 );
 a19812a <=( A199  and  a19811a );
 a19813a <=( a19812a  and  a19807a );
 a19817a <=( A267  and  A266 );
 a19818a <=( (not A203)  and  a19817a );
 a19822a <=( (not A301)  and  (not A299) );
 a19823a <=( (not A298)  and  a19822a );
 a19824a <=( a19823a  and  a19818a );
 a19827a <=( (not A166)  and  A167 );
 a19831a <=( A202  and  A200 );
 a19832a <=( A199  and  a19831a );
 a19833a <=( a19832a  and  a19827a );
 a19837a <=( A267  and  A266 );
 a19838a <=( (not A203)  and  a19837a );
 a19842a <=( A302  and  (not A299) );
 a19843a <=( (not A298)  and  a19842a );
 a19844a <=( a19843a  and  a19838a );
 a19847a <=( (not A166)  and  A167 );
 a19851a <=( (not A201)  and  A200 );
 a19852a <=( A199  and  a19851a );
 a19853a <=( a19852a  and  a19847a );
 a19857a <=( (not A266)  and  (not A265) );
 a19858a <=( (not A202)  and  a19857a );
 a19862a <=( A300  and  A299 );
 a19863a <=( (not A268)  and  a19862a );
 a19864a <=( a19863a  and  a19858a );
 a19867a <=( (not A166)  and  A167 );
 a19871a <=( (not A201)  and  A200 );
 a19872a <=( A199  and  a19871a );
 a19873a <=( a19872a  and  a19867a );
 a19877a <=( (not A266)  and  (not A265) );
 a19878a <=( (not A202)  and  a19877a );
 a19882a <=( A300  and  A298 );
 a19883a <=( (not A268)  and  a19882a );
 a19884a <=( a19883a  and  a19878a );
 a19887a <=( (not A166)  and  A167 );
 a19891a <=( (not A201)  and  A200 );
 a19892a <=( A199  and  a19891a );
 a19893a <=( a19892a  and  a19887a );
 a19897a <=( (not A266)  and  (not A265) );
 a19898a <=( (not A202)  and  a19897a );
 a19902a <=( A300  and  A299 );
 a19903a <=( A269  and  a19902a );
 a19904a <=( a19903a  and  a19898a );
 a19907a <=( (not A166)  and  A167 );
 a19911a <=( (not A201)  and  A200 );
 a19912a <=( A199  and  a19911a );
 a19913a <=( a19912a  and  a19907a );
 a19917a <=( (not A266)  and  (not A265) );
 a19918a <=( (not A202)  and  a19917a );
 a19922a <=( A300  and  A298 );
 a19923a <=( A269  and  a19922a );
 a19924a <=( a19923a  and  a19918a );
 a19927a <=( (not A166)  and  A167 );
 a19931a <=( (not A201)  and  A200 );
 a19932a <=( A199  and  a19931a );
 a19933a <=( a19932a  and  a19927a );
 a19937a <=( (not A266)  and  (not A265) );
 a19938a <=( A203  and  a19937a );
 a19942a <=( A300  and  A299 );
 a19943a <=( (not A268)  and  a19942a );
 a19944a <=( a19943a  and  a19938a );
 a19947a <=( (not A166)  and  A167 );
 a19951a <=( (not A201)  and  A200 );
 a19952a <=( A199  and  a19951a );
 a19953a <=( a19952a  and  a19947a );
 a19957a <=( (not A266)  and  (not A265) );
 a19958a <=( A203  and  a19957a );
 a19962a <=( A300  and  A298 );
 a19963a <=( (not A268)  and  a19962a );
 a19964a <=( a19963a  and  a19958a );
 a19967a <=( (not A166)  and  A167 );
 a19971a <=( (not A201)  and  A200 );
 a19972a <=( A199  and  a19971a );
 a19973a <=( a19972a  and  a19967a );
 a19977a <=( (not A266)  and  (not A265) );
 a19978a <=( A203  and  a19977a );
 a19982a <=( A300  and  A299 );
 a19983a <=( A269  and  a19982a );
 a19984a <=( a19983a  and  a19978a );
 a19987a <=( (not A166)  and  A167 );
 a19991a <=( (not A201)  and  A200 );
 a19992a <=( A199  and  a19991a );
 a19993a <=( a19992a  and  a19987a );
 a19997a <=( (not A266)  and  (not A265) );
 a19998a <=( A203  and  a19997a );
 a20002a <=( A300  and  A298 );
 a20003a <=( A269  and  a20002a );
 a20004a <=( a20003a  and  a19998a );
 a20007a <=( (not A166)  and  A167 );
 a20011a <=( (not A202)  and  A200 );
 a20012a <=( (not A199)  and  a20011a );
 a20013a <=( a20012a  and  a20007a );
 a20017a <=( A267  and  A265 );
 a20018a <=( A203  and  a20017a );
 a20022a <=( (not A301)  and  (not A299) );
 a20023a <=( (not A298)  and  a20022a );
 a20024a <=( a20023a  and  a20018a );
 a20027a <=( (not A166)  and  A167 );
 a20031a <=( (not A202)  and  A200 );
 a20032a <=( (not A199)  and  a20031a );
 a20033a <=( a20032a  and  a20027a );
 a20037a <=( A267  and  A265 );
 a20038a <=( A203  and  a20037a );
 a20042a <=( A302  and  (not A299) );
 a20043a <=( (not A298)  and  a20042a );
 a20044a <=( a20043a  and  a20038a );
 a20047a <=( (not A166)  and  A167 );
 a20051a <=( (not A202)  and  A200 );
 a20052a <=( (not A199)  and  a20051a );
 a20053a <=( a20052a  and  a20047a );
 a20057a <=( A267  and  A266 );
 a20058a <=( A203  and  a20057a );
 a20062a <=( (not A301)  and  (not A299) );
 a20063a <=( (not A298)  and  a20062a );
 a20064a <=( a20063a  and  a20058a );
 a20067a <=( (not A166)  and  A167 );
 a20071a <=( (not A202)  and  A200 );
 a20072a <=( (not A199)  and  a20071a );
 a20073a <=( a20072a  and  a20067a );
 a20077a <=( A267  and  A266 );
 a20078a <=( A203  and  a20077a );
 a20082a <=( A302  and  (not A299) );
 a20083a <=( (not A298)  and  a20082a );
 a20084a <=( a20083a  and  a20078a );
 a20087a <=( (not A166)  and  A167 );
 a20091a <=( (not A201)  and  A200 );
 a20092a <=( (not A199)  and  a20091a );
 a20093a <=( a20092a  and  a20087a );
 a20097a <=( (not A266)  and  (not A265) );
 a20098a <=( A202  and  a20097a );
 a20102a <=( A300  and  A299 );
 a20103a <=( (not A268)  and  a20102a );
 a20104a <=( a20103a  and  a20098a );
 a20107a <=( (not A166)  and  A167 );
 a20111a <=( (not A201)  and  A200 );
 a20112a <=( (not A199)  and  a20111a );
 a20113a <=( a20112a  and  a20107a );
 a20117a <=( (not A266)  and  (not A265) );
 a20118a <=( A202  and  a20117a );
 a20122a <=( A300  and  A298 );
 a20123a <=( (not A268)  and  a20122a );
 a20124a <=( a20123a  and  a20118a );
 a20127a <=( (not A166)  and  A167 );
 a20131a <=( (not A201)  and  A200 );
 a20132a <=( (not A199)  and  a20131a );
 a20133a <=( a20132a  and  a20127a );
 a20137a <=( (not A266)  and  (not A265) );
 a20138a <=( A202  and  a20137a );
 a20142a <=( A300  and  A299 );
 a20143a <=( A269  and  a20142a );
 a20144a <=( a20143a  and  a20138a );
 a20147a <=( (not A166)  and  A167 );
 a20151a <=( (not A201)  and  A200 );
 a20152a <=( (not A199)  and  a20151a );
 a20153a <=( a20152a  and  a20147a );
 a20157a <=( (not A266)  and  (not A265) );
 a20158a <=( A202  and  a20157a );
 a20162a <=( A300  and  A298 );
 a20163a <=( A269  and  a20162a );
 a20164a <=( a20163a  and  a20158a );
 a20167a <=( (not A166)  and  A167 );
 a20171a <=( (not A201)  and  A200 );
 a20172a <=( (not A199)  and  a20171a );
 a20173a <=( a20172a  and  a20167a );
 a20177a <=( (not A266)  and  (not A265) );
 a20178a <=( (not A203)  and  a20177a );
 a20182a <=( A300  and  A299 );
 a20183a <=( (not A268)  and  a20182a );
 a20184a <=( a20183a  and  a20178a );
 a20187a <=( (not A166)  and  A167 );
 a20191a <=( (not A201)  and  A200 );
 a20192a <=( (not A199)  and  a20191a );
 a20193a <=( a20192a  and  a20187a );
 a20197a <=( (not A266)  and  (not A265) );
 a20198a <=( (not A203)  and  a20197a );
 a20202a <=( A300  and  A298 );
 a20203a <=( (not A268)  and  a20202a );
 a20204a <=( a20203a  and  a20198a );
 a20207a <=( (not A166)  and  A167 );
 a20211a <=( (not A201)  and  A200 );
 a20212a <=( (not A199)  and  a20211a );
 a20213a <=( a20212a  and  a20207a );
 a20217a <=( (not A266)  and  (not A265) );
 a20218a <=( (not A203)  and  a20217a );
 a20222a <=( A300  and  A299 );
 a20223a <=( A269  and  a20222a );
 a20224a <=( a20223a  and  a20218a );
 a20227a <=( (not A166)  and  A167 );
 a20231a <=( (not A201)  and  A200 );
 a20232a <=( (not A199)  and  a20231a );
 a20233a <=( a20232a  and  a20227a );
 a20237a <=( (not A266)  and  (not A265) );
 a20238a <=( (not A203)  and  a20237a );
 a20242a <=( A300  and  A298 );
 a20243a <=( A269  and  a20242a );
 a20244a <=( a20243a  and  a20238a );
 a20247a <=( (not A166)  and  A167 );
 a20251a <=( (not A202)  and  (not A200) );
 a20252a <=( A199  and  a20251a );
 a20253a <=( a20252a  and  a20247a );
 a20257a <=( A267  and  A265 );
 a20258a <=( A203  and  a20257a );
 a20262a <=( (not A301)  and  (not A299) );
 a20263a <=( (not A298)  and  a20262a );
 a20264a <=( a20263a  and  a20258a );
 a20267a <=( (not A166)  and  A167 );
 a20271a <=( (not A202)  and  (not A200) );
 a20272a <=( A199  and  a20271a );
 a20273a <=( a20272a  and  a20267a );
 a20277a <=( A267  and  A265 );
 a20278a <=( A203  and  a20277a );
 a20282a <=( A302  and  (not A299) );
 a20283a <=( (not A298)  and  a20282a );
 a20284a <=( a20283a  and  a20278a );
 a20287a <=( (not A166)  and  A167 );
 a20291a <=( (not A202)  and  (not A200) );
 a20292a <=( A199  and  a20291a );
 a20293a <=( a20292a  and  a20287a );
 a20297a <=( A267  and  A266 );
 a20298a <=( A203  and  a20297a );
 a20302a <=( (not A301)  and  (not A299) );
 a20303a <=( (not A298)  and  a20302a );
 a20304a <=( a20303a  and  a20298a );
 a20307a <=( (not A166)  and  A167 );
 a20311a <=( (not A202)  and  (not A200) );
 a20312a <=( A199  and  a20311a );
 a20313a <=( a20312a  and  a20307a );
 a20317a <=( A267  and  A266 );
 a20318a <=( A203  and  a20317a );
 a20322a <=( A302  and  (not A299) );
 a20323a <=( (not A298)  and  a20322a );
 a20324a <=( a20323a  and  a20318a );
 a20327a <=( (not A166)  and  A167 );
 a20331a <=( (not A201)  and  (not A200) );
 a20332a <=( A199  and  a20331a );
 a20333a <=( a20332a  and  a20327a );
 a20337a <=( (not A266)  and  (not A265) );
 a20338a <=( A202  and  a20337a );
 a20342a <=( A300  and  A299 );
 a20343a <=( (not A268)  and  a20342a );
 a20344a <=( a20343a  and  a20338a );
 a20347a <=( (not A166)  and  A167 );
 a20351a <=( (not A201)  and  (not A200) );
 a20352a <=( A199  and  a20351a );
 a20353a <=( a20352a  and  a20347a );
 a20357a <=( (not A266)  and  (not A265) );
 a20358a <=( A202  and  a20357a );
 a20362a <=( A300  and  A298 );
 a20363a <=( (not A268)  and  a20362a );
 a20364a <=( a20363a  and  a20358a );
 a20367a <=( (not A166)  and  A167 );
 a20371a <=( (not A201)  and  (not A200) );
 a20372a <=( A199  and  a20371a );
 a20373a <=( a20372a  and  a20367a );
 a20377a <=( (not A266)  and  (not A265) );
 a20378a <=( A202  and  a20377a );
 a20382a <=( A300  and  A299 );
 a20383a <=( A269  and  a20382a );
 a20384a <=( a20383a  and  a20378a );
 a20387a <=( (not A166)  and  A167 );
 a20391a <=( (not A201)  and  (not A200) );
 a20392a <=( A199  and  a20391a );
 a20393a <=( a20392a  and  a20387a );
 a20397a <=( (not A266)  and  (not A265) );
 a20398a <=( A202  and  a20397a );
 a20402a <=( A300  and  A298 );
 a20403a <=( A269  and  a20402a );
 a20404a <=( a20403a  and  a20398a );
 a20407a <=( (not A166)  and  A167 );
 a20411a <=( (not A201)  and  (not A200) );
 a20412a <=( A199  and  a20411a );
 a20413a <=( a20412a  and  a20407a );
 a20417a <=( (not A266)  and  (not A265) );
 a20418a <=( (not A203)  and  a20417a );
 a20422a <=( A300  and  A299 );
 a20423a <=( (not A268)  and  a20422a );
 a20424a <=( a20423a  and  a20418a );
 a20427a <=( (not A166)  and  A167 );
 a20431a <=( (not A201)  and  (not A200) );
 a20432a <=( A199  and  a20431a );
 a20433a <=( a20432a  and  a20427a );
 a20437a <=( (not A266)  and  (not A265) );
 a20438a <=( (not A203)  and  a20437a );
 a20442a <=( A300  and  A298 );
 a20443a <=( (not A268)  and  a20442a );
 a20444a <=( a20443a  and  a20438a );
 a20447a <=( (not A166)  and  A167 );
 a20451a <=( (not A201)  and  (not A200) );
 a20452a <=( A199  and  a20451a );
 a20453a <=( a20452a  and  a20447a );
 a20457a <=( (not A266)  and  (not A265) );
 a20458a <=( (not A203)  and  a20457a );
 a20462a <=( A300  and  A299 );
 a20463a <=( A269  and  a20462a );
 a20464a <=( a20463a  and  a20458a );
 a20467a <=( (not A166)  and  A167 );
 a20471a <=( (not A201)  and  (not A200) );
 a20472a <=( A199  and  a20471a );
 a20473a <=( a20472a  and  a20467a );
 a20477a <=( (not A266)  and  (not A265) );
 a20478a <=( (not A203)  and  a20477a );
 a20482a <=( A300  and  A298 );
 a20483a <=( A269  and  a20482a );
 a20484a <=( a20483a  and  a20478a );
 a20487a <=( (not A166)  and  A167 );
 a20491a <=( (not A202)  and  (not A200) );
 a20492a <=( (not A199)  and  a20491a );
 a20493a <=( a20492a  and  a20487a );
 a20497a <=( (not A267)  and  A266 );
 a20498a <=( A265  and  a20497a );
 a20502a <=( A300  and  A299 );
 a20503a <=( (not A268)  and  a20502a );
 a20504a <=( a20503a  and  a20498a );
 a20507a <=( (not A166)  and  A167 );
 a20511a <=( (not A202)  and  (not A200) );
 a20512a <=( (not A199)  and  a20511a );
 a20513a <=( a20512a  and  a20507a );
 a20517a <=( (not A267)  and  A266 );
 a20518a <=( A265  and  a20517a );
 a20522a <=( A300  and  A298 );
 a20523a <=( (not A268)  and  a20522a );
 a20524a <=( a20523a  and  a20518a );
 a20527a <=( (not A166)  and  A167 );
 a20531a <=( (not A202)  and  (not A200) );
 a20532a <=( (not A199)  and  a20531a );
 a20533a <=( a20532a  and  a20527a );
 a20537a <=( (not A267)  and  A266 );
 a20538a <=( A265  and  a20537a );
 a20542a <=( A300  and  A299 );
 a20543a <=( A269  and  a20542a );
 a20544a <=( a20543a  and  a20538a );
 a20547a <=( (not A166)  and  A167 );
 a20551a <=( (not A202)  and  (not A200) );
 a20552a <=( (not A199)  and  a20551a );
 a20553a <=( a20552a  and  a20547a );
 a20557a <=( (not A267)  and  A266 );
 a20558a <=( A265  and  a20557a );
 a20562a <=( A300  and  A298 );
 a20563a <=( A269  and  a20562a );
 a20564a <=( a20563a  and  a20558a );
 a20567a <=( (not A166)  and  A167 );
 a20571a <=( (not A202)  and  (not A200) );
 a20572a <=( (not A199)  and  a20571a );
 a20573a <=( a20572a  and  a20567a );
 a20577a <=( (not A267)  and  A266 );
 a20578a <=( (not A265)  and  a20577a );
 a20582a <=( A300  and  A299 );
 a20583a <=( A268  and  a20582a );
 a20584a <=( a20583a  and  a20578a );
 a20587a <=( (not A166)  and  A167 );
 a20591a <=( (not A202)  and  (not A200) );
 a20592a <=( (not A199)  and  a20591a );
 a20593a <=( a20592a  and  a20587a );
 a20597a <=( (not A267)  and  A266 );
 a20598a <=( (not A265)  and  a20597a );
 a20602a <=( A300  and  A298 );
 a20603a <=( A268  and  a20602a );
 a20604a <=( a20603a  and  a20598a );
 a20607a <=( (not A166)  and  A167 );
 a20611a <=( (not A202)  and  (not A200) );
 a20612a <=( (not A199)  and  a20611a );
 a20613a <=( a20612a  and  a20607a );
 a20617a <=( (not A267)  and  A266 );
 a20618a <=( (not A265)  and  a20617a );
 a20622a <=( A300  and  A299 );
 a20623a <=( (not A269)  and  a20622a );
 a20624a <=( a20623a  and  a20618a );
 a20627a <=( (not A166)  and  A167 );
 a20631a <=( (not A202)  and  (not A200) );
 a20632a <=( (not A199)  and  a20631a );
 a20633a <=( a20632a  and  a20627a );
 a20637a <=( (not A267)  and  A266 );
 a20638a <=( (not A265)  and  a20637a );
 a20642a <=( A300  and  A298 );
 a20643a <=( (not A269)  and  a20642a );
 a20644a <=( a20643a  and  a20638a );
 a20647a <=( (not A166)  and  A167 );
 a20651a <=( (not A202)  and  (not A200) );
 a20652a <=( (not A199)  and  a20651a );
 a20653a <=( a20652a  and  a20647a );
 a20657a <=( (not A267)  and  (not A266) );
 a20658a <=( A265  and  a20657a );
 a20662a <=( A300  and  A299 );
 a20663a <=( A268  and  a20662a );
 a20664a <=( a20663a  and  a20658a );
 a20667a <=( (not A166)  and  A167 );
 a20671a <=( (not A202)  and  (not A200) );
 a20672a <=( (not A199)  and  a20671a );
 a20673a <=( a20672a  and  a20667a );
 a20677a <=( (not A267)  and  (not A266) );
 a20678a <=( A265  and  a20677a );
 a20682a <=( A300  and  A298 );
 a20683a <=( A268  and  a20682a );
 a20684a <=( a20683a  and  a20678a );
 a20687a <=( (not A166)  and  A167 );
 a20691a <=( (not A202)  and  (not A200) );
 a20692a <=( (not A199)  and  a20691a );
 a20693a <=( a20692a  and  a20687a );
 a20697a <=( (not A267)  and  (not A266) );
 a20698a <=( A265  and  a20697a );
 a20702a <=( A300  and  A299 );
 a20703a <=( (not A269)  and  a20702a );
 a20704a <=( a20703a  and  a20698a );
 a20707a <=( (not A166)  and  A167 );
 a20711a <=( (not A202)  and  (not A200) );
 a20712a <=( (not A199)  and  a20711a );
 a20713a <=( a20712a  and  a20707a );
 a20717a <=( (not A267)  and  (not A266) );
 a20718a <=( A265  and  a20717a );
 a20722a <=( A300  and  A298 );
 a20723a <=( (not A269)  and  a20722a );
 a20724a <=( a20723a  and  a20718a );
 a20727a <=( (not A166)  and  A167 );
 a20731a <=( A203  and  (not A200) );
 a20732a <=( (not A199)  and  a20731a );
 a20733a <=( a20732a  and  a20727a );
 a20737a <=( (not A267)  and  A266 );
 a20738a <=( A265  and  a20737a );
 a20742a <=( A300  and  A299 );
 a20743a <=( (not A268)  and  a20742a );
 a20744a <=( a20743a  and  a20738a );
 a20747a <=( (not A166)  and  A167 );
 a20751a <=( A203  and  (not A200) );
 a20752a <=( (not A199)  and  a20751a );
 a20753a <=( a20752a  and  a20747a );
 a20757a <=( (not A267)  and  A266 );
 a20758a <=( A265  and  a20757a );
 a20762a <=( A300  and  A298 );
 a20763a <=( (not A268)  and  a20762a );
 a20764a <=( a20763a  and  a20758a );
 a20767a <=( (not A166)  and  A167 );
 a20771a <=( A203  and  (not A200) );
 a20772a <=( (not A199)  and  a20771a );
 a20773a <=( a20772a  and  a20767a );
 a20777a <=( (not A267)  and  A266 );
 a20778a <=( A265  and  a20777a );
 a20782a <=( A300  and  A299 );
 a20783a <=( A269  and  a20782a );
 a20784a <=( a20783a  and  a20778a );
 a20787a <=( (not A166)  and  A167 );
 a20791a <=( A203  and  (not A200) );
 a20792a <=( (not A199)  and  a20791a );
 a20793a <=( a20792a  and  a20787a );
 a20797a <=( (not A267)  and  A266 );
 a20798a <=( A265  and  a20797a );
 a20802a <=( A300  and  A298 );
 a20803a <=( A269  and  a20802a );
 a20804a <=( a20803a  and  a20798a );
 a20807a <=( (not A166)  and  A167 );
 a20811a <=( A203  and  (not A200) );
 a20812a <=( (not A199)  and  a20811a );
 a20813a <=( a20812a  and  a20807a );
 a20817a <=( (not A267)  and  A266 );
 a20818a <=( (not A265)  and  a20817a );
 a20822a <=( A300  and  A299 );
 a20823a <=( A268  and  a20822a );
 a20824a <=( a20823a  and  a20818a );
 a20827a <=( (not A166)  and  A167 );
 a20831a <=( A203  and  (not A200) );
 a20832a <=( (not A199)  and  a20831a );
 a20833a <=( a20832a  and  a20827a );
 a20837a <=( (not A267)  and  A266 );
 a20838a <=( (not A265)  and  a20837a );
 a20842a <=( A300  and  A298 );
 a20843a <=( A268  and  a20842a );
 a20844a <=( a20843a  and  a20838a );
 a20847a <=( (not A166)  and  A167 );
 a20851a <=( A203  and  (not A200) );
 a20852a <=( (not A199)  and  a20851a );
 a20853a <=( a20852a  and  a20847a );
 a20857a <=( (not A267)  and  A266 );
 a20858a <=( (not A265)  and  a20857a );
 a20862a <=( A300  and  A299 );
 a20863a <=( (not A269)  and  a20862a );
 a20864a <=( a20863a  and  a20858a );
 a20867a <=( (not A166)  and  A167 );
 a20871a <=( A203  and  (not A200) );
 a20872a <=( (not A199)  and  a20871a );
 a20873a <=( a20872a  and  a20867a );
 a20877a <=( (not A267)  and  A266 );
 a20878a <=( (not A265)  and  a20877a );
 a20882a <=( A300  and  A298 );
 a20883a <=( (not A269)  and  a20882a );
 a20884a <=( a20883a  and  a20878a );
 a20887a <=( (not A166)  and  A167 );
 a20891a <=( A203  and  (not A200) );
 a20892a <=( (not A199)  and  a20891a );
 a20893a <=( a20892a  and  a20887a );
 a20897a <=( (not A267)  and  (not A266) );
 a20898a <=( A265  and  a20897a );
 a20902a <=( A300  and  A299 );
 a20903a <=( A268  and  a20902a );
 a20904a <=( a20903a  and  a20898a );
 a20907a <=( (not A166)  and  A167 );
 a20911a <=( A203  and  (not A200) );
 a20912a <=( (not A199)  and  a20911a );
 a20913a <=( a20912a  and  a20907a );
 a20917a <=( (not A267)  and  (not A266) );
 a20918a <=( A265  and  a20917a );
 a20922a <=( A300  and  A298 );
 a20923a <=( A268  and  a20922a );
 a20924a <=( a20923a  and  a20918a );
 a20927a <=( (not A166)  and  A167 );
 a20931a <=( A203  and  (not A200) );
 a20932a <=( (not A199)  and  a20931a );
 a20933a <=( a20932a  and  a20927a );
 a20937a <=( (not A267)  and  (not A266) );
 a20938a <=( A265  and  a20937a );
 a20942a <=( A300  and  A299 );
 a20943a <=( (not A269)  and  a20942a );
 a20944a <=( a20943a  and  a20938a );
 a20947a <=( (not A166)  and  A167 );
 a20951a <=( A203  and  (not A200) );
 a20952a <=( (not A199)  and  a20951a );
 a20953a <=( a20952a  and  a20947a );
 a20957a <=( (not A267)  and  (not A266) );
 a20958a <=( A265  and  a20957a );
 a20962a <=( A300  and  A298 );
 a20963a <=( (not A269)  and  a20962a );
 a20964a <=( a20963a  and  a20958a );
 a20967a <=( (not A166)  and  A167 );
 a20971a <=( A202  and  (not A200) );
 a20972a <=( (not A199)  and  a20971a );
 a20973a <=( a20972a  and  a20967a );
 a20977a <=( A267  and  A265 );
 a20978a <=( (not A203)  and  a20977a );
 a20982a <=( (not A301)  and  (not A299) );
 a20983a <=( (not A298)  and  a20982a );
 a20984a <=( a20983a  and  a20978a );
 a20987a <=( (not A166)  and  A167 );
 a20991a <=( A202  and  (not A200) );
 a20992a <=( (not A199)  and  a20991a );
 a20993a <=( a20992a  and  a20987a );
 a20997a <=( A267  and  A265 );
 a20998a <=( (not A203)  and  a20997a );
 a21002a <=( A302  and  (not A299) );
 a21003a <=( (not A298)  and  a21002a );
 a21004a <=( a21003a  and  a20998a );
 a21007a <=( (not A166)  and  A167 );
 a21011a <=( A202  and  (not A200) );
 a21012a <=( (not A199)  and  a21011a );
 a21013a <=( a21012a  and  a21007a );
 a21017a <=( A267  and  A266 );
 a21018a <=( (not A203)  and  a21017a );
 a21022a <=( (not A301)  and  (not A299) );
 a21023a <=( (not A298)  and  a21022a );
 a21024a <=( a21023a  and  a21018a );
 a21027a <=( (not A166)  and  A167 );
 a21031a <=( A202  and  (not A200) );
 a21032a <=( (not A199)  and  a21031a );
 a21033a <=( a21032a  and  a21027a );
 a21037a <=( A267  and  A266 );
 a21038a <=( (not A203)  and  a21037a );
 a21042a <=( A302  and  (not A299) );
 a21043a <=( (not A298)  and  a21042a );
 a21044a <=( a21043a  and  a21038a );
 a21047a <=( (not A166)  and  (not A167) );
 a21051a <=( (not A265)  and  A201 );
 a21052a <=( A199  and  a21051a );
 a21053a <=( a21052a  and  a21047a );
 a21057a <=( A298  and  (not A268) );
 a21058a <=( (not A266)  and  a21057a );
 a21062a <=( (not A302)  and  A301 );
 a21063a <=( A299  and  a21062a );
 a21064a <=( a21063a  and  a21058a );
 a21067a <=( (not A166)  and  (not A167) );
 a21071a <=( (not A265)  and  A201 );
 a21072a <=( A199  and  a21071a );
 a21073a <=( a21072a  and  a21067a );
 a21077a <=( A298  and  (not A268) );
 a21078a <=( (not A266)  and  a21077a );
 a21082a <=( A302  and  (not A301) );
 a21083a <=( (not A299)  and  a21082a );
 a21084a <=( a21083a  and  a21078a );
 a21087a <=( (not A166)  and  (not A167) );
 a21091a <=( (not A265)  and  A201 );
 a21092a <=( A199  and  a21091a );
 a21093a <=( a21092a  and  a21087a );
 a21097a <=( (not A298)  and  (not A268) );
 a21098a <=( (not A266)  and  a21097a );
 a21102a <=( A302  and  (not A301) );
 a21103a <=( A299  and  a21102a );
 a21104a <=( a21103a  and  a21098a );
 a21107a <=( (not A166)  and  (not A167) );
 a21111a <=( (not A265)  and  A201 );
 a21112a <=( A199  and  a21111a );
 a21113a <=( a21112a  and  a21107a );
 a21117a <=( (not A298)  and  (not A268) );
 a21118a <=( (not A266)  and  a21117a );
 a21122a <=( (not A302)  and  A301 );
 a21123a <=( (not A299)  and  a21122a );
 a21124a <=( a21123a  and  a21118a );
 a21127a <=( (not A166)  and  (not A167) );
 a21131a <=( (not A265)  and  A201 );
 a21132a <=( A199  and  a21131a );
 a21133a <=( a21132a  and  a21127a );
 a21137a <=( A298  and  A269 );
 a21138a <=( (not A266)  and  a21137a );
 a21142a <=( (not A302)  and  A301 );
 a21143a <=( A299  and  a21142a );
 a21144a <=( a21143a  and  a21138a );
 a21147a <=( (not A166)  and  (not A167) );
 a21151a <=( (not A265)  and  A201 );
 a21152a <=( A199  and  a21151a );
 a21153a <=( a21152a  and  a21147a );
 a21157a <=( A298  and  A269 );
 a21158a <=( (not A266)  and  a21157a );
 a21162a <=( A302  and  (not A301) );
 a21163a <=( (not A299)  and  a21162a );
 a21164a <=( a21163a  and  a21158a );
 a21167a <=( (not A166)  and  (not A167) );
 a21171a <=( (not A265)  and  A201 );
 a21172a <=( A199  and  a21171a );
 a21173a <=( a21172a  and  a21167a );
 a21177a <=( (not A298)  and  A269 );
 a21178a <=( (not A266)  and  a21177a );
 a21182a <=( A302  and  (not A301) );
 a21183a <=( A299  and  a21182a );
 a21184a <=( a21183a  and  a21178a );
 a21187a <=( (not A166)  and  (not A167) );
 a21191a <=( (not A265)  and  A201 );
 a21192a <=( A199  and  a21191a );
 a21193a <=( a21192a  and  a21187a );
 a21197a <=( (not A298)  and  A269 );
 a21198a <=( (not A266)  and  a21197a );
 a21202a <=( (not A302)  and  A301 );
 a21203a <=( (not A299)  and  a21202a );
 a21204a <=( a21203a  and  a21198a );
 a21207a <=( (not A166)  and  (not A167) );
 a21211a <=( (not A265)  and  A201 );
 a21212a <=( A200  and  a21211a );
 a21213a <=( a21212a  and  a21207a );
 a21217a <=( A298  and  (not A268) );
 a21218a <=( (not A266)  and  a21217a );
 a21222a <=( (not A302)  and  A301 );
 a21223a <=( A299  and  a21222a );
 a21224a <=( a21223a  and  a21218a );
 a21227a <=( (not A166)  and  (not A167) );
 a21231a <=( (not A265)  and  A201 );
 a21232a <=( A200  and  a21231a );
 a21233a <=( a21232a  and  a21227a );
 a21237a <=( A298  and  (not A268) );
 a21238a <=( (not A266)  and  a21237a );
 a21242a <=( A302  and  (not A301) );
 a21243a <=( (not A299)  and  a21242a );
 a21244a <=( a21243a  and  a21238a );
 a21247a <=( (not A166)  and  (not A167) );
 a21251a <=( (not A265)  and  A201 );
 a21252a <=( A200  and  a21251a );
 a21253a <=( a21252a  and  a21247a );
 a21257a <=( (not A298)  and  (not A268) );
 a21258a <=( (not A266)  and  a21257a );
 a21262a <=( A302  and  (not A301) );
 a21263a <=( A299  and  a21262a );
 a21264a <=( a21263a  and  a21258a );
 a21267a <=( (not A166)  and  (not A167) );
 a21271a <=( (not A265)  and  A201 );
 a21272a <=( A200  and  a21271a );
 a21273a <=( a21272a  and  a21267a );
 a21277a <=( (not A298)  and  (not A268) );
 a21278a <=( (not A266)  and  a21277a );
 a21282a <=( (not A302)  and  A301 );
 a21283a <=( (not A299)  and  a21282a );
 a21284a <=( a21283a  and  a21278a );
 a21287a <=( (not A166)  and  (not A167) );
 a21291a <=( (not A265)  and  A201 );
 a21292a <=( A200  and  a21291a );
 a21293a <=( a21292a  and  a21287a );
 a21297a <=( A298  and  A269 );
 a21298a <=( (not A266)  and  a21297a );
 a21302a <=( (not A302)  and  A301 );
 a21303a <=( A299  and  a21302a );
 a21304a <=( a21303a  and  a21298a );
 a21307a <=( (not A166)  and  (not A167) );
 a21311a <=( (not A265)  and  A201 );
 a21312a <=( A200  and  a21311a );
 a21313a <=( a21312a  and  a21307a );
 a21317a <=( A298  and  A269 );
 a21318a <=( (not A266)  and  a21317a );
 a21322a <=( A302  and  (not A301) );
 a21323a <=( (not A299)  and  a21322a );
 a21324a <=( a21323a  and  a21318a );
 a21327a <=( (not A166)  and  (not A167) );
 a21331a <=( (not A265)  and  A201 );
 a21332a <=( A200  and  a21331a );
 a21333a <=( a21332a  and  a21327a );
 a21337a <=( (not A298)  and  A269 );
 a21338a <=( (not A266)  and  a21337a );
 a21342a <=( A302  and  (not A301) );
 a21343a <=( A299  and  a21342a );
 a21344a <=( a21343a  and  a21338a );
 a21347a <=( (not A166)  and  (not A167) );
 a21351a <=( (not A265)  and  A201 );
 a21352a <=( A200  and  a21351a );
 a21353a <=( a21352a  and  a21347a );
 a21357a <=( (not A298)  and  A269 );
 a21358a <=( (not A266)  and  a21357a );
 a21362a <=( (not A302)  and  A301 );
 a21363a <=( (not A299)  and  a21362a );
 a21364a <=( a21363a  and  a21358a );
 a21367a <=( (not A166)  and  (not A167) );
 a21371a <=( A202  and  A200 );
 a21372a <=( A199  and  a21371a );
 a21373a <=( a21372a  and  a21367a );
 a21377a <=( (not A266)  and  (not A265) );
 a21378a <=( (not A203)  and  a21377a );
 a21382a <=( A300  and  A299 );
 a21383a <=( (not A268)  and  a21382a );
 a21384a <=( a21383a  and  a21378a );
 a21387a <=( (not A166)  and  (not A167) );
 a21391a <=( A202  and  A200 );
 a21392a <=( A199  and  a21391a );
 a21393a <=( a21392a  and  a21387a );
 a21397a <=( (not A266)  and  (not A265) );
 a21398a <=( (not A203)  and  a21397a );
 a21402a <=( A300  and  A298 );
 a21403a <=( (not A268)  and  a21402a );
 a21404a <=( a21403a  and  a21398a );
 a21407a <=( (not A166)  and  (not A167) );
 a21411a <=( A202  and  A200 );
 a21412a <=( A199  and  a21411a );
 a21413a <=( a21412a  and  a21407a );
 a21417a <=( (not A266)  and  (not A265) );
 a21418a <=( (not A203)  and  a21417a );
 a21422a <=( A300  and  A299 );
 a21423a <=( A269  and  a21422a );
 a21424a <=( a21423a  and  a21418a );
 a21427a <=( (not A166)  and  (not A167) );
 a21431a <=( A202  and  A200 );
 a21432a <=( A199  and  a21431a );
 a21433a <=( a21432a  and  a21427a );
 a21437a <=( (not A266)  and  (not A265) );
 a21438a <=( (not A203)  and  a21437a );
 a21442a <=( A300  and  A298 );
 a21443a <=( A269  and  a21442a );
 a21444a <=( a21443a  and  a21438a );
 a21447a <=( (not A166)  and  (not A167) );
 a21451a <=( (not A201)  and  A200 );
 a21452a <=( A199  and  a21451a );
 a21453a <=( a21452a  and  a21447a );
 a21457a <=( A267  and  A265 );
 a21458a <=( (not A202)  and  a21457a );
 a21462a <=( (not A301)  and  (not A299) );
 a21463a <=( (not A298)  and  a21462a );
 a21464a <=( a21463a  and  a21458a );
 a21467a <=( (not A166)  and  (not A167) );
 a21471a <=( (not A201)  and  A200 );
 a21472a <=( A199  and  a21471a );
 a21473a <=( a21472a  and  a21467a );
 a21477a <=( A267  and  A265 );
 a21478a <=( (not A202)  and  a21477a );
 a21482a <=( A302  and  (not A299) );
 a21483a <=( (not A298)  and  a21482a );
 a21484a <=( a21483a  and  a21478a );
 a21487a <=( (not A166)  and  (not A167) );
 a21491a <=( (not A201)  and  A200 );
 a21492a <=( A199  and  a21491a );
 a21493a <=( a21492a  and  a21487a );
 a21497a <=( A267  and  A266 );
 a21498a <=( (not A202)  and  a21497a );
 a21502a <=( (not A301)  and  (not A299) );
 a21503a <=( (not A298)  and  a21502a );
 a21504a <=( a21503a  and  a21498a );
 a21507a <=( (not A166)  and  (not A167) );
 a21511a <=( (not A201)  and  A200 );
 a21512a <=( A199  and  a21511a );
 a21513a <=( a21512a  and  a21507a );
 a21517a <=( A267  and  A266 );
 a21518a <=( (not A202)  and  a21517a );
 a21522a <=( A302  and  (not A299) );
 a21523a <=( (not A298)  and  a21522a );
 a21524a <=( a21523a  and  a21518a );
 a21527a <=( (not A166)  and  (not A167) );
 a21531a <=( (not A201)  and  A200 );
 a21532a <=( A199  and  a21531a );
 a21533a <=( a21532a  and  a21527a );
 a21537a <=( A267  and  A265 );
 a21538a <=( A203  and  a21537a );
 a21542a <=( (not A301)  and  (not A299) );
 a21543a <=( (not A298)  and  a21542a );
 a21544a <=( a21543a  and  a21538a );
 a21547a <=( (not A166)  and  (not A167) );
 a21551a <=( (not A201)  and  A200 );
 a21552a <=( A199  and  a21551a );
 a21553a <=( a21552a  and  a21547a );
 a21557a <=( A267  and  A265 );
 a21558a <=( A203  and  a21557a );
 a21562a <=( A302  and  (not A299) );
 a21563a <=( (not A298)  and  a21562a );
 a21564a <=( a21563a  and  a21558a );
 a21567a <=( (not A166)  and  (not A167) );
 a21571a <=( (not A201)  and  A200 );
 a21572a <=( A199  and  a21571a );
 a21573a <=( a21572a  and  a21567a );
 a21577a <=( A267  and  A266 );
 a21578a <=( A203  and  a21577a );
 a21582a <=( (not A301)  and  (not A299) );
 a21583a <=( (not A298)  and  a21582a );
 a21584a <=( a21583a  and  a21578a );
 a21587a <=( (not A166)  and  (not A167) );
 a21591a <=( (not A201)  and  A200 );
 a21592a <=( A199  and  a21591a );
 a21593a <=( a21592a  and  a21587a );
 a21597a <=( A267  and  A266 );
 a21598a <=( A203  and  a21597a );
 a21602a <=( A302  and  (not A299) );
 a21603a <=( (not A298)  and  a21602a );
 a21604a <=( a21603a  and  a21598a );
 a21607a <=( (not A166)  and  (not A167) );
 a21611a <=( (not A202)  and  A200 );
 a21612a <=( (not A199)  and  a21611a );
 a21613a <=( a21612a  and  a21607a );
 a21617a <=( (not A266)  and  (not A265) );
 a21618a <=( A203  and  a21617a );
 a21622a <=( A300  and  A299 );
 a21623a <=( (not A268)  and  a21622a );
 a21624a <=( a21623a  and  a21618a );
 a21627a <=( (not A166)  and  (not A167) );
 a21631a <=( (not A202)  and  A200 );
 a21632a <=( (not A199)  and  a21631a );
 a21633a <=( a21632a  and  a21627a );
 a21637a <=( (not A266)  and  (not A265) );
 a21638a <=( A203  and  a21637a );
 a21642a <=( A300  and  A298 );
 a21643a <=( (not A268)  and  a21642a );
 a21644a <=( a21643a  and  a21638a );
 a21647a <=( (not A166)  and  (not A167) );
 a21651a <=( (not A202)  and  A200 );
 a21652a <=( (not A199)  and  a21651a );
 a21653a <=( a21652a  and  a21647a );
 a21657a <=( (not A266)  and  (not A265) );
 a21658a <=( A203  and  a21657a );
 a21662a <=( A300  and  A299 );
 a21663a <=( A269  and  a21662a );
 a21664a <=( a21663a  and  a21658a );
 a21667a <=( (not A166)  and  (not A167) );
 a21671a <=( (not A202)  and  A200 );
 a21672a <=( (not A199)  and  a21671a );
 a21673a <=( a21672a  and  a21667a );
 a21677a <=( (not A266)  and  (not A265) );
 a21678a <=( A203  and  a21677a );
 a21682a <=( A300  and  A298 );
 a21683a <=( A269  and  a21682a );
 a21684a <=( a21683a  and  a21678a );
 a21687a <=( (not A166)  and  (not A167) );
 a21691a <=( (not A201)  and  A200 );
 a21692a <=( (not A199)  and  a21691a );
 a21693a <=( a21692a  and  a21687a );
 a21697a <=( A267  and  A265 );
 a21698a <=( A202  and  a21697a );
 a21702a <=( (not A301)  and  (not A299) );
 a21703a <=( (not A298)  and  a21702a );
 a21704a <=( a21703a  and  a21698a );
 a21707a <=( (not A166)  and  (not A167) );
 a21711a <=( (not A201)  and  A200 );
 a21712a <=( (not A199)  and  a21711a );
 a21713a <=( a21712a  and  a21707a );
 a21717a <=( A267  and  A265 );
 a21718a <=( A202  and  a21717a );
 a21722a <=( A302  and  (not A299) );
 a21723a <=( (not A298)  and  a21722a );
 a21724a <=( a21723a  and  a21718a );
 a21727a <=( (not A166)  and  (not A167) );
 a21731a <=( (not A201)  and  A200 );
 a21732a <=( (not A199)  and  a21731a );
 a21733a <=( a21732a  and  a21727a );
 a21737a <=( A267  and  A266 );
 a21738a <=( A202  and  a21737a );
 a21742a <=( (not A301)  and  (not A299) );
 a21743a <=( (not A298)  and  a21742a );
 a21744a <=( a21743a  and  a21738a );
 a21747a <=( (not A166)  and  (not A167) );
 a21751a <=( (not A201)  and  A200 );
 a21752a <=( (not A199)  and  a21751a );
 a21753a <=( a21752a  and  a21747a );
 a21757a <=( A267  and  A266 );
 a21758a <=( A202  and  a21757a );
 a21762a <=( A302  and  (not A299) );
 a21763a <=( (not A298)  and  a21762a );
 a21764a <=( a21763a  and  a21758a );
 a21767a <=( (not A166)  and  (not A167) );
 a21771a <=( (not A201)  and  A200 );
 a21772a <=( (not A199)  and  a21771a );
 a21773a <=( a21772a  and  a21767a );
 a21777a <=( A267  and  A265 );
 a21778a <=( (not A203)  and  a21777a );
 a21782a <=( (not A301)  and  (not A299) );
 a21783a <=( (not A298)  and  a21782a );
 a21784a <=( a21783a  and  a21778a );
 a21787a <=( (not A166)  and  (not A167) );
 a21791a <=( (not A201)  and  A200 );
 a21792a <=( (not A199)  and  a21791a );
 a21793a <=( a21792a  and  a21787a );
 a21797a <=( A267  and  A265 );
 a21798a <=( (not A203)  and  a21797a );
 a21802a <=( A302  and  (not A299) );
 a21803a <=( (not A298)  and  a21802a );
 a21804a <=( a21803a  and  a21798a );
 a21807a <=( (not A166)  and  (not A167) );
 a21811a <=( (not A201)  and  A200 );
 a21812a <=( (not A199)  and  a21811a );
 a21813a <=( a21812a  and  a21807a );
 a21817a <=( A267  and  A266 );
 a21818a <=( (not A203)  and  a21817a );
 a21822a <=( (not A301)  and  (not A299) );
 a21823a <=( (not A298)  and  a21822a );
 a21824a <=( a21823a  and  a21818a );
 a21827a <=( (not A166)  and  (not A167) );
 a21831a <=( (not A201)  and  A200 );
 a21832a <=( (not A199)  and  a21831a );
 a21833a <=( a21832a  and  a21827a );
 a21837a <=( A267  and  A266 );
 a21838a <=( (not A203)  and  a21837a );
 a21842a <=( A302  and  (not A299) );
 a21843a <=( (not A298)  and  a21842a );
 a21844a <=( a21843a  and  a21838a );
 a21847a <=( (not A166)  and  (not A167) );
 a21851a <=( (not A202)  and  (not A200) );
 a21852a <=( A199  and  a21851a );
 a21853a <=( a21852a  and  a21847a );
 a21857a <=( (not A266)  and  (not A265) );
 a21858a <=( A203  and  a21857a );
 a21862a <=( A300  and  A299 );
 a21863a <=( (not A268)  and  a21862a );
 a21864a <=( a21863a  and  a21858a );
 a21867a <=( (not A166)  and  (not A167) );
 a21871a <=( (not A202)  and  (not A200) );
 a21872a <=( A199  and  a21871a );
 a21873a <=( a21872a  and  a21867a );
 a21877a <=( (not A266)  and  (not A265) );
 a21878a <=( A203  and  a21877a );
 a21882a <=( A300  and  A298 );
 a21883a <=( (not A268)  and  a21882a );
 a21884a <=( a21883a  and  a21878a );
 a21887a <=( (not A166)  and  (not A167) );
 a21891a <=( (not A202)  and  (not A200) );
 a21892a <=( A199  and  a21891a );
 a21893a <=( a21892a  and  a21887a );
 a21897a <=( (not A266)  and  (not A265) );
 a21898a <=( A203  and  a21897a );
 a21902a <=( A300  and  A299 );
 a21903a <=( A269  and  a21902a );
 a21904a <=( a21903a  and  a21898a );
 a21907a <=( (not A166)  and  (not A167) );
 a21911a <=( (not A202)  and  (not A200) );
 a21912a <=( A199  and  a21911a );
 a21913a <=( a21912a  and  a21907a );
 a21917a <=( (not A266)  and  (not A265) );
 a21918a <=( A203  and  a21917a );
 a21922a <=( A300  and  A298 );
 a21923a <=( A269  and  a21922a );
 a21924a <=( a21923a  and  a21918a );
 a21927a <=( (not A166)  and  (not A167) );
 a21931a <=( (not A201)  and  (not A200) );
 a21932a <=( A199  and  a21931a );
 a21933a <=( a21932a  and  a21927a );
 a21937a <=( A267  and  A265 );
 a21938a <=( A202  and  a21937a );
 a21942a <=( (not A301)  and  (not A299) );
 a21943a <=( (not A298)  and  a21942a );
 a21944a <=( a21943a  and  a21938a );
 a21947a <=( (not A166)  and  (not A167) );
 a21951a <=( (not A201)  and  (not A200) );
 a21952a <=( A199  and  a21951a );
 a21953a <=( a21952a  and  a21947a );
 a21957a <=( A267  and  A265 );
 a21958a <=( A202  and  a21957a );
 a21962a <=( A302  and  (not A299) );
 a21963a <=( (not A298)  and  a21962a );
 a21964a <=( a21963a  and  a21958a );
 a21967a <=( (not A166)  and  (not A167) );
 a21971a <=( (not A201)  and  (not A200) );
 a21972a <=( A199  and  a21971a );
 a21973a <=( a21972a  and  a21967a );
 a21977a <=( A267  and  A266 );
 a21978a <=( A202  and  a21977a );
 a21982a <=( (not A301)  and  (not A299) );
 a21983a <=( (not A298)  and  a21982a );
 a21984a <=( a21983a  and  a21978a );
 a21987a <=( (not A166)  and  (not A167) );
 a21991a <=( (not A201)  and  (not A200) );
 a21992a <=( A199  and  a21991a );
 a21993a <=( a21992a  and  a21987a );
 a21997a <=( A267  and  A266 );
 a21998a <=( A202  and  a21997a );
 a22002a <=( A302  and  (not A299) );
 a22003a <=( (not A298)  and  a22002a );
 a22004a <=( a22003a  and  a21998a );
 a22007a <=( (not A166)  and  (not A167) );
 a22011a <=( (not A201)  and  (not A200) );
 a22012a <=( A199  and  a22011a );
 a22013a <=( a22012a  and  a22007a );
 a22017a <=( A267  and  A265 );
 a22018a <=( (not A203)  and  a22017a );
 a22022a <=( (not A301)  and  (not A299) );
 a22023a <=( (not A298)  and  a22022a );
 a22024a <=( a22023a  and  a22018a );
 a22027a <=( (not A166)  and  (not A167) );
 a22031a <=( (not A201)  and  (not A200) );
 a22032a <=( A199  and  a22031a );
 a22033a <=( a22032a  and  a22027a );
 a22037a <=( A267  and  A265 );
 a22038a <=( (not A203)  and  a22037a );
 a22042a <=( A302  and  (not A299) );
 a22043a <=( (not A298)  and  a22042a );
 a22044a <=( a22043a  and  a22038a );
 a22047a <=( (not A166)  and  (not A167) );
 a22051a <=( (not A201)  and  (not A200) );
 a22052a <=( A199  and  a22051a );
 a22053a <=( a22052a  and  a22047a );
 a22057a <=( A267  and  A266 );
 a22058a <=( (not A203)  and  a22057a );
 a22062a <=( (not A301)  and  (not A299) );
 a22063a <=( (not A298)  and  a22062a );
 a22064a <=( a22063a  and  a22058a );
 a22067a <=( (not A166)  and  (not A167) );
 a22071a <=( (not A201)  and  (not A200) );
 a22072a <=( A199  and  a22071a );
 a22073a <=( a22072a  and  a22067a );
 a22077a <=( A267  and  A266 );
 a22078a <=( (not A203)  and  a22077a );
 a22082a <=( A302  and  (not A299) );
 a22083a <=( (not A298)  and  a22082a );
 a22084a <=( a22083a  and  a22078a );
 a22087a <=( (not A166)  and  (not A167) );
 a22091a <=( (not A202)  and  (not A200) );
 a22092a <=( (not A199)  and  a22091a );
 a22093a <=( a22092a  and  a22087a );
 a22097a <=( A298  and  A267 );
 a22098a <=( A265  and  a22097a );
 a22102a <=( (not A301)  and  (not A300) );
 a22103a <=( A299  and  a22102a );
 a22104a <=( a22103a  and  a22098a );
 a22107a <=( (not A166)  and  (not A167) );
 a22111a <=( (not A202)  and  (not A200) );
 a22112a <=( (not A199)  and  a22111a );
 a22113a <=( a22112a  and  a22107a );
 a22117a <=( A298  and  A267 );
 a22118a <=( A265  and  a22117a );
 a22122a <=( A302  and  (not A300) );
 a22123a <=( A299  and  a22122a );
 a22124a <=( a22123a  and  a22118a );
 a22127a <=( (not A166)  and  (not A167) );
 a22131a <=( (not A202)  and  (not A200) );
 a22132a <=( (not A199)  and  a22131a );
 a22133a <=( a22132a  and  a22127a );
 a22137a <=( A298  and  A267 );
 a22138a <=( A265  and  a22137a );
 a22142a <=( A301  and  (not A300) );
 a22143a <=( (not A299)  and  a22142a );
 a22144a <=( a22143a  and  a22138a );
 a22147a <=( (not A166)  and  (not A167) );
 a22151a <=( (not A202)  and  (not A200) );
 a22152a <=( (not A199)  and  a22151a );
 a22153a <=( a22152a  and  a22147a );
 a22157a <=( A298  and  A267 );
 a22158a <=( A265  and  a22157a );
 a22162a <=( (not A302)  and  (not A300) );
 a22163a <=( (not A299)  and  a22162a );
 a22164a <=( a22163a  and  a22158a );
 a22167a <=( (not A166)  and  (not A167) );
 a22171a <=( (not A202)  and  (not A200) );
 a22172a <=( (not A199)  and  a22171a );
 a22173a <=( a22172a  and  a22167a );
 a22177a <=( (not A298)  and  A267 );
 a22178a <=( A265  and  a22177a );
 a22182a <=( A301  and  (not A300) );
 a22183a <=( A299  and  a22182a );
 a22184a <=( a22183a  and  a22178a );
 a22187a <=( (not A166)  and  (not A167) );
 a22191a <=( (not A202)  and  (not A200) );
 a22192a <=( (not A199)  and  a22191a );
 a22193a <=( a22192a  and  a22187a );
 a22197a <=( (not A298)  and  A267 );
 a22198a <=( A265  and  a22197a );
 a22202a <=( (not A302)  and  (not A300) );
 a22203a <=( A299  and  a22202a );
 a22204a <=( a22203a  and  a22198a );
 a22207a <=( (not A166)  and  (not A167) );
 a22211a <=( (not A202)  and  (not A200) );
 a22212a <=( (not A199)  and  a22211a );
 a22213a <=( a22212a  and  a22207a );
 a22217a <=( A298  and  A267 );
 a22218a <=( A266  and  a22217a );
 a22222a <=( (not A301)  and  (not A300) );
 a22223a <=( A299  and  a22222a );
 a22224a <=( a22223a  and  a22218a );
 a22227a <=( (not A166)  and  (not A167) );
 a22231a <=( (not A202)  and  (not A200) );
 a22232a <=( (not A199)  and  a22231a );
 a22233a <=( a22232a  and  a22227a );
 a22237a <=( A298  and  A267 );
 a22238a <=( A266  and  a22237a );
 a22242a <=( A302  and  (not A300) );
 a22243a <=( A299  and  a22242a );
 a22244a <=( a22243a  and  a22238a );
 a22247a <=( (not A166)  and  (not A167) );
 a22251a <=( (not A202)  and  (not A200) );
 a22252a <=( (not A199)  and  a22251a );
 a22253a <=( a22252a  and  a22247a );
 a22257a <=( A298  and  A267 );
 a22258a <=( A266  and  a22257a );
 a22262a <=( A301  and  (not A300) );
 a22263a <=( (not A299)  and  a22262a );
 a22264a <=( a22263a  and  a22258a );
 a22267a <=( (not A166)  and  (not A167) );
 a22271a <=( (not A202)  and  (not A200) );
 a22272a <=( (not A199)  and  a22271a );
 a22273a <=( a22272a  and  a22267a );
 a22277a <=( A298  and  A267 );
 a22278a <=( A266  and  a22277a );
 a22282a <=( (not A302)  and  (not A300) );
 a22283a <=( (not A299)  and  a22282a );
 a22284a <=( a22283a  and  a22278a );
 a22287a <=( (not A166)  and  (not A167) );
 a22291a <=( (not A202)  and  (not A200) );
 a22292a <=( (not A199)  and  a22291a );
 a22293a <=( a22292a  and  a22287a );
 a22297a <=( (not A298)  and  A267 );
 a22298a <=( A266  and  a22297a );
 a22302a <=( A301  and  (not A300) );
 a22303a <=( A299  and  a22302a );
 a22304a <=( a22303a  and  a22298a );
 a22307a <=( (not A166)  and  (not A167) );
 a22311a <=( (not A202)  and  (not A200) );
 a22312a <=( (not A199)  and  a22311a );
 a22313a <=( a22312a  and  a22307a );
 a22317a <=( (not A298)  and  A267 );
 a22318a <=( A266  and  a22317a );
 a22322a <=( (not A302)  and  (not A300) );
 a22323a <=( A299  and  a22322a );
 a22324a <=( a22323a  and  a22318a );
 a22327a <=( (not A166)  and  (not A167) );
 a22331a <=( A203  and  (not A200) );
 a22332a <=( (not A199)  and  a22331a );
 a22333a <=( a22332a  and  a22327a );
 a22337a <=( A298  and  A267 );
 a22338a <=( A265  and  a22337a );
 a22342a <=( (not A301)  and  (not A300) );
 a22343a <=( A299  and  a22342a );
 a22344a <=( a22343a  and  a22338a );
 a22347a <=( (not A166)  and  (not A167) );
 a22351a <=( A203  and  (not A200) );
 a22352a <=( (not A199)  and  a22351a );
 a22353a <=( a22352a  and  a22347a );
 a22357a <=( A298  and  A267 );
 a22358a <=( A265  and  a22357a );
 a22362a <=( A302  and  (not A300) );
 a22363a <=( A299  and  a22362a );
 a22364a <=( a22363a  and  a22358a );
 a22367a <=( (not A166)  and  (not A167) );
 a22371a <=( A203  and  (not A200) );
 a22372a <=( (not A199)  and  a22371a );
 a22373a <=( a22372a  and  a22367a );
 a22377a <=( A298  and  A267 );
 a22378a <=( A265  and  a22377a );
 a22382a <=( A301  and  (not A300) );
 a22383a <=( (not A299)  and  a22382a );
 a22384a <=( a22383a  and  a22378a );
 a22387a <=( (not A166)  and  (not A167) );
 a22391a <=( A203  and  (not A200) );
 a22392a <=( (not A199)  and  a22391a );
 a22393a <=( a22392a  and  a22387a );
 a22397a <=( A298  and  A267 );
 a22398a <=( A265  and  a22397a );
 a22402a <=( (not A302)  and  (not A300) );
 a22403a <=( (not A299)  and  a22402a );
 a22404a <=( a22403a  and  a22398a );
 a22407a <=( (not A166)  and  (not A167) );
 a22411a <=( A203  and  (not A200) );
 a22412a <=( (not A199)  and  a22411a );
 a22413a <=( a22412a  and  a22407a );
 a22417a <=( (not A298)  and  A267 );
 a22418a <=( A265  and  a22417a );
 a22422a <=( A301  and  (not A300) );
 a22423a <=( A299  and  a22422a );
 a22424a <=( a22423a  and  a22418a );
 a22427a <=( (not A166)  and  (not A167) );
 a22431a <=( A203  and  (not A200) );
 a22432a <=( (not A199)  and  a22431a );
 a22433a <=( a22432a  and  a22427a );
 a22437a <=( (not A298)  and  A267 );
 a22438a <=( A265  and  a22437a );
 a22442a <=( (not A302)  and  (not A300) );
 a22443a <=( A299  and  a22442a );
 a22444a <=( a22443a  and  a22438a );
 a22447a <=( (not A166)  and  (not A167) );
 a22451a <=( A203  and  (not A200) );
 a22452a <=( (not A199)  and  a22451a );
 a22453a <=( a22452a  and  a22447a );
 a22457a <=( A298  and  A267 );
 a22458a <=( A266  and  a22457a );
 a22462a <=( (not A301)  and  (not A300) );
 a22463a <=( A299  and  a22462a );
 a22464a <=( a22463a  and  a22458a );
 a22467a <=( (not A166)  and  (not A167) );
 a22471a <=( A203  and  (not A200) );
 a22472a <=( (not A199)  and  a22471a );
 a22473a <=( a22472a  and  a22467a );
 a22477a <=( A298  and  A267 );
 a22478a <=( A266  and  a22477a );
 a22482a <=( A302  and  (not A300) );
 a22483a <=( A299  and  a22482a );
 a22484a <=( a22483a  and  a22478a );
 a22487a <=( (not A166)  and  (not A167) );
 a22491a <=( A203  and  (not A200) );
 a22492a <=( (not A199)  and  a22491a );
 a22493a <=( a22492a  and  a22487a );
 a22497a <=( A298  and  A267 );
 a22498a <=( A266  and  a22497a );
 a22502a <=( A301  and  (not A300) );
 a22503a <=( (not A299)  and  a22502a );
 a22504a <=( a22503a  and  a22498a );
 a22507a <=( (not A166)  and  (not A167) );
 a22511a <=( A203  and  (not A200) );
 a22512a <=( (not A199)  and  a22511a );
 a22513a <=( a22512a  and  a22507a );
 a22517a <=( A298  and  A267 );
 a22518a <=( A266  and  a22517a );
 a22522a <=( (not A302)  and  (not A300) );
 a22523a <=( (not A299)  and  a22522a );
 a22524a <=( a22523a  and  a22518a );
 a22527a <=( (not A166)  and  (not A167) );
 a22531a <=( A203  and  (not A200) );
 a22532a <=( (not A199)  and  a22531a );
 a22533a <=( a22532a  and  a22527a );
 a22537a <=( (not A298)  and  A267 );
 a22538a <=( A266  and  a22537a );
 a22542a <=( A301  and  (not A300) );
 a22543a <=( A299  and  a22542a );
 a22544a <=( a22543a  and  a22538a );
 a22547a <=( (not A166)  and  (not A167) );
 a22551a <=( A203  and  (not A200) );
 a22552a <=( (not A199)  and  a22551a );
 a22553a <=( a22552a  and  a22547a );
 a22557a <=( (not A298)  and  A267 );
 a22558a <=( A266  and  a22557a );
 a22562a <=( (not A302)  and  (not A300) );
 a22563a <=( A299  and  a22562a );
 a22564a <=( a22563a  and  a22558a );
 a22567a <=( (not A166)  and  (not A167) );
 a22571a <=( A202  and  (not A200) );
 a22572a <=( (not A199)  and  a22571a );
 a22573a <=( a22572a  and  a22567a );
 a22577a <=( (not A266)  and  (not A265) );
 a22578a <=( (not A203)  and  a22577a );
 a22582a <=( A300  and  A299 );
 a22583a <=( (not A268)  and  a22582a );
 a22584a <=( a22583a  and  a22578a );
 a22587a <=( (not A166)  and  (not A167) );
 a22591a <=( A202  and  (not A200) );
 a22592a <=( (not A199)  and  a22591a );
 a22593a <=( a22592a  and  a22587a );
 a22597a <=( (not A266)  and  (not A265) );
 a22598a <=( (not A203)  and  a22597a );
 a22602a <=( A300  and  A298 );
 a22603a <=( (not A268)  and  a22602a );
 a22604a <=( a22603a  and  a22598a );
 a22607a <=( (not A166)  and  (not A167) );
 a22611a <=( A202  and  (not A200) );
 a22612a <=( (not A199)  and  a22611a );
 a22613a <=( a22612a  and  a22607a );
 a22617a <=( (not A266)  and  (not A265) );
 a22618a <=( (not A203)  and  a22617a );
 a22622a <=( A300  and  A299 );
 a22623a <=( A269  and  a22622a );
 a22624a <=( a22623a  and  a22618a );
 a22627a <=( (not A166)  and  (not A167) );
 a22631a <=( A202  and  (not A200) );
 a22632a <=( (not A199)  and  a22631a );
 a22633a <=( a22632a  and  a22627a );
 a22637a <=( (not A266)  and  (not A265) );
 a22638a <=( (not A203)  and  a22637a );
 a22642a <=( A300  and  A298 );
 a22643a <=( A269  and  a22642a );
 a22644a <=( a22643a  and  a22638a );
 a22647a <=( (not A167)  and  (not A168) );
 a22651a <=( (not A265)  and  A201 );
 a22652a <=( A199  and  a22651a );
 a22653a <=( a22652a  and  a22647a );
 a22657a <=( A298  and  (not A268) );
 a22658a <=( (not A266)  and  a22657a );
 a22662a <=( (not A302)  and  A301 );
 a22663a <=( A299  and  a22662a );
 a22664a <=( a22663a  and  a22658a );
 a22667a <=( (not A167)  and  (not A168) );
 a22671a <=( (not A265)  and  A201 );
 a22672a <=( A199  and  a22671a );
 a22673a <=( a22672a  and  a22667a );
 a22677a <=( A298  and  (not A268) );
 a22678a <=( (not A266)  and  a22677a );
 a22682a <=( A302  and  (not A301) );
 a22683a <=( (not A299)  and  a22682a );
 a22684a <=( a22683a  and  a22678a );
 a22687a <=( (not A167)  and  (not A168) );
 a22691a <=( (not A265)  and  A201 );
 a22692a <=( A199  and  a22691a );
 a22693a <=( a22692a  and  a22687a );
 a22697a <=( (not A298)  and  (not A268) );
 a22698a <=( (not A266)  and  a22697a );
 a22702a <=( A302  and  (not A301) );
 a22703a <=( A299  and  a22702a );
 a22704a <=( a22703a  and  a22698a );
 a22707a <=( (not A167)  and  (not A168) );
 a22711a <=( (not A265)  and  A201 );
 a22712a <=( A199  and  a22711a );
 a22713a <=( a22712a  and  a22707a );
 a22717a <=( (not A298)  and  (not A268) );
 a22718a <=( (not A266)  and  a22717a );
 a22722a <=( (not A302)  and  A301 );
 a22723a <=( (not A299)  and  a22722a );
 a22724a <=( a22723a  and  a22718a );
 a22727a <=( (not A167)  and  (not A168) );
 a22731a <=( (not A265)  and  A201 );
 a22732a <=( A199  and  a22731a );
 a22733a <=( a22732a  and  a22727a );
 a22737a <=( A298  and  A269 );
 a22738a <=( (not A266)  and  a22737a );
 a22742a <=( (not A302)  and  A301 );
 a22743a <=( A299  and  a22742a );
 a22744a <=( a22743a  and  a22738a );
 a22747a <=( (not A167)  and  (not A168) );
 a22751a <=( (not A265)  and  A201 );
 a22752a <=( A199  and  a22751a );
 a22753a <=( a22752a  and  a22747a );
 a22757a <=( A298  and  A269 );
 a22758a <=( (not A266)  and  a22757a );
 a22762a <=( A302  and  (not A301) );
 a22763a <=( (not A299)  and  a22762a );
 a22764a <=( a22763a  and  a22758a );
 a22767a <=( (not A167)  and  (not A168) );
 a22771a <=( (not A265)  and  A201 );
 a22772a <=( A199  and  a22771a );
 a22773a <=( a22772a  and  a22767a );
 a22777a <=( (not A298)  and  A269 );
 a22778a <=( (not A266)  and  a22777a );
 a22782a <=( A302  and  (not A301) );
 a22783a <=( A299  and  a22782a );
 a22784a <=( a22783a  and  a22778a );
 a22787a <=( (not A167)  and  (not A168) );
 a22791a <=( (not A265)  and  A201 );
 a22792a <=( A199  and  a22791a );
 a22793a <=( a22792a  and  a22787a );
 a22797a <=( (not A298)  and  A269 );
 a22798a <=( (not A266)  and  a22797a );
 a22802a <=( (not A302)  and  A301 );
 a22803a <=( (not A299)  and  a22802a );
 a22804a <=( a22803a  and  a22798a );
 a22807a <=( (not A167)  and  (not A168) );
 a22811a <=( (not A265)  and  A201 );
 a22812a <=( A200  and  a22811a );
 a22813a <=( a22812a  and  a22807a );
 a22817a <=( A298  and  (not A268) );
 a22818a <=( (not A266)  and  a22817a );
 a22822a <=( (not A302)  and  A301 );
 a22823a <=( A299  and  a22822a );
 a22824a <=( a22823a  and  a22818a );
 a22827a <=( (not A167)  and  (not A168) );
 a22831a <=( (not A265)  and  A201 );
 a22832a <=( A200  and  a22831a );
 a22833a <=( a22832a  and  a22827a );
 a22837a <=( A298  and  (not A268) );
 a22838a <=( (not A266)  and  a22837a );
 a22842a <=( A302  and  (not A301) );
 a22843a <=( (not A299)  and  a22842a );
 a22844a <=( a22843a  and  a22838a );
 a22847a <=( (not A167)  and  (not A168) );
 a22851a <=( (not A265)  and  A201 );
 a22852a <=( A200  and  a22851a );
 a22853a <=( a22852a  and  a22847a );
 a22857a <=( (not A298)  and  (not A268) );
 a22858a <=( (not A266)  and  a22857a );
 a22862a <=( A302  and  (not A301) );
 a22863a <=( A299  and  a22862a );
 a22864a <=( a22863a  and  a22858a );
 a22867a <=( (not A167)  and  (not A168) );
 a22871a <=( (not A265)  and  A201 );
 a22872a <=( A200  and  a22871a );
 a22873a <=( a22872a  and  a22867a );
 a22877a <=( (not A298)  and  (not A268) );
 a22878a <=( (not A266)  and  a22877a );
 a22882a <=( (not A302)  and  A301 );
 a22883a <=( (not A299)  and  a22882a );
 a22884a <=( a22883a  and  a22878a );
 a22887a <=( (not A167)  and  (not A168) );
 a22891a <=( (not A265)  and  A201 );
 a22892a <=( A200  and  a22891a );
 a22893a <=( a22892a  and  a22887a );
 a22897a <=( A298  and  A269 );
 a22898a <=( (not A266)  and  a22897a );
 a22902a <=( (not A302)  and  A301 );
 a22903a <=( A299  and  a22902a );
 a22904a <=( a22903a  and  a22898a );
 a22907a <=( (not A167)  and  (not A168) );
 a22911a <=( (not A265)  and  A201 );
 a22912a <=( A200  and  a22911a );
 a22913a <=( a22912a  and  a22907a );
 a22917a <=( A298  and  A269 );
 a22918a <=( (not A266)  and  a22917a );
 a22922a <=( A302  and  (not A301) );
 a22923a <=( (not A299)  and  a22922a );
 a22924a <=( a22923a  and  a22918a );
 a22927a <=( (not A167)  and  (not A168) );
 a22931a <=( (not A265)  and  A201 );
 a22932a <=( A200  and  a22931a );
 a22933a <=( a22932a  and  a22927a );
 a22937a <=( (not A298)  and  A269 );
 a22938a <=( (not A266)  and  a22937a );
 a22942a <=( A302  and  (not A301) );
 a22943a <=( A299  and  a22942a );
 a22944a <=( a22943a  and  a22938a );
 a22947a <=( (not A167)  and  (not A168) );
 a22951a <=( (not A265)  and  A201 );
 a22952a <=( A200  and  a22951a );
 a22953a <=( a22952a  and  a22947a );
 a22957a <=( (not A298)  and  A269 );
 a22958a <=( (not A266)  and  a22957a );
 a22962a <=( (not A302)  and  A301 );
 a22963a <=( (not A299)  and  a22962a );
 a22964a <=( a22963a  and  a22958a );
 a22967a <=( (not A167)  and  (not A168) );
 a22971a <=( A202  and  A200 );
 a22972a <=( A199  and  a22971a );
 a22973a <=( a22972a  and  a22967a );
 a22977a <=( (not A266)  and  (not A265) );
 a22978a <=( (not A203)  and  a22977a );
 a22982a <=( A300  and  A299 );
 a22983a <=( (not A268)  and  a22982a );
 a22984a <=( a22983a  and  a22978a );
 a22987a <=( (not A167)  and  (not A168) );
 a22991a <=( A202  and  A200 );
 a22992a <=( A199  and  a22991a );
 a22993a <=( a22992a  and  a22987a );
 a22997a <=( (not A266)  and  (not A265) );
 a22998a <=( (not A203)  and  a22997a );
 a23002a <=( A300  and  A298 );
 a23003a <=( (not A268)  and  a23002a );
 a23004a <=( a23003a  and  a22998a );
 a23007a <=( (not A167)  and  (not A168) );
 a23011a <=( A202  and  A200 );
 a23012a <=( A199  and  a23011a );
 a23013a <=( a23012a  and  a23007a );
 a23017a <=( (not A266)  and  (not A265) );
 a23018a <=( (not A203)  and  a23017a );
 a23022a <=( A300  and  A299 );
 a23023a <=( A269  and  a23022a );
 a23024a <=( a23023a  and  a23018a );
 a23027a <=( (not A167)  and  (not A168) );
 a23031a <=( A202  and  A200 );
 a23032a <=( A199  and  a23031a );
 a23033a <=( a23032a  and  a23027a );
 a23037a <=( (not A266)  and  (not A265) );
 a23038a <=( (not A203)  and  a23037a );
 a23042a <=( A300  and  A298 );
 a23043a <=( A269  and  a23042a );
 a23044a <=( a23043a  and  a23038a );
 a23047a <=( (not A167)  and  (not A168) );
 a23051a <=( (not A201)  and  A200 );
 a23052a <=( A199  and  a23051a );
 a23053a <=( a23052a  and  a23047a );
 a23057a <=( A267  and  A265 );
 a23058a <=( (not A202)  and  a23057a );
 a23062a <=( (not A301)  and  (not A299) );
 a23063a <=( (not A298)  and  a23062a );
 a23064a <=( a23063a  and  a23058a );
 a23067a <=( (not A167)  and  (not A168) );
 a23071a <=( (not A201)  and  A200 );
 a23072a <=( A199  and  a23071a );
 a23073a <=( a23072a  and  a23067a );
 a23077a <=( A267  and  A265 );
 a23078a <=( (not A202)  and  a23077a );
 a23082a <=( A302  and  (not A299) );
 a23083a <=( (not A298)  and  a23082a );
 a23084a <=( a23083a  and  a23078a );
 a23087a <=( (not A167)  and  (not A168) );
 a23091a <=( (not A201)  and  A200 );
 a23092a <=( A199  and  a23091a );
 a23093a <=( a23092a  and  a23087a );
 a23097a <=( A267  and  A266 );
 a23098a <=( (not A202)  and  a23097a );
 a23102a <=( (not A301)  and  (not A299) );
 a23103a <=( (not A298)  and  a23102a );
 a23104a <=( a23103a  and  a23098a );
 a23107a <=( (not A167)  and  (not A168) );
 a23111a <=( (not A201)  and  A200 );
 a23112a <=( A199  and  a23111a );
 a23113a <=( a23112a  and  a23107a );
 a23117a <=( A267  and  A266 );
 a23118a <=( (not A202)  and  a23117a );
 a23122a <=( A302  and  (not A299) );
 a23123a <=( (not A298)  and  a23122a );
 a23124a <=( a23123a  and  a23118a );
 a23127a <=( (not A167)  and  (not A168) );
 a23131a <=( (not A201)  and  A200 );
 a23132a <=( A199  and  a23131a );
 a23133a <=( a23132a  and  a23127a );
 a23137a <=( A267  and  A265 );
 a23138a <=( A203  and  a23137a );
 a23142a <=( (not A301)  and  (not A299) );
 a23143a <=( (not A298)  and  a23142a );
 a23144a <=( a23143a  and  a23138a );
 a23147a <=( (not A167)  and  (not A168) );
 a23151a <=( (not A201)  and  A200 );
 a23152a <=( A199  and  a23151a );
 a23153a <=( a23152a  and  a23147a );
 a23157a <=( A267  and  A265 );
 a23158a <=( A203  and  a23157a );
 a23162a <=( A302  and  (not A299) );
 a23163a <=( (not A298)  and  a23162a );
 a23164a <=( a23163a  and  a23158a );
 a23167a <=( (not A167)  and  (not A168) );
 a23171a <=( (not A201)  and  A200 );
 a23172a <=( A199  and  a23171a );
 a23173a <=( a23172a  and  a23167a );
 a23177a <=( A267  and  A266 );
 a23178a <=( A203  and  a23177a );
 a23182a <=( (not A301)  and  (not A299) );
 a23183a <=( (not A298)  and  a23182a );
 a23184a <=( a23183a  and  a23178a );
 a23187a <=( (not A167)  and  (not A168) );
 a23191a <=( (not A201)  and  A200 );
 a23192a <=( A199  and  a23191a );
 a23193a <=( a23192a  and  a23187a );
 a23197a <=( A267  and  A266 );
 a23198a <=( A203  and  a23197a );
 a23202a <=( A302  and  (not A299) );
 a23203a <=( (not A298)  and  a23202a );
 a23204a <=( a23203a  and  a23198a );
 a23207a <=( (not A167)  and  (not A168) );
 a23211a <=( (not A202)  and  A200 );
 a23212a <=( (not A199)  and  a23211a );
 a23213a <=( a23212a  and  a23207a );
 a23217a <=( (not A266)  and  (not A265) );
 a23218a <=( A203  and  a23217a );
 a23222a <=( A300  and  A299 );
 a23223a <=( (not A268)  and  a23222a );
 a23224a <=( a23223a  and  a23218a );
 a23227a <=( (not A167)  and  (not A168) );
 a23231a <=( (not A202)  and  A200 );
 a23232a <=( (not A199)  and  a23231a );
 a23233a <=( a23232a  and  a23227a );
 a23237a <=( (not A266)  and  (not A265) );
 a23238a <=( A203  and  a23237a );
 a23242a <=( A300  and  A298 );
 a23243a <=( (not A268)  and  a23242a );
 a23244a <=( a23243a  and  a23238a );
 a23247a <=( (not A167)  and  (not A168) );
 a23251a <=( (not A202)  and  A200 );
 a23252a <=( (not A199)  and  a23251a );
 a23253a <=( a23252a  and  a23247a );
 a23257a <=( (not A266)  and  (not A265) );
 a23258a <=( A203  and  a23257a );
 a23262a <=( A300  and  A299 );
 a23263a <=( A269  and  a23262a );
 a23264a <=( a23263a  and  a23258a );
 a23267a <=( (not A167)  and  (not A168) );
 a23271a <=( (not A202)  and  A200 );
 a23272a <=( (not A199)  and  a23271a );
 a23273a <=( a23272a  and  a23267a );
 a23277a <=( (not A266)  and  (not A265) );
 a23278a <=( A203  and  a23277a );
 a23282a <=( A300  and  A298 );
 a23283a <=( A269  and  a23282a );
 a23284a <=( a23283a  and  a23278a );
 a23287a <=( (not A167)  and  (not A168) );
 a23291a <=( (not A201)  and  A200 );
 a23292a <=( (not A199)  and  a23291a );
 a23293a <=( a23292a  and  a23287a );
 a23297a <=( A267  and  A265 );
 a23298a <=( A202  and  a23297a );
 a23302a <=( (not A301)  and  (not A299) );
 a23303a <=( (not A298)  and  a23302a );
 a23304a <=( a23303a  and  a23298a );
 a23307a <=( (not A167)  and  (not A168) );
 a23311a <=( (not A201)  and  A200 );
 a23312a <=( (not A199)  and  a23311a );
 a23313a <=( a23312a  and  a23307a );
 a23317a <=( A267  and  A265 );
 a23318a <=( A202  and  a23317a );
 a23322a <=( A302  and  (not A299) );
 a23323a <=( (not A298)  and  a23322a );
 a23324a <=( a23323a  and  a23318a );
 a23327a <=( (not A167)  and  (not A168) );
 a23331a <=( (not A201)  and  A200 );
 a23332a <=( (not A199)  and  a23331a );
 a23333a <=( a23332a  and  a23327a );
 a23337a <=( A267  and  A266 );
 a23338a <=( A202  and  a23337a );
 a23342a <=( (not A301)  and  (not A299) );
 a23343a <=( (not A298)  and  a23342a );
 a23344a <=( a23343a  and  a23338a );
 a23347a <=( (not A167)  and  (not A168) );
 a23351a <=( (not A201)  and  A200 );
 a23352a <=( (not A199)  and  a23351a );
 a23353a <=( a23352a  and  a23347a );
 a23357a <=( A267  and  A266 );
 a23358a <=( A202  and  a23357a );
 a23362a <=( A302  and  (not A299) );
 a23363a <=( (not A298)  and  a23362a );
 a23364a <=( a23363a  and  a23358a );
 a23367a <=( (not A167)  and  (not A168) );
 a23371a <=( (not A201)  and  A200 );
 a23372a <=( (not A199)  and  a23371a );
 a23373a <=( a23372a  and  a23367a );
 a23377a <=( A267  and  A265 );
 a23378a <=( (not A203)  and  a23377a );
 a23382a <=( (not A301)  and  (not A299) );
 a23383a <=( (not A298)  and  a23382a );
 a23384a <=( a23383a  and  a23378a );
 a23387a <=( (not A167)  and  (not A168) );
 a23391a <=( (not A201)  and  A200 );
 a23392a <=( (not A199)  and  a23391a );
 a23393a <=( a23392a  and  a23387a );
 a23397a <=( A267  and  A265 );
 a23398a <=( (not A203)  and  a23397a );
 a23402a <=( A302  and  (not A299) );
 a23403a <=( (not A298)  and  a23402a );
 a23404a <=( a23403a  and  a23398a );
 a23407a <=( (not A167)  and  (not A168) );
 a23411a <=( (not A201)  and  A200 );
 a23412a <=( (not A199)  and  a23411a );
 a23413a <=( a23412a  and  a23407a );
 a23417a <=( A267  and  A266 );
 a23418a <=( (not A203)  and  a23417a );
 a23422a <=( (not A301)  and  (not A299) );
 a23423a <=( (not A298)  and  a23422a );
 a23424a <=( a23423a  and  a23418a );
 a23427a <=( (not A167)  and  (not A168) );
 a23431a <=( (not A201)  and  A200 );
 a23432a <=( (not A199)  and  a23431a );
 a23433a <=( a23432a  and  a23427a );
 a23437a <=( A267  and  A266 );
 a23438a <=( (not A203)  and  a23437a );
 a23442a <=( A302  and  (not A299) );
 a23443a <=( (not A298)  and  a23442a );
 a23444a <=( a23443a  and  a23438a );
 a23447a <=( (not A167)  and  (not A168) );
 a23451a <=( (not A202)  and  (not A200) );
 a23452a <=( A199  and  a23451a );
 a23453a <=( a23452a  and  a23447a );
 a23457a <=( (not A266)  and  (not A265) );
 a23458a <=( A203  and  a23457a );
 a23462a <=( A300  and  A299 );
 a23463a <=( (not A268)  and  a23462a );
 a23464a <=( a23463a  and  a23458a );
 a23467a <=( (not A167)  and  (not A168) );
 a23471a <=( (not A202)  and  (not A200) );
 a23472a <=( A199  and  a23471a );
 a23473a <=( a23472a  and  a23467a );
 a23477a <=( (not A266)  and  (not A265) );
 a23478a <=( A203  and  a23477a );
 a23482a <=( A300  and  A298 );
 a23483a <=( (not A268)  and  a23482a );
 a23484a <=( a23483a  and  a23478a );
 a23487a <=( (not A167)  and  (not A168) );
 a23491a <=( (not A202)  and  (not A200) );
 a23492a <=( A199  and  a23491a );
 a23493a <=( a23492a  and  a23487a );
 a23497a <=( (not A266)  and  (not A265) );
 a23498a <=( A203  and  a23497a );
 a23502a <=( A300  and  A299 );
 a23503a <=( A269  and  a23502a );
 a23504a <=( a23503a  and  a23498a );
 a23507a <=( (not A167)  and  (not A168) );
 a23511a <=( (not A202)  and  (not A200) );
 a23512a <=( A199  and  a23511a );
 a23513a <=( a23512a  and  a23507a );
 a23517a <=( (not A266)  and  (not A265) );
 a23518a <=( A203  and  a23517a );
 a23522a <=( A300  and  A298 );
 a23523a <=( A269  and  a23522a );
 a23524a <=( a23523a  and  a23518a );
 a23527a <=( (not A167)  and  (not A168) );
 a23531a <=( (not A201)  and  (not A200) );
 a23532a <=( A199  and  a23531a );
 a23533a <=( a23532a  and  a23527a );
 a23537a <=( A267  and  A265 );
 a23538a <=( A202  and  a23537a );
 a23542a <=( (not A301)  and  (not A299) );
 a23543a <=( (not A298)  and  a23542a );
 a23544a <=( a23543a  and  a23538a );
 a23547a <=( (not A167)  and  (not A168) );
 a23551a <=( (not A201)  and  (not A200) );
 a23552a <=( A199  and  a23551a );
 a23553a <=( a23552a  and  a23547a );
 a23557a <=( A267  and  A265 );
 a23558a <=( A202  and  a23557a );
 a23562a <=( A302  and  (not A299) );
 a23563a <=( (not A298)  and  a23562a );
 a23564a <=( a23563a  and  a23558a );
 a23567a <=( (not A167)  and  (not A168) );
 a23571a <=( (not A201)  and  (not A200) );
 a23572a <=( A199  and  a23571a );
 a23573a <=( a23572a  and  a23567a );
 a23577a <=( A267  and  A266 );
 a23578a <=( A202  and  a23577a );
 a23582a <=( (not A301)  and  (not A299) );
 a23583a <=( (not A298)  and  a23582a );
 a23584a <=( a23583a  and  a23578a );
 a23587a <=( (not A167)  and  (not A168) );
 a23591a <=( (not A201)  and  (not A200) );
 a23592a <=( A199  and  a23591a );
 a23593a <=( a23592a  and  a23587a );
 a23597a <=( A267  and  A266 );
 a23598a <=( A202  and  a23597a );
 a23602a <=( A302  and  (not A299) );
 a23603a <=( (not A298)  and  a23602a );
 a23604a <=( a23603a  and  a23598a );
 a23607a <=( (not A167)  and  (not A168) );
 a23611a <=( (not A201)  and  (not A200) );
 a23612a <=( A199  and  a23611a );
 a23613a <=( a23612a  and  a23607a );
 a23617a <=( A267  and  A265 );
 a23618a <=( (not A203)  and  a23617a );
 a23622a <=( (not A301)  and  (not A299) );
 a23623a <=( (not A298)  and  a23622a );
 a23624a <=( a23623a  and  a23618a );
 a23627a <=( (not A167)  and  (not A168) );
 a23631a <=( (not A201)  and  (not A200) );
 a23632a <=( A199  and  a23631a );
 a23633a <=( a23632a  and  a23627a );
 a23637a <=( A267  and  A265 );
 a23638a <=( (not A203)  and  a23637a );
 a23642a <=( A302  and  (not A299) );
 a23643a <=( (not A298)  and  a23642a );
 a23644a <=( a23643a  and  a23638a );
 a23647a <=( (not A167)  and  (not A168) );
 a23651a <=( (not A201)  and  (not A200) );
 a23652a <=( A199  and  a23651a );
 a23653a <=( a23652a  and  a23647a );
 a23657a <=( A267  and  A266 );
 a23658a <=( (not A203)  and  a23657a );
 a23662a <=( (not A301)  and  (not A299) );
 a23663a <=( (not A298)  and  a23662a );
 a23664a <=( a23663a  and  a23658a );
 a23667a <=( (not A167)  and  (not A168) );
 a23671a <=( (not A201)  and  (not A200) );
 a23672a <=( A199  and  a23671a );
 a23673a <=( a23672a  and  a23667a );
 a23677a <=( A267  and  A266 );
 a23678a <=( (not A203)  and  a23677a );
 a23682a <=( A302  and  (not A299) );
 a23683a <=( (not A298)  and  a23682a );
 a23684a <=( a23683a  and  a23678a );
 a23687a <=( (not A167)  and  (not A168) );
 a23691a <=( (not A202)  and  (not A200) );
 a23692a <=( (not A199)  and  a23691a );
 a23693a <=( a23692a  and  a23687a );
 a23697a <=( A298  and  A267 );
 a23698a <=( A265  and  a23697a );
 a23702a <=( (not A301)  and  (not A300) );
 a23703a <=( A299  and  a23702a );
 a23704a <=( a23703a  and  a23698a );
 a23707a <=( (not A167)  and  (not A168) );
 a23711a <=( (not A202)  and  (not A200) );
 a23712a <=( (not A199)  and  a23711a );
 a23713a <=( a23712a  and  a23707a );
 a23717a <=( A298  and  A267 );
 a23718a <=( A265  and  a23717a );
 a23722a <=( A302  and  (not A300) );
 a23723a <=( A299  and  a23722a );
 a23724a <=( a23723a  and  a23718a );
 a23727a <=( (not A167)  and  (not A168) );
 a23731a <=( (not A202)  and  (not A200) );
 a23732a <=( (not A199)  and  a23731a );
 a23733a <=( a23732a  and  a23727a );
 a23737a <=( A298  and  A267 );
 a23738a <=( A265  and  a23737a );
 a23742a <=( A301  and  (not A300) );
 a23743a <=( (not A299)  and  a23742a );
 a23744a <=( a23743a  and  a23738a );
 a23747a <=( (not A167)  and  (not A168) );
 a23751a <=( (not A202)  and  (not A200) );
 a23752a <=( (not A199)  and  a23751a );
 a23753a <=( a23752a  and  a23747a );
 a23757a <=( A298  and  A267 );
 a23758a <=( A265  and  a23757a );
 a23762a <=( (not A302)  and  (not A300) );
 a23763a <=( (not A299)  and  a23762a );
 a23764a <=( a23763a  and  a23758a );
 a23767a <=( (not A167)  and  (not A168) );
 a23771a <=( (not A202)  and  (not A200) );
 a23772a <=( (not A199)  and  a23771a );
 a23773a <=( a23772a  and  a23767a );
 a23777a <=( (not A298)  and  A267 );
 a23778a <=( A265  and  a23777a );
 a23782a <=( A301  and  (not A300) );
 a23783a <=( A299  and  a23782a );
 a23784a <=( a23783a  and  a23778a );
 a23787a <=( (not A167)  and  (not A168) );
 a23791a <=( (not A202)  and  (not A200) );
 a23792a <=( (not A199)  and  a23791a );
 a23793a <=( a23792a  and  a23787a );
 a23797a <=( (not A298)  and  A267 );
 a23798a <=( A265  and  a23797a );
 a23802a <=( (not A302)  and  (not A300) );
 a23803a <=( A299  and  a23802a );
 a23804a <=( a23803a  and  a23798a );
 a23807a <=( (not A167)  and  (not A168) );
 a23811a <=( (not A202)  and  (not A200) );
 a23812a <=( (not A199)  and  a23811a );
 a23813a <=( a23812a  and  a23807a );
 a23817a <=( A298  and  A267 );
 a23818a <=( A266  and  a23817a );
 a23822a <=( (not A301)  and  (not A300) );
 a23823a <=( A299  and  a23822a );
 a23824a <=( a23823a  and  a23818a );
 a23827a <=( (not A167)  and  (not A168) );
 a23831a <=( (not A202)  and  (not A200) );
 a23832a <=( (not A199)  and  a23831a );
 a23833a <=( a23832a  and  a23827a );
 a23837a <=( A298  and  A267 );
 a23838a <=( A266  and  a23837a );
 a23842a <=( A302  and  (not A300) );
 a23843a <=( A299  and  a23842a );
 a23844a <=( a23843a  and  a23838a );
 a23847a <=( (not A167)  and  (not A168) );
 a23851a <=( (not A202)  and  (not A200) );
 a23852a <=( (not A199)  and  a23851a );
 a23853a <=( a23852a  and  a23847a );
 a23857a <=( A298  and  A267 );
 a23858a <=( A266  and  a23857a );
 a23862a <=( A301  and  (not A300) );
 a23863a <=( (not A299)  and  a23862a );
 a23864a <=( a23863a  and  a23858a );
 a23867a <=( (not A167)  and  (not A168) );
 a23871a <=( (not A202)  and  (not A200) );
 a23872a <=( (not A199)  and  a23871a );
 a23873a <=( a23872a  and  a23867a );
 a23877a <=( A298  and  A267 );
 a23878a <=( A266  and  a23877a );
 a23882a <=( (not A302)  and  (not A300) );
 a23883a <=( (not A299)  and  a23882a );
 a23884a <=( a23883a  and  a23878a );
 a23887a <=( (not A167)  and  (not A168) );
 a23891a <=( (not A202)  and  (not A200) );
 a23892a <=( (not A199)  and  a23891a );
 a23893a <=( a23892a  and  a23887a );
 a23897a <=( (not A298)  and  A267 );
 a23898a <=( A266  and  a23897a );
 a23902a <=( A301  and  (not A300) );
 a23903a <=( A299  and  a23902a );
 a23904a <=( a23903a  and  a23898a );
 a23907a <=( (not A167)  and  (not A168) );
 a23911a <=( (not A202)  and  (not A200) );
 a23912a <=( (not A199)  and  a23911a );
 a23913a <=( a23912a  and  a23907a );
 a23917a <=( (not A298)  and  A267 );
 a23918a <=( A266  and  a23917a );
 a23922a <=( (not A302)  and  (not A300) );
 a23923a <=( A299  and  a23922a );
 a23924a <=( a23923a  and  a23918a );
 a23927a <=( (not A167)  and  (not A168) );
 a23931a <=( A203  and  (not A200) );
 a23932a <=( (not A199)  and  a23931a );
 a23933a <=( a23932a  and  a23927a );
 a23937a <=( A298  and  A267 );
 a23938a <=( A265  and  a23937a );
 a23942a <=( (not A301)  and  (not A300) );
 a23943a <=( A299  and  a23942a );
 a23944a <=( a23943a  and  a23938a );
 a23947a <=( (not A167)  and  (not A168) );
 a23951a <=( A203  and  (not A200) );
 a23952a <=( (not A199)  and  a23951a );
 a23953a <=( a23952a  and  a23947a );
 a23957a <=( A298  and  A267 );
 a23958a <=( A265  and  a23957a );
 a23962a <=( A302  and  (not A300) );
 a23963a <=( A299  and  a23962a );
 a23964a <=( a23963a  and  a23958a );
 a23967a <=( (not A167)  and  (not A168) );
 a23971a <=( A203  and  (not A200) );
 a23972a <=( (not A199)  and  a23971a );
 a23973a <=( a23972a  and  a23967a );
 a23977a <=( A298  and  A267 );
 a23978a <=( A265  and  a23977a );
 a23982a <=( A301  and  (not A300) );
 a23983a <=( (not A299)  and  a23982a );
 a23984a <=( a23983a  and  a23978a );
 a23987a <=( (not A167)  and  (not A168) );
 a23991a <=( A203  and  (not A200) );
 a23992a <=( (not A199)  and  a23991a );
 a23993a <=( a23992a  and  a23987a );
 a23997a <=( A298  and  A267 );
 a23998a <=( A265  and  a23997a );
 a24002a <=( (not A302)  and  (not A300) );
 a24003a <=( (not A299)  and  a24002a );
 a24004a <=( a24003a  and  a23998a );
 a24007a <=( (not A167)  and  (not A168) );
 a24011a <=( A203  and  (not A200) );
 a24012a <=( (not A199)  and  a24011a );
 a24013a <=( a24012a  and  a24007a );
 a24017a <=( (not A298)  and  A267 );
 a24018a <=( A265  and  a24017a );
 a24022a <=( A301  and  (not A300) );
 a24023a <=( A299  and  a24022a );
 a24024a <=( a24023a  and  a24018a );
 a24027a <=( (not A167)  and  (not A168) );
 a24031a <=( A203  and  (not A200) );
 a24032a <=( (not A199)  and  a24031a );
 a24033a <=( a24032a  and  a24027a );
 a24037a <=( (not A298)  and  A267 );
 a24038a <=( A265  and  a24037a );
 a24042a <=( (not A302)  and  (not A300) );
 a24043a <=( A299  and  a24042a );
 a24044a <=( a24043a  and  a24038a );
 a24047a <=( (not A167)  and  (not A168) );
 a24051a <=( A203  and  (not A200) );
 a24052a <=( (not A199)  and  a24051a );
 a24053a <=( a24052a  and  a24047a );
 a24057a <=( A298  and  A267 );
 a24058a <=( A266  and  a24057a );
 a24062a <=( (not A301)  and  (not A300) );
 a24063a <=( A299  and  a24062a );
 a24064a <=( a24063a  and  a24058a );
 a24067a <=( (not A167)  and  (not A168) );
 a24071a <=( A203  and  (not A200) );
 a24072a <=( (not A199)  and  a24071a );
 a24073a <=( a24072a  and  a24067a );
 a24077a <=( A298  and  A267 );
 a24078a <=( A266  and  a24077a );
 a24082a <=( A302  and  (not A300) );
 a24083a <=( A299  and  a24082a );
 a24084a <=( a24083a  and  a24078a );
 a24087a <=( (not A167)  and  (not A168) );
 a24091a <=( A203  and  (not A200) );
 a24092a <=( (not A199)  and  a24091a );
 a24093a <=( a24092a  and  a24087a );
 a24097a <=( A298  and  A267 );
 a24098a <=( A266  and  a24097a );
 a24102a <=( A301  and  (not A300) );
 a24103a <=( (not A299)  and  a24102a );
 a24104a <=( a24103a  and  a24098a );
 a24107a <=( (not A167)  and  (not A168) );
 a24111a <=( A203  and  (not A200) );
 a24112a <=( (not A199)  and  a24111a );
 a24113a <=( a24112a  and  a24107a );
 a24117a <=( A298  and  A267 );
 a24118a <=( A266  and  a24117a );
 a24122a <=( (not A302)  and  (not A300) );
 a24123a <=( (not A299)  and  a24122a );
 a24124a <=( a24123a  and  a24118a );
 a24127a <=( (not A167)  and  (not A168) );
 a24131a <=( A203  and  (not A200) );
 a24132a <=( (not A199)  and  a24131a );
 a24133a <=( a24132a  and  a24127a );
 a24137a <=( (not A298)  and  A267 );
 a24138a <=( A266  and  a24137a );
 a24142a <=( A301  and  (not A300) );
 a24143a <=( A299  and  a24142a );
 a24144a <=( a24143a  and  a24138a );
 a24147a <=( (not A167)  and  (not A168) );
 a24151a <=( A203  and  (not A200) );
 a24152a <=( (not A199)  and  a24151a );
 a24153a <=( a24152a  and  a24147a );
 a24157a <=( (not A298)  and  A267 );
 a24158a <=( A266  and  a24157a );
 a24162a <=( (not A302)  and  (not A300) );
 a24163a <=( A299  and  a24162a );
 a24164a <=( a24163a  and  a24158a );
 a24167a <=( (not A167)  and  (not A168) );
 a24171a <=( A202  and  (not A200) );
 a24172a <=( (not A199)  and  a24171a );
 a24173a <=( a24172a  and  a24167a );
 a24177a <=( (not A266)  and  (not A265) );
 a24178a <=( (not A203)  and  a24177a );
 a24182a <=( A300  and  A299 );
 a24183a <=( (not A268)  and  a24182a );
 a24184a <=( a24183a  and  a24178a );
 a24187a <=( (not A167)  and  (not A168) );
 a24191a <=( A202  and  (not A200) );
 a24192a <=( (not A199)  and  a24191a );
 a24193a <=( a24192a  and  a24187a );
 a24197a <=( (not A266)  and  (not A265) );
 a24198a <=( (not A203)  and  a24197a );
 a24202a <=( A300  and  A298 );
 a24203a <=( (not A268)  and  a24202a );
 a24204a <=( a24203a  and  a24198a );
 a24207a <=( (not A167)  and  (not A168) );
 a24211a <=( A202  and  (not A200) );
 a24212a <=( (not A199)  and  a24211a );
 a24213a <=( a24212a  and  a24207a );
 a24217a <=( (not A266)  and  (not A265) );
 a24218a <=( (not A203)  and  a24217a );
 a24222a <=( A300  and  A299 );
 a24223a <=( A269  and  a24222a );
 a24224a <=( a24223a  and  a24218a );
 a24227a <=( (not A167)  and  (not A168) );
 a24231a <=( A202  and  (not A200) );
 a24232a <=( (not A199)  and  a24231a );
 a24233a <=( a24232a  and  a24227a );
 a24237a <=( (not A266)  and  (not A265) );
 a24238a <=( (not A203)  and  a24237a );
 a24242a <=( A300  and  A298 );
 a24243a <=( A269  and  a24242a );
 a24244a <=( a24243a  and  a24238a );
 a24247a <=( A168  and  A170 );
 a24251a <=( A199  and  A166 );
 a24252a <=( (not A167)  and  a24251a );
 a24253a <=( a24252a  and  a24247a );
 a24257a <=( A267  and  A265 );
 a24258a <=( A201  and  a24257a );
 a24262a <=( (not A301)  and  (not A299) );
 a24263a <=( (not A298)  and  a24262a );
 a24264a <=( a24263a  and  a24258a );
 a24267a <=( A168  and  A170 );
 a24271a <=( A199  and  A166 );
 a24272a <=( (not A167)  and  a24271a );
 a24273a <=( a24272a  and  a24267a );
 a24277a <=( A267  and  A265 );
 a24278a <=( A201  and  a24277a );
 a24282a <=( A302  and  (not A299) );
 a24283a <=( (not A298)  and  a24282a );
 a24284a <=( a24283a  and  a24278a );
 a24287a <=( A168  and  A170 );
 a24291a <=( A199  and  A166 );
 a24292a <=( (not A167)  and  a24291a );
 a24293a <=( a24292a  and  a24287a );
 a24297a <=( A267  and  A266 );
 a24298a <=( A201  and  a24297a );
 a24302a <=( (not A301)  and  (not A299) );
 a24303a <=( (not A298)  and  a24302a );
 a24304a <=( a24303a  and  a24298a );
 a24307a <=( A168  and  A170 );
 a24311a <=( A199  and  A166 );
 a24312a <=( (not A167)  and  a24311a );
 a24313a <=( a24312a  and  a24307a );
 a24317a <=( A267  and  A266 );
 a24318a <=( A201  and  a24317a );
 a24322a <=( A302  and  (not A299) );
 a24323a <=( (not A298)  and  a24322a );
 a24324a <=( a24323a  and  a24318a );
 a24327a <=( A168  and  A170 );
 a24331a <=( A200  and  A166 );
 a24332a <=( (not A167)  and  a24331a );
 a24333a <=( a24332a  and  a24327a );
 a24337a <=( A267  and  A265 );
 a24338a <=( A201  and  a24337a );
 a24342a <=( (not A301)  and  (not A299) );
 a24343a <=( (not A298)  and  a24342a );
 a24344a <=( a24343a  and  a24338a );
 a24347a <=( A168  and  A170 );
 a24351a <=( A200  and  A166 );
 a24352a <=( (not A167)  and  a24351a );
 a24353a <=( a24352a  and  a24347a );
 a24357a <=( A267  and  A265 );
 a24358a <=( A201  and  a24357a );
 a24362a <=( A302  and  (not A299) );
 a24363a <=( (not A298)  and  a24362a );
 a24364a <=( a24363a  and  a24358a );
 a24367a <=( A168  and  A170 );
 a24371a <=( A200  and  A166 );
 a24372a <=( (not A167)  and  a24371a );
 a24373a <=( a24372a  and  a24367a );
 a24377a <=( A267  and  A266 );
 a24378a <=( A201  and  a24377a );
 a24382a <=( (not A301)  and  (not A299) );
 a24383a <=( (not A298)  and  a24382a );
 a24384a <=( a24383a  and  a24378a );
 a24387a <=( A168  and  A170 );
 a24391a <=( A200  and  A166 );
 a24392a <=( (not A167)  and  a24391a );
 a24393a <=( a24392a  and  a24387a );
 a24397a <=( A267  and  A266 );
 a24398a <=( A201  and  a24397a );
 a24402a <=( A302  and  (not A299) );
 a24403a <=( (not A298)  and  a24402a );
 a24404a <=( a24403a  and  a24398a );
 a24407a <=( A168  and  A169 );
 a24411a <=( A199  and  A166 );
 a24412a <=( (not A167)  and  a24411a );
 a24413a <=( a24412a  and  a24407a );
 a24417a <=( A267  and  A265 );
 a24418a <=( A201  and  a24417a );
 a24422a <=( (not A301)  and  (not A299) );
 a24423a <=( (not A298)  and  a24422a );
 a24424a <=( a24423a  and  a24418a );
 a24427a <=( A168  and  A169 );
 a24431a <=( A199  and  A166 );
 a24432a <=( (not A167)  and  a24431a );
 a24433a <=( a24432a  and  a24427a );
 a24437a <=( A267  and  A265 );
 a24438a <=( A201  and  a24437a );
 a24442a <=( A302  and  (not A299) );
 a24443a <=( (not A298)  and  a24442a );
 a24444a <=( a24443a  and  a24438a );
 a24447a <=( A168  and  A169 );
 a24451a <=( A199  and  A166 );
 a24452a <=( (not A167)  and  a24451a );
 a24453a <=( a24452a  and  a24447a );
 a24457a <=( A267  and  A266 );
 a24458a <=( A201  and  a24457a );
 a24462a <=( (not A301)  and  (not A299) );
 a24463a <=( (not A298)  and  a24462a );
 a24464a <=( a24463a  and  a24458a );
 a24467a <=( A168  and  A169 );
 a24471a <=( A199  and  A166 );
 a24472a <=( (not A167)  and  a24471a );
 a24473a <=( a24472a  and  a24467a );
 a24477a <=( A267  and  A266 );
 a24478a <=( A201  and  a24477a );
 a24482a <=( A302  and  (not A299) );
 a24483a <=( (not A298)  and  a24482a );
 a24484a <=( a24483a  and  a24478a );
 a24487a <=( A168  and  A169 );
 a24491a <=( A200  and  A166 );
 a24492a <=( (not A167)  and  a24491a );
 a24493a <=( a24492a  and  a24487a );
 a24497a <=( A267  and  A265 );
 a24498a <=( A201  and  a24497a );
 a24502a <=( (not A301)  and  (not A299) );
 a24503a <=( (not A298)  and  a24502a );
 a24504a <=( a24503a  and  a24498a );
 a24507a <=( A168  and  A169 );
 a24511a <=( A200  and  A166 );
 a24512a <=( (not A167)  and  a24511a );
 a24513a <=( a24512a  and  a24507a );
 a24517a <=( A267  and  A265 );
 a24518a <=( A201  and  a24517a );
 a24522a <=( A302  and  (not A299) );
 a24523a <=( (not A298)  and  a24522a );
 a24524a <=( a24523a  and  a24518a );
 a24527a <=( A168  and  A169 );
 a24531a <=( A200  and  A166 );
 a24532a <=( (not A167)  and  a24531a );
 a24533a <=( a24532a  and  a24527a );
 a24537a <=( A267  and  A266 );
 a24538a <=( A201  and  a24537a );
 a24542a <=( (not A301)  and  (not A299) );
 a24543a <=( (not A298)  and  a24542a );
 a24544a <=( a24543a  and  a24538a );
 a24547a <=( A168  and  A169 );
 a24551a <=( A200  and  A166 );
 a24552a <=( (not A167)  and  a24551a );
 a24553a <=( a24552a  and  a24547a );
 a24557a <=( A267  and  A266 );
 a24558a <=( A201  and  a24557a );
 a24562a <=( A302  and  (not A299) );
 a24563a <=( (not A298)  and  a24562a );
 a24564a <=( a24563a  and  a24558a );
 a24567a <=( (not A169)  and  (not A170) );
 a24571a <=( A201  and  A199 );
 a24572a <=( (not A167)  and  a24571a );
 a24573a <=( a24572a  and  a24567a );
 a24577a <=( (not A267)  and  A266 );
 a24578a <=( A265  and  a24577a );
 a24582a <=( A300  and  A299 );
 a24583a <=( (not A268)  and  a24582a );
 a24584a <=( a24583a  and  a24578a );
 a24587a <=( (not A169)  and  (not A170) );
 a24591a <=( A201  and  A199 );
 a24592a <=( (not A167)  and  a24591a );
 a24593a <=( a24592a  and  a24587a );
 a24597a <=( (not A267)  and  A266 );
 a24598a <=( A265  and  a24597a );
 a24602a <=( A300  and  A298 );
 a24603a <=( (not A268)  and  a24602a );
 a24604a <=( a24603a  and  a24598a );
 a24607a <=( (not A169)  and  (not A170) );
 a24611a <=( A201  and  A199 );
 a24612a <=( (not A167)  and  a24611a );
 a24613a <=( a24612a  and  a24607a );
 a24617a <=( (not A267)  and  A266 );
 a24618a <=( A265  and  a24617a );
 a24622a <=( A300  and  A299 );
 a24623a <=( A269  and  a24622a );
 a24624a <=( a24623a  and  a24618a );
 a24627a <=( (not A169)  and  (not A170) );
 a24631a <=( A201  and  A199 );
 a24632a <=( (not A167)  and  a24631a );
 a24633a <=( a24632a  and  a24627a );
 a24637a <=( (not A267)  and  A266 );
 a24638a <=( A265  and  a24637a );
 a24642a <=( A300  and  A298 );
 a24643a <=( A269  and  a24642a );
 a24644a <=( a24643a  and  a24638a );
 a24647a <=( (not A169)  and  (not A170) );
 a24651a <=( A201  and  A199 );
 a24652a <=( (not A167)  and  a24651a );
 a24653a <=( a24652a  and  a24647a );
 a24657a <=( (not A267)  and  A266 );
 a24658a <=( (not A265)  and  a24657a );
 a24662a <=( A300  and  A299 );
 a24663a <=( A268  and  a24662a );
 a24664a <=( a24663a  and  a24658a );
 a24667a <=( (not A169)  and  (not A170) );
 a24671a <=( A201  and  A199 );
 a24672a <=( (not A167)  and  a24671a );
 a24673a <=( a24672a  and  a24667a );
 a24677a <=( (not A267)  and  A266 );
 a24678a <=( (not A265)  and  a24677a );
 a24682a <=( A300  and  A298 );
 a24683a <=( A268  and  a24682a );
 a24684a <=( a24683a  and  a24678a );
 a24687a <=( (not A169)  and  (not A170) );
 a24691a <=( A201  and  A199 );
 a24692a <=( (not A167)  and  a24691a );
 a24693a <=( a24692a  and  a24687a );
 a24697a <=( (not A267)  and  A266 );
 a24698a <=( (not A265)  and  a24697a );
 a24702a <=( A300  and  A299 );
 a24703a <=( (not A269)  and  a24702a );
 a24704a <=( a24703a  and  a24698a );
 a24707a <=( (not A169)  and  (not A170) );
 a24711a <=( A201  and  A199 );
 a24712a <=( (not A167)  and  a24711a );
 a24713a <=( a24712a  and  a24707a );
 a24717a <=( (not A267)  and  A266 );
 a24718a <=( (not A265)  and  a24717a );
 a24722a <=( A300  and  A298 );
 a24723a <=( (not A269)  and  a24722a );
 a24724a <=( a24723a  and  a24718a );
 a24727a <=( (not A169)  and  (not A170) );
 a24731a <=( A201  and  A199 );
 a24732a <=( (not A167)  and  a24731a );
 a24733a <=( a24732a  and  a24727a );
 a24737a <=( (not A267)  and  (not A266) );
 a24738a <=( A265  and  a24737a );
 a24742a <=( A300  and  A299 );
 a24743a <=( A268  and  a24742a );
 a24744a <=( a24743a  and  a24738a );
 a24747a <=( (not A169)  and  (not A170) );
 a24751a <=( A201  and  A199 );
 a24752a <=( (not A167)  and  a24751a );
 a24753a <=( a24752a  and  a24747a );
 a24757a <=( (not A267)  and  (not A266) );
 a24758a <=( A265  and  a24757a );
 a24762a <=( A300  and  A298 );
 a24763a <=( A268  and  a24762a );
 a24764a <=( a24763a  and  a24758a );
 a24767a <=( (not A169)  and  (not A170) );
 a24771a <=( A201  and  A199 );
 a24772a <=( (not A167)  and  a24771a );
 a24773a <=( a24772a  and  a24767a );
 a24777a <=( (not A267)  and  (not A266) );
 a24778a <=( A265  and  a24777a );
 a24782a <=( A300  and  A299 );
 a24783a <=( (not A269)  and  a24782a );
 a24784a <=( a24783a  and  a24778a );
 a24787a <=( (not A169)  and  (not A170) );
 a24791a <=( A201  and  A199 );
 a24792a <=( (not A167)  and  a24791a );
 a24793a <=( a24792a  and  a24787a );
 a24797a <=( (not A267)  and  (not A266) );
 a24798a <=( A265  and  a24797a );
 a24802a <=( A300  and  A298 );
 a24803a <=( (not A269)  and  a24802a );
 a24804a <=( a24803a  and  a24798a );
 a24807a <=( (not A169)  and  (not A170) );
 a24811a <=( A201  and  A200 );
 a24812a <=( (not A167)  and  a24811a );
 a24813a <=( a24812a  and  a24807a );
 a24817a <=( (not A267)  and  A266 );
 a24818a <=( A265  and  a24817a );
 a24822a <=( A300  and  A299 );
 a24823a <=( (not A268)  and  a24822a );
 a24824a <=( a24823a  and  a24818a );
 a24827a <=( (not A169)  and  (not A170) );
 a24831a <=( A201  and  A200 );
 a24832a <=( (not A167)  and  a24831a );
 a24833a <=( a24832a  and  a24827a );
 a24837a <=( (not A267)  and  A266 );
 a24838a <=( A265  and  a24837a );
 a24842a <=( A300  and  A298 );
 a24843a <=( (not A268)  and  a24842a );
 a24844a <=( a24843a  and  a24838a );
 a24847a <=( (not A169)  and  (not A170) );
 a24851a <=( A201  and  A200 );
 a24852a <=( (not A167)  and  a24851a );
 a24853a <=( a24852a  and  a24847a );
 a24857a <=( (not A267)  and  A266 );
 a24858a <=( A265  and  a24857a );
 a24862a <=( A300  and  A299 );
 a24863a <=( A269  and  a24862a );
 a24864a <=( a24863a  and  a24858a );
 a24867a <=( (not A169)  and  (not A170) );
 a24871a <=( A201  and  A200 );
 a24872a <=( (not A167)  and  a24871a );
 a24873a <=( a24872a  and  a24867a );
 a24877a <=( (not A267)  and  A266 );
 a24878a <=( A265  and  a24877a );
 a24882a <=( A300  and  A298 );
 a24883a <=( A269  and  a24882a );
 a24884a <=( a24883a  and  a24878a );
 a24887a <=( (not A169)  and  (not A170) );
 a24891a <=( A201  and  A200 );
 a24892a <=( (not A167)  and  a24891a );
 a24893a <=( a24892a  and  a24887a );
 a24897a <=( (not A267)  and  A266 );
 a24898a <=( (not A265)  and  a24897a );
 a24902a <=( A300  and  A299 );
 a24903a <=( A268  and  a24902a );
 a24904a <=( a24903a  and  a24898a );
 a24907a <=( (not A169)  and  (not A170) );
 a24911a <=( A201  and  A200 );
 a24912a <=( (not A167)  and  a24911a );
 a24913a <=( a24912a  and  a24907a );
 a24917a <=( (not A267)  and  A266 );
 a24918a <=( (not A265)  and  a24917a );
 a24922a <=( A300  and  A298 );
 a24923a <=( A268  and  a24922a );
 a24924a <=( a24923a  and  a24918a );
 a24927a <=( (not A169)  and  (not A170) );
 a24931a <=( A201  and  A200 );
 a24932a <=( (not A167)  and  a24931a );
 a24933a <=( a24932a  and  a24927a );
 a24937a <=( (not A267)  and  A266 );
 a24938a <=( (not A265)  and  a24937a );
 a24942a <=( A300  and  A299 );
 a24943a <=( (not A269)  and  a24942a );
 a24944a <=( a24943a  and  a24938a );
 a24947a <=( (not A169)  and  (not A170) );
 a24951a <=( A201  and  A200 );
 a24952a <=( (not A167)  and  a24951a );
 a24953a <=( a24952a  and  a24947a );
 a24957a <=( (not A267)  and  A266 );
 a24958a <=( (not A265)  and  a24957a );
 a24962a <=( A300  and  A298 );
 a24963a <=( (not A269)  and  a24962a );
 a24964a <=( a24963a  and  a24958a );
 a24967a <=( (not A169)  and  (not A170) );
 a24971a <=( A201  and  A200 );
 a24972a <=( (not A167)  and  a24971a );
 a24973a <=( a24972a  and  a24967a );
 a24977a <=( (not A267)  and  (not A266) );
 a24978a <=( A265  and  a24977a );
 a24982a <=( A300  and  A299 );
 a24983a <=( A268  and  a24982a );
 a24984a <=( a24983a  and  a24978a );
 a24987a <=( (not A169)  and  (not A170) );
 a24991a <=( A201  and  A200 );
 a24992a <=( (not A167)  and  a24991a );
 a24993a <=( a24992a  and  a24987a );
 a24997a <=( (not A267)  and  (not A266) );
 a24998a <=( A265  and  a24997a );
 a25002a <=( A300  and  A298 );
 a25003a <=( A268  and  a25002a );
 a25004a <=( a25003a  and  a24998a );
 a25007a <=( (not A169)  and  (not A170) );
 a25011a <=( A201  and  A200 );
 a25012a <=( (not A167)  and  a25011a );
 a25013a <=( a25012a  and  a25007a );
 a25017a <=( (not A267)  and  (not A266) );
 a25018a <=( A265  and  a25017a );
 a25022a <=( A300  and  A299 );
 a25023a <=( (not A269)  and  a25022a );
 a25024a <=( a25023a  and  a25018a );
 a25027a <=( (not A169)  and  (not A170) );
 a25031a <=( A201  and  A200 );
 a25032a <=( (not A167)  and  a25031a );
 a25033a <=( a25032a  and  a25027a );
 a25037a <=( (not A267)  and  (not A266) );
 a25038a <=( A265  and  a25037a );
 a25042a <=( A300  and  A298 );
 a25043a <=( (not A269)  and  a25042a );
 a25044a <=( a25043a  and  a25038a );
 a25047a <=( (not A169)  and  (not A170) );
 a25051a <=( (not A200)  and  (not A199) );
 a25052a <=( (not A167)  and  a25051a );
 a25053a <=( a25052a  and  a25047a );
 a25057a <=( A267  and  A265 );
 a25058a <=( (not A202)  and  a25057a );
 a25062a <=( (not A301)  and  (not A299) );
 a25063a <=( (not A298)  and  a25062a );
 a25064a <=( a25063a  and  a25058a );
 a25067a <=( (not A169)  and  (not A170) );
 a25071a <=( (not A200)  and  (not A199) );
 a25072a <=( (not A167)  and  a25071a );
 a25073a <=( a25072a  and  a25067a );
 a25077a <=( A267  and  A265 );
 a25078a <=( (not A202)  and  a25077a );
 a25082a <=( A302  and  (not A299) );
 a25083a <=( (not A298)  and  a25082a );
 a25084a <=( a25083a  and  a25078a );
 a25087a <=( (not A169)  and  (not A170) );
 a25091a <=( (not A200)  and  (not A199) );
 a25092a <=( (not A167)  and  a25091a );
 a25093a <=( a25092a  and  a25087a );
 a25097a <=( A267  and  A266 );
 a25098a <=( (not A202)  and  a25097a );
 a25102a <=( (not A301)  and  (not A299) );
 a25103a <=( (not A298)  and  a25102a );
 a25104a <=( a25103a  and  a25098a );
 a25107a <=( (not A169)  and  (not A170) );
 a25111a <=( (not A200)  and  (not A199) );
 a25112a <=( (not A167)  and  a25111a );
 a25113a <=( a25112a  and  a25107a );
 a25117a <=( A267  and  A266 );
 a25118a <=( (not A202)  and  a25117a );
 a25122a <=( A302  and  (not A299) );
 a25123a <=( (not A298)  and  a25122a );
 a25124a <=( a25123a  and  a25118a );
 a25127a <=( (not A169)  and  (not A170) );
 a25131a <=( (not A200)  and  (not A199) );
 a25132a <=( (not A167)  and  a25131a );
 a25133a <=( a25132a  and  a25127a );
 a25137a <=( A267  and  A265 );
 a25138a <=( A203  and  a25137a );
 a25142a <=( (not A301)  and  (not A299) );
 a25143a <=( (not A298)  and  a25142a );
 a25144a <=( a25143a  and  a25138a );
 a25147a <=( (not A169)  and  (not A170) );
 a25151a <=( (not A200)  and  (not A199) );
 a25152a <=( (not A167)  and  a25151a );
 a25153a <=( a25152a  and  a25147a );
 a25157a <=( A267  and  A265 );
 a25158a <=( A203  and  a25157a );
 a25162a <=( A302  and  (not A299) );
 a25163a <=( (not A298)  and  a25162a );
 a25164a <=( a25163a  and  a25158a );
 a25167a <=( (not A169)  and  (not A170) );
 a25171a <=( (not A200)  and  (not A199) );
 a25172a <=( (not A167)  and  a25171a );
 a25173a <=( a25172a  and  a25167a );
 a25177a <=( A267  and  A266 );
 a25178a <=( A203  and  a25177a );
 a25182a <=( (not A301)  and  (not A299) );
 a25183a <=( (not A298)  and  a25182a );
 a25184a <=( a25183a  and  a25178a );
 a25187a <=( (not A169)  and  (not A170) );
 a25191a <=( (not A200)  and  (not A199) );
 a25192a <=( (not A167)  and  a25191a );
 a25193a <=( a25192a  and  a25187a );
 a25197a <=( A267  and  A266 );
 a25198a <=( A203  and  a25197a );
 a25202a <=( A302  and  (not A299) );
 a25203a <=( (not A298)  and  a25202a );
 a25204a <=( a25203a  and  a25198a );
 a25208a <=( A199  and  A166 );
 a25209a <=( A167  and  a25208a );
 a25213a <=( A266  and  A265 );
 a25214a <=( A201  and  a25213a );
 a25215a <=( a25214a  and  a25209a );
 a25219a <=( A298  and  (not A268) );
 a25220a <=( (not A267)  and  a25219a );
 a25224a <=( (not A302)  and  A301 );
 a25225a <=( A299  and  a25224a );
 a25226a <=( a25225a  and  a25220a );
 a25230a <=( A199  and  A166 );
 a25231a <=( A167  and  a25230a );
 a25235a <=( A266  and  A265 );
 a25236a <=( A201  and  a25235a );
 a25237a <=( a25236a  and  a25231a );
 a25241a <=( A298  and  (not A268) );
 a25242a <=( (not A267)  and  a25241a );
 a25246a <=( A302  and  (not A301) );
 a25247a <=( (not A299)  and  a25246a );
 a25248a <=( a25247a  and  a25242a );
 a25252a <=( A199  and  A166 );
 a25253a <=( A167  and  a25252a );
 a25257a <=( A266  and  A265 );
 a25258a <=( A201  and  a25257a );
 a25259a <=( a25258a  and  a25253a );
 a25263a <=( (not A298)  and  (not A268) );
 a25264a <=( (not A267)  and  a25263a );
 a25268a <=( A302  and  (not A301) );
 a25269a <=( A299  and  a25268a );
 a25270a <=( a25269a  and  a25264a );
 a25274a <=( A199  and  A166 );
 a25275a <=( A167  and  a25274a );
 a25279a <=( A266  and  A265 );
 a25280a <=( A201  and  a25279a );
 a25281a <=( a25280a  and  a25275a );
 a25285a <=( (not A298)  and  (not A268) );
 a25286a <=( (not A267)  and  a25285a );
 a25290a <=( (not A302)  and  A301 );
 a25291a <=( (not A299)  and  a25290a );
 a25292a <=( a25291a  and  a25286a );
 a25296a <=( A199  and  A166 );
 a25297a <=( A167  and  a25296a );
 a25301a <=( A266  and  A265 );
 a25302a <=( A201  and  a25301a );
 a25303a <=( a25302a  and  a25297a );
 a25307a <=( A298  and  A269 );
 a25308a <=( (not A267)  and  a25307a );
 a25312a <=( (not A302)  and  A301 );
 a25313a <=( A299  and  a25312a );
 a25314a <=( a25313a  and  a25308a );
 a25318a <=( A199  and  A166 );
 a25319a <=( A167  and  a25318a );
 a25323a <=( A266  and  A265 );
 a25324a <=( A201  and  a25323a );
 a25325a <=( a25324a  and  a25319a );
 a25329a <=( A298  and  A269 );
 a25330a <=( (not A267)  and  a25329a );
 a25334a <=( A302  and  (not A301) );
 a25335a <=( (not A299)  and  a25334a );
 a25336a <=( a25335a  and  a25330a );
 a25340a <=( A199  and  A166 );
 a25341a <=( A167  and  a25340a );
 a25345a <=( A266  and  A265 );
 a25346a <=( A201  and  a25345a );
 a25347a <=( a25346a  and  a25341a );
 a25351a <=( (not A298)  and  A269 );
 a25352a <=( (not A267)  and  a25351a );
 a25356a <=( A302  and  (not A301) );
 a25357a <=( A299  and  a25356a );
 a25358a <=( a25357a  and  a25352a );
 a25362a <=( A199  and  A166 );
 a25363a <=( A167  and  a25362a );
 a25367a <=( A266  and  A265 );
 a25368a <=( A201  and  a25367a );
 a25369a <=( a25368a  and  a25363a );
 a25373a <=( (not A298)  and  A269 );
 a25374a <=( (not A267)  and  a25373a );
 a25378a <=( (not A302)  and  A301 );
 a25379a <=( (not A299)  and  a25378a );
 a25380a <=( a25379a  and  a25374a );
 a25384a <=( A199  and  A166 );
 a25385a <=( A167  and  a25384a );
 a25389a <=( A266  and  (not A265) );
 a25390a <=( A201  and  a25389a );
 a25391a <=( a25390a  and  a25385a );
 a25395a <=( A298  and  A268 );
 a25396a <=( (not A267)  and  a25395a );
 a25400a <=( (not A302)  and  A301 );
 a25401a <=( A299  and  a25400a );
 a25402a <=( a25401a  and  a25396a );
 a25406a <=( A199  and  A166 );
 a25407a <=( A167  and  a25406a );
 a25411a <=( A266  and  (not A265) );
 a25412a <=( A201  and  a25411a );
 a25413a <=( a25412a  and  a25407a );
 a25417a <=( A298  and  A268 );
 a25418a <=( (not A267)  and  a25417a );
 a25422a <=( A302  and  (not A301) );
 a25423a <=( (not A299)  and  a25422a );
 a25424a <=( a25423a  and  a25418a );
 a25428a <=( A199  and  A166 );
 a25429a <=( A167  and  a25428a );
 a25433a <=( A266  and  (not A265) );
 a25434a <=( A201  and  a25433a );
 a25435a <=( a25434a  and  a25429a );
 a25439a <=( (not A298)  and  A268 );
 a25440a <=( (not A267)  and  a25439a );
 a25444a <=( A302  and  (not A301) );
 a25445a <=( A299  and  a25444a );
 a25446a <=( a25445a  and  a25440a );
 a25450a <=( A199  and  A166 );
 a25451a <=( A167  and  a25450a );
 a25455a <=( A266  and  (not A265) );
 a25456a <=( A201  and  a25455a );
 a25457a <=( a25456a  and  a25451a );
 a25461a <=( (not A298)  and  A268 );
 a25462a <=( (not A267)  and  a25461a );
 a25466a <=( (not A302)  and  A301 );
 a25467a <=( (not A299)  and  a25466a );
 a25468a <=( a25467a  and  a25462a );
 a25472a <=( A199  and  A166 );
 a25473a <=( A167  and  a25472a );
 a25477a <=( A266  and  (not A265) );
 a25478a <=( A201  and  a25477a );
 a25479a <=( a25478a  and  a25473a );
 a25483a <=( A298  and  (not A269) );
 a25484a <=( (not A267)  and  a25483a );
 a25488a <=( (not A302)  and  A301 );
 a25489a <=( A299  and  a25488a );
 a25490a <=( a25489a  and  a25484a );
 a25494a <=( A199  and  A166 );
 a25495a <=( A167  and  a25494a );
 a25499a <=( A266  and  (not A265) );
 a25500a <=( A201  and  a25499a );
 a25501a <=( a25500a  and  a25495a );
 a25505a <=( A298  and  (not A269) );
 a25506a <=( (not A267)  and  a25505a );
 a25510a <=( A302  and  (not A301) );
 a25511a <=( (not A299)  and  a25510a );
 a25512a <=( a25511a  and  a25506a );
 a25516a <=( A199  and  A166 );
 a25517a <=( A167  and  a25516a );
 a25521a <=( A266  and  (not A265) );
 a25522a <=( A201  and  a25521a );
 a25523a <=( a25522a  and  a25517a );
 a25527a <=( (not A298)  and  (not A269) );
 a25528a <=( (not A267)  and  a25527a );
 a25532a <=( A302  and  (not A301) );
 a25533a <=( A299  and  a25532a );
 a25534a <=( a25533a  and  a25528a );
 a25538a <=( A199  and  A166 );
 a25539a <=( A167  and  a25538a );
 a25543a <=( A266  and  (not A265) );
 a25544a <=( A201  and  a25543a );
 a25545a <=( a25544a  and  a25539a );
 a25549a <=( (not A298)  and  (not A269) );
 a25550a <=( (not A267)  and  a25549a );
 a25554a <=( (not A302)  and  A301 );
 a25555a <=( (not A299)  and  a25554a );
 a25556a <=( a25555a  and  a25550a );
 a25560a <=( A199  and  A166 );
 a25561a <=( A167  and  a25560a );
 a25565a <=( (not A266)  and  A265 );
 a25566a <=( A201  and  a25565a );
 a25567a <=( a25566a  and  a25561a );
 a25571a <=( A298  and  A268 );
 a25572a <=( (not A267)  and  a25571a );
 a25576a <=( (not A302)  and  A301 );
 a25577a <=( A299  and  a25576a );
 a25578a <=( a25577a  and  a25572a );
 a25582a <=( A199  and  A166 );
 a25583a <=( A167  and  a25582a );
 a25587a <=( (not A266)  and  A265 );
 a25588a <=( A201  and  a25587a );
 a25589a <=( a25588a  and  a25583a );
 a25593a <=( A298  and  A268 );
 a25594a <=( (not A267)  and  a25593a );
 a25598a <=( A302  and  (not A301) );
 a25599a <=( (not A299)  and  a25598a );
 a25600a <=( a25599a  and  a25594a );
 a25604a <=( A199  and  A166 );
 a25605a <=( A167  and  a25604a );
 a25609a <=( (not A266)  and  A265 );
 a25610a <=( A201  and  a25609a );
 a25611a <=( a25610a  and  a25605a );
 a25615a <=( (not A298)  and  A268 );
 a25616a <=( (not A267)  and  a25615a );
 a25620a <=( A302  and  (not A301) );
 a25621a <=( A299  and  a25620a );
 a25622a <=( a25621a  and  a25616a );
 a25626a <=( A199  and  A166 );
 a25627a <=( A167  and  a25626a );
 a25631a <=( (not A266)  and  A265 );
 a25632a <=( A201  and  a25631a );
 a25633a <=( a25632a  and  a25627a );
 a25637a <=( (not A298)  and  A268 );
 a25638a <=( (not A267)  and  a25637a );
 a25642a <=( (not A302)  and  A301 );
 a25643a <=( (not A299)  and  a25642a );
 a25644a <=( a25643a  and  a25638a );
 a25648a <=( A199  and  A166 );
 a25649a <=( A167  and  a25648a );
 a25653a <=( (not A266)  and  A265 );
 a25654a <=( A201  and  a25653a );
 a25655a <=( a25654a  and  a25649a );
 a25659a <=( A298  and  (not A269) );
 a25660a <=( (not A267)  and  a25659a );
 a25664a <=( (not A302)  and  A301 );
 a25665a <=( A299  and  a25664a );
 a25666a <=( a25665a  and  a25660a );
 a25670a <=( A199  and  A166 );
 a25671a <=( A167  and  a25670a );
 a25675a <=( (not A266)  and  A265 );
 a25676a <=( A201  and  a25675a );
 a25677a <=( a25676a  and  a25671a );
 a25681a <=( A298  and  (not A269) );
 a25682a <=( (not A267)  and  a25681a );
 a25686a <=( A302  and  (not A301) );
 a25687a <=( (not A299)  and  a25686a );
 a25688a <=( a25687a  and  a25682a );
 a25692a <=( A199  and  A166 );
 a25693a <=( A167  and  a25692a );
 a25697a <=( (not A266)  and  A265 );
 a25698a <=( A201  and  a25697a );
 a25699a <=( a25698a  and  a25693a );
 a25703a <=( (not A298)  and  (not A269) );
 a25704a <=( (not A267)  and  a25703a );
 a25708a <=( A302  and  (not A301) );
 a25709a <=( A299  and  a25708a );
 a25710a <=( a25709a  and  a25704a );
 a25714a <=( A199  and  A166 );
 a25715a <=( A167  and  a25714a );
 a25719a <=( (not A266)  and  A265 );
 a25720a <=( A201  and  a25719a );
 a25721a <=( a25720a  and  a25715a );
 a25725a <=( (not A298)  and  (not A269) );
 a25726a <=( (not A267)  and  a25725a );
 a25730a <=( (not A302)  and  A301 );
 a25731a <=( (not A299)  and  a25730a );
 a25732a <=( a25731a  and  a25726a );
 a25736a <=( A200  and  A166 );
 a25737a <=( A167  and  a25736a );
 a25741a <=( A266  and  A265 );
 a25742a <=( A201  and  a25741a );
 a25743a <=( a25742a  and  a25737a );
 a25747a <=( A298  and  (not A268) );
 a25748a <=( (not A267)  and  a25747a );
 a25752a <=( (not A302)  and  A301 );
 a25753a <=( A299  and  a25752a );
 a25754a <=( a25753a  and  a25748a );
 a25758a <=( A200  and  A166 );
 a25759a <=( A167  and  a25758a );
 a25763a <=( A266  and  A265 );
 a25764a <=( A201  and  a25763a );
 a25765a <=( a25764a  and  a25759a );
 a25769a <=( A298  and  (not A268) );
 a25770a <=( (not A267)  and  a25769a );
 a25774a <=( A302  and  (not A301) );
 a25775a <=( (not A299)  and  a25774a );
 a25776a <=( a25775a  and  a25770a );
 a25780a <=( A200  and  A166 );
 a25781a <=( A167  and  a25780a );
 a25785a <=( A266  and  A265 );
 a25786a <=( A201  and  a25785a );
 a25787a <=( a25786a  and  a25781a );
 a25791a <=( (not A298)  and  (not A268) );
 a25792a <=( (not A267)  and  a25791a );
 a25796a <=( A302  and  (not A301) );
 a25797a <=( A299  and  a25796a );
 a25798a <=( a25797a  and  a25792a );
 a25802a <=( A200  and  A166 );
 a25803a <=( A167  and  a25802a );
 a25807a <=( A266  and  A265 );
 a25808a <=( A201  and  a25807a );
 a25809a <=( a25808a  and  a25803a );
 a25813a <=( (not A298)  and  (not A268) );
 a25814a <=( (not A267)  and  a25813a );
 a25818a <=( (not A302)  and  A301 );
 a25819a <=( (not A299)  and  a25818a );
 a25820a <=( a25819a  and  a25814a );
 a25824a <=( A200  and  A166 );
 a25825a <=( A167  and  a25824a );
 a25829a <=( A266  and  A265 );
 a25830a <=( A201  and  a25829a );
 a25831a <=( a25830a  and  a25825a );
 a25835a <=( A298  and  A269 );
 a25836a <=( (not A267)  and  a25835a );
 a25840a <=( (not A302)  and  A301 );
 a25841a <=( A299  and  a25840a );
 a25842a <=( a25841a  and  a25836a );
 a25846a <=( A200  and  A166 );
 a25847a <=( A167  and  a25846a );
 a25851a <=( A266  and  A265 );
 a25852a <=( A201  and  a25851a );
 a25853a <=( a25852a  and  a25847a );
 a25857a <=( A298  and  A269 );
 a25858a <=( (not A267)  and  a25857a );
 a25862a <=( A302  and  (not A301) );
 a25863a <=( (not A299)  and  a25862a );
 a25864a <=( a25863a  and  a25858a );
 a25868a <=( A200  and  A166 );
 a25869a <=( A167  and  a25868a );
 a25873a <=( A266  and  A265 );
 a25874a <=( A201  and  a25873a );
 a25875a <=( a25874a  and  a25869a );
 a25879a <=( (not A298)  and  A269 );
 a25880a <=( (not A267)  and  a25879a );
 a25884a <=( A302  and  (not A301) );
 a25885a <=( A299  and  a25884a );
 a25886a <=( a25885a  and  a25880a );
 a25890a <=( A200  and  A166 );
 a25891a <=( A167  and  a25890a );
 a25895a <=( A266  and  A265 );
 a25896a <=( A201  and  a25895a );
 a25897a <=( a25896a  and  a25891a );
 a25901a <=( (not A298)  and  A269 );
 a25902a <=( (not A267)  and  a25901a );
 a25906a <=( (not A302)  and  A301 );
 a25907a <=( (not A299)  and  a25906a );
 a25908a <=( a25907a  and  a25902a );
 a25912a <=( A200  and  A166 );
 a25913a <=( A167  and  a25912a );
 a25917a <=( A266  and  (not A265) );
 a25918a <=( A201  and  a25917a );
 a25919a <=( a25918a  and  a25913a );
 a25923a <=( A298  and  A268 );
 a25924a <=( (not A267)  and  a25923a );
 a25928a <=( (not A302)  and  A301 );
 a25929a <=( A299  and  a25928a );
 a25930a <=( a25929a  and  a25924a );
 a25934a <=( A200  and  A166 );
 a25935a <=( A167  and  a25934a );
 a25939a <=( A266  and  (not A265) );
 a25940a <=( A201  and  a25939a );
 a25941a <=( a25940a  and  a25935a );
 a25945a <=( A298  and  A268 );
 a25946a <=( (not A267)  and  a25945a );
 a25950a <=( A302  and  (not A301) );
 a25951a <=( (not A299)  and  a25950a );
 a25952a <=( a25951a  and  a25946a );
 a25956a <=( A200  and  A166 );
 a25957a <=( A167  and  a25956a );
 a25961a <=( A266  and  (not A265) );
 a25962a <=( A201  and  a25961a );
 a25963a <=( a25962a  and  a25957a );
 a25967a <=( (not A298)  and  A268 );
 a25968a <=( (not A267)  and  a25967a );
 a25972a <=( A302  and  (not A301) );
 a25973a <=( A299  and  a25972a );
 a25974a <=( a25973a  and  a25968a );
 a25978a <=( A200  and  A166 );
 a25979a <=( A167  and  a25978a );
 a25983a <=( A266  and  (not A265) );
 a25984a <=( A201  and  a25983a );
 a25985a <=( a25984a  and  a25979a );
 a25989a <=( (not A298)  and  A268 );
 a25990a <=( (not A267)  and  a25989a );
 a25994a <=( (not A302)  and  A301 );
 a25995a <=( (not A299)  and  a25994a );
 a25996a <=( a25995a  and  a25990a );
 a26000a <=( A200  and  A166 );
 a26001a <=( A167  and  a26000a );
 a26005a <=( A266  and  (not A265) );
 a26006a <=( A201  and  a26005a );
 a26007a <=( a26006a  and  a26001a );
 a26011a <=( A298  and  (not A269) );
 a26012a <=( (not A267)  and  a26011a );
 a26016a <=( (not A302)  and  A301 );
 a26017a <=( A299  and  a26016a );
 a26018a <=( a26017a  and  a26012a );
 a26022a <=( A200  and  A166 );
 a26023a <=( A167  and  a26022a );
 a26027a <=( A266  and  (not A265) );
 a26028a <=( A201  and  a26027a );
 a26029a <=( a26028a  and  a26023a );
 a26033a <=( A298  and  (not A269) );
 a26034a <=( (not A267)  and  a26033a );
 a26038a <=( A302  and  (not A301) );
 a26039a <=( (not A299)  and  a26038a );
 a26040a <=( a26039a  and  a26034a );
 a26044a <=( A200  and  A166 );
 a26045a <=( A167  and  a26044a );
 a26049a <=( A266  and  (not A265) );
 a26050a <=( A201  and  a26049a );
 a26051a <=( a26050a  and  a26045a );
 a26055a <=( (not A298)  and  (not A269) );
 a26056a <=( (not A267)  and  a26055a );
 a26060a <=( A302  and  (not A301) );
 a26061a <=( A299  and  a26060a );
 a26062a <=( a26061a  and  a26056a );
 a26066a <=( A200  and  A166 );
 a26067a <=( A167  and  a26066a );
 a26071a <=( A266  and  (not A265) );
 a26072a <=( A201  and  a26071a );
 a26073a <=( a26072a  and  a26067a );
 a26077a <=( (not A298)  and  (not A269) );
 a26078a <=( (not A267)  and  a26077a );
 a26082a <=( (not A302)  and  A301 );
 a26083a <=( (not A299)  and  a26082a );
 a26084a <=( a26083a  and  a26078a );
 a26088a <=( A200  and  A166 );
 a26089a <=( A167  and  a26088a );
 a26093a <=( (not A266)  and  A265 );
 a26094a <=( A201  and  a26093a );
 a26095a <=( a26094a  and  a26089a );
 a26099a <=( A298  and  A268 );
 a26100a <=( (not A267)  and  a26099a );
 a26104a <=( (not A302)  and  A301 );
 a26105a <=( A299  and  a26104a );
 a26106a <=( a26105a  and  a26100a );
 a26110a <=( A200  and  A166 );
 a26111a <=( A167  and  a26110a );
 a26115a <=( (not A266)  and  A265 );
 a26116a <=( A201  and  a26115a );
 a26117a <=( a26116a  and  a26111a );
 a26121a <=( A298  and  A268 );
 a26122a <=( (not A267)  and  a26121a );
 a26126a <=( A302  and  (not A301) );
 a26127a <=( (not A299)  and  a26126a );
 a26128a <=( a26127a  and  a26122a );
 a26132a <=( A200  and  A166 );
 a26133a <=( A167  and  a26132a );
 a26137a <=( (not A266)  and  A265 );
 a26138a <=( A201  and  a26137a );
 a26139a <=( a26138a  and  a26133a );
 a26143a <=( (not A298)  and  A268 );
 a26144a <=( (not A267)  and  a26143a );
 a26148a <=( A302  and  (not A301) );
 a26149a <=( A299  and  a26148a );
 a26150a <=( a26149a  and  a26144a );
 a26154a <=( A200  and  A166 );
 a26155a <=( A167  and  a26154a );
 a26159a <=( (not A266)  and  A265 );
 a26160a <=( A201  and  a26159a );
 a26161a <=( a26160a  and  a26155a );
 a26165a <=( (not A298)  and  A268 );
 a26166a <=( (not A267)  and  a26165a );
 a26170a <=( (not A302)  and  A301 );
 a26171a <=( (not A299)  and  a26170a );
 a26172a <=( a26171a  and  a26166a );
 a26176a <=( A200  and  A166 );
 a26177a <=( A167  and  a26176a );
 a26181a <=( (not A266)  and  A265 );
 a26182a <=( A201  and  a26181a );
 a26183a <=( a26182a  and  a26177a );
 a26187a <=( A298  and  (not A269) );
 a26188a <=( (not A267)  and  a26187a );
 a26192a <=( (not A302)  and  A301 );
 a26193a <=( A299  and  a26192a );
 a26194a <=( a26193a  and  a26188a );
 a26198a <=( A200  and  A166 );
 a26199a <=( A167  and  a26198a );
 a26203a <=( (not A266)  and  A265 );
 a26204a <=( A201  and  a26203a );
 a26205a <=( a26204a  and  a26199a );
 a26209a <=( A298  and  (not A269) );
 a26210a <=( (not A267)  and  a26209a );
 a26214a <=( A302  and  (not A301) );
 a26215a <=( (not A299)  and  a26214a );
 a26216a <=( a26215a  and  a26210a );
 a26220a <=( A200  and  A166 );
 a26221a <=( A167  and  a26220a );
 a26225a <=( (not A266)  and  A265 );
 a26226a <=( A201  and  a26225a );
 a26227a <=( a26226a  and  a26221a );
 a26231a <=( (not A298)  and  (not A269) );
 a26232a <=( (not A267)  and  a26231a );
 a26236a <=( A302  and  (not A301) );
 a26237a <=( A299  and  a26236a );
 a26238a <=( a26237a  and  a26232a );
 a26242a <=( A200  and  A166 );
 a26243a <=( A167  and  a26242a );
 a26247a <=( (not A266)  and  A265 );
 a26248a <=( A201  and  a26247a );
 a26249a <=( a26248a  and  a26243a );
 a26253a <=( (not A298)  and  (not A269) );
 a26254a <=( (not A267)  and  a26253a );
 a26258a <=( (not A302)  and  A301 );
 a26259a <=( (not A299)  and  a26258a );
 a26260a <=( a26259a  and  a26254a );
 a26264a <=( A199  and  A166 );
 a26265a <=( A167  and  a26264a );
 a26269a <=( (not A203)  and  A202 );
 a26270a <=( A200  and  a26269a );
 a26271a <=( a26270a  and  a26265a );
 a26275a <=( (not A267)  and  A266 );
 a26276a <=( A265  and  a26275a );
 a26280a <=( A300  and  A299 );
 a26281a <=( (not A268)  and  a26280a );
 a26282a <=( a26281a  and  a26276a );
 a26286a <=( A199  and  A166 );
 a26287a <=( A167  and  a26286a );
 a26291a <=( (not A203)  and  A202 );
 a26292a <=( A200  and  a26291a );
 a26293a <=( a26292a  and  a26287a );
 a26297a <=( (not A267)  and  A266 );
 a26298a <=( A265  and  a26297a );
 a26302a <=( A300  and  A298 );
 a26303a <=( (not A268)  and  a26302a );
 a26304a <=( a26303a  and  a26298a );
 a26308a <=( A199  and  A166 );
 a26309a <=( A167  and  a26308a );
 a26313a <=( (not A203)  and  A202 );
 a26314a <=( A200  and  a26313a );
 a26315a <=( a26314a  and  a26309a );
 a26319a <=( (not A267)  and  A266 );
 a26320a <=( A265  and  a26319a );
 a26324a <=( A300  and  A299 );
 a26325a <=( A269  and  a26324a );
 a26326a <=( a26325a  and  a26320a );
 a26330a <=( A199  and  A166 );
 a26331a <=( A167  and  a26330a );
 a26335a <=( (not A203)  and  A202 );
 a26336a <=( A200  and  a26335a );
 a26337a <=( a26336a  and  a26331a );
 a26341a <=( (not A267)  and  A266 );
 a26342a <=( A265  and  a26341a );
 a26346a <=( A300  and  A298 );
 a26347a <=( A269  and  a26346a );
 a26348a <=( a26347a  and  a26342a );
 a26352a <=( A199  and  A166 );
 a26353a <=( A167  and  a26352a );
 a26357a <=( (not A203)  and  A202 );
 a26358a <=( A200  and  a26357a );
 a26359a <=( a26358a  and  a26353a );
 a26363a <=( (not A267)  and  A266 );
 a26364a <=( (not A265)  and  a26363a );
 a26368a <=( A300  and  A299 );
 a26369a <=( A268  and  a26368a );
 a26370a <=( a26369a  and  a26364a );
 a26374a <=( A199  and  A166 );
 a26375a <=( A167  and  a26374a );
 a26379a <=( (not A203)  and  A202 );
 a26380a <=( A200  and  a26379a );
 a26381a <=( a26380a  and  a26375a );
 a26385a <=( (not A267)  and  A266 );
 a26386a <=( (not A265)  and  a26385a );
 a26390a <=( A300  and  A298 );
 a26391a <=( A268  and  a26390a );
 a26392a <=( a26391a  and  a26386a );
 a26396a <=( A199  and  A166 );
 a26397a <=( A167  and  a26396a );
 a26401a <=( (not A203)  and  A202 );
 a26402a <=( A200  and  a26401a );
 a26403a <=( a26402a  and  a26397a );
 a26407a <=( (not A267)  and  A266 );
 a26408a <=( (not A265)  and  a26407a );
 a26412a <=( A300  and  A299 );
 a26413a <=( (not A269)  and  a26412a );
 a26414a <=( a26413a  and  a26408a );
 a26418a <=( A199  and  A166 );
 a26419a <=( A167  and  a26418a );
 a26423a <=( (not A203)  and  A202 );
 a26424a <=( A200  and  a26423a );
 a26425a <=( a26424a  and  a26419a );
 a26429a <=( (not A267)  and  A266 );
 a26430a <=( (not A265)  and  a26429a );
 a26434a <=( A300  and  A298 );
 a26435a <=( (not A269)  and  a26434a );
 a26436a <=( a26435a  and  a26430a );
 a26440a <=( A199  and  A166 );
 a26441a <=( A167  and  a26440a );
 a26445a <=( (not A203)  and  A202 );
 a26446a <=( A200  and  a26445a );
 a26447a <=( a26446a  and  a26441a );
 a26451a <=( (not A267)  and  (not A266) );
 a26452a <=( A265  and  a26451a );
 a26456a <=( A300  and  A299 );
 a26457a <=( A268  and  a26456a );
 a26458a <=( a26457a  and  a26452a );
 a26462a <=( A199  and  A166 );
 a26463a <=( A167  and  a26462a );
 a26467a <=( (not A203)  and  A202 );
 a26468a <=( A200  and  a26467a );
 a26469a <=( a26468a  and  a26463a );
 a26473a <=( (not A267)  and  (not A266) );
 a26474a <=( A265  and  a26473a );
 a26478a <=( A300  and  A298 );
 a26479a <=( A268  and  a26478a );
 a26480a <=( a26479a  and  a26474a );
 a26484a <=( A199  and  A166 );
 a26485a <=( A167  and  a26484a );
 a26489a <=( (not A203)  and  A202 );
 a26490a <=( A200  and  a26489a );
 a26491a <=( a26490a  and  a26485a );
 a26495a <=( (not A267)  and  (not A266) );
 a26496a <=( A265  and  a26495a );
 a26500a <=( A300  and  A299 );
 a26501a <=( (not A269)  and  a26500a );
 a26502a <=( a26501a  and  a26496a );
 a26506a <=( A199  and  A166 );
 a26507a <=( A167  and  a26506a );
 a26511a <=( (not A203)  and  A202 );
 a26512a <=( A200  and  a26511a );
 a26513a <=( a26512a  and  a26507a );
 a26517a <=( (not A267)  and  (not A266) );
 a26518a <=( A265  and  a26517a );
 a26522a <=( A300  and  A298 );
 a26523a <=( (not A269)  and  a26522a );
 a26524a <=( a26523a  and  a26518a );
 a26528a <=( A199  and  A166 );
 a26529a <=( A167  and  a26528a );
 a26533a <=( (not A202)  and  (not A201) );
 a26534a <=( A200  and  a26533a );
 a26535a <=( a26534a  and  a26529a );
 a26539a <=( A298  and  A267 );
 a26540a <=( A265  and  a26539a );
 a26544a <=( (not A301)  and  (not A300) );
 a26545a <=( A299  and  a26544a );
 a26546a <=( a26545a  and  a26540a );
 a26550a <=( A199  and  A166 );
 a26551a <=( A167  and  a26550a );
 a26555a <=( (not A202)  and  (not A201) );
 a26556a <=( A200  and  a26555a );
 a26557a <=( a26556a  and  a26551a );
 a26561a <=( A298  and  A267 );
 a26562a <=( A265  and  a26561a );
 a26566a <=( A302  and  (not A300) );
 a26567a <=( A299  and  a26566a );
 a26568a <=( a26567a  and  a26562a );
 a26572a <=( A199  and  A166 );
 a26573a <=( A167  and  a26572a );
 a26577a <=( (not A202)  and  (not A201) );
 a26578a <=( A200  and  a26577a );
 a26579a <=( a26578a  and  a26573a );
 a26583a <=( A298  and  A267 );
 a26584a <=( A265  and  a26583a );
 a26588a <=( A301  and  (not A300) );
 a26589a <=( (not A299)  and  a26588a );
 a26590a <=( a26589a  and  a26584a );
 a26594a <=( A199  and  A166 );
 a26595a <=( A167  and  a26594a );
 a26599a <=( (not A202)  and  (not A201) );
 a26600a <=( A200  and  a26599a );
 a26601a <=( a26600a  and  a26595a );
 a26605a <=( A298  and  A267 );
 a26606a <=( A265  and  a26605a );
 a26610a <=( (not A302)  and  (not A300) );
 a26611a <=( (not A299)  and  a26610a );
 a26612a <=( a26611a  and  a26606a );
 a26616a <=( A199  and  A166 );
 a26617a <=( A167  and  a26616a );
 a26621a <=( (not A202)  and  (not A201) );
 a26622a <=( A200  and  a26621a );
 a26623a <=( a26622a  and  a26617a );
 a26627a <=( (not A298)  and  A267 );
 a26628a <=( A265  and  a26627a );
 a26632a <=( A301  and  (not A300) );
 a26633a <=( A299  and  a26632a );
 a26634a <=( a26633a  and  a26628a );
 a26638a <=( A199  and  A166 );
 a26639a <=( A167  and  a26638a );
 a26643a <=( (not A202)  and  (not A201) );
 a26644a <=( A200  and  a26643a );
 a26645a <=( a26644a  and  a26639a );
 a26649a <=( (not A298)  and  A267 );
 a26650a <=( A265  and  a26649a );
 a26654a <=( (not A302)  and  (not A300) );
 a26655a <=( A299  and  a26654a );
 a26656a <=( a26655a  and  a26650a );
 a26660a <=( A199  and  A166 );
 a26661a <=( A167  and  a26660a );
 a26665a <=( (not A202)  and  (not A201) );
 a26666a <=( A200  and  a26665a );
 a26667a <=( a26666a  and  a26661a );
 a26671a <=( A298  and  A267 );
 a26672a <=( A266  and  a26671a );
 a26676a <=( (not A301)  and  (not A300) );
 a26677a <=( A299  and  a26676a );
 a26678a <=( a26677a  and  a26672a );
 a26682a <=( A199  and  A166 );
 a26683a <=( A167  and  a26682a );
 a26687a <=( (not A202)  and  (not A201) );
 a26688a <=( A200  and  a26687a );
 a26689a <=( a26688a  and  a26683a );
 a26693a <=( A298  and  A267 );
 a26694a <=( A266  and  a26693a );
 a26698a <=( A302  and  (not A300) );
 a26699a <=( A299  and  a26698a );
 a26700a <=( a26699a  and  a26694a );
 a26704a <=( A199  and  A166 );
 a26705a <=( A167  and  a26704a );
 a26709a <=( (not A202)  and  (not A201) );
 a26710a <=( A200  and  a26709a );
 a26711a <=( a26710a  and  a26705a );
 a26715a <=( A298  and  A267 );
 a26716a <=( A266  and  a26715a );
 a26720a <=( A301  and  (not A300) );
 a26721a <=( (not A299)  and  a26720a );
 a26722a <=( a26721a  and  a26716a );
 a26726a <=( A199  and  A166 );
 a26727a <=( A167  and  a26726a );
 a26731a <=( (not A202)  and  (not A201) );
 a26732a <=( A200  and  a26731a );
 a26733a <=( a26732a  and  a26727a );
 a26737a <=( A298  and  A267 );
 a26738a <=( A266  and  a26737a );
 a26742a <=( (not A302)  and  (not A300) );
 a26743a <=( (not A299)  and  a26742a );
 a26744a <=( a26743a  and  a26738a );
 a26748a <=( A199  and  A166 );
 a26749a <=( A167  and  a26748a );
 a26753a <=( (not A202)  and  (not A201) );
 a26754a <=( A200  and  a26753a );
 a26755a <=( a26754a  and  a26749a );
 a26759a <=( (not A298)  and  A267 );
 a26760a <=( A266  and  a26759a );
 a26764a <=( A301  and  (not A300) );
 a26765a <=( A299  and  a26764a );
 a26766a <=( a26765a  and  a26760a );
 a26770a <=( A199  and  A166 );
 a26771a <=( A167  and  a26770a );
 a26775a <=( (not A202)  and  (not A201) );
 a26776a <=( A200  and  a26775a );
 a26777a <=( a26776a  and  a26771a );
 a26781a <=( (not A298)  and  A267 );
 a26782a <=( A266  and  a26781a );
 a26786a <=( (not A302)  and  (not A300) );
 a26787a <=( A299  and  a26786a );
 a26788a <=( a26787a  and  a26782a );
 a26792a <=( A199  and  A166 );
 a26793a <=( A167  and  a26792a );
 a26797a <=( A203  and  (not A201) );
 a26798a <=( A200  and  a26797a );
 a26799a <=( a26798a  and  a26793a );
 a26803a <=( A298  and  A267 );
 a26804a <=( A265  and  a26803a );
 a26808a <=( (not A301)  and  (not A300) );
 a26809a <=( A299  and  a26808a );
 a26810a <=( a26809a  and  a26804a );
 a26814a <=( A199  and  A166 );
 a26815a <=( A167  and  a26814a );
 a26819a <=( A203  and  (not A201) );
 a26820a <=( A200  and  a26819a );
 a26821a <=( a26820a  and  a26815a );
 a26825a <=( A298  and  A267 );
 a26826a <=( A265  and  a26825a );
 a26830a <=( A302  and  (not A300) );
 a26831a <=( A299  and  a26830a );
 a26832a <=( a26831a  and  a26826a );
 a26836a <=( A199  and  A166 );
 a26837a <=( A167  and  a26836a );
 a26841a <=( A203  and  (not A201) );
 a26842a <=( A200  and  a26841a );
 a26843a <=( a26842a  and  a26837a );
 a26847a <=( A298  and  A267 );
 a26848a <=( A265  and  a26847a );
 a26852a <=( A301  and  (not A300) );
 a26853a <=( (not A299)  and  a26852a );
 a26854a <=( a26853a  and  a26848a );
 a26858a <=( A199  and  A166 );
 a26859a <=( A167  and  a26858a );
 a26863a <=( A203  and  (not A201) );
 a26864a <=( A200  and  a26863a );
 a26865a <=( a26864a  and  a26859a );
 a26869a <=( A298  and  A267 );
 a26870a <=( A265  and  a26869a );
 a26874a <=( (not A302)  and  (not A300) );
 a26875a <=( (not A299)  and  a26874a );
 a26876a <=( a26875a  and  a26870a );
 a26880a <=( A199  and  A166 );
 a26881a <=( A167  and  a26880a );
 a26885a <=( A203  and  (not A201) );
 a26886a <=( A200  and  a26885a );
 a26887a <=( a26886a  and  a26881a );
 a26891a <=( (not A298)  and  A267 );
 a26892a <=( A265  and  a26891a );
 a26896a <=( A301  and  (not A300) );
 a26897a <=( A299  and  a26896a );
 a26898a <=( a26897a  and  a26892a );
 a26902a <=( A199  and  A166 );
 a26903a <=( A167  and  a26902a );
 a26907a <=( A203  and  (not A201) );
 a26908a <=( A200  and  a26907a );
 a26909a <=( a26908a  and  a26903a );
 a26913a <=( (not A298)  and  A267 );
 a26914a <=( A265  and  a26913a );
 a26918a <=( (not A302)  and  (not A300) );
 a26919a <=( A299  and  a26918a );
 a26920a <=( a26919a  and  a26914a );
 a26924a <=( A199  and  A166 );
 a26925a <=( A167  and  a26924a );
 a26929a <=( A203  and  (not A201) );
 a26930a <=( A200  and  a26929a );
 a26931a <=( a26930a  and  a26925a );
 a26935a <=( A298  and  A267 );
 a26936a <=( A266  and  a26935a );
 a26940a <=( (not A301)  and  (not A300) );
 a26941a <=( A299  and  a26940a );
 a26942a <=( a26941a  and  a26936a );
 a26946a <=( A199  and  A166 );
 a26947a <=( A167  and  a26946a );
 a26951a <=( A203  and  (not A201) );
 a26952a <=( A200  and  a26951a );
 a26953a <=( a26952a  and  a26947a );
 a26957a <=( A298  and  A267 );
 a26958a <=( A266  and  a26957a );
 a26962a <=( A302  and  (not A300) );
 a26963a <=( A299  and  a26962a );
 a26964a <=( a26963a  and  a26958a );
 a26968a <=( A199  and  A166 );
 a26969a <=( A167  and  a26968a );
 a26973a <=( A203  and  (not A201) );
 a26974a <=( A200  and  a26973a );
 a26975a <=( a26974a  and  a26969a );
 a26979a <=( A298  and  A267 );
 a26980a <=( A266  and  a26979a );
 a26984a <=( A301  and  (not A300) );
 a26985a <=( (not A299)  and  a26984a );
 a26986a <=( a26985a  and  a26980a );
 a26990a <=( A199  and  A166 );
 a26991a <=( A167  and  a26990a );
 a26995a <=( A203  and  (not A201) );
 a26996a <=( A200  and  a26995a );
 a26997a <=( a26996a  and  a26991a );
 a27001a <=( A298  and  A267 );
 a27002a <=( A266  and  a27001a );
 a27006a <=( (not A302)  and  (not A300) );
 a27007a <=( (not A299)  and  a27006a );
 a27008a <=( a27007a  and  a27002a );
 a27012a <=( A199  and  A166 );
 a27013a <=( A167  and  a27012a );
 a27017a <=( A203  and  (not A201) );
 a27018a <=( A200  and  a27017a );
 a27019a <=( a27018a  and  a27013a );
 a27023a <=( (not A298)  and  A267 );
 a27024a <=( A266  and  a27023a );
 a27028a <=( A301  and  (not A300) );
 a27029a <=( A299  and  a27028a );
 a27030a <=( a27029a  and  a27024a );
 a27034a <=( A199  and  A166 );
 a27035a <=( A167  and  a27034a );
 a27039a <=( A203  and  (not A201) );
 a27040a <=( A200  and  a27039a );
 a27041a <=( a27040a  and  a27035a );
 a27045a <=( (not A298)  and  A267 );
 a27046a <=( A266  and  a27045a );
 a27050a <=( (not A302)  and  (not A300) );
 a27051a <=( A299  and  a27050a );
 a27052a <=( a27051a  and  a27046a );
 a27056a <=( (not A199)  and  A166 );
 a27057a <=( A167  and  a27056a );
 a27061a <=( A203  and  (not A202) );
 a27062a <=( A200  and  a27061a );
 a27063a <=( a27062a  and  a27057a );
 a27067a <=( (not A267)  and  A266 );
 a27068a <=( A265  and  a27067a );
 a27072a <=( A300  and  A299 );
 a27073a <=( (not A268)  and  a27072a );
 a27074a <=( a27073a  and  a27068a );
 a27078a <=( (not A199)  and  A166 );
 a27079a <=( A167  and  a27078a );
 a27083a <=( A203  and  (not A202) );
 a27084a <=( A200  and  a27083a );
 a27085a <=( a27084a  and  a27079a );
 a27089a <=( (not A267)  and  A266 );
 a27090a <=( A265  and  a27089a );
 a27094a <=( A300  and  A298 );
 a27095a <=( (not A268)  and  a27094a );
 a27096a <=( a27095a  and  a27090a );
 a27100a <=( (not A199)  and  A166 );
 a27101a <=( A167  and  a27100a );
 a27105a <=( A203  and  (not A202) );
 a27106a <=( A200  and  a27105a );
 a27107a <=( a27106a  and  a27101a );
 a27111a <=( (not A267)  and  A266 );
 a27112a <=( A265  and  a27111a );
 a27116a <=( A300  and  A299 );
 a27117a <=( A269  and  a27116a );
 a27118a <=( a27117a  and  a27112a );
 a27122a <=( (not A199)  and  A166 );
 a27123a <=( A167  and  a27122a );
 a27127a <=( A203  and  (not A202) );
 a27128a <=( A200  and  a27127a );
 a27129a <=( a27128a  and  a27123a );
 a27133a <=( (not A267)  and  A266 );
 a27134a <=( A265  and  a27133a );
 a27138a <=( A300  and  A298 );
 a27139a <=( A269  and  a27138a );
 a27140a <=( a27139a  and  a27134a );
 a27144a <=( (not A199)  and  A166 );
 a27145a <=( A167  and  a27144a );
 a27149a <=( A203  and  (not A202) );
 a27150a <=( A200  and  a27149a );
 a27151a <=( a27150a  and  a27145a );
 a27155a <=( (not A267)  and  A266 );
 a27156a <=( (not A265)  and  a27155a );
 a27160a <=( A300  and  A299 );
 a27161a <=( A268  and  a27160a );
 a27162a <=( a27161a  and  a27156a );
 a27166a <=( (not A199)  and  A166 );
 a27167a <=( A167  and  a27166a );
 a27171a <=( A203  and  (not A202) );
 a27172a <=( A200  and  a27171a );
 a27173a <=( a27172a  and  a27167a );
 a27177a <=( (not A267)  and  A266 );
 a27178a <=( (not A265)  and  a27177a );
 a27182a <=( A300  and  A298 );
 a27183a <=( A268  and  a27182a );
 a27184a <=( a27183a  and  a27178a );
 a27188a <=( (not A199)  and  A166 );
 a27189a <=( A167  and  a27188a );
 a27193a <=( A203  and  (not A202) );
 a27194a <=( A200  and  a27193a );
 a27195a <=( a27194a  and  a27189a );
 a27199a <=( (not A267)  and  A266 );
 a27200a <=( (not A265)  and  a27199a );
 a27204a <=( A300  and  A299 );
 a27205a <=( (not A269)  and  a27204a );
 a27206a <=( a27205a  and  a27200a );
 a27210a <=( (not A199)  and  A166 );
 a27211a <=( A167  and  a27210a );
 a27215a <=( A203  and  (not A202) );
 a27216a <=( A200  and  a27215a );
 a27217a <=( a27216a  and  a27211a );
 a27221a <=( (not A267)  and  A266 );
 a27222a <=( (not A265)  and  a27221a );
 a27226a <=( A300  and  A298 );
 a27227a <=( (not A269)  and  a27226a );
 a27228a <=( a27227a  and  a27222a );
 a27232a <=( (not A199)  and  A166 );
 a27233a <=( A167  and  a27232a );
 a27237a <=( A203  and  (not A202) );
 a27238a <=( A200  and  a27237a );
 a27239a <=( a27238a  and  a27233a );
 a27243a <=( (not A267)  and  (not A266) );
 a27244a <=( A265  and  a27243a );
 a27248a <=( A300  and  A299 );
 a27249a <=( A268  and  a27248a );
 a27250a <=( a27249a  and  a27244a );
 a27254a <=( (not A199)  and  A166 );
 a27255a <=( A167  and  a27254a );
 a27259a <=( A203  and  (not A202) );
 a27260a <=( A200  and  a27259a );
 a27261a <=( a27260a  and  a27255a );
 a27265a <=( (not A267)  and  (not A266) );
 a27266a <=( A265  and  a27265a );
 a27270a <=( A300  and  A298 );
 a27271a <=( A268  and  a27270a );
 a27272a <=( a27271a  and  a27266a );
 a27276a <=( (not A199)  and  A166 );
 a27277a <=( A167  and  a27276a );
 a27281a <=( A203  and  (not A202) );
 a27282a <=( A200  and  a27281a );
 a27283a <=( a27282a  and  a27277a );
 a27287a <=( (not A267)  and  (not A266) );
 a27288a <=( A265  and  a27287a );
 a27292a <=( A300  and  A299 );
 a27293a <=( (not A269)  and  a27292a );
 a27294a <=( a27293a  and  a27288a );
 a27298a <=( (not A199)  and  A166 );
 a27299a <=( A167  and  a27298a );
 a27303a <=( A203  and  (not A202) );
 a27304a <=( A200  and  a27303a );
 a27305a <=( a27304a  and  a27299a );
 a27309a <=( (not A267)  and  (not A266) );
 a27310a <=( A265  and  a27309a );
 a27314a <=( A300  and  A298 );
 a27315a <=( (not A269)  and  a27314a );
 a27316a <=( a27315a  and  a27310a );
 a27320a <=( (not A199)  and  A166 );
 a27321a <=( A167  and  a27320a );
 a27325a <=( A202  and  (not A201) );
 a27326a <=( A200  and  a27325a );
 a27327a <=( a27326a  and  a27321a );
 a27331a <=( A298  and  A267 );
 a27332a <=( A265  and  a27331a );
 a27336a <=( (not A301)  and  (not A300) );
 a27337a <=( A299  and  a27336a );
 a27338a <=( a27337a  and  a27332a );
 a27342a <=( (not A199)  and  A166 );
 a27343a <=( A167  and  a27342a );
 a27347a <=( A202  and  (not A201) );
 a27348a <=( A200  and  a27347a );
 a27349a <=( a27348a  and  a27343a );
 a27353a <=( A298  and  A267 );
 a27354a <=( A265  and  a27353a );
 a27358a <=( A302  and  (not A300) );
 a27359a <=( A299  and  a27358a );
 a27360a <=( a27359a  and  a27354a );
 a27364a <=( (not A199)  and  A166 );
 a27365a <=( A167  and  a27364a );
 a27369a <=( A202  and  (not A201) );
 a27370a <=( A200  and  a27369a );
 a27371a <=( a27370a  and  a27365a );
 a27375a <=( A298  and  A267 );
 a27376a <=( A265  and  a27375a );
 a27380a <=( A301  and  (not A300) );
 a27381a <=( (not A299)  and  a27380a );
 a27382a <=( a27381a  and  a27376a );
 a27386a <=( (not A199)  and  A166 );
 a27387a <=( A167  and  a27386a );
 a27391a <=( A202  and  (not A201) );
 a27392a <=( A200  and  a27391a );
 a27393a <=( a27392a  and  a27387a );
 a27397a <=( A298  and  A267 );
 a27398a <=( A265  and  a27397a );
 a27402a <=( (not A302)  and  (not A300) );
 a27403a <=( (not A299)  and  a27402a );
 a27404a <=( a27403a  and  a27398a );
 a27408a <=( (not A199)  and  A166 );
 a27409a <=( A167  and  a27408a );
 a27413a <=( A202  and  (not A201) );
 a27414a <=( A200  and  a27413a );
 a27415a <=( a27414a  and  a27409a );
 a27419a <=( (not A298)  and  A267 );
 a27420a <=( A265  and  a27419a );
 a27424a <=( A301  and  (not A300) );
 a27425a <=( A299  and  a27424a );
 a27426a <=( a27425a  and  a27420a );
 a27430a <=( (not A199)  and  A166 );
 a27431a <=( A167  and  a27430a );
 a27435a <=( A202  and  (not A201) );
 a27436a <=( A200  and  a27435a );
 a27437a <=( a27436a  and  a27431a );
 a27441a <=( (not A298)  and  A267 );
 a27442a <=( A265  and  a27441a );
 a27446a <=( (not A302)  and  (not A300) );
 a27447a <=( A299  and  a27446a );
 a27448a <=( a27447a  and  a27442a );
 a27452a <=( (not A199)  and  A166 );
 a27453a <=( A167  and  a27452a );
 a27457a <=( A202  and  (not A201) );
 a27458a <=( A200  and  a27457a );
 a27459a <=( a27458a  and  a27453a );
 a27463a <=( A298  and  A267 );
 a27464a <=( A266  and  a27463a );
 a27468a <=( (not A301)  and  (not A300) );
 a27469a <=( A299  and  a27468a );
 a27470a <=( a27469a  and  a27464a );
 a27474a <=( (not A199)  and  A166 );
 a27475a <=( A167  and  a27474a );
 a27479a <=( A202  and  (not A201) );
 a27480a <=( A200  and  a27479a );
 a27481a <=( a27480a  and  a27475a );
 a27485a <=( A298  and  A267 );
 a27486a <=( A266  and  a27485a );
 a27490a <=( A302  and  (not A300) );
 a27491a <=( A299  and  a27490a );
 a27492a <=( a27491a  and  a27486a );
 a27496a <=( (not A199)  and  A166 );
 a27497a <=( A167  and  a27496a );
 a27501a <=( A202  and  (not A201) );
 a27502a <=( A200  and  a27501a );
 a27503a <=( a27502a  and  a27497a );
 a27507a <=( A298  and  A267 );
 a27508a <=( A266  and  a27507a );
 a27512a <=( A301  and  (not A300) );
 a27513a <=( (not A299)  and  a27512a );
 a27514a <=( a27513a  and  a27508a );
 a27518a <=( (not A199)  and  A166 );
 a27519a <=( A167  and  a27518a );
 a27523a <=( A202  and  (not A201) );
 a27524a <=( A200  and  a27523a );
 a27525a <=( a27524a  and  a27519a );
 a27529a <=( A298  and  A267 );
 a27530a <=( A266  and  a27529a );
 a27534a <=( (not A302)  and  (not A300) );
 a27535a <=( (not A299)  and  a27534a );
 a27536a <=( a27535a  and  a27530a );
 a27540a <=( (not A199)  and  A166 );
 a27541a <=( A167  and  a27540a );
 a27545a <=( A202  and  (not A201) );
 a27546a <=( A200  and  a27545a );
 a27547a <=( a27546a  and  a27541a );
 a27551a <=( (not A298)  and  A267 );
 a27552a <=( A266  and  a27551a );
 a27556a <=( A301  and  (not A300) );
 a27557a <=( A299  and  a27556a );
 a27558a <=( a27557a  and  a27552a );
 a27562a <=( (not A199)  and  A166 );
 a27563a <=( A167  and  a27562a );
 a27567a <=( A202  and  (not A201) );
 a27568a <=( A200  and  a27567a );
 a27569a <=( a27568a  and  a27563a );
 a27573a <=( (not A298)  and  A267 );
 a27574a <=( A266  and  a27573a );
 a27578a <=( (not A302)  and  (not A300) );
 a27579a <=( A299  and  a27578a );
 a27580a <=( a27579a  and  a27574a );
 a27584a <=( (not A199)  and  A166 );
 a27585a <=( A167  and  a27584a );
 a27589a <=( (not A203)  and  (not A201) );
 a27590a <=( A200  and  a27589a );
 a27591a <=( a27590a  and  a27585a );
 a27595a <=( A298  and  A267 );
 a27596a <=( A265  and  a27595a );
 a27600a <=( (not A301)  and  (not A300) );
 a27601a <=( A299  and  a27600a );
 a27602a <=( a27601a  and  a27596a );
 a27606a <=( (not A199)  and  A166 );
 a27607a <=( A167  and  a27606a );
 a27611a <=( (not A203)  and  (not A201) );
 a27612a <=( A200  and  a27611a );
 a27613a <=( a27612a  and  a27607a );
 a27617a <=( A298  and  A267 );
 a27618a <=( A265  and  a27617a );
 a27622a <=( A302  and  (not A300) );
 a27623a <=( A299  and  a27622a );
 a27624a <=( a27623a  and  a27618a );
 a27628a <=( (not A199)  and  A166 );
 a27629a <=( A167  and  a27628a );
 a27633a <=( (not A203)  and  (not A201) );
 a27634a <=( A200  and  a27633a );
 a27635a <=( a27634a  and  a27629a );
 a27639a <=( A298  and  A267 );
 a27640a <=( A265  and  a27639a );
 a27644a <=( A301  and  (not A300) );
 a27645a <=( (not A299)  and  a27644a );
 a27646a <=( a27645a  and  a27640a );
 a27650a <=( (not A199)  and  A166 );
 a27651a <=( A167  and  a27650a );
 a27655a <=( (not A203)  and  (not A201) );
 a27656a <=( A200  and  a27655a );
 a27657a <=( a27656a  and  a27651a );
 a27661a <=( A298  and  A267 );
 a27662a <=( A265  and  a27661a );
 a27666a <=( (not A302)  and  (not A300) );
 a27667a <=( (not A299)  and  a27666a );
 a27668a <=( a27667a  and  a27662a );
 a27672a <=( (not A199)  and  A166 );
 a27673a <=( A167  and  a27672a );
 a27677a <=( (not A203)  and  (not A201) );
 a27678a <=( A200  and  a27677a );
 a27679a <=( a27678a  and  a27673a );
 a27683a <=( (not A298)  and  A267 );
 a27684a <=( A265  and  a27683a );
 a27688a <=( A301  and  (not A300) );
 a27689a <=( A299  and  a27688a );
 a27690a <=( a27689a  and  a27684a );
 a27694a <=( (not A199)  and  A166 );
 a27695a <=( A167  and  a27694a );
 a27699a <=( (not A203)  and  (not A201) );
 a27700a <=( A200  and  a27699a );
 a27701a <=( a27700a  and  a27695a );
 a27705a <=( (not A298)  and  A267 );
 a27706a <=( A265  and  a27705a );
 a27710a <=( (not A302)  and  (not A300) );
 a27711a <=( A299  and  a27710a );
 a27712a <=( a27711a  and  a27706a );
 a27716a <=( (not A199)  and  A166 );
 a27717a <=( A167  and  a27716a );
 a27721a <=( (not A203)  and  (not A201) );
 a27722a <=( A200  and  a27721a );
 a27723a <=( a27722a  and  a27717a );
 a27727a <=( A298  and  A267 );
 a27728a <=( A266  and  a27727a );
 a27732a <=( (not A301)  and  (not A300) );
 a27733a <=( A299  and  a27732a );
 a27734a <=( a27733a  and  a27728a );
 a27738a <=( (not A199)  and  A166 );
 a27739a <=( A167  and  a27738a );
 a27743a <=( (not A203)  and  (not A201) );
 a27744a <=( A200  and  a27743a );
 a27745a <=( a27744a  and  a27739a );
 a27749a <=( A298  and  A267 );
 a27750a <=( A266  and  a27749a );
 a27754a <=( A302  and  (not A300) );
 a27755a <=( A299  and  a27754a );
 a27756a <=( a27755a  and  a27750a );
 a27760a <=( (not A199)  and  A166 );
 a27761a <=( A167  and  a27760a );
 a27765a <=( (not A203)  and  (not A201) );
 a27766a <=( A200  and  a27765a );
 a27767a <=( a27766a  and  a27761a );
 a27771a <=( A298  and  A267 );
 a27772a <=( A266  and  a27771a );
 a27776a <=( A301  and  (not A300) );
 a27777a <=( (not A299)  and  a27776a );
 a27778a <=( a27777a  and  a27772a );
 a27782a <=( (not A199)  and  A166 );
 a27783a <=( A167  and  a27782a );
 a27787a <=( (not A203)  and  (not A201) );
 a27788a <=( A200  and  a27787a );
 a27789a <=( a27788a  and  a27783a );
 a27793a <=( A298  and  A267 );
 a27794a <=( A266  and  a27793a );
 a27798a <=( (not A302)  and  (not A300) );
 a27799a <=( (not A299)  and  a27798a );
 a27800a <=( a27799a  and  a27794a );
 a27804a <=( (not A199)  and  A166 );
 a27805a <=( A167  and  a27804a );
 a27809a <=( (not A203)  and  (not A201) );
 a27810a <=( A200  and  a27809a );
 a27811a <=( a27810a  and  a27805a );
 a27815a <=( (not A298)  and  A267 );
 a27816a <=( A266  and  a27815a );
 a27820a <=( A301  and  (not A300) );
 a27821a <=( A299  and  a27820a );
 a27822a <=( a27821a  and  a27816a );
 a27826a <=( (not A199)  and  A166 );
 a27827a <=( A167  and  a27826a );
 a27831a <=( (not A203)  and  (not A201) );
 a27832a <=( A200  and  a27831a );
 a27833a <=( a27832a  and  a27827a );
 a27837a <=( (not A298)  and  A267 );
 a27838a <=( A266  and  a27837a );
 a27842a <=( (not A302)  and  (not A300) );
 a27843a <=( A299  and  a27842a );
 a27844a <=( a27843a  and  a27838a );
 a27848a <=( A199  and  A166 );
 a27849a <=( A167  and  a27848a );
 a27853a <=( A203  and  (not A202) );
 a27854a <=( (not A200)  and  a27853a );
 a27855a <=( a27854a  and  a27849a );
 a27859a <=( (not A267)  and  A266 );
 a27860a <=( A265  and  a27859a );
 a27864a <=( A300  and  A299 );
 a27865a <=( (not A268)  and  a27864a );
 a27866a <=( a27865a  and  a27860a );
 a27870a <=( A199  and  A166 );
 a27871a <=( A167  and  a27870a );
 a27875a <=( A203  and  (not A202) );
 a27876a <=( (not A200)  and  a27875a );
 a27877a <=( a27876a  and  a27871a );
 a27881a <=( (not A267)  and  A266 );
 a27882a <=( A265  and  a27881a );
 a27886a <=( A300  and  A298 );
 a27887a <=( (not A268)  and  a27886a );
 a27888a <=( a27887a  and  a27882a );
 a27892a <=( A199  and  A166 );
 a27893a <=( A167  and  a27892a );
 a27897a <=( A203  and  (not A202) );
 a27898a <=( (not A200)  and  a27897a );
 a27899a <=( a27898a  and  a27893a );
 a27903a <=( (not A267)  and  A266 );
 a27904a <=( A265  and  a27903a );
 a27908a <=( A300  and  A299 );
 a27909a <=( A269  and  a27908a );
 a27910a <=( a27909a  and  a27904a );
 a27914a <=( A199  and  A166 );
 a27915a <=( A167  and  a27914a );
 a27919a <=( A203  and  (not A202) );
 a27920a <=( (not A200)  and  a27919a );
 a27921a <=( a27920a  and  a27915a );
 a27925a <=( (not A267)  and  A266 );
 a27926a <=( A265  and  a27925a );
 a27930a <=( A300  and  A298 );
 a27931a <=( A269  and  a27930a );
 a27932a <=( a27931a  and  a27926a );
 a27936a <=( A199  and  A166 );
 a27937a <=( A167  and  a27936a );
 a27941a <=( A203  and  (not A202) );
 a27942a <=( (not A200)  and  a27941a );
 a27943a <=( a27942a  and  a27937a );
 a27947a <=( (not A267)  and  A266 );
 a27948a <=( (not A265)  and  a27947a );
 a27952a <=( A300  and  A299 );
 a27953a <=( A268  and  a27952a );
 a27954a <=( a27953a  and  a27948a );
 a27958a <=( A199  and  A166 );
 a27959a <=( A167  and  a27958a );
 a27963a <=( A203  and  (not A202) );
 a27964a <=( (not A200)  and  a27963a );
 a27965a <=( a27964a  and  a27959a );
 a27969a <=( (not A267)  and  A266 );
 a27970a <=( (not A265)  and  a27969a );
 a27974a <=( A300  and  A298 );
 a27975a <=( A268  and  a27974a );
 a27976a <=( a27975a  and  a27970a );
 a27980a <=( A199  and  A166 );
 a27981a <=( A167  and  a27980a );
 a27985a <=( A203  and  (not A202) );
 a27986a <=( (not A200)  and  a27985a );
 a27987a <=( a27986a  and  a27981a );
 a27991a <=( (not A267)  and  A266 );
 a27992a <=( (not A265)  and  a27991a );
 a27996a <=( A300  and  A299 );
 a27997a <=( (not A269)  and  a27996a );
 a27998a <=( a27997a  and  a27992a );
 a28002a <=( A199  and  A166 );
 a28003a <=( A167  and  a28002a );
 a28007a <=( A203  and  (not A202) );
 a28008a <=( (not A200)  and  a28007a );
 a28009a <=( a28008a  and  a28003a );
 a28013a <=( (not A267)  and  A266 );
 a28014a <=( (not A265)  and  a28013a );
 a28018a <=( A300  and  A298 );
 a28019a <=( (not A269)  and  a28018a );
 a28020a <=( a28019a  and  a28014a );
 a28024a <=( A199  and  A166 );
 a28025a <=( A167  and  a28024a );
 a28029a <=( A203  and  (not A202) );
 a28030a <=( (not A200)  and  a28029a );
 a28031a <=( a28030a  and  a28025a );
 a28035a <=( (not A267)  and  (not A266) );
 a28036a <=( A265  and  a28035a );
 a28040a <=( A300  and  A299 );
 a28041a <=( A268  and  a28040a );
 a28042a <=( a28041a  and  a28036a );
 a28046a <=( A199  and  A166 );
 a28047a <=( A167  and  a28046a );
 a28051a <=( A203  and  (not A202) );
 a28052a <=( (not A200)  and  a28051a );
 a28053a <=( a28052a  and  a28047a );
 a28057a <=( (not A267)  and  (not A266) );
 a28058a <=( A265  and  a28057a );
 a28062a <=( A300  and  A298 );
 a28063a <=( A268  and  a28062a );
 a28064a <=( a28063a  and  a28058a );
 a28068a <=( A199  and  A166 );
 a28069a <=( A167  and  a28068a );
 a28073a <=( A203  and  (not A202) );
 a28074a <=( (not A200)  and  a28073a );
 a28075a <=( a28074a  and  a28069a );
 a28079a <=( (not A267)  and  (not A266) );
 a28080a <=( A265  and  a28079a );
 a28084a <=( A300  and  A299 );
 a28085a <=( (not A269)  and  a28084a );
 a28086a <=( a28085a  and  a28080a );
 a28090a <=( A199  and  A166 );
 a28091a <=( A167  and  a28090a );
 a28095a <=( A203  and  (not A202) );
 a28096a <=( (not A200)  and  a28095a );
 a28097a <=( a28096a  and  a28091a );
 a28101a <=( (not A267)  and  (not A266) );
 a28102a <=( A265  and  a28101a );
 a28106a <=( A300  and  A298 );
 a28107a <=( (not A269)  and  a28106a );
 a28108a <=( a28107a  and  a28102a );
 a28112a <=( A199  and  A166 );
 a28113a <=( A167  and  a28112a );
 a28117a <=( A202  and  (not A201) );
 a28118a <=( (not A200)  and  a28117a );
 a28119a <=( a28118a  and  a28113a );
 a28123a <=( A298  and  A267 );
 a28124a <=( A265  and  a28123a );
 a28128a <=( (not A301)  and  (not A300) );
 a28129a <=( A299  and  a28128a );
 a28130a <=( a28129a  and  a28124a );
 a28134a <=( A199  and  A166 );
 a28135a <=( A167  and  a28134a );
 a28139a <=( A202  and  (not A201) );
 a28140a <=( (not A200)  and  a28139a );
 a28141a <=( a28140a  and  a28135a );
 a28145a <=( A298  and  A267 );
 a28146a <=( A265  and  a28145a );
 a28150a <=( A302  and  (not A300) );
 a28151a <=( A299  and  a28150a );
 a28152a <=( a28151a  and  a28146a );
 a28156a <=( A199  and  A166 );
 a28157a <=( A167  and  a28156a );
 a28161a <=( A202  and  (not A201) );
 a28162a <=( (not A200)  and  a28161a );
 a28163a <=( a28162a  and  a28157a );
 a28167a <=( A298  and  A267 );
 a28168a <=( A265  and  a28167a );
 a28172a <=( A301  and  (not A300) );
 a28173a <=( (not A299)  and  a28172a );
 a28174a <=( a28173a  and  a28168a );
 a28178a <=( A199  and  A166 );
 a28179a <=( A167  and  a28178a );
 a28183a <=( A202  and  (not A201) );
 a28184a <=( (not A200)  and  a28183a );
 a28185a <=( a28184a  and  a28179a );
 a28189a <=( A298  and  A267 );
 a28190a <=( A265  and  a28189a );
 a28194a <=( (not A302)  and  (not A300) );
 a28195a <=( (not A299)  and  a28194a );
 a28196a <=( a28195a  and  a28190a );
 a28200a <=( A199  and  A166 );
 a28201a <=( A167  and  a28200a );
 a28205a <=( A202  and  (not A201) );
 a28206a <=( (not A200)  and  a28205a );
 a28207a <=( a28206a  and  a28201a );
 a28211a <=( (not A298)  and  A267 );
 a28212a <=( A265  and  a28211a );
 a28216a <=( A301  and  (not A300) );
 a28217a <=( A299  and  a28216a );
 a28218a <=( a28217a  and  a28212a );
 a28222a <=( A199  and  A166 );
 a28223a <=( A167  and  a28222a );
 a28227a <=( A202  and  (not A201) );
 a28228a <=( (not A200)  and  a28227a );
 a28229a <=( a28228a  and  a28223a );
 a28233a <=( (not A298)  and  A267 );
 a28234a <=( A265  and  a28233a );
 a28238a <=( (not A302)  and  (not A300) );
 a28239a <=( A299  and  a28238a );
 a28240a <=( a28239a  and  a28234a );
 a28244a <=( A199  and  A166 );
 a28245a <=( A167  and  a28244a );
 a28249a <=( A202  and  (not A201) );
 a28250a <=( (not A200)  and  a28249a );
 a28251a <=( a28250a  and  a28245a );
 a28255a <=( A298  and  A267 );
 a28256a <=( A266  and  a28255a );
 a28260a <=( (not A301)  and  (not A300) );
 a28261a <=( A299  and  a28260a );
 a28262a <=( a28261a  and  a28256a );
 a28266a <=( A199  and  A166 );
 a28267a <=( A167  and  a28266a );
 a28271a <=( A202  and  (not A201) );
 a28272a <=( (not A200)  and  a28271a );
 a28273a <=( a28272a  and  a28267a );
 a28277a <=( A298  and  A267 );
 a28278a <=( A266  and  a28277a );
 a28282a <=( A302  and  (not A300) );
 a28283a <=( A299  and  a28282a );
 a28284a <=( a28283a  and  a28278a );
 a28288a <=( A199  and  A166 );
 a28289a <=( A167  and  a28288a );
 a28293a <=( A202  and  (not A201) );
 a28294a <=( (not A200)  and  a28293a );
 a28295a <=( a28294a  and  a28289a );
 a28299a <=( A298  and  A267 );
 a28300a <=( A266  and  a28299a );
 a28304a <=( A301  and  (not A300) );
 a28305a <=( (not A299)  and  a28304a );
 a28306a <=( a28305a  and  a28300a );
 a28310a <=( A199  and  A166 );
 a28311a <=( A167  and  a28310a );
 a28315a <=( A202  and  (not A201) );
 a28316a <=( (not A200)  and  a28315a );
 a28317a <=( a28316a  and  a28311a );
 a28321a <=( A298  and  A267 );
 a28322a <=( A266  and  a28321a );
 a28326a <=( (not A302)  and  (not A300) );
 a28327a <=( (not A299)  and  a28326a );
 a28328a <=( a28327a  and  a28322a );
 a28332a <=( A199  and  A166 );
 a28333a <=( A167  and  a28332a );
 a28337a <=( A202  and  (not A201) );
 a28338a <=( (not A200)  and  a28337a );
 a28339a <=( a28338a  and  a28333a );
 a28343a <=( (not A298)  and  A267 );
 a28344a <=( A266  and  a28343a );
 a28348a <=( A301  and  (not A300) );
 a28349a <=( A299  and  a28348a );
 a28350a <=( a28349a  and  a28344a );
 a28354a <=( A199  and  A166 );
 a28355a <=( A167  and  a28354a );
 a28359a <=( A202  and  (not A201) );
 a28360a <=( (not A200)  and  a28359a );
 a28361a <=( a28360a  and  a28355a );
 a28365a <=( (not A298)  and  A267 );
 a28366a <=( A266  and  a28365a );
 a28370a <=( (not A302)  and  (not A300) );
 a28371a <=( A299  and  a28370a );
 a28372a <=( a28371a  and  a28366a );
 a28376a <=( A199  and  A166 );
 a28377a <=( A167  and  a28376a );
 a28381a <=( (not A203)  and  (not A201) );
 a28382a <=( (not A200)  and  a28381a );
 a28383a <=( a28382a  and  a28377a );
 a28387a <=( A298  and  A267 );
 a28388a <=( A265  and  a28387a );
 a28392a <=( (not A301)  and  (not A300) );
 a28393a <=( A299  and  a28392a );
 a28394a <=( a28393a  and  a28388a );
 a28398a <=( A199  and  A166 );
 a28399a <=( A167  and  a28398a );
 a28403a <=( (not A203)  and  (not A201) );
 a28404a <=( (not A200)  and  a28403a );
 a28405a <=( a28404a  and  a28399a );
 a28409a <=( A298  and  A267 );
 a28410a <=( A265  and  a28409a );
 a28414a <=( A302  and  (not A300) );
 a28415a <=( A299  and  a28414a );
 a28416a <=( a28415a  and  a28410a );
 a28420a <=( A199  and  A166 );
 a28421a <=( A167  and  a28420a );
 a28425a <=( (not A203)  and  (not A201) );
 a28426a <=( (not A200)  and  a28425a );
 a28427a <=( a28426a  and  a28421a );
 a28431a <=( A298  and  A267 );
 a28432a <=( A265  and  a28431a );
 a28436a <=( A301  and  (not A300) );
 a28437a <=( (not A299)  and  a28436a );
 a28438a <=( a28437a  and  a28432a );
 a28442a <=( A199  and  A166 );
 a28443a <=( A167  and  a28442a );
 a28447a <=( (not A203)  and  (not A201) );
 a28448a <=( (not A200)  and  a28447a );
 a28449a <=( a28448a  and  a28443a );
 a28453a <=( A298  and  A267 );
 a28454a <=( A265  and  a28453a );
 a28458a <=( (not A302)  and  (not A300) );
 a28459a <=( (not A299)  and  a28458a );
 a28460a <=( a28459a  and  a28454a );
 a28464a <=( A199  and  A166 );
 a28465a <=( A167  and  a28464a );
 a28469a <=( (not A203)  and  (not A201) );
 a28470a <=( (not A200)  and  a28469a );
 a28471a <=( a28470a  and  a28465a );
 a28475a <=( (not A298)  and  A267 );
 a28476a <=( A265  and  a28475a );
 a28480a <=( A301  and  (not A300) );
 a28481a <=( A299  and  a28480a );
 a28482a <=( a28481a  and  a28476a );
 a28486a <=( A199  and  A166 );
 a28487a <=( A167  and  a28486a );
 a28491a <=( (not A203)  and  (not A201) );
 a28492a <=( (not A200)  and  a28491a );
 a28493a <=( a28492a  and  a28487a );
 a28497a <=( (not A298)  and  A267 );
 a28498a <=( A265  and  a28497a );
 a28502a <=( (not A302)  and  (not A300) );
 a28503a <=( A299  and  a28502a );
 a28504a <=( a28503a  and  a28498a );
 a28508a <=( A199  and  A166 );
 a28509a <=( A167  and  a28508a );
 a28513a <=( (not A203)  and  (not A201) );
 a28514a <=( (not A200)  and  a28513a );
 a28515a <=( a28514a  and  a28509a );
 a28519a <=( A298  and  A267 );
 a28520a <=( A266  and  a28519a );
 a28524a <=( (not A301)  and  (not A300) );
 a28525a <=( A299  and  a28524a );
 a28526a <=( a28525a  and  a28520a );
 a28530a <=( A199  and  A166 );
 a28531a <=( A167  and  a28530a );
 a28535a <=( (not A203)  and  (not A201) );
 a28536a <=( (not A200)  and  a28535a );
 a28537a <=( a28536a  and  a28531a );
 a28541a <=( A298  and  A267 );
 a28542a <=( A266  and  a28541a );
 a28546a <=( A302  and  (not A300) );
 a28547a <=( A299  and  a28546a );
 a28548a <=( a28547a  and  a28542a );
 a28552a <=( A199  and  A166 );
 a28553a <=( A167  and  a28552a );
 a28557a <=( (not A203)  and  (not A201) );
 a28558a <=( (not A200)  and  a28557a );
 a28559a <=( a28558a  and  a28553a );
 a28563a <=( A298  and  A267 );
 a28564a <=( A266  and  a28563a );
 a28568a <=( A301  and  (not A300) );
 a28569a <=( (not A299)  and  a28568a );
 a28570a <=( a28569a  and  a28564a );
 a28574a <=( A199  and  A166 );
 a28575a <=( A167  and  a28574a );
 a28579a <=( (not A203)  and  (not A201) );
 a28580a <=( (not A200)  and  a28579a );
 a28581a <=( a28580a  and  a28575a );
 a28585a <=( A298  and  A267 );
 a28586a <=( A266  and  a28585a );
 a28590a <=( (not A302)  and  (not A300) );
 a28591a <=( (not A299)  and  a28590a );
 a28592a <=( a28591a  and  a28586a );
 a28596a <=( A199  and  A166 );
 a28597a <=( A167  and  a28596a );
 a28601a <=( (not A203)  and  (not A201) );
 a28602a <=( (not A200)  and  a28601a );
 a28603a <=( a28602a  and  a28597a );
 a28607a <=( (not A298)  and  A267 );
 a28608a <=( A266  and  a28607a );
 a28612a <=( A301  and  (not A300) );
 a28613a <=( A299  and  a28612a );
 a28614a <=( a28613a  and  a28608a );
 a28618a <=( A199  and  A166 );
 a28619a <=( A167  and  a28618a );
 a28623a <=( (not A203)  and  (not A201) );
 a28624a <=( (not A200)  and  a28623a );
 a28625a <=( a28624a  and  a28619a );
 a28629a <=( (not A298)  and  A267 );
 a28630a <=( A266  and  a28629a );
 a28634a <=( (not A302)  and  (not A300) );
 a28635a <=( A299  and  a28634a );
 a28636a <=( a28635a  and  a28630a );
 a28640a <=( (not A199)  and  A166 );
 a28641a <=( A167  and  a28640a );
 a28645a <=( A265  and  (not A202) );
 a28646a <=( (not A200)  and  a28645a );
 a28647a <=( a28646a  and  a28641a );
 a28651a <=( (not A269)  and  A268 );
 a28652a <=( A266  and  a28651a );
 a28656a <=( (not A301)  and  (not A299) );
 a28657a <=( (not A298)  and  a28656a );
 a28658a <=( a28657a  and  a28652a );
 a28662a <=( (not A199)  and  A166 );
 a28663a <=( A167  and  a28662a );
 a28667a <=( A265  and  (not A202) );
 a28668a <=( (not A200)  and  a28667a );
 a28669a <=( a28668a  and  a28663a );
 a28673a <=( (not A269)  and  A268 );
 a28674a <=( A266  and  a28673a );
 a28678a <=( A302  and  (not A299) );
 a28679a <=( (not A298)  and  a28678a );
 a28680a <=( a28679a  and  a28674a );
 a28684a <=( (not A199)  and  A166 );
 a28685a <=( A167  and  a28684a );
 a28689a <=( (not A265)  and  (not A202) );
 a28690a <=( (not A200)  and  a28689a );
 a28691a <=( a28690a  and  a28685a );
 a28695a <=( A269  and  (not A268) );
 a28696a <=( A266  and  a28695a );
 a28700a <=( (not A301)  and  (not A299) );
 a28701a <=( (not A298)  and  a28700a );
 a28702a <=( a28701a  and  a28696a );
 a28706a <=( (not A199)  and  A166 );
 a28707a <=( A167  and  a28706a );
 a28711a <=( (not A265)  and  (not A202) );
 a28712a <=( (not A200)  and  a28711a );
 a28713a <=( a28712a  and  a28707a );
 a28717a <=( A269  and  (not A268) );
 a28718a <=( A266  and  a28717a );
 a28722a <=( A302  and  (not A299) );
 a28723a <=( (not A298)  and  a28722a );
 a28724a <=( a28723a  and  a28718a );
 a28728a <=( (not A199)  and  A166 );
 a28729a <=( A167  and  a28728a );
 a28733a <=( A265  and  (not A202) );
 a28734a <=( (not A200)  and  a28733a );
 a28735a <=( a28734a  and  a28729a );
 a28739a <=( A269  and  (not A268) );
 a28740a <=( (not A266)  and  a28739a );
 a28744a <=( (not A301)  and  (not A299) );
 a28745a <=( (not A298)  and  a28744a );
 a28746a <=( a28745a  and  a28740a );
 a28750a <=( (not A199)  and  A166 );
 a28751a <=( A167  and  a28750a );
 a28755a <=( A265  and  (not A202) );
 a28756a <=( (not A200)  and  a28755a );
 a28757a <=( a28756a  and  a28751a );
 a28761a <=( A269  and  (not A268) );
 a28762a <=( (not A266)  and  a28761a );
 a28766a <=( A302  and  (not A299) );
 a28767a <=( (not A298)  and  a28766a );
 a28768a <=( a28767a  and  a28762a );
 a28772a <=( (not A199)  and  A166 );
 a28773a <=( A167  and  a28772a );
 a28777a <=( (not A265)  and  (not A202) );
 a28778a <=( (not A200)  and  a28777a );
 a28779a <=( a28778a  and  a28773a );
 a28783a <=( (not A269)  and  A268 );
 a28784a <=( (not A266)  and  a28783a );
 a28788a <=( (not A301)  and  (not A299) );
 a28789a <=( (not A298)  and  a28788a );
 a28790a <=( a28789a  and  a28784a );
 a28794a <=( (not A199)  and  A166 );
 a28795a <=( A167  and  a28794a );
 a28799a <=( (not A265)  and  (not A202) );
 a28800a <=( (not A200)  and  a28799a );
 a28801a <=( a28800a  and  a28795a );
 a28805a <=( (not A269)  and  A268 );
 a28806a <=( (not A266)  and  a28805a );
 a28810a <=( A302  and  (not A299) );
 a28811a <=( (not A298)  and  a28810a );
 a28812a <=( a28811a  and  a28806a );
 a28816a <=( (not A199)  and  A166 );
 a28817a <=( A167  and  a28816a );
 a28821a <=( A265  and  A203 );
 a28822a <=( (not A200)  and  a28821a );
 a28823a <=( a28822a  and  a28817a );
 a28827a <=( (not A269)  and  A268 );
 a28828a <=( A266  and  a28827a );
 a28832a <=( (not A301)  and  (not A299) );
 a28833a <=( (not A298)  and  a28832a );
 a28834a <=( a28833a  and  a28828a );
 a28838a <=( (not A199)  and  A166 );
 a28839a <=( A167  and  a28838a );
 a28843a <=( A265  and  A203 );
 a28844a <=( (not A200)  and  a28843a );
 a28845a <=( a28844a  and  a28839a );
 a28849a <=( (not A269)  and  A268 );
 a28850a <=( A266  and  a28849a );
 a28854a <=( A302  and  (not A299) );
 a28855a <=( (not A298)  and  a28854a );
 a28856a <=( a28855a  and  a28850a );
 a28860a <=( (not A199)  and  A166 );
 a28861a <=( A167  and  a28860a );
 a28865a <=( (not A265)  and  A203 );
 a28866a <=( (not A200)  and  a28865a );
 a28867a <=( a28866a  and  a28861a );
 a28871a <=( A269  and  (not A268) );
 a28872a <=( A266  and  a28871a );
 a28876a <=( (not A301)  and  (not A299) );
 a28877a <=( (not A298)  and  a28876a );
 a28878a <=( a28877a  and  a28872a );
 a28882a <=( (not A199)  and  A166 );
 a28883a <=( A167  and  a28882a );
 a28887a <=( (not A265)  and  A203 );
 a28888a <=( (not A200)  and  a28887a );
 a28889a <=( a28888a  and  a28883a );
 a28893a <=( A269  and  (not A268) );
 a28894a <=( A266  and  a28893a );
 a28898a <=( A302  and  (not A299) );
 a28899a <=( (not A298)  and  a28898a );
 a28900a <=( a28899a  and  a28894a );
 a28904a <=( (not A199)  and  A166 );
 a28905a <=( A167  and  a28904a );
 a28909a <=( A265  and  A203 );
 a28910a <=( (not A200)  and  a28909a );
 a28911a <=( a28910a  and  a28905a );
 a28915a <=( A269  and  (not A268) );
 a28916a <=( (not A266)  and  a28915a );
 a28920a <=( (not A301)  and  (not A299) );
 a28921a <=( (not A298)  and  a28920a );
 a28922a <=( a28921a  and  a28916a );
 a28926a <=( (not A199)  and  A166 );
 a28927a <=( A167  and  a28926a );
 a28931a <=( A265  and  A203 );
 a28932a <=( (not A200)  and  a28931a );
 a28933a <=( a28932a  and  a28927a );
 a28937a <=( A269  and  (not A268) );
 a28938a <=( (not A266)  and  a28937a );
 a28942a <=( A302  and  (not A299) );
 a28943a <=( (not A298)  and  a28942a );
 a28944a <=( a28943a  and  a28938a );
 a28948a <=( (not A199)  and  A166 );
 a28949a <=( A167  and  a28948a );
 a28953a <=( (not A265)  and  A203 );
 a28954a <=( (not A200)  and  a28953a );
 a28955a <=( a28954a  and  a28949a );
 a28959a <=( (not A269)  and  A268 );
 a28960a <=( (not A266)  and  a28959a );
 a28964a <=( (not A301)  and  (not A299) );
 a28965a <=( (not A298)  and  a28964a );
 a28966a <=( a28965a  and  a28960a );
 a28970a <=( (not A199)  and  A166 );
 a28971a <=( A167  and  a28970a );
 a28975a <=( (not A265)  and  A203 );
 a28976a <=( (not A200)  and  a28975a );
 a28977a <=( a28976a  and  a28971a );
 a28981a <=( (not A269)  and  A268 );
 a28982a <=( (not A266)  and  a28981a );
 a28986a <=( A302  and  (not A299) );
 a28987a <=( (not A298)  and  a28986a );
 a28988a <=( a28987a  and  a28982a );
 a28992a <=( (not A199)  and  A166 );
 a28993a <=( A167  and  a28992a );
 a28997a <=( (not A203)  and  A202 );
 a28998a <=( (not A200)  and  a28997a );
 a28999a <=( a28998a  and  a28993a );
 a29003a <=( (not A267)  and  A266 );
 a29004a <=( A265  and  a29003a );
 a29008a <=( A300  and  A299 );
 a29009a <=( (not A268)  and  a29008a );
 a29010a <=( a29009a  and  a29004a );
 a29014a <=( (not A199)  and  A166 );
 a29015a <=( A167  and  a29014a );
 a29019a <=( (not A203)  and  A202 );
 a29020a <=( (not A200)  and  a29019a );
 a29021a <=( a29020a  and  a29015a );
 a29025a <=( (not A267)  and  A266 );
 a29026a <=( A265  and  a29025a );
 a29030a <=( A300  and  A298 );
 a29031a <=( (not A268)  and  a29030a );
 a29032a <=( a29031a  and  a29026a );
 a29036a <=( (not A199)  and  A166 );
 a29037a <=( A167  and  a29036a );
 a29041a <=( (not A203)  and  A202 );
 a29042a <=( (not A200)  and  a29041a );
 a29043a <=( a29042a  and  a29037a );
 a29047a <=( (not A267)  and  A266 );
 a29048a <=( A265  and  a29047a );
 a29052a <=( A300  and  A299 );
 a29053a <=( A269  and  a29052a );
 a29054a <=( a29053a  and  a29048a );
 a29058a <=( (not A199)  and  A166 );
 a29059a <=( A167  and  a29058a );
 a29063a <=( (not A203)  and  A202 );
 a29064a <=( (not A200)  and  a29063a );
 a29065a <=( a29064a  and  a29059a );
 a29069a <=( (not A267)  and  A266 );
 a29070a <=( A265  and  a29069a );
 a29074a <=( A300  and  A298 );
 a29075a <=( A269  and  a29074a );
 a29076a <=( a29075a  and  a29070a );
 a29080a <=( (not A199)  and  A166 );
 a29081a <=( A167  and  a29080a );
 a29085a <=( (not A203)  and  A202 );
 a29086a <=( (not A200)  and  a29085a );
 a29087a <=( a29086a  and  a29081a );
 a29091a <=( (not A267)  and  A266 );
 a29092a <=( (not A265)  and  a29091a );
 a29096a <=( A300  and  A299 );
 a29097a <=( A268  and  a29096a );
 a29098a <=( a29097a  and  a29092a );
 a29102a <=( (not A199)  and  A166 );
 a29103a <=( A167  and  a29102a );
 a29107a <=( (not A203)  and  A202 );
 a29108a <=( (not A200)  and  a29107a );
 a29109a <=( a29108a  and  a29103a );
 a29113a <=( (not A267)  and  A266 );
 a29114a <=( (not A265)  and  a29113a );
 a29118a <=( A300  and  A298 );
 a29119a <=( A268  and  a29118a );
 a29120a <=( a29119a  and  a29114a );
 a29124a <=( (not A199)  and  A166 );
 a29125a <=( A167  and  a29124a );
 a29129a <=( (not A203)  and  A202 );
 a29130a <=( (not A200)  and  a29129a );
 a29131a <=( a29130a  and  a29125a );
 a29135a <=( (not A267)  and  A266 );
 a29136a <=( (not A265)  and  a29135a );
 a29140a <=( A300  and  A299 );
 a29141a <=( (not A269)  and  a29140a );
 a29142a <=( a29141a  and  a29136a );
 a29146a <=( (not A199)  and  A166 );
 a29147a <=( A167  and  a29146a );
 a29151a <=( (not A203)  and  A202 );
 a29152a <=( (not A200)  and  a29151a );
 a29153a <=( a29152a  and  a29147a );
 a29157a <=( (not A267)  and  A266 );
 a29158a <=( (not A265)  and  a29157a );
 a29162a <=( A300  and  A298 );
 a29163a <=( (not A269)  and  a29162a );
 a29164a <=( a29163a  and  a29158a );
 a29168a <=( (not A199)  and  A166 );
 a29169a <=( A167  and  a29168a );
 a29173a <=( (not A203)  and  A202 );
 a29174a <=( (not A200)  and  a29173a );
 a29175a <=( a29174a  and  a29169a );
 a29179a <=( (not A267)  and  (not A266) );
 a29180a <=( A265  and  a29179a );
 a29184a <=( A300  and  A299 );
 a29185a <=( A268  and  a29184a );
 a29186a <=( a29185a  and  a29180a );
 a29190a <=( (not A199)  and  A166 );
 a29191a <=( A167  and  a29190a );
 a29195a <=( (not A203)  and  A202 );
 a29196a <=( (not A200)  and  a29195a );
 a29197a <=( a29196a  and  a29191a );
 a29201a <=( (not A267)  and  (not A266) );
 a29202a <=( A265  and  a29201a );
 a29206a <=( A300  and  A298 );
 a29207a <=( A268  and  a29206a );
 a29208a <=( a29207a  and  a29202a );
 a29212a <=( (not A199)  and  A166 );
 a29213a <=( A167  and  a29212a );
 a29217a <=( (not A203)  and  A202 );
 a29218a <=( (not A200)  and  a29217a );
 a29219a <=( a29218a  and  a29213a );
 a29223a <=( (not A267)  and  (not A266) );
 a29224a <=( A265  and  a29223a );
 a29228a <=( A300  and  A299 );
 a29229a <=( (not A269)  and  a29228a );
 a29230a <=( a29229a  and  a29224a );
 a29234a <=( (not A199)  and  A166 );
 a29235a <=( A167  and  a29234a );
 a29239a <=( (not A203)  and  A202 );
 a29240a <=( (not A200)  and  a29239a );
 a29241a <=( a29240a  and  a29235a );
 a29245a <=( (not A267)  and  (not A266) );
 a29246a <=( A265  and  a29245a );
 a29250a <=( A300  and  A298 );
 a29251a <=( (not A269)  and  a29250a );
 a29252a <=( a29251a  and  a29246a );
 a29256a <=( A199  and  (not A166) );
 a29257a <=( A167  and  a29256a );
 a29261a <=( A266  and  A265 );
 a29262a <=( A201  and  a29261a );
 a29263a <=( a29262a  and  a29257a );
 a29267a <=( A298  and  (not A269) );
 a29268a <=( A268  and  a29267a );
 a29272a <=( (not A301)  and  (not A300) );
 a29273a <=( A299  and  a29272a );
 a29274a <=( a29273a  and  a29268a );
 a29278a <=( A199  and  (not A166) );
 a29279a <=( A167  and  a29278a );
 a29283a <=( A266  and  A265 );
 a29284a <=( A201  and  a29283a );
 a29285a <=( a29284a  and  a29279a );
 a29289a <=( A298  and  (not A269) );
 a29290a <=( A268  and  a29289a );
 a29294a <=( A302  and  (not A300) );
 a29295a <=( A299  and  a29294a );
 a29296a <=( a29295a  and  a29290a );
 a29300a <=( A199  and  (not A166) );
 a29301a <=( A167  and  a29300a );
 a29305a <=( A266  and  A265 );
 a29306a <=( A201  and  a29305a );
 a29307a <=( a29306a  and  a29301a );
 a29311a <=( A298  and  (not A269) );
 a29312a <=( A268  and  a29311a );
 a29316a <=( A301  and  (not A300) );
 a29317a <=( (not A299)  and  a29316a );
 a29318a <=( a29317a  and  a29312a );
 a29322a <=( A199  and  (not A166) );
 a29323a <=( A167  and  a29322a );
 a29327a <=( A266  and  A265 );
 a29328a <=( A201  and  a29327a );
 a29329a <=( a29328a  and  a29323a );
 a29333a <=( A298  and  (not A269) );
 a29334a <=( A268  and  a29333a );
 a29338a <=( (not A302)  and  (not A300) );
 a29339a <=( (not A299)  and  a29338a );
 a29340a <=( a29339a  and  a29334a );
 a29344a <=( A199  and  (not A166) );
 a29345a <=( A167  and  a29344a );
 a29349a <=( A266  and  A265 );
 a29350a <=( A201  and  a29349a );
 a29351a <=( a29350a  and  a29345a );
 a29355a <=( (not A298)  and  (not A269) );
 a29356a <=( A268  and  a29355a );
 a29360a <=( A301  and  (not A300) );
 a29361a <=( A299  and  a29360a );
 a29362a <=( a29361a  and  a29356a );
 a29366a <=( A199  and  (not A166) );
 a29367a <=( A167  and  a29366a );
 a29371a <=( A266  and  A265 );
 a29372a <=( A201  and  a29371a );
 a29373a <=( a29372a  and  a29367a );
 a29377a <=( (not A298)  and  (not A269) );
 a29378a <=( A268  and  a29377a );
 a29382a <=( (not A302)  and  (not A300) );
 a29383a <=( A299  and  a29382a );
 a29384a <=( a29383a  and  a29378a );
 a29388a <=( A199  and  (not A166) );
 a29389a <=( A167  and  a29388a );
 a29393a <=( A266  and  (not A265) );
 a29394a <=( A201  and  a29393a );
 a29395a <=( a29394a  and  a29389a );
 a29399a <=( A298  and  A269 );
 a29400a <=( (not A268)  and  a29399a );
 a29404a <=( (not A301)  and  (not A300) );
 a29405a <=( A299  and  a29404a );
 a29406a <=( a29405a  and  a29400a );
 a29410a <=( A199  and  (not A166) );
 a29411a <=( A167  and  a29410a );
 a29415a <=( A266  and  (not A265) );
 a29416a <=( A201  and  a29415a );
 a29417a <=( a29416a  and  a29411a );
 a29421a <=( A298  and  A269 );
 a29422a <=( (not A268)  and  a29421a );
 a29426a <=( A302  and  (not A300) );
 a29427a <=( A299  and  a29426a );
 a29428a <=( a29427a  and  a29422a );
 a29432a <=( A199  and  (not A166) );
 a29433a <=( A167  and  a29432a );
 a29437a <=( A266  and  (not A265) );
 a29438a <=( A201  and  a29437a );
 a29439a <=( a29438a  and  a29433a );
 a29443a <=( A298  and  A269 );
 a29444a <=( (not A268)  and  a29443a );
 a29448a <=( A301  and  (not A300) );
 a29449a <=( (not A299)  and  a29448a );
 a29450a <=( a29449a  and  a29444a );
 a29454a <=( A199  and  (not A166) );
 a29455a <=( A167  and  a29454a );
 a29459a <=( A266  and  (not A265) );
 a29460a <=( A201  and  a29459a );
 a29461a <=( a29460a  and  a29455a );
 a29465a <=( A298  and  A269 );
 a29466a <=( (not A268)  and  a29465a );
 a29470a <=( (not A302)  and  (not A300) );
 a29471a <=( (not A299)  and  a29470a );
 a29472a <=( a29471a  and  a29466a );
 a29476a <=( A199  and  (not A166) );
 a29477a <=( A167  and  a29476a );
 a29481a <=( A266  and  (not A265) );
 a29482a <=( A201  and  a29481a );
 a29483a <=( a29482a  and  a29477a );
 a29487a <=( (not A298)  and  A269 );
 a29488a <=( (not A268)  and  a29487a );
 a29492a <=( A301  and  (not A300) );
 a29493a <=( A299  and  a29492a );
 a29494a <=( a29493a  and  a29488a );
 a29498a <=( A199  and  (not A166) );
 a29499a <=( A167  and  a29498a );
 a29503a <=( A266  and  (not A265) );
 a29504a <=( A201  and  a29503a );
 a29505a <=( a29504a  and  a29499a );
 a29509a <=( (not A298)  and  A269 );
 a29510a <=( (not A268)  and  a29509a );
 a29514a <=( (not A302)  and  (not A300) );
 a29515a <=( A299  and  a29514a );
 a29516a <=( a29515a  and  a29510a );
 a29520a <=( A199  and  (not A166) );
 a29521a <=( A167  and  a29520a );
 a29525a <=( (not A266)  and  A265 );
 a29526a <=( A201  and  a29525a );
 a29527a <=( a29526a  and  a29521a );
 a29531a <=( A298  and  A269 );
 a29532a <=( (not A268)  and  a29531a );
 a29536a <=( (not A301)  and  (not A300) );
 a29537a <=( A299  and  a29536a );
 a29538a <=( a29537a  and  a29532a );
 a29542a <=( A199  and  (not A166) );
 a29543a <=( A167  and  a29542a );
 a29547a <=( (not A266)  and  A265 );
 a29548a <=( A201  and  a29547a );
 a29549a <=( a29548a  and  a29543a );
 a29553a <=( A298  and  A269 );
 a29554a <=( (not A268)  and  a29553a );
 a29558a <=( A302  and  (not A300) );
 a29559a <=( A299  and  a29558a );
 a29560a <=( a29559a  and  a29554a );
 a29564a <=( A199  and  (not A166) );
 a29565a <=( A167  and  a29564a );
 a29569a <=( (not A266)  and  A265 );
 a29570a <=( A201  and  a29569a );
 a29571a <=( a29570a  and  a29565a );
 a29575a <=( A298  and  A269 );
 a29576a <=( (not A268)  and  a29575a );
 a29580a <=( A301  and  (not A300) );
 a29581a <=( (not A299)  and  a29580a );
 a29582a <=( a29581a  and  a29576a );
 a29586a <=( A199  and  (not A166) );
 a29587a <=( A167  and  a29586a );
 a29591a <=( (not A266)  and  A265 );
 a29592a <=( A201  and  a29591a );
 a29593a <=( a29592a  and  a29587a );
 a29597a <=( A298  and  A269 );
 a29598a <=( (not A268)  and  a29597a );
 a29602a <=( (not A302)  and  (not A300) );
 a29603a <=( (not A299)  and  a29602a );
 a29604a <=( a29603a  and  a29598a );
 a29608a <=( A199  and  (not A166) );
 a29609a <=( A167  and  a29608a );
 a29613a <=( (not A266)  and  A265 );
 a29614a <=( A201  and  a29613a );
 a29615a <=( a29614a  and  a29609a );
 a29619a <=( (not A298)  and  A269 );
 a29620a <=( (not A268)  and  a29619a );
 a29624a <=( A301  and  (not A300) );
 a29625a <=( A299  and  a29624a );
 a29626a <=( a29625a  and  a29620a );
 a29630a <=( A199  and  (not A166) );
 a29631a <=( A167  and  a29630a );
 a29635a <=( (not A266)  and  A265 );
 a29636a <=( A201  and  a29635a );
 a29637a <=( a29636a  and  a29631a );
 a29641a <=( (not A298)  and  A269 );
 a29642a <=( (not A268)  and  a29641a );
 a29646a <=( (not A302)  and  (not A300) );
 a29647a <=( A299  and  a29646a );
 a29648a <=( a29647a  and  a29642a );
 a29652a <=( A199  and  (not A166) );
 a29653a <=( A167  and  a29652a );
 a29657a <=( (not A266)  and  (not A265) );
 a29658a <=( A201  and  a29657a );
 a29659a <=( a29658a  and  a29653a );
 a29663a <=( A298  and  (not A269) );
 a29664a <=( A268  and  a29663a );
 a29668a <=( (not A301)  and  (not A300) );
 a29669a <=( A299  and  a29668a );
 a29670a <=( a29669a  and  a29664a );
 a29674a <=( A199  and  (not A166) );
 a29675a <=( A167  and  a29674a );
 a29679a <=( (not A266)  and  (not A265) );
 a29680a <=( A201  and  a29679a );
 a29681a <=( a29680a  and  a29675a );
 a29685a <=( A298  and  (not A269) );
 a29686a <=( A268  and  a29685a );
 a29690a <=( A302  and  (not A300) );
 a29691a <=( A299  and  a29690a );
 a29692a <=( a29691a  and  a29686a );
 a29696a <=( A199  and  (not A166) );
 a29697a <=( A167  and  a29696a );
 a29701a <=( (not A266)  and  (not A265) );
 a29702a <=( A201  and  a29701a );
 a29703a <=( a29702a  and  a29697a );
 a29707a <=( A298  and  (not A269) );
 a29708a <=( A268  and  a29707a );
 a29712a <=( A301  and  (not A300) );
 a29713a <=( (not A299)  and  a29712a );
 a29714a <=( a29713a  and  a29708a );
 a29718a <=( A199  and  (not A166) );
 a29719a <=( A167  and  a29718a );
 a29723a <=( (not A266)  and  (not A265) );
 a29724a <=( A201  and  a29723a );
 a29725a <=( a29724a  and  a29719a );
 a29729a <=( A298  and  (not A269) );
 a29730a <=( A268  and  a29729a );
 a29734a <=( (not A302)  and  (not A300) );
 a29735a <=( (not A299)  and  a29734a );
 a29736a <=( a29735a  and  a29730a );
 a29740a <=( A199  and  (not A166) );
 a29741a <=( A167  and  a29740a );
 a29745a <=( (not A266)  and  (not A265) );
 a29746a <=( A201  and  a29745a );
 a29747a <=( a29746a  and  a29741a );
 a29751a <=( (not A298)  and  (not A269) );
 a29752a <=( A268  and  a29751a );
 a29756a <=( A301  and  (not A300) );
 a29757a <=( A299  and  a29756a );
 a29758a <=( a29757a  and  a29752a );
 a29762a <=( A199  and  (not A166) );
 a29763a <=( A167  and  a29762a );
 a29767a <=( (not A266)  and  (not A265) );
 a29768a <=( A201  and  a29767a );
 a29769a <=( a29768a  and  a29763a );
 a29773a <=( (not A298)  and  (not A269) );
 a29774a <=( A268  and  a29773a );
 a29778a <=( (not A302)  and  (not A300) );
 a29779a <=( A299  and  a29778a );
 a29780a <=( a29779a  and  a29774a );
 a29784a <=( A200  and  (not A166) );
 a29785a <=( A167  and  a29784a );
 a29789a <=( A266  and  A265 );
 a29790a <=( A201  and  a29789a );
 a29791a <=( a29790a  and  a29785a );
 a29795a <=( A298  and  (not A269) );
 a29796a <=( A268  and  a29795a );
 a29800a <=( (not A301)  and  (not A300) );
 a29801a <=( A299  and  a29800a );
 a29802a <=( a29801a  and  a29796a );
 a29806a <=( A200  and  (not A166) );
 a29807a <=( A167  and  a29806a );
 a29811a <=( A266  and  A265 );
 a29812a <=( A201  and  a29811a );
 a29813a <=( a29812a  and  a29807a );
 a29817a <=( A298  and  (not A269) );
 a29818a <=( A268  and  a29817a );
 a29822a <=( A302  and  (not A300) );
 a29823a <=( A299  and  a29822a );
 a29824a <=( a29823a  and  a29818a );
 a29828a <=( A200  and  (not A166) );
 a29829a <=( A167  and  a29828a );
 a29833a <=( A266  and  A265 );
 a29834a <=( A201  and  a29833a );
 a29835a <=( a29834a  and  a29829a );
 a29839a <=( A298  and  (not A269) );
 a29840a <=( A268  and  a29839a );
 a29844a <=( A301  and  (not A300) );
 a29845a <=( (not A299)  and  a29844a );
 a29846a <=( a29845a  and  a29840a );
 a29850a <=( A200  and  (not A166) );
 a29851a <=( A167  and  a29850a );
 a29855a <=( A266  and  A265 );
 a29856a <=( A201  and  a29855a );
 a29857a <=( a29856a  and  a29851a );
 a29861a <=( A298  and  (not A269) );
 a29862a <=( A268  and  a29861a );
 a29866a <=( (not A302)  and  (not A300) );
 a29867a <=( (not A299)  and  a29866a );
 a29868a <=( a29867a  and  a29862a );
 a29872a <=( A200  and  (not A166) );
 a29873a <=( A167  and  a29872a );
 a29877a <=( A266  and  A265 );
 a29878a <=( A201  and  a29877a );
 a29879a <=( a29878a  and  a29873a );
 a29883a <=( (not A298)  and  (not A269) );
 a29884a <=( A268  and  a29883a );
 a29888a <=( A301  and  (not A300) );
 a29889a <=( A299  and  a29888a );
 a29890a <=( a29889a  and  a29884a );
 a29894a <=( A200  and  (not A166) );
 a29895a <=( A167  and  a29894a );
 a29899a <=( A266  and  A265 );
 a29900a <=( A201  and  a29899a );
 a29901a <=( a29900a  and  a29895a );
 a29905a <=( (not A298)  and  (not A269) );
 a29906a <=( A268  and  a29905a );
 a29910a <=( (not A302)  and  (not A300) );
 a29911a <=( A299  and  a29910a );
 a29912a <=( a29911a  and  a29906a );
 a29916a <=( A200  and  (not A166) );
 a29917a <=( A167  and  a29916a );
 a29921a <=( A266  and  (not A265) );
 a29922a <=( A201  and  a29921a );
 a29923a <=( a29922a  and  a29917a );
 a29927a <=( A298  and  A269 );
 a29928a <=( (not A268)  and  a29927a );
 a29932a <=( (not A301)  and  (not A300) );
 a29933a <=( A299  and  a29932a );
 a29934a <=( a29933a  and  a29928a );
 a29938a <=( A200  and  (not A166) );
 a29939a <=( A167  and  a29938a );
 a29943a <=( A266  and  (not A265) );
 a29944a <=( A201  and  a29943a );
 a29945a <=( a29944a  and  a29939a );
 a29949a <=( A298  and  A269 );
 a29950a <=( (not A268)  and  a29949a );
 a29954a <=( A302  and  (not A300) );
 a29955a <=( A299  and  a29954a );
 a29956a <=( a29955a  and  a29950a );
 a29960a <=( A200  and  (not A166) );
 a29961a <=( A167  and  a29960a );
 a29965a <=( A266  and  (not A265) );
 a29966a <=( A201  and  a29965a );
 a29967a <=( a29966a  and  a29961a );
 a29971a <=( A298  and  A269 );
 a29972a <=( (not A268)  and  a29971a );
 a29976a <=( A301  and  (not A300) );
 a29977a <=( (not A299)  and  a29976a );
 a29978a <=( a29977a  and  a29972a );
 a29982a <=( A200  and  (not A166) );
 a29983a <=( A167  and  a29982a );
 a29987a <=( A266  and  (not A265) );
 a29988a <=( A201  and  a29987a );
 a29989a <=( a29988a  and  a29983a );
 a29993a <=( A298  and  A269 );
 a29994a <=( (not A268)  and  a29993a );
 a29998a <=( (not A302)  and  (not A300) );
 a29999a <=( (not A299)  and  a29998a );
 a30000a <=( a29999a  and  a29994a );
 a30004a <=( A200  and  (not A166) );
 a30005a <=( A167  and  a30004a );
 a30009a <=( A266  and  (not A265) );
 a30010a <=( A201  and  a30009a );
 a30011a <=( a30010a  and  a30005a );
 a30015a <=( (not A298)  and  A269 );
 a30016a <=( (not A268)  and  a30015a );
 a30020a <=( A301  and  (not A300) );
 a30021a <=( A299  and  a30020a );
 a30022a <=( a30021a  and  a30016a );
 a30026a <=( A200  and  (not A166) );
 a30027a <=( A167  and  a30026a );
 a30031a <=( A266  and  (not A265) );
 a30032a <=( A201  and  a30031a );
 a30033a <=( a30032a  and  a30027a );
 a30037a <=( (not A298)  and  A269 );
 a30038a <=( (not A268)  and  a30037a );
 a30042a <=( (not A302)  and  (not A300) );
 a30043a <=( A299  and  a30042a );
 a30044a <=( a30043a  and  a30038a );
 a30048a <=( A200  and  (not A166) );
 a30049a <=( A167  and  a30048a );
 a30053a <=( (not A266)  and  A265 );
 a30054a <=( A201  and  a30053a );
 a30055a <=( a30054a  and  a30049a );
 a30059a <=( A298  and  A269 );
 a30060a <=( (not A268)  and  a30059a );
 a30064a <=( (not A301)  and  (not A300) );
 a30065a <=( A299  and  a30064a );
 a30066a <=( a30065a  and  a30060a );
 a30070a <=( A200  and  (not A166) );
 a30071a <=( A167  and  a30070a );
 a30075a <=( (not A266)  and  A265 );
 a30076a <=( A201  and  a30075a );
 a30077a <=( a30076a  and  a30071a );
 a30081a <=( A298  and  A269 );
 a30082a <=( (not A268)  and  a30081a );
 a30086a <=( A302  and  (not A300) );
 a30087a <=( A299  and  a30086a );
 a30088a <=( a30087a  and  a30082a );
 a30092a <=( A200  and  (not A166) );
 a30093a <=( A167  and  a30092a );
 a30097a <=( (not A266)  and  A265 );
 a30098a <=( A201  and  a30097a );
 a30099a <=( a30098a  and  a30093a );
 a30103a <=( A298  and  A269 );
 a30104a <=( (not A268)  and  a30103a );
 a30108a <=( A301  and  (not A300) );
 a30109a <=( (not A299)  and  a30108a );
 a30110a <=( a30109a  and  a30104a );
 a30114a <=( A200  and  (not A166) );
 a30115a <=( A167  and  a30114a );
 a30119a <=( (not A266)  and  A265 );
 a30120a <=( A201  and  a30119a );
 a30121a <=( a30120a  and  a30115a );
 a30125a <=( A298  and  A269 );
 a30126a <=( (not A268)  and  a30125a );
 a30130a <=( (not A302)  and  (not A300) );
 a30131a <=( (not A299)  and  a30130a );
 a30132a <=( a30131a  and  a30126a );
 a30136a <=( A200  and  (not A166) );
 a30137a <=( A167  and  a30136a );
 a30141a <=( (not A266)  and  A265 );
 a30142a <=( A201  and  a30141a );
 a30143a <=( a30142a  and  a30137a );
 a30147a <=( (not A298)  and  A269 );
 a30148a <=( (not A268)  and  a30147a );
 a30152a <=( A301  and  (not A300) );
 a30153a <=( A299  and  a30152a );
 a30154a <=( a30153a  and  a30148a );
 a30158a <=( A200  and  (not A166) );
 a30159a <=( A167  and  a30158a );
 a30163a <=( (not A266)  and  A265 );
 a30164a <=( A201  and  a30163a );
 a30165a <=( a30164a  and  a30159a );
 a30169a <=( (not A298)  and  A269 );
 a30170a <=( (not A268)  and  a30169a );
 a30174a <=( (not A302)  and  (not A300) );
 a30175a <=( A299  and  a30174a );
 a30176a <=( a30175a  and  a30170a );
 a30180a <=( A200  and  (not A166) );
 a30181a <=( A167  and  a30180a );
 a30185a <=( (not A266)  and  (not A265) );
 a30186a <=( A201  and  a30185a );
 a30187a <=( a30186a  and  a30181a );
 a30191a <=( A298  and  (not A269) );
 a30192a <=( A268  and  a30191a );
 a30196a <=( (not A301)  and  (not A300) );
 a30197a <=( A299  and  a30196a );
 a30198a <=( a30197a  and  a30192a );
 a30202a <=( A200  and  (not A166) );
 a30203a <=( A167  and  a30202a );
 a30207a <=( (not A266)  and  (not A265) );
 a30208a <=( A201  and  a30207a );
 a30209a <=( a30208a  and  a30203a );
 a30213a <=( A298  and  (not A269) );
 a30214a <=( A268  and  a30213a );
 a30218a <=( A302  and  (not A300) );
 a30219a <=( A299  and  a30218a );
 a30220a <=( a30219a  and  a30214a );
 a30224a <=( A200  and  (not A166) );
 a30225a <=( A167  and  a30224a );
 a30229a <=( (not A266)  and  (not A265) );
 a30230a <=( A201  and  a30229a );
 a30231a <=( a30230a  and  a30225a );
 a30235a <=( A298  and  (not A269) );
 a30236a <=( A268  and  a30235a );
 a30240a <=( A301  and  (not A300) );
 a30241a <=( (not A299)  and  a30240a );
 a30242a <=( a30241a  and  a30236a );
 a30246a <=( A200  and  (not A166) );
 a30247a <=( A167  and  a30246a );
 a30251a <=( (not A266)  and  (not A265) );
 a30252a <=( A201  and  a30251a );
 a30253a <=( a30252a  and  a30247a );
 a30257a <=( A298  and  (not A269) );
 a30258a <=( A268  and  a30257a );
 a30262a <=( (not A302)  and  (not A300) );
 a30263a <=( (not A299)  and  a30262a );
 a30264a <=( a30263a  and  a30258a );
 a30268a <=( A200  and  (not A166) );
 a30269a <=( A167  and  a30268a );
 a30273a <=( (not A266)  and  (not A265) );
 a30274a <=( A201  and  a30273a );
 a30275a <=( a30274a  and  a30269a );
 a30279a <=( (not A298)  and  (not A269) );
 a30280a <=( A268  and  a30279a );
 a30284a <=( A301  and  (not A300) );
 a30285a <=( A299  and  a30284a );
 a30286a <=( a30285a  and  a30280a );
 a30290a <=( A200  and  (not A166) );
 a30291a <=( A167  and  a30290a );
 a30295a <=( (not A266)  and  (not A265) );
 a30296a <=( A201  and  a30295a );
 a30297a <=( a30296a  and  a30291a );
 a30301a <=( (not A298)  and  (not A269) );
 a30302a <=( A268  and  a30301a );
 a30306a <=( (not A302)  and  (not A300) );
 a30307a <=( A299  and  a30306a );
 a30308a <=( a30307a  and  a30302a );
 a30312a <=( A199  and  (not A166) );
 a30313a <=( A167  and  a30312a );
 a30317a <=( (not A203)  and  A202 );
 a30318a <=( A200  and  a30317a );
 a30319a <=( a30318a  and  a30313a );
 a30323a <=( A298  and  A267 );
 a30324a <=( A265  and  a30323a );
 a30328a <=( (not A301)  and  (not A300) );
 a30329a <=( A299  and  a30328a );
 a30330a <=( a30329a  and  a30324a );
 a30334a <=( A199  and  (not A166) );
 a30335a <=( A167  and  a30334a );
 a30339a <=( (not A203)  and  A202 );
 a30340a <=( A200  and  a30339a );
 a30341a <=( a30340a  and  a30335a );
 a30345a <=( A298  and  A267 );
 a30346a <=( A265  and  a30345a );
 a30350a <=( A302  and  (not A300) );
 a30351a <=( A299  and  a30350a );
 a30352a <=( a30351a  and  a30346a );
 a30356a <=( A199  and  (not A166) );
 a30357a <=( A167  and  a30356a );
 a30361a <=( (not A203)  and  A202 );
 a30362a <=( A200  and  a30361a );
 a30363a <=( a30362a  and  a30357a );
 a30367a <=( A298  and  A267 );
 a30368a <=( A265  and  a30367a );
 a30372a <=( A301  and  (not A300) );
 a30373a <=( (not A299)  and  a30372a );
 a30374a <=( a30373a  and  a30368a );
 a30378a <=( A199  and  (not A166) );
 a30379a <=( A167  and  a30378a );
 a30383a <=( (not A203)  and  A202 );
 a30384a <=( A200  and  a30383a );
 a30385a <=( a30384a  and  a30379a );
 a30389a <=( A298  and  A267 );
 a30390a <=( A265  and  a30389a );
 a30394a <=( (not A302)  and  (not A300) );
 a30395a <=( (not A299)  and  a30394a );
 a30396a <=( a30395a  and  a30390a );
 a30400a <=( A199  and  (not A166) );
 a30401a <=( A167  and  a30400a );
 a30405a <=( (not A203)  and  A202 );
 a30406a <=( A200  and  a30405a );
 a30407a <=( a30406a  and  a30401a );
 a30411a <=( (not A298)  and  A267 );
 a30412a <=( A265  and  a30411a );
 a30416a <=( A301  and  (not A300) );
 a30417a <=( A299  and  a30416a );
 a30418a <=( a30417a  and  a30412a );
 a30422a <=( A199  and  (not A166) );
 a30423a <=( A167  and  a30422a );
 a30427a <=( (not A203)  and  A202 );
 a30428a <=( A200  and  a30427a );
 a30429a <=( a30428a  and  a30423a );
 a30433a <=( (not A298)  and  A267 );
 a30434a <=( A265  and  a30433a );
 a30438a <=( (not A302)  and  (not A300) );
 a30439a <=( A299  and  a30438a );
 a30440a <=( a30439a  and  a30434a );
 a30444a <=( A199  and  (not A166) );
 a30445a <=( A167  and  a30444a );
 a30449a <=( (not A203)  and  A202 );
 a30450a <=( A200  and  a30449a );
 a30451a <=( a30450a  and  a30445a );
 a30455a <=( A298  and  A267 );
 a30456a <=( A266  and  a30455a );
 a30460a <=( (not A301)  and  (not A300) );
 a30461a <=( A299  and  a30460a );
 a30462a <=( a30461a  and  a30456a );
 a30466a <=( A199  and  (not A166) );
 a30467a <=( A167  and  a30466a );
 a30471a <=( (not A203)  and  A202 );
 a30472a <=( A200  and  a30471a );
 a30473a <=( a30472a  and  a30467a );
 a30477a <=( A298  and  A267 );
 a30478a <=( A266  and  a30477a );
 a30482a <=( A302  and  (not A300) );
 a30483a <=( A299  and  a30482a );
 a30484a <=( a30483a  and  a30478a );
 a30488a <=( A199  and  (not A166) );
 a30489a <=( A167  and  a30488a );
 a30493a <=( (not A203)  and  A202 );
 a30494a <=( A200  and  a30493a );
 a30495a <=( a30494a  and  a30489a );
 a30499a <=( A298  and  A267 );
 a30500a <=( A266  and  a30499a );
 a30504a <=( A301  and  (not A300) );
 a30505a <=( (not A299)  and  a30504a );
 a30506a <=( a30505a  and  a30500a );
 a30510a <=( A199  and  (not A166) );
 a30511a <=( A167  and  a30510a );
 a30515a <=( (not A203)  and  A202 );
 a30516a <=( A200  and  a30515a );
 a30517a <=( a30516a  and  a30511a );
 a30521a <=( A298  and  A267 );
 a30522a <=( A266  and  a30521a );
 a30526a <=( (not A302)  and  (not A300) );
 a30527a <=( (not A299)  and  a30526a );
 a30528a <=( a30527a  and  a30522a );
 a30532a <=( A199  and  (not A166) );
 a30533a <=( A167  and  a30532a );
 a30537a <=( (not A203)  and  A202 );
 a30538a <=( A200  and  a30537a );
 a30539a <=( a30538a  and  a30533a );
 a30543a <=( (not A298)  and  A267 );
 a30544a <=( A266  and  a30543a );
 a30548a <=( A301  and  (not A300) );
 a30549a <=( A299  and  a30548a );
 a30550a <=( a30549a  and  a30544a );
 a30554a <=( A199  and  (not A166) );
 a30555a <=( A167  and  a30554a );
 a30559a <=( (not A203)  and  A202 );
 a30560a <=( A200  and  a30559a );
 a30561a <=( a30560a  and  a30555a );
 a30565a <=( (not A298)  and  A267 );
 a30566a <=( A266  and  a30565a );
 a30570a <=( (not A302)  and  (not A300) );
 a30571a <=( A299  and  a30570a );
 a30572a <=( a30571a  and  a30566a );
 a30576a <=( A199  and  (not A166) );
 a30577a <=( A167  and  a30576a );
 a30581a <=( (not A202)  and  (not A201) );
 a30582a <=( A200  and  a30581a );
 a30583a <=( a30582a  and  a30577a );
 a30587a <=( (not A267)  and  A266 );
 a30588a <=( A265  and  a30587a );
 a30592a <=( A300  and  A299 );
 a30593a <=( (not A268)  and  a30592a );
 a30594a <=( a30593a  and  a30588a );
 a30598a <=( A199  and  (not A166) );
 a30599a <=( A167  and  a30598a );
 a30603a <=( (not A202)  and  (not A201) );
 a30604a <=( A200  and  a30603a );
 a30605a <=( a30604a  and  a30599a );
 a30609a <=( (not A267)  and  A266 );
 a30610a <=( A265  and  a30609a );
 a30614a <=( A300  and  A298 );
 a30615a <=( (not A268)  and  a30614a );
 a30616a <=( a30615a  and  a30610a );
 a30620a <=( A199  and  (not A166) );
 a30621a <=( A167  and  a30620a );
 a30625a <=( (not A202)  and  (not A201) );
 a30626a <=( A200  and  a30625a );
 a30627a <=( a30626a  and  a30621a );
 a30631a <=( (not A267)  and  A266 );
 a30632a <=( A265  and  a30631a );
 a30636a <=( A300  and  A299 );
 a30637a <=( A269  and  a30636a );
 a30638a <=( a30637a  and  a30632a );
 a30642a <=( A199  and  (not A166) );
 a30643a <=( A167  and  a30642a );
 a30647a <=( (not A202)  and  (not A201) );
 a30648a <=( A200  and  a30647a );
 a30649a <=( a30648a  and  a30643a );
 a30653a <=( (not A267)  and  A266 );
 a30654a <=( A265  and  a30653a );
 a30658a <=( A300  and  A298 );
 a30659a <=( A269  and  a30658a );
 a30660a <=( a30659a  and  a30654a );
 a30664a <=( A199  and  (not A166) );
 a30665a <=( A167  and  a30664a );
 a30669a <=( (not A202)  and  (not A201) );
 a30670a <=( A200  and  a30669a );
 a30671a <=( a30670a  and  a30665a );
 a30675a <=( (not A267)  and  A266 );
 a30676a <=( (not A265)  and  a30675a );
 a30680a <=( A300  and  A299 );
 a30681a <=( A268  and  a30680a );
 a30682a <=( a30681a  and  a30676a );
 a30686a <=( A199  and  (not A166) );
 a30687a <=( A167  and  a30686a );
 a30691a <=( (not A202)  and  (not A201) );
 a30692a <=( A200  and  a30691a );
 a30693a <=( a30692a  and  a30687a );
 a30697a <=( (not A267)  and  A266 );
 a30698a <=( (not A265)  and  a30697a );
 a30702a <=( A300  and  A298 );
 a30703a <=( A268  and  a30702a );
 a30704a <=( a30703a  and  a30698a );
 a30708a <=( A199  and  (not A166) );
 a30709a <=( A167  and  a30708a );
 a30713a <=( (not A202)  and  (not A201) );
 a30714a <=( A200  and  a30713a );
 a30715a <=( a30714a  and  a30709a );
 a30719a <=( (not A267)  and  A266 );
 a30720a <=( (not A265)  and  a30719a );
 a30724a <=( A300  and  A299 );
 a30725a <=( (not A269)  and  a30724a );
 a30726a <=( a30725a  and  a30720a );
 a30730a <=( A199  and  (not A166) );
 a30731a <=( A167  and  a30730a );
 a30735a <=( (not A202)  and  (not A201) );
 a30736a <=( A200  and  a30735a );
 a30737a <=( a30736a  and  a30731a );
 a30741a <=( (not A267)  and  A266 );
 a30742a <=( (not A265)  and  a30741a );
 a30746a <=( A300  and  A298 );
 a30747a <=( (not A269)  and  a30746a );
 a30748a <=( a30747a  and  a30742a );
 a30752a <=( A199  and  (not A166) );
 a30753a <=( A167  and  a30752a );
 a30757a <=( (not A202)  and  (not A201) );
 a30758a <=( A200  and  a30757a );
 a30759a <=( a30758a  and  a30753a );
 a30763a <=( (not A267)  and  (not A266) );
 a30764a <=( A265  and  a30763a );
 a30768a <=( A300  and  A299 );
 a30769a <=( A268  and  a30768a );
 a30770a <=( a30769a  and  a30764a );
 a30774a <=( A199  and  (not A166) );
 a30775a <=( A167  and  a30774a );
 a30779a <=( (not A202)  and  (not A201) );
 a30780a <=( A200  and  a30779a );
 a30781a <=( a30780a  and  a30775a );
 a30785a <=( (not A267)  and  (not A266) );
 a30786a <=( A265  and  a30785a );
 a30790a <=( A300  and  A298 );
 a30791a <=( A268  and  a30790a );
 a30792a <=( a30791a  and  a30786a );
 a30796a <=( A199  and  (not A166) );
 a30797a <=( A167  and  a30796a );
 a30801a <=( (not A202)  and  (not A201) );
 a30802a <=( A200  and  a30801a );
 a30803a <=( a30802a  and  a30797a );
 a30807a <=( (not A267)  and  (not A266) );
 a30808a <=( A265  and  a30807a );
 a30812a <=( A300  and  A299 );
 a30813a <=( (not A269)  and  a30812a );
 a30814a <=( a30813a  and  a30808a );
 a30818a <=( A199  and  (not A166) );
 a30819a <=( A167  and  a30818a );
 a30823a <=( (not A202)  and  (not A201) );
 a30824a <=( A200  and  a30823a );
 a30825a <=( a30824a  and  a30819a );
 a30829a <=( (not A267)  and  (not A266) );
 a30830a <=( A265  and  a30829a );
 a30834a <=( A300  and  A298 );
 a30835a <=( (not A269)  and  a30834a );
 a30836a <=( a30835a  and  a30830a );
 a30840a <=( A199  and  (not A166) );
 a30841a <=( A167  and  a30840a );
 a30845a <=( A203  and  (not A201) );
 a30846a <=( A200  and  a30845a );
 a30847a <=( a30846a  and  a30841a );
 a30851a <=( (not A267)  and  A266 );
 a30852a <=( A265  and  a30851a );
 a30856a <=( A300  and  A299 );
 a30857a <=( (not A268)  and  a30856a );
 a30858a <=( a30857a  and  a30852a );
 a30862a <=( A199  and  (not A166) );
 a30863a <=( A167  and  a30862a );
 a30867a <=( A203  and  (not A201) );
 a30868a <=( A200  and  a30867a );
 a30869a <=( a30868a  and  a30863a );
 a30873a <=( (not A267)  and  A266 );
 a30874a <=( A265  and  a30873a );
 a30878a <=( A300  and  A298 );
 a30879a <=( (not A268)  and  a30878a );
 a30880a <=( a30879a  and  a30874a );
 a30884a <=( A199  and  (not A166) );
 a30885a <=( A167  and  a30884a );
 a30889a <=( A203  and  (not A201) );
 a30890a <=( A200  and  a30889a );
 a30891a <=( a30890a  and  a30885a );
 a30895a <=( (not A267)  and  A266 );
 a30896a <=( A265  and  a30895a );
 a30900a <=( A300  and  A299 );
 a30901a <=( A269  and  a30900a );
 a30902a <=( a30901a  and  a30896a );
 a30906a <=( A199  and  (not A166) );
 a30907a <=( A167  and  a30906a );
 a30911a <=( A203  and  (not A201) );
 a30912a <=( A200  and  a30911a );
 a30913a <=( a30912a  and  a30907a );
 a30917a <=( (not A267)  and  A266 );
 a30918a <=( A265  and  a30917a );
 a30922a <=( A300  and  A298 );
 a30923a <=( A269  and  a30922a );
 a30924a <=( a30923a  and  a30918a );
 a30928a <=( A199  and  (not A166) );
 a30929a <=( A167  and  a30928a );
 a30933a <=( A203  and  (not A201) );
 a30934a <=( A200  and  a30933a );
 a30935a <=( a30934a  and  a30929a );
 a30939a <=( (not A267)  and  A266 );
 a30940a <=( (not A265)  and  a30939a );
 a30944a <=( A300  and  A299 );
 a30945a <=( A268  and  a30944a );
 a30946a <=( a30945a  and  a30940a );
 a30950a <=( A199  and  (not A166) );
 a30951a <=( A167  and  a30950a );
 a30955a <=( A203  and  (not A201) );
 a30956a <=( A200  and  a30955a );
 a30957a <=( a30956a  and  a30951a );
 a30961a <=( (not A267)  and  A266 );
 a30962a <=( (not A265)  and  a30961a );
 a30966a <=( A300  and  A298 );
 a30967a <=( A268  and  a30966a );
 a30968a <=( a30967a  and  a30962a );
 a30972a <=( A199  and  (not A166) );
 a30973a <=( A167  and  a30972a );
 a30977a <=( A203  and  (not A201) );
 a30978a <=( A200  and  a30977a );
 a30979a <=( a30978a  and  a30973a );
 a30983a <=( (not A267)  and  A266 );
 a30984a <=( (not A265)  and  a30983a );
 a30988a <=( A300  and  A299 );
 a30989a <=( (not A269)  and  a30988a );
 a30990a <=( a30989a  and  a30984a );
 a30994a <=( A199  and  (not A166) );
 a30995a <=( A167  and  a30994a );
 a30999a <=( A203  and  (not A201) );
 a31000a <=( A200  and  a30999a );
 a31001a <=( a31000a  and  a30995a );
 a31005a <=( (not A267)  and  A266 );
 a31006a <=( (not A265)  and  a31005a );
 a31010a <=( A300  and  A298 );
 a31011a <=( (not A269)  and  a31010a );
 a31012a <=( a31011a  and  a31006a );
 a31016a <=( A199  and  (not A166) );
 a31017a <=( A167  and  a31016a );
 a31021a <=( A203  and  (not A201) );
 a31022a <=( A200  and  a31021a );
 a31023a <=( a31022a  and  a31017a );
 a31027a <=( (not A267)  and  (not A266) );
 a31028a <=( A265  and  a31027a );
 a31032a <=( A300  and  A299 );
 a31033a <=( A268  and  a31032a );
 a31034a <=( a31033a  and  a31028a );
 a31038a <=( A199  and  (not A166) );
 a31039a <=( A167  and  a31038a );
 a31043a <=( A203  and  (not A201) );
 a31044a <=( A200  and  a31043a );
 a31045a <=( a31044a  and  a31039a );
 a31049a <=( (not A267)  and  (not A266) );
 a31050a <=( A265  and  a31049a );
 a31054a <=( A300  and  A298 );
 a31055a <=( A268  and  a31054a );
 a31056a <=( a31055a  and  a31050a );
 a31060a <=( A199  and  (not A166) );
 a31061a <=( A167  and  a31060a );
 a31065a <=( A203  and  (not A201) );
 a31066a <=( A200  and  a31065a );
 a31067a <=( a31066a  and  a31061a );
 a31071a <=( (not A267)  and  (not A266) );
 a31072a <=( A265  and  a31071a );
 a31076a <=( A300  and  A299 );
 a31077a <=( (not A269)  and  a31076a );
 a31078a <=( a31077a  and  a31072a );
 a31082a <=( A199  and  (not A166) );
 a31083a <=( A167  and  a31082a );
 a31087a <=( A203  and  (not A201) );
 a31088a <=( A200  and  a31087a );
 a31089a <=( a31088a  and  a31083a );
 a31093a <=( (not A267)  and  (not A266) );
 a31094a <=( A265  and  a31093a );
 a31098a <=( A300  and  A298 );
 a31099a <=( (not A269)  and  a31098a );
 a31100a <=( a31099a  and  a31094a );
 a31104a <=( (not A199)  and  (not A166) );
 a31105a <=( A167  and  a31104a );
 a31109a <=( A203  and  (not A202) );
 a31110a <=( A200  and  a31109a );
 a31111a <=( a31110a  and  a31105a );
 a31115a <=( A298  and  A267 );
 a31116a <=( A265  and  a31115a );
 a31120a <=( (not A301)  and  (not A300) );
 a31121a <=( A299  and  a31120a );
 a31122a <=( a31121a  and  a31116a );
 a31126a <=( (not A199)  and  (not A166) );
 a31127a <=( A167  and  a31126a );
 a31131a <=( A203  and  (not A202) );
 a31132a <=( A200  and  a31131a );
 a31133a <=( a31132a  and  a31127a );
 a31137a <=( A298  and  A267 );
 a31138a <=( A265  and  a31137a );
 a31142a <=( A302  and  (not A300) );
 a31143a <=( A299  and  a31142a );
 a31144a <=( a31143a  and  a31138a );
 a31148a <=( (not A199)  and  (not A166) );
 a31149a <=( A167  and  a31148a );
 a31153a <=( A203  and  (not A202) );
 a31154a <=( A200  and  a31153a );
 a31155a <=( a31154a  and  a31149a );
 a31159a <=( A298  and  A267 );
 a31160a <=( A265  and  a31159a );
 a31164a <=( A301  and  (not A300) );
 a31165a <=( (not A299)  and  a31164a );
 a31166a <=( a31165a  and  a31160a );
 a31170a <=( (not A199)  and  (not A166) );
 a31171a <=( A167  and  a31170a );
 a31175a <=( A203  and  (not A202) );
 a31176a <=( A200  and  a31175a );
 a31177a <=( a31176a  and  a31171a );
 a31181a <=( A298  and  A267 );
 a31182a <=( A265  and  a31181a );
 a31186a <=( (not A302)  and  (not A300) );
 a31187a <=( (not A299)  and  a31186a );
 a31188a <=( a31187a  and  a31182a );
 a31192a <=( (not A199)  and  (not A166) );
 a31193a <=( A167  and  a31192a );
 a31197a <=( A203  and  (not A202) );
 a31198a <=( A200  and  a31197a );
 a31199a <=( a31198a  and  a31193a );
 a31203a <=( (not A298)  and  A267 );
 a31204a <=( A265  and  a31203a );
 a31208a <=( A301  and  (not A300) );
 a31209a <=( A299  and  a31208a );
 a31210a <=( a31209a  and  a31204a );
 a31214a <=( (not A199)  and  (not A166) );
 a31215a <=( A167  and  a31214a );
 a31219a <=( A203  and  (not A202) );
 a31220a <=( A200  and  a31219a );
 a31221a <=( a31220a  and  a31215a );
 a31225a <=( (not A298)  and  A267 );
 a31226a <=( A265  and  a31225a );
 a31230a <=( (not A302)  and  (not A300) );
 a31231a <=( A299  and  a31230a );
 a31232a <=( a31231a  and  a31226a );
 a31236a <=( (not A199)  and  (not A166) );
 a31237a <=( A167  and  a31236a );
 a31241a <=( A203  and  (not A202) );
 a31242a <=( A200  and  a31241a );
 a31243a <=( a31242a  and  a31237a );
 a31247a <=( A298  and  A267 );
 a31248a <=( A266  and  a31247a );
 a31252a <=( (not A301)  and  (not A300) );
 a31253a <=( A299  and  a31252a );
 a31254a <=( a31253a  and  a31248a );
 a31258a <=( (not A199)  and  (not A166) );
 a31259a <=( A167  and  a31258a );
 a31263a <=( A203  and  (not A202) );
 a31264a <=( A200  and  a31263a );
 a31265a <=( a31264a  and  a31259a );
 a31269a <=( A298  and  A267 );
 a31270a <=( A266  and  a31269a );
 a31274a <=( A302  and  (not A300) );
 a31275a <=( A299  and  a31274a );
 a31276a <=( a31275a  and  a31270a );
 a31280a <=( (not A199)  and  (not A166) );
 a31281a <=( A167  and  a31280a );
 a31285a <=( A203  and  (not A202) );
 a31286a <=( A200  and  a31285a );
 a31287a <=( a31286a  and  a31281a );
 a31291a <=( A298  and  A267 );
 a31292a <=( A266  and  a31291a );
 a31296a <=( A301  and  (not A300) );
 a31297a <=( (not A299)  and  a31296a );
 a31298a <=( a31297a  and  a31292a );
 a31302a <=( (not A199)  and  (not A166) );
 a31303a <=( A167  and  a31302a );
 a31307a <=( A203  and  (not A202) );
 a31308a <=( A200  and  a31307a );
 a31309a <=( a31308a  and  a31303a );
 a31313a <=( A298  and  A267 );
 a31314a <=( A266  and  a31313a );
 a31318a <=( (not A302)  and  (not A300) );
 a31319a <=( (not A299)  and  a31318a );
 a31320a <=( a31319a  and  a31314a );
 a31324a <=( (not A199)  and  (not A166) );
 a31325a <=( A167  and  a31324a );
 a31329a <=( A203  and  (not A202) );
 a31330a <=( A200  and  a31329a );
 a31331a <=( a31330a  and  a31325a );
 a31335a <=( (not A298)  and  A267 );
 a31336a <=( A266  and  a31335a );
 a31340a <=( A301  and  (not A300) );
 a31341a <=( A299  and  a31340a );
 a31342a <=( a31341a  and  a31336a );
 a31346a <=( (not A199)  and  (not A166) );
 a31347a <=( A167  and  a31346a );
 a31351a <=( A203  and  (not A202) );
 a31352a <=( A200  and  a31351a );
 a31353a <=( a31352a  and  a31347a );
 a31357a <=( (not A298)  and  A267 );
 a31358a <=( A266  and  a31357a );
 a31362a <=( (not A302)  and  (not A300) );
 a31363a <=( A299  and  a31362a );
 a31364a <=( a31363a  and  a31358a );
 a31368a <=( (not A199)  and  (not A166) );
 a31369a <=( A167  and  a31368a );
 a31373a <=( A202  and  (not A201) );
 a31374a <=( A200  and  a31373a );
 a31375a <=( a31374a  and  a31369a );
 a31379a <=( (not A267)  and  A266 );
 a31380a <=( A265  and  a31379a );
 a31384a <=( A300  and  A299 );
 a31385a <=( (not A268)  and  a31384a );
 a31386a <=( a31385a  and  a31380a );
 a31390a <=( (not A199)  and  (not A166) );
 a31391a <=( A167  and  a31390a );
 a31395a <=( A202  and  (not A201) );
 a31396a <=( A200  and  a31395a );
 a31397a <=( a31396a  and  a31391a );
 a31401a <=( (not A267)  and  A266 );
 a31402a <=( A265  and  a31401a );
 a31406a <=( A300  and  A298 );
 a31407a <=( (not A268)  and  a31406a );
 a31408a <=( a31407a  and  a31402a );
 a31412a <=( (not A199)  and  (not A166) );
 a31413a <=( A167  and  a31412a );
 a31417a <=( A202  and  (not A201) );
 a31418a <=( A200  and  a31417a );
 a31419a <=( a31418a  and  a31413a );
 a31423a <=( (not A267)  and  A266 );
 a31424a <=( A265  and  a31423a );
 a31428a <=( A300  and  A299 );
 a31429a <=( A269  and  a31428a );
 a31430a <=( a31429a  and  a31424a );
 a31434a <=( (not A199)  and  (not A166) );
 a31435a <=( A167  and  a31434a );
 a31439a <=( A202  and  (not A201) );
 a31440a <=( A200  and  a31439a );
 a31441a <=( a31440a  and  a31435a );
 a31445a <=( (not A267)  and  A266 );
 a31446a <=( A265  and  a31445a );
 a31450a <=( A300  and  A298 );
 a31451a <=( A269  and  a31450a );
 a31452a <=( a31451a  and  a31446a );
 a31456a <=( (not A199)  and  (not A166) );
 a31457a <=( A167  and  a31456a );
 a31461a <=( A202  and  (not A201) );
 a31462a <=( A200  and  a31461a );
 a31463a <=( a31462a  and  a31457a );
 a31467a <=( (not A267)  and  A266 );
 a31468a <=( (not A265)  and  a31467a );
 a31472a <=( A300  and  A299 );
 a31473a <=( A268  and  a31472a );
 a31474a <=( a31473a  and  a31468a );
 a31478a <=( (not A199)  and  (not A166) );
 a31479a <=( A167  and  a31478a );
 a31483a <=( A202  and  (not A201) );
 a31484a <=( A200  and  a31483a );
 a31485a <=( a31484a  and  a31479a );
 a31489a <=( (not A267)  and  A266 );
 a31490a <=( (not A265)  and  a31489a );
 a31494a <=( A300  and  A298 );
 a31495a <=( A268  and  a31494a );
 a31496a <=( a31495a  and  a31490a );
 a31500a <=( (not A199)  and  (not A166) );
 a31501a <=( A167  and  a31500a );
 a31505a <=( A202  and  (not A201) );
 a31506a <=( A200  and  a31505a );
 a31507a <=( a31506a  and  a31501a );
 a31511a <=( (not A267)  and  A266 );
 a31512a <=( (not A265)  and  a31511a );
 a31516a <=( A300  and  A299 );
 a31517a <=( (not A269)  and  a31516a );
 a31518a <=( a31517a  and  a31512a );
 a31522a <=( (not A199)  and  (not A166) );
 a31523a <=( A167  and  a31522a );
 a31527a <=( A202  and  (not A201) );
 a31528a <=( A200  and  a31527a );
 a31529a <=( a31528a  and  a31523a );
 a31533a <=( (not A267)  and  A266 );
 a31534a <=( (not A265)  and  a31533a );
 a31538a <=( A300  and  A298 );
 a31539a <=( (not A269)  and  a31538a );
 a31540a <=( a31539a  and  a31534a );
 a31544a <=( (not A199)  and  (not A166) );
 a31545a <=( A167  and  a31544a );
 a31549a <=( A202  and  (not A201) );
 a31550a <=( A200  and  a31549a );
 a31551a <=( a31550a  and  a31545a );
 a31555a <=( (not A267)  and  (not A266) );
 a31556a <=( A265  and  a31555a );
 a31560a <=( A300  and  A299 );
 a31561a <=( A268  and  a31560a );
 a31562a <=( a31561a  and  a31556a );
 a31566a <=( (not A199)  and  (not A166) );
 a31567a <=( A167  and  a31566a );
 a31571a <=( A202  and  (not A201) );
 a31572a <=( A200  and  a31571a );
 a31573a <=( a31572a  and  a31567a );
 a31577a <=( (not A267)  and  (not A266) );
 a31578a <=( A265  and  a31577a );
 a31582a <=( A300  and  A298 );
 a31583a <=( A268  and  a31582a );
 a31584a <=( a31583a  and  a31578a );
 a31588a <=( (not A199)  and  (not A166) );
 a31589a <=( A167  and  a31588a );
 a31593a <=( A202  and  (not A201) );
 a31594a <=( A200  and  a31593a );
 a31595a <=( a31594a  and  a31589a );
 a31599a <=( (not A267)  and  (not A266) );
 a31600a <=( A265  and  a31599a );
 a31604a <=( A300  and  A299 );
 a31605a <=( (not A269)  and  a31604a );
 a31606a <=( a31605a  and  a31600a );
 a31610a <=( (not A199)  and  (not A166) );
 a31611a <=( A167  and  a31610a );
 a31615a <=( A202  and  (not A201) );
 a31616a <=( A200  and  a31615a );
 a31617a <=( a31616a  and  a31611a );
 a31621a <=( (not A267)  and  (not A266) );
 a31622a <=( A265  and  a31621a );
 a31626a <=( A300  and  A298 );
 a31627a <=( (not A269)  and  a31626a );
 a31628a <=( a31627a  and  a31622a );
 a31632a <=( (not A199)  and  (not A166) );
 a31633a <=( A167  and  a31632a );
 a31637a <=( (not A203)  and  (not A201) );
 a31638a <=( A200  and  a31637a );
 a31639a <=( a31638a  and  a31633a );
 a31643a <=( (not A267)  and  A266 );
 a31644a <=( A265  and  a31643a );
 a31648a <=( A300  and  A299 );
 a31649a <=( (not A268)  and  a31648a );
 a31650a <=( a31649a  and  a31644a );
 a31654a <=( (not A199)  and  (not A166) );
 a31655a <=( A167  and  a31654a );
 a31659a <=( (not A203)  and  (not A201) );
 a31660a <=( A200  and  a31659a );
 a31661a <=( a31660a  and  a31655a );
 a31665a <=( (not A267)  and  A266 );
 a31666a <=( A265  and  a31665a );
 a31670a <=( A300  and  A298 );
 a31671a <=( (not A268)  and  a31670a );
 a31672a <=( a31671a  and  a31666a );
 a31676a <=( (not A199)  and  (not A166) );
 a31677a <=( A167  and  a31676a );
 a31681a <=( (not A203)  and  (not A201) );
 a31682a <=( A200  and  a31681a );
 a31683a <=( a31682a  and  a31677a );
 a31687a <=( (not A267)  and  A266 );
 a31688a <=( A265  and  a31687a );
 a31692a <=( A300  and  A299 );
 a31693a <=( A269  and  a31692a );
 a31694a <=( a31693a  and  a31688a );
 a31698a <=( (not A199)  and  (not A166) );
 a31699a <=( A167  and  a31698a );
 a31703a <=( (not A203)  and  (not A201) );
 a31704a <=( A200  and  a31703a );
 a31705a <=( a31704a  and  a31699a );
 a31709a <=( (not A267)  and  A266 );
 a31710a <=( A265  and  a31709a );
 a31714a <=( A300  and  A298 );
 a31715a <=( A269  and  a31714a );
 a31716a <=( a31715a  and  a31710a );
 a31720a <=( (not A199)  and  (not A166) );
 a31721a <=( A167  and  a31720a );
 a31725a <=( (not A203)  and  (not A201) );
 a31726a <=( A200  and  a31725a );
 a31727a <=( a31726a  and  a31721a );
 a31731a <=( (not A267)  and  A266 );
 a31732a <=( (not A265)  and  a31731a );
 a31736a <=( A300  and  A299 );
 a31737a <=( A268  and  a31736a );
 a31738a <=( a31737a  and  a31732a );
 a31742a <=( (not A199)  and  (not A166) );
 a31743a <=( A167  and  a31742a );
 a31747a <=( (not A203)  and  (not A201) );
 a31748a <=( A200  and  a31747a );
 a31749a <=( a31748a  and  a31743a );
 a31753a <=( (not A267)  and  A266 );
 a31754a <=( (not A265)  and  a31753a );
 a31758a <=( A300  and  A298 );
 a31759a <=( A268  and  a31758a );
 a31760a <=( a31759a  and  a31754a );
 a31764a <=( (not A199)  and  (not A166) );
 a31765a <=( A167  and  a31764a );
 a31769a <=( (not A203)  and  (not A201) );
 a31770a <=( A200  and  a31769a );
 a31771a <=( a31770a  and  a31765a );
 a31775a <=( (not A267)  and  A266 );
 a31776a <=( (not A265)  and  a31775a );
 a31780a <=( A300  and  A299 );
 a31781a <=( (not A269)  and  a31780a );
 a31782a <=( a31781a  and  a31776a );
 a31786a <=( (not A199)  and  (not A166) );
 a31787a <=( A167  and  a31786a );
 a31791a <=( (not A203)  and  (not A201) );
 a31792a <=( A200  and  a31791a );
 a31793a <=( a31792a  and  a31787a );
 a31797a <=( (not A267)  and  A266 );
 a31798a <=( (not A265)  and  a31797a );
 a31802a <=( A300  and  A298 );
 a31803a <=( (not A269)  and  a31802a );
 a31804a <=( a31803a  and  a31798a );
 a31808a <=( (not A199)  and  (not A166) );
 a31809a <=( A167  and  a31808a );
 a31813a <=( (not A203)  and  (not A201) );
 a31814a <=( A200  and  a31813a );
 a31815a <=( a31814a  and  a31809a );
 a31819a <=( (not A267)  and  (not A266) );
 a31820a <=( A265  and  a31819a );
 a31824a <=( A300  and  A299 );
 a31825a <=( A268  and  a31824a );
 a31826a <=( a31825a  and  a31820a );
 a31830a <=( (not A199)  and  (not A166) );
 a31831a <=( A167  and  a31830a );
 a31835a <=( (not A203)  and  (not A201) );
 a31836a <=( A200  and  a31835a );
 a31837a <=( a31836a  and  a31831a );
 a31841a <=( (not A267)  and  (not A266) );
 a31842a <=( A265  and  a31841a );
 a31846a <=( A300  and  A298 );
 a31847a <=( A268  and  a31846a );
 a31848a <=( a31847a  and  a31842a );
 a31852a <=( (not A199)  and  (not A166) );
 a31853a <=( A167  and  a31852a );
 a31857a <=( (not A203)  and  (not A201) );
 a31858a <=( A200  and  a31857a );
 a31859a <=( a31858a  and  a31853a );
 a31863a <=( (not A267)  and  (not A266) );
 a31864a <=( A265  and  a31863a );
 a31868a <=( A300  and  A299 );
 a31869a <=( (not A269)  and  a31868a );
 a31870a <=( a31869a  and  a31864a );
 a31874a <=( (not A199)  and  (not A166) );
 a31875a <=( A167  and  a31874a );
 a31879a <=( (not A203)  and  (not A201) );
 a31880a <=( A200  and  a31879a );
 a31881a <=( a31880a  and  a31875a );
 a31885a <=( (not A267)  and  (not A266) );
 a31886a <=( A265  and  a31885a );
 a31890a <=( A300  and  A298 );
 a31891a <=( (not A269)  and  a31890a );
 a31892a <=( a31891a  and  a31886a );
 a31896a <=( A199  and  (not A166) );
 a31897a <=( A167  and  a31896a );
 a31901a <=( A203  and  (not A202) );
 a31902a <=( (not A200)  and  a31901a );
 a31903a <=( a31902a  and  a31897a );
 a31907a <=( A298  and  A267 );
 a31908a <=( A265  and  a31907a );
 a31912a <=( (not A301)  and  (not A300) );
 a31913a <=( A299  and  a31912a );
 a31914a <=( a31913a  and  a31908a );
 a31918a <=( A199  and  (not A166) );
 a31919a <=( A167  and  a31918a );
 a31923a <=( A203  and  (not A202) );
 a31924a <=( (not A200)  and  a31923a );
 a31925a <=( a31924a  and  a31919a );
 a31929a <=( A298  and  A267 );
 a31930a <=( A265  and  a31929a );
 a31934a <=( A302  and  (not A300) );
 a31935a <=( A299  and  a31934a );
 a31936a <=( a31935a  and  a31930a );
 a31940a <=( A199  and  (not A166) );
 a31941a <=( A167  and  a31940a );
 a31945a <=( A203  and  (not A202) );
 a31946a <=( (not A200)  and  a31945a );
 a31947a <=( a31946a  and  a31941a );
 a31951a <=( A298  and  A267 );
 a31952a <=( A265  and  a31951a );
 a31956a <=( A301  and  (not A300) );
 a31957a <=( (not A299)  and  a31956a );
 a31958a <=( a31957a  and  a31952a );
 a31962a <=( A199  and  (not A166) );
 a31963a <=( A167  and  a31962a );
 a31967a <=( A203  and  (not A202) );
 a31968a <=( (not A200)  and  a31967a );
 a31969a <=( a31968a  and  a31963a );
 a31973a <=( A298  and  A267 );
 a31974a <=( A265  and  a31973a );
 a31978a <=( (not A302)  and  (not A300) );
 a31979a <=( (not A299)  and  a31978a );
 a31980a <=( a31979a  and  a31974a );
 a31984a <=( A199  and  (not A166) );
 a31985a <=( A167  and  a31984a );
 a31989a <=( A203  and  (not A202) );
 a31990a <=( (not A200)  and  a31989a );
 a31991a <=( a31990a  and  a31985a );
 a31995a <=( (not A298)  and  A267 );
 a31996a <=( A265  and  a31995a );
 a32000a <=( A301  and  (not A300) );
 a32001a <=( A299  and  a32000a );
 a32002a <=( a32001a  and  a31996a );
 a32006a <=( A199  and  (not A166) );
 a32007a <=( A167  and  a32006a );
 a32011a <=( A203  and  (not A202) );
 a32012a <=( (not A200)  and  a32011a );
 a32013a <=( a32012a  and  a32007a );
 a32017a <=( (not A298)  and  A267 );
 a32018a <=( A265  and  a32017a );
 a32022a <=( (not A302)  and  (not A300) );
 a32023a <=( A299  and  a32022a );
 a32024a <=( a32023a  and  a32018a );
 a32028a <=( A199  and  (not A166) );
 a32029a <=( A167  and  a32028a );
 a32033a <=( A203  and  (not A202) );
 a32034a <=( (not A200)  and  a32033a );
 a32035a <=( a32034a  and  a32029a );
 a32039a <=( A298  and  A267 );
 a32040a <=( A266  and  a32039a );
 a32044a <=( (not A301)  and  (not A300) );
 a32045a <=( A299  and  a32044a );
 a32046a <=( a32045a  and  a32040a );
 a32050a <=( A199  and  (not A166) );
 a32051a <=( A167  and  a32050a );
 a32055a <=( A203  and  (not A202) );
 a32056a <=( (not A200)  and  a32055a );
 a32057a <=( a32056a  and  a32051a );
 a32061a <=( A298  and  A267 );
 a32062a <=( A266  and  a32061a );
 a32066a <=( A302  and  (not A300) );
 a32067a <=( A299  and  a32066a );
 a32068a <=( a32067a  and  a32062a );
 a32072a <=( A199  and  (not A166) );
 a32073a <=( A167  and  a32072a );
 a32077a <=( A203  and  (not A202) );
 a32078a <=( (not A200)  and  a32077a );
 a32079a <=( a32078a  and  a32073a );
 a32083a <=( A298  and  A267 );
 a32084a <=( A266  and  a32083a );
 a32088a <=( A301  and  (not A300) );
 a32089a <=( (not A299)  and  a32088a );
 a32090a <=( a32089a  and  a32084a );
 a32094a <=( A199  and  (not A166) );
 a32095a <=( A167  and  a32094a );
 a32099a <=( A203  and  (not A202) );
 a32100a <=( (not A200)  and  a32099a );
 a32101a <=( a32100a  and  a32095a );
 a32105a <=( A298  and  A267 );
 a32106a <=( A266  and  a32105a );
 a32110a <=( (not A302)  and  (not A300) );
 a32111a <=( (not A299)  and  a32110a );
 a32112a <=( a32111a  and  a32106a );
 a32116a <=( A199  and  (not A166) );
 a32117a <=( A167  and  a32116a );
 a32121a <=( A203  and  (not A202) );
 a32122a <=( (not A200)  and  a32121a );
 a32123a <=( a32122a  and  a32117a );
 a32127a <=( (not A298)  and  A267 );
 a32128a <=( A266  and  a32127a );
 a32132a <=( A301  and  (not A300) );
 a32133a <=( A299  and  a32132a );
 a32134a <=( a32133a  and  a32128a );
 a32138a <=( A199  and  (not A166) );
 a32139a <=( A167  and  a32138a );
 a32143a <=( A203  and  (not A202) );
 a32144a <=( (not A200)  and  a32143a );
 a32145a <=( a32144a  and  a32139a );
 a32149a <=( (not A298)  and  A267 );
 a32150a <=( A266  and  a32149a );
 a32154a <=( (not A302)  and  (not A300) );
 a32155a <=( A299  and  a32154a );
 a32156a <=( a32155a  and  a32150a );
 a32160a <=( A199  and  (not A166) );
 a32161a <=( A167  and  a32160a );
 a32165a <=( A202  and  (not A201) );
 a32166a <=( (not A200)  and  a32165a );
 a32167a <=( a32166a  and  a32161a );
 a32171a <=( (not A267)  and  A266 );
 a32172a <=( A265  and  a32171a );
 a32176a <=( A300  and  A299 );
 a32177a <=( (not A268)  and  a32176a );
 a32178a <=( a32177a  and  a32172a );
 a32182a <=( A199  and  (not A166) );
 a32183a <=( A167  and  a32182a );
 a32187a <=( A202  and  (not A201) );
 a32188a <=( (not A200)  and  a32187a );
 a32189a <=( a32188a  and  a32183a );
 a32193a <=( (not A267)  and  A266 );
 a32194a <=( A265  and  a32193a );
 a32198a <=( A300  and  A298 );
 a32199a <=( (not A268)  and  a32198a );
 a32200a <=( a32199a  and  a32194a );
 a32204a <=( A199  and  (not A166) );
 a32205a <=( A167  and  a32204a );
 a32209a <=( A202  and  (not A201) );
 a32210a <=( (not A200)  and  a32209a );
 a32211a <=( a32210a  and  a32205a );
 a32215a <=( (not A267)  and  A266 );
 a32216a <=( A265  and  a32215a );
 a32220a <=( A300  and  A299 );
 a32221a <=( A269  and  a32220a );
 a32222a <=( a32221a  and  a32216a );
 a32226a <=( A199  and  (not A166) );
 a32227a <=( A167  and  a32226a );
 a32231a <=( A202  and  (not A201) );
 a32232a <=( (not A200)  and  a32231a );
 a32233a <=( a32232a  and  a32227a );
 a32237a <=( (not A267)  and  A266 );
 a32238a <=( A265  and  a32237a );
 a32242a <=( A300  and  A298 );
 a32243a <=( A269  and  a32242a );
 a32244a <=( a32243a  and  a32238a );
 a32248a <=( A199  and  (not A166) );
 a32249a <=( A167  and  a32248a );
 a32253a <=( A202  and  (not A201) );
 a32254a <=( (not A200)  and  a32253a );
 a32255a <=( a32254a  and  a32249a );
 a32259a <=( (not A267)  and  A266 );
 a32260a <=( (not A265)  and  a32259a );
 a32264a <=( A300  and  A299 );
 a32265a <=( A268  and  a32264a );
 a32266a <=( a32265a  and  a32260a );
 a32270a <=( A199  and  (not A166) );
 a32271a <=( A167  and  a32270a );
 a32275a <=( A202  and  (not A201) );
 a32276a <=( (not A200)  and  a32275a );
 a32277a <=( a32276a  and  a32271a );
 a32281a <=( (not A267)  and  A266 );
 a32282a <=( (not A265)  and  a32281a );
 a32286a <=( A300  and  A298 );
 a32287a <=( A268  and  a32286a );
 a32288a <=( a32287a  and  a32282a );
 a32292a <=( A199  and  (not A166) );
 a32293a <=( A167  and  a32292a );
 a32297a <=( A202  and  (not A201) );
 a32298a <=( (not A200)  and  a32297a );
 a32299a <=( a32298a  and  a32293a );
 a32303a <=( (not A267)  and  A266 );
 a32304a <=( (not A265)  and  a32303a );
 a32308a <=( A300  and  A299 );
 a32309a <=( (not A269)  and  a32308a );
 a32310a <=( a32309a  and  a32304a );
 a32314a <=( A199  and  (not A166) );
 a32315a <=( A167  and  a32314a );
 a32319a <=( A202  and  (not A201) );
 a32320a <=( (not A200)  and  a32319a );
 a32321a <=( a32320a  and  a32315a );
 a32325a <=( (not A267)  and  A266 );
 a32326a <=( (not A265)  and  a32325a );
 a32330a <=( A300  and  A298 );
 a32331a <=( (not A269)  and  a32330a );
 a32332a <=( a32331a  and  a32326a );
 a32336a <=( A199  and  (not A166) );
 a32337a <=( A167  and  a32336a );
 a32341a <=( A202  and  (not A201) );
 a32342a <=( (not A200)  and  a32341a );
 a32343a <=( a32342a  and  a32337a );
 a32347a <=( (not A267)  and  (not A266) );
 a32348a <=( A265  and  a32347a );
 a32352a <=( A300  and  A299 );
 a32353a <=( A268  and  a32352a );
 a32354a <=( a32353a  and  a32348a );
 a32358a <=( A199  and  (not A166) );
 a32359a <=( A167  and  a32358a );
 a32363a <=( A202  and  (not A201) );
 a32364a <=( (not A200)  and  a32363a );
 a32365a <=( a32364a  and  a32359a );
 a32369a <=( (not A267)  and  (not A266) );
 a32370a <=( A265  and  a32369a );
 a32374a <=( A300  and  A298 );
 a32375a <=( A268  and  a32374a );
 a32376a <=( a32375a  and  a32370a );
 a32380a <=( A199  and  (not A166) );
 a32381a <=( A167  and  a32380a );
 a32385a <=( A202  and  (not A201) );
 a32386a <=( (not A200)  and  a32385a );
 a32387a <=( a32386a  and  a32381a );
 a32391a <=( (not A267)  and  (not A266) );
 a32392a <=( A265  and  a32391a );
 a32396a <=( A300  and  A299 );
 a32397a <=( (not A269)  and  a32396a );
 a32398a <=( a32397a  and  a32392a );
 a32402a <=( A199  and  (not A166) );
 a32403a <=( A167  and  a32402a );
 a32407a <=( A202  and  (not A201) );
 a32408a <=( (not A200)  and  a32407a );
 a32409a <=( a32408a  and  a32403a );
 a32413a <=( (not A267)  and  (not A266) );
 a32414a <=( A265  and  a32413a );
 a32418a <=( A300  and  A298 );
 a32419a <=( (not A269)  and  a32418a );
 a32420a <=( a32419a  and  a32414a );
 a32424a <=( A199  and  (not A166) );
 a32425a <=( A167  and  a32424a );
 a32429a <=( (not A203)  and  (not A201) );
 a32430a <=( (not A200)  and  a32429a );
 a32431a <=( a32430a  and  a32425a );
 a32435a <=( (not A267)  and  A266 );
 a32436a <=( A265  and  a32435a );
 a32440a <=( A300  and  A299 );
 a32441a <=( (not A268)  and  a32440a );
 a32442a <=( a32441a  and  a32436a );
 a32446a <=( A199  and  (not A166) );
 a32447a <=( A167  and  a32446a );
 a32451a <=( (not A203)  and  (not A201) );
 a32452a <=( (not A200)  and  a32451a );
 a32453a <=( a32452a  and  a32447a );
 a32457a <=( (not A267)  and  A266 );
 a32458a <=( A265  and  a32457a );
 a32462a <=( A300  and  A298 );
 a32463a <=( (not A268)  and  a32462a );
 a32464a <=( a32463a  and  a32458a );
 a32468a <=( A199  and  (not A166) );
 a32469a <=( A167  and  a32468a );
 a32473a <=( (not A203)  and  (not A201) );
 a32474a <=( (not A200)  and  a32473a );
 a32475a <=( a32474a  and  a32469a );
 a32479a <=( (not A267)  and  A266 );
 a32480a <=( A265  and  a32479a );
 a32484a <=( A300  and  A299 );
 a32485a <=( A269  and  a32484a );
 a32486a <=( a32485a  and  a32480a );
 a32490a <=( A199  and  (not A166) );
 a32491a <=( A167  and  a32490a );
 a32495a <=( (not A203)  and  (not A201) );
 a32496a <=( (not A200)  and  a32495a );
 a32497a <=( a32496a  and  a32491a );
 a32501a <=( (not A267)  and  A266 );
 a32502a <=( A265  and  a32501a );
 a32506a <=( A300  and  A298 );
 a32507a <=( A269  and  a32506a );
 a32508a <=( a32507a  and  a32502a );
 a32512a <=( A199  and  (not A166) );
 a32513a <=( A167  and  a32512a );
 a32517a <=( (not A203)  and  (not A201) );
 a32518a <=( (not A200)  and  a32517a );
 a32519a <=( a32518a  and  a32513a );
 a32523a <=( (not A267)  and  A266 );
 a32524a <=( (not A265)  and  a32523a );
 a32528a <=( A300  and  A299 );
 a32529a <=( A268  and  a32528a );
 a32530a <=( a32529a  and  a32524a );
 a32534a <=( A199  and  (not A166) );
 a32535a <=( A167  and  a32534a );
 a32539a <=( (not A203)  and  (not A201) );
 a32540a <=( (not A200)  and  a32539a );
 a32541a <=( a32540a  and  a32535a );
 a32545a <=( (not A267)  and  A266 );
 a32546a <=( (not A265)  and  a32545a );
 a32550a <=( A300  and  A298 );
 a32551a <=( A268  and  a32550a );
 a32552a <=( a32551a  and  a32546a );
 a32556a <=( A199  and  (not A166) );
 a32557a <=( A167  and  a32556a );
 a32561a <=( (not A203)  and  (not A201) );
 a32562a <=( (not A200)  and  a32561a );
 a32563a <=( a32562a  and  a32557a );
 a32567a <=( (not A267)  and  A266 );
 a32568a <=( (not A265)  and  a32567a );
 a32572a <=( A300  and  A299 );
 a32573a <=( (not A269)  and  a32572a );
 a32574a <=( a32573a  and  a32568a );
 a32578a <=( A199  and  (not A166) );
 a32579a <=( A167  and  a32578a );
 a32583a <=( (not A203)  and  (not A201) );
 a32584a <=( (not A200)  and  a32583a );
 a32585a <=( a32584a  and  a32579a );
 a32589a <=( (not A267)  and  A266 );
 a32590a <=( (not A265)  and  a32589a );
 a32594a <=( A300  and  A298 );
 a32595a <=( (not A269)  and  a32594a );
 a32596a <=( a32595a  and  a32590a );
 a32600a <=( A199  and  (not A166) );
 a32601a <=( A167  and  a32600a );
 a32605a <=( (not A203)  and  (not A201) );
 a32606a <=( (not A200)  and  a32605a );
 a32607a <=( a32606a  and  a32601a );
 a32611a <=( (not A267)  and  (not A266) );
 a32612a <=( A265  and  a32611a );
 a32616a <=( A300  and  A299 );
 a32617a <=( A268  and  a32616a );
 a32618a <=( a32617a  and  a32612a );
 a32622a <=( A199  and  (not A166) );
 a32623a <=( A167  and  a32622a );
 a32627a <=( (not A203)  and  (not A201) );
 a32628a <=( (not A200)  and  a32627a );
 a32629a <=( a32628a  and  a32623a );
 a32633a <=( (not A267)  and  (not A266) );
 a32634a <=( A265  and  a32633a );
 a32638a <=( A300  and  A298 );
 a32639a <=( A268  and  a32638a );
 a32640a <=( a32639a  and  a32634a );
 a32644a <=( A199  and  (not A166) );
 a32645a <=( A167  and  a32644a );
 a32649a <=( (not A203)  and  (not A201) );
 a32650a <=( (not A200)  and  a32649a );
 a32651a <=( a32650a  and  a32645a );
 a32655a <=( (not A267)  and  (not A266) );
 a32656a <=( A265  and  a32655a );
 a32660a <=( A300  and  A299 );
 a32661a <=( (not A269)  and  a32660a );
 a32662a <=( a32661a  and  a32656a );
 a32666a <=( A199  and  (not A166) );
 a32667a <=( A167  and  a32666a );
 a32671a <=( (not A203)  and  (not A201) );
 a32672a <=( (not A200)  and  a32671a );
 a32673a <=( a32672a  and  a32667a );
 a32677a <=( (not A267)  and  (not A266) );
 a32678a <=( A265  and  a32677a );
 a32682a <=( A300  and  A298 );
 a32683a <=( (not A269)  and  a32682a );
 a32684a <=( a32683a  and  a32678a );
 a32688a <=( (not A199)  and  (not A166) );
 a32689a <=( A167  and  a32688a );
 a32693a <=( (not A265)  and  (not A202) );
 a32694a <=( (not A200)  and  a32693a );
 a32695a <=( a32694a  and  a32689a );
 a32699a <=( A298  and  (not A268) );
 a32700a <=( (not A266)  and  a32699a );
 a32704a <=( (not A302)  and  A301 );
 a32705a <=( A299  and  a32704a );
 a32706a <=( a32705a  and  a32700a );
 a32710a <=( (not A199)  and  (not A166) );
 a32711a <=( A167  and  a32710a );
 a32715a <=( (not A265)  and  (not A202) );
 a32716a <=( (not A200)  and  a32715a );
 a32717a <=( a32716a  and  a32711a );
 a32721a <=( A298  and  (not A268) );
 a32722a <=( (not A266)  and  a32721a );
 a32726a <=( A302  and  (not A301) );
 a32727a <=( (not A299)  and  a32726a );
 a32728a <=( a32727a  and  a32722a );
 a32732a <=( (not A199)  and  (not A166) );
 a32733a <=( A167  and  a32732a );
 a32737a <=( (not A265)  and  (not A202) );
 a32738a <=( (not A200)  and  a32737a );
 a32739a <=( a32738a  and  a32733a );
 a32743a <=( (not A298)  and  (not A268) );
 a32744a <=( (not A266)  and  a32743a );
 a32748a <=( A302  and  (not A301) );
 a32749a <=( A299  and  a32748a );
 a32750a <=( a32749a  and  a32744a );
 a32754a <=( (not A199)  and  (not A166) );
 a32755a <=( A167  and  a32754a );
 a32759a <=( (not A265)  and  (not A202) );
 a32760a <=( (not A200)  and  a32759a );
 a32761a <=( a32760a  and  a32755a );
 a32765a <=( (not A298)  and  (not A268) );
 a32766a <=( (not A266)  and  a32765a );
 a32770a <=( (not A302)  and  A301 );
 a32771a <=( (not A299)  and  a32770a );
 a32772a <=( a32771a  and  a32766a );
 a32776a <=( (not A199)  and  (not A166) );
 a32777a <=( A167  and  a32776a );
 a32781a <=( (not A265)  and  (not A202) );
 a32782a <=( (not A200)  and  a32781a );
 a32783a <=( a32782a  and  a32777a );
 a32787a <=( A298  and  A269 );
 a32788a <=( (not A266)  and  a32787a );
 a32792a <=( (not A302)  and  A301 );
 a32793a <=( A299  and  a32792a );
 a32794a <=( a32793a  and  a32788a );
 a32798a <=( (not A199)  and  (not A166) );
 a32799a <=( A167  and  a32798a );
 a32803a <=( (not A265)  and  (not A202) );
 a32804a <=( (not A200)  and  a32803a );
 a32805a <=( a32804a  and  a32799a );
 a32809a <=( A298  and  A269 );
 a32810a <=( (not A266)  and  a32809a );
 a32814a <=( A302  and  (not A301) );
 a32815a <=( (not A299)  and  a32814a );
 a32816a <=( a32815a  and  a32810a );
 a32820a <=( (not A199)  and  (not A166) );
 a32821a <=( A167  and  a32820a );
 a32825a <=( (not A265)  and  (not A202) );
 a32826a <=( (not A200)  and  a32825a );
 a32827a <=( a32826a  and  a32821a );
 a32831a <=( (not A298)  and  A269 );
 a32832a <=( (not A266)  and  a32831a );
 a32836a <=( A302  and  (not A301) );
 a32837a <=( A299  and  a32836a );
 a32838a <=( a32837a  and  a32832a );
 a32842a <=( (not A199)  and  (not A166) );
 a32843a <=( A167  and  a32842a );
 a32847a <=( (not A265)  and  (not A202) );
 a32848a <=( (not A200)  and  a32847a );
 a32849a <=( a32848a  and  a32843a );
 a32853a <=( (not A298)  and  A269 );
 a32854a <=( (not A266)  and  a32853a );
 a32858a <=( (not A302)  and  A301 );
 a32859a <=( (not A299)  and  a32858a );
 a32860a <=( a32859a  and  a32854a );
 a32864a <=( (not A199)  and  (not A166) );
 a32865a <=( A167  and  a32864a );
 a32869a <=( (not A265)  and  A203 );
 a32870a <=( (not A200)  and  a32869a );
 a32871a <=( a32870a  and  a32865a );
 a32875a <=( A298  and  (not A268) );
 a32876a <=( (not A266)  and  a32875a );
 a32880a <=( (not A302)  and  A301 );
 a32881a <=( A299  and  a32880a );
 a32882a <=( a32881a  and  a32876a );
 a32886a <=( (not A199)  and  (not A166) );
 a32887a <=( A167  and  a32886a );
 a32891a <=( (not A265)  and  A203 );
 a32892a <=( (not A200)  and  a32891a );
 a32893a <=( a32892a  and  a32887a );
 a32897a <=( A298  and  (not A268) );
 a32898a <=( (not A266)  and  a32897a );
 a32902a <=( A302  and  (not A301) );
 a32903a <=( (not A299)  and  a32902a );
 a32904a <=( a32903a  and  a32898a );
 a32908a <=( (not A199)  and  (not A166) );
 a32909a <=( A167  and  a32908a );
 a32913a <=( (not A265)  and  A203 );
 a32914a <=( (not A200)  and  a32913a );
 a32915a <=( a32914a  and  a32909a );
 a32919a <=( (not A298)  and  (not A268) );
 a32920a <=( (not A266)  and  a32919a );
 a32924a <=( A302  and  (not A301) );
 a32925a <=( A299  and  a32924a );
 a32926a <=( a32925a  and  a32920a );
 a32930a <=( (not A199)  and  (not A166) );
 a32931a <=( A167  and  a32930a );
 a32935a <=( (not A265)  and  A203 );
 a32936a <=( (not A200)  and  a32935a );
 a32937a <=( a32936a  and  a32931a );
 a32941a <=( (not A298)  and  (not A268) );
 a32942a <=( (not A266)  and  a32941a );
 a32946a <=( (not A302)  and  A301 );
 a32947a <=( (not A299)  and  a32946a );
 a32948a <=( a32947a  and  a32942a );
 a32952a <=( (not A199)  and  (not A166) );
 a32953a <=( A167  and  a32952a );
 a32957a <=( (not A265)  and  A203 );
 a32958a <=( (not A200)  and  a32957a );
 a32959a <=( a32958a  and  a32953a );
 a32963a <=( A298  and  A269 );
 a32964a <=( (not A266)  and  a32963a );
 a32968a <=( (not A302)  and  A301 );
 a32969a <=( A299  and  a32968a );
 a32970a <=( a32969a  and  a32964a );
 a32974a <=( (not A199)  and  (not A166) );
 a32975a <=( A167  and  a32974a );
 a32979a <=( (not A265)  and  A203 );
 a32980a <=( (not A200)  and  a32979a );
 a32981a <=( a32980a  and  a32975a );
 a32985a <=( A298  and  A269 );
 a32986a <=( (not A266)  and  a32985a );
 a32990a <=( A302  and  (not A301) );
 a32991a <=( (not A299)  and  a32990a );
 a32992a <=( a32991a  and  a32986a );
 a32996a <=( (not A199)  and  (not A166) );
 a32997a <=( A167  and  a32996a );
 a33001a <=( (not A265)  and  A203 );
 a33002a <=( (not A200)  and  a33001a );
 a33003a <=( a33002a  and  a32997a );
 a33007a <=( (not A298)  and  A269 );
 a33008a <=( (not A266)  and  a33007a );
 a33012a <=( A302  and  (not A301) );
 a33013a <=( A299  and  a33012a );
 a33014a <=( a33013a  and  a33008a );
 a33018a <=( (not A199)  and  (not A166) );
 a33019a <=( A167  and  a33018a );
 a33023a <=( (not A265)  and  A203 );
 a33024a <=( (not A200)  and  a33023a );
 a33025a <=( a33024a  and  a33019a );
 a33029a <=( (not A298)  and  A269 );
 a33030a <=( (not A266)  and  a33029a );
 a33034a <=( (not A302)  and  A301 );
 a33035a <=( (not A299)  and  a33034a );
 a33036a <=( a33035a  and  a33030a );
 a33040a <=( (not A199)  and  (not A166) );
 a33041a <=( A167  and  a33040a );
 a33045a <=( (not A203)  and  A202 );
 a33046a <=( (not A200)  and  a33045a );
 a33047a <=( a33046a  and  a33041a );
 a33051a <=( A298  and  A267 );
 a33052a <=( A265  and  a33051a );
 a33056a <=( (not A301)  and  (not A300) );
 a33057a <=( A299  and  a33056a );
 a33058a <=( a33057a  and  a33052a );
 a33062a <=( (not A199)  and  (not A166) );
 a33063a <=( A167  and  a33062a );
 a33067a <=( (not A203)  and  A202 );
 a33068a <=( (not A200)  and  a33067a );
 a33069a <=( a33068a  and  a33063a );
 a33073a <=( A298  and  A267 );
 a33074a <=( A265  and  a33073a );
 a33078a <=( A302  and  (not A300) );
 a33079a <=( A299  and  a33078a );
 a33080a <=( a33079a  and  a33074a );
 a33084a <=( (not A199)  and  (not A166) );
 a33085a <=( A167  and  a33084a );
 a33089a <=( (not A203)  and  A202 );
 a33090a <=( (not A200)  and  a33089a );
 a33091a <=( a33090a  and  a33085a );
 a33095a <=( A298  and  A267 );
 a33096a <=( A265  and  a33095a );
 a33100a <=( A301  and  (not A300) );
 a33101a <=( (not A299)  and  a33100a );
 a33102a <=( a33101a  and  a33096a );
 a33106a <=( (not A199)  and  (not A166) );
 a33107a <=( A167  and  a33106a );
 a33111a <=( (not A203)  and  A202 );
 a33112a <=( (not A200)  and  a33111a );
 a33113a <=( a33112a  and  a33107a );
 a33117a <=( A298  and  A267 );
 a33118a <=( A265  and  a33117a );
 a33122a <=( (not A302)  and  (not A300) );
 a33123a <=( (not A299)  and  a33122a );
 a33124a <=( a33123a  and  a33118a );
 a33128a <=( (not A199)  and  (not A166) );
 a33129a <=( A167  and  a33128a );
 a33133a <=( (not A203)  and  A202 );
 a33134a <=( (not A200)  and  a33133a );
 a33135a <=( a33134a  and  a33129a );
 a33139a <=( (not A298)  and  A267 );
 a33140a <=( A265  and  a33139a );
 a33144a <=( A301  and  (not A300) );
 a33145a <=( A299  and  a33144a );
 a33146a <=( a33145a  and  a33140a );
 a33150a <=( (not A199)  and  (not A166) );
 a33151a <=( A167  and  a33150a );
 a33155a <=( (not A203)  and  A202 );
 a33156a <=( (not A200)  and  a33155a );
 a33157a <=( a33156a  and  a33151a );
 a33161a <=( (not A298)  and  A267 );
 a33162a <=( A265  and  a33161a );
 a33166a <=( (not A302)  and  (not A300) );
 a33167a <=( A299  and  a33166a );
 a33168a <=( a33167a  and  a33162a );
 a33172a <=( (not A199)  and  (not A166) );
 a33173a <=( A167  and  a33172a );
 a33177a <=( (not A203)  and  A202 );
 a33178a <=( (not A200)  and  a33177a );
 a33179a <=( a33178a  and  a33173a );
 a33183a <=( A298  and  A267 );
 a33184a <=( A266  and  a33183a );
 a33188a <=( (not A301)  and  (not A300) );
 a33189a <=( A299  and  a33188a );
 a33190a <=( a33189a  and  a33184a );
 a33194a <=( (not A199)  and  (not A166) );
 a33195a <=( A167  and  a33194a );
 a33199a <=( (not A203)  and  A202 );
 a33200a <=( (not A200)  and  a33199a );
 a33201a <=( a33200a  and  a33195a );
 a33205a <=( A298  and  A267 );
 a33206a <=( A266  and  a33205a );
 a33210a <=( A302  and  (not A300) );
 a33211a <=( A299  and  a33210a );
 a33212a <=( a33211a  and  a33206a );
 a33216a <=( (not A199)  and  (not A166) );
 a33217a <=( A167  and  a33216a );
 a33221a <=( (not A203)  and  A202 );
 a33222a <=( (not A200)  and  a33221a );
 a33223a <=( a33222a  and  a33217a );
 a33227a <=( A298  and  A267 );
 a33228a <=( A266  and  a33227a );
 a33232a <=( A301  and  (not A300) );
 a33233a <=( (not A299)  and  a33232a );
 a33234a <=( a33233a  and  a33228a );
 a33238a <=( (not A199)  and  (not A166) );
 a33239a <=( A167  and  a33238a );
 a33243a <=( (not A203)  and  A202 );
 a33244a <=( (not A200)  and  a33243a );
 a33245a <=( a33244a  and  a33239a );
 a33249a <=( A298  and  A267 );
 a33250a <=( A266  and  a33249a );
 a33254a <=( (not A302)  and  (not A300) );
 a33255a <=( (not A299)  and  a33254a );
 a33256a <=( a33255a  and  a33250a );
 a33260a <=( (not A199)  and  (not A166) );
 a33261a <=( A167  and  a33260a );
 a33265a <=( (not A203)  and  A202 );
 a33266a <=( (not A200)  and  a33265a );
 a33267a <=( a33266a  and  a33261a );
 a33271a <=( (not A298)  and  A267 );
 a33272a <=( A266  and  a33271a );
 a33276a <=( A301  and  (not A300) );
 a33277a <=( A299  and  a33276a );
 a33278a <=( a33277a  and  a33272a );
 a33282a <=( (not A199)  and  (not A166) );
 a33283a <=( A167  and  a33282a );
 a33287a <=( (not A203)  and  A202 );
 a33288a <=( (not A200)  and  a33287a );
 a33289a <=( a33288a  and  a33283a );
 a33293a <=( (not A298)  and  A267 );
 a33294a <=( A266  and  a33293a );
 a33298a <=( (not A302)  and  (not A300) );
 a33299a <=( A299  and  a33298a );
 a33300a <=( a33299a  and  a33294a );
 a33304a <=( A199  and  (not A166) );
 a33305a <=( (not A167)  and  a33304a );
 a33309a <=( A266  and  A265 );
 a33310a <=( A201  and  a33309a );
 a33311a <=( a33310a  and  a33305a );
 a33315a <=( A298  and  (not A268) );
 a33316a <=( (not A267)  and  a33315a );
 a33320a <=( (not A302)  and  A301 );
 a33321a <=( A299  and  a33320a );
 a33322a <=( a33321a  and  a33316a );
 a33326a <=( A199  and  (not A166) );
 a33327a <=( (not A167)  and  a33326a );
 a33331a <=( A266  and  A265 );
 a33332a <=( A201  and  a33331a );
 a33333a <=( a33332a  and  a33327a );
 a33337a <=( A298  and  (not A268) );
 a33338a <=( (not A267)  and  a33337a );
 a33342a <=( A302  and  (not A301) );
 a33343a <=( (not A299)  and  a33342a );
 a33344a <=( a33343a  and  a33338a );
 a33348a <=( A199  and  (not A166) );
 a33349a <=( (not A167)  and  a33348a );
 a33353a <=( A266  and  A265 );
 a33354a <=( A201  and  a33353a );
 a33355a <=( a33354a  and  a33349a );
 a33359a <=( (not A298)  and  (not A268) );
 a33360a <=( (not A267)  and  a33359a );
 a33364a <=( A302  and  (not A301) );
 a33365a <=( A299  and  a33364a );
 a33366a <=( a33365a  and  a33360a );
 a33370a <=( A199  and  (not A166) );
 a33371a <=( (not A167)  and  a33370a );
 a33375a <=( A266  and  A265 );
 a33376a <=( A201  and  a33375a );
 a33377a <=( a33376a  and  a33371a );
 a33381a <=( (not A298)  and  (not A268) );
 a33382a <=( (not A267)  and  a33381a );
 a33386a <=( (not A302)  and  A301 );
 a33387a <=( (not A299)  and  a33386a );
 a33388a <=( a33387a  and  a33382a );
 a33392a <=( A199  and  (not A166) );
 a33393a <=( (not A167)  and  a33392a );
 a33397a <=( A266  and  A265 );
 a33398a <=( A201  and  a33397a );
 a33399a <=( a33398a  and  a33393a );
 a33403a <=( A298  and  A269 );
 a33404a <=( (not A267)  and  a33403a );
 a33408a <=( (not A302)  and  A301 );
 a33409a <=( A299  and  a33408a );
 a33410a <=( a33409a  and  a33404a );
 a33414a <=( A199  and  (not A166) );
 a33415a <=( (not A167)  and  a33414a );
 a33419a <=( A266  and  A265 );
 a33420a <=( A201  and  a33419a );
 a33421a <=( a33420a  and  a33415a );
 a33425a <=( A298  and  A269 );
 a33426a <=( (not A267)  and  a33425a );
 a33430a <=( A302  and  (not A301) );
 a33431a <=( (not A299)  and  a33430a );
 a33432a <=( a33431a  and  a33426a );
 a33436a <=( A199  and  (not A166) );
 a33437a <=( (not A167)  and  a33436a );
 a33441a <=( A266  and  A265 );
 a33442a <=( A201  and  a33441a );
 a33443a <=( a33442a  and  a33437a );
 a33447a <=( (not A298)  and  A269 );
 a33448a <=( (not A267)  and  a33447a );
 a33452a <=( A302  and  (not A301) );
 a33453a <=( A299  and  a33452a );
 a33454a <=( a33453a  and  a33448a );
 a33458a <=( A199  and  (not A166) );
 a33459a <=( (not A167)  and  a33458a );
 a33463a <=( A266  and  A265 );
 a33464a <=( A201  and  a33463a );
 a33465a <=( a33464a  and  a33459a );
 a33469a <=( (not A298)  and  A269 );
 a33470a <=( (not A267)  and  a33469a );
 a33474a <=( (not A302)  and  A301 );
 a33475a <=( (not A299)  and  a33474a );
 a33476a <=( a33475a  and  a33470a );
 a33480a <=( A199  and  (not A166) );
 a33481a <=( (not A167)  and  a33480a );
 a33485a <=( A266  and  (not A265) );
 a33486a <=( A201  and  a33485a );
 a33487a <=( a33486a  and  a33481a );
 a33491a <=( A298  and  A268 );
 a33492a <=( (not A267)  and  a33491a );
 a33496a <=( (not A302)  and  A301 );
 a33497a <=( A299  and  a33496a );
 a33498a <=( a33497a  and  a33492a );
 a33502a <=( A199  and  (not A166) );
 a33503a <=( (not A167)  and  a33502a );
 a33507a <=( A266  and  (not A265) );
 a33508a <=( A201  and  a33507a );
 a33509a <=( a33508a  and  a33503a );
 a33513a <=( A298  and  A268 );
 a33514a <=( (not A267)  and  a33513a );
 a33518a <=( A302  and  (not A301) );
 a33519a <=( (not A299)  and  a33518a );
 a33520a <=( a33519a  and  a33514a );
 a33524a <=( A199  and  (not A166) );
 a33525a <=( (not A167)  and  a33524a );
 a33529a <=( A266  and  (not A265) );
 a33530a <=( A201  and  a33529a );
 a33531a <=( a33530a  and  a33525a );
 a33535a <=( (not A298)  and  A268 );
 a33536a <=( (not A267)  and  a33535a );
 a33540a <=( A302  and  (not A301) );
 a33541a <=( A299  and  a33540a );
 a33542a <=( a33541a  and  a33536a );
 a33546a <=( A199  and  (not A166) );
 a33547a <=( (not A167)  and  a33546a );
 a33551a <=( A266  and  (not A265) );
 a33552a <=( A201  and  a33551a );
 a33553a <=( a33552a  and  a33547a );
 a33557a <=( (not A298)  and  A268 );
 a33558a <=( (not A267)  and  a33557a );
 a33562a <=( (not A302)  and  A301 );
 a33563a <=( (not A299)  and  a33562a );
 a33564a <=( a33563a  and  a33558a );
 a33568a <=( A199  and  (not A166) );
 a33569a <=( (not A167)  and  a33568a );
 a33573a <=( A266  and  (not A265) );
 a33574a <=( A201  and  a33573a );
 a33575a <=( a33574a  and  a33569a );
 a33579a <=( A298  and  (not A269) );
 a33580a <=( (not A267)  and  a33579a );
 a33584a <=( (not A302)  and  A301 );
 a33585a <=( A299  and  a33584a );
 a33586a <=( a33585a  and  a33580a );
 a33590a <=( A199  and  (not A166) );
 a33591a <=( (not A167)  and  a33590a );
 a33595a <=( A266  and  (not A265) );
 a33596a <=( A201  and  a33595a );
 a33597a <=( a33596a  and  a33591a );
 a33601a <=( A298  and  (not A269) );
 a33602a <=( (not A267)  and  a33601a );
 a33606a <=( A302  and  (not A301) );
 a33607a <=( (not A299)  and  a33606a );
 a33608a <=( a33607a  and  a33602a );
 a33612a <=( A199  and  (not A166) );
 a33613a <=( (not A167)  and  a33612a );
 a33617a <=( A266  and  (not A265) );
 a33618a <=( A201  and  a33617a );
 a33619a <=( a33618a  and  a33613a );
 a33623a <=( (not A298)  and  (not A269) );
 a33624a <=( (not A267)  and  a33623a );
 a33628a <=( A302  and  (not A301) );
 a33629a <=( A299  and  a33628a );
 a33630a <=( a33629a  and  a33624a );
 a33634a <=( A199  and  (not A166) );
 a33635a <=( (not A167)  and  a33634a );
 a33639a <=( A266  and  (not A265) );
 a33640a <=( A201  and  a33639a );
 a33641a <=( a33640a  and  a33635a );
 a33645a <=( (not A298)  and  (not A269) );
 a33646a <=( (not A267)  and  a33645a );
 a33650a <=( (not A302)  and  A301 );
 a33651a <=( (not A299)  and  a33650a );
 a33652a <=( a33651a  and  a33646a );
 a33656a <=( A199  and  (not A166) );
 a33657a <=( (not A167)  and  a33656a );
 a33661a <=( (not A266)  and  A265 );
 a33662a <=( A201  and  a33661a );
 a33663a <=( a33662a  and  a33657a );
 a33667a <=( A298  and  A268 );
 a33668a <=( (not A267)  and  a33667a );
 a33672a <=( (not A302)  and  A301 );
 a33673a <=( A299  and  a33672a );
 a33674a <=( a33673a  and  a33668a );
 a33678a <=( A199  and  (not A166) );
 a33679a <=( (not A167)  and  a33678a );
 a33683a <=( (not A266)  and  A265 );
 a33684a <=( A201  and  a33683a );
 a33685a <=( a33684a  and  a33679a );
 a33689a <=( A298  and  A268 );
 a33690a <=( (not A267)  and  a33689a );
 a33694a <=( A302  and  (not A301) );
 a33695a <=( (not A299)  and  a33694a );
 a33696a <=( a33695a  and  a33690a );
 a33700a <=( A199  and  (not A166) );
 a33701a <=( (not A167)  and  a33700a );
 a33705a <=( (not A266)  and  A265 );
 a33706a <=( A201  and  a33705a );
 a33707a <=( a33706a  and  a33701a );
 a33711a <=( (not A298)  and  A268 );
 a33712a <=( (not A267)  and  a33711a );
 a33716a <=( A302  and  (not A301) );
 a33717a <=( A299  and  a33716a );
 a33718a <=( a33717a  and  a33712a );
 a33722a <=( A199  and  (not A166) );
 a33723a <=( (not A167)  and  a33722a );
 a33727a <=( (not A266)  and  A265 );
 a33728a <=( A201  and  a33727a );
 a33729a <=( a33728a  and  a33723a );
 a33733a <=( (not A298)  and  A268 );
 a33734a <=( (not A267)  and  a33733a );
 a33738a <=( (not A302)  and  A301 );
 a33739a <=( (not A299)  and  a33738a );
 a33740a <=( a33739a  and  a33734a );
 a33744a <=( A199  and  (not A166) );
 a33745a <=( (not A167)  and  a33744a );
 a33749a <=( (not A266)  and  A265 );
 a33750a <=( A201  and  a33749a );
 a33751a <=( a33750a  and  a33745a );
 a33755a <=( A298  and  (not A269) );
 a33756a <=( (not A267)  and  a33755a );
 a33760a <=( (not A302)  and  A301 );
 a33761a <=( A299  and  a33760a );
 a33762a <=( a33761a  and  a33756a );
 a33766a <=( A199  and  (not A166) );
 a33767a <=( (not A167)  and  a33766a );
 a33771a <=( (not A266)  and  A265 );
 a33772a <=( A201  and  a33771a );
 a33773a <=( a33772a  and  a33767a );
 a33777a <=( A298  and  (not A269) );
 a33778a <=( (not A267)  and  a33777a );
 a33782a <=( A302  and  (not A301) );
 a33783a <=( (not A299)  and  a33782a );
 a33784a <=( a33783a  and  a33778a );
 a33788a <=( A199  and  (not A166) );
 a33789a <=( (not A167)  and  a33788a );
 a33793a <=( (not A266)  and  A265 );
 a33794a <=( A201  and  a33793a );
 a33795a <=( a33794a  and  a33789a );
 a33799a <=( (not A298)  and  (not A269) );
 a33800a <=( (not A267)  and  a33799a );
 a33804a <=( A302  and  (not A301) );
 a33805a <=( A299  and  a33804a );
 a33806a <=( a33805a  and  a33800a );
 a33810a <=( A199  and  (not A166) );
 a33811a <=( (not A167)  and  a33810a );
 a33815a <=( (not A266)  and  A265 );
 a33816a <=( A201  and  a33815a );
 a33817a <=( a33816a  and  a33811a );
 a33821a <=( (not A298)  and  (not A269) );
 a33822a <=( (not A267)  and  a33821a );
 a33826a <=( (not A302)  and  A301 );
 a33827a <=( (not A299)  and  a33826a );
 a33828a <=( a33827a  and  a33822a );
 a33832a <=( A200  and  (not A166) );
 a33833a <=( (not A167)  and  a33832a );
 a33837a <=( A266  and  A265 );
 a33838a <=( A201  and  a33837a );
 a33839a <=( a33838a  and  a33833a );
 a33843a <=( A298  and  (not A268) );
 a33844a <=( (not A267)  and  a33843a );
 a33848a <=( (not A302)  and  A301 );
 a33849a <=( A299  and  a33848a );
 a33850a <=( a33849a  and  a33844a );
 a33854a <=( A200  and  (not A166) );
 a33855a <=( (not A167)  and  a33854a );
 a33859a <=( A266  and  A265 );
 a33860a <=( A201  and  a33859a );
 a33861a <=( a33860a  and  a33855a );
 a33865a <=( A298  and  (not A268) );
 a33866a <=( (not A267)  and  a33865a );
 a33870a <=( A302  and  (not A301) );
 a33871a <=( (not A299)  and  a33870a );
 a33872a <=( a33871a  and  a33866a );
 a33876a <=( A200  and  (not A166) );
 a33877a <=( (not A167)  and  a33876a );
 a33881a <=( A266  and  A265 );
 a33882a <=( A201  and  a33881a );
 a33883a <=( a33882a  and  a33877a );
 a33887a <=( (not A298)  and  (not A268) );
 a33888a <=( (not A267)  and  a33887a );
 a33892a <=( A302  and  (not A301) );
 a33893a <=( A299  and  a33892a );
 a33894a <=( a33893a  and  a33888a );
 a33898a <=( A200  and  (not A166) );
 a33899a <=( (not A167)  and  a33898a );
 a33903a <=( A266  and  A265 );
 a33904a <=( A201  and  a33903a );
 a33905a <=( a33904a  and  a33899a );
 a33909a <=( (not A298)  and  (not A268) );
 a33910a <=( (not A267)  and  a33909a );
 a33914a <=( (not A302)  and  A301 );
 a33915a <=( (not A299)  and  a33914a );
 a33916a <=( a33915a  and  a33910a );
 a33920a <=( A200  and  (not A166) );
 a33921a <=( (not A167)  and  a33920a );
 a33925a <=( A266  and  A265 );
 a33926a <=( A201  and  a33925a );
 a33927a <=( a33926a  and  a33921a );
 a33931a <=( A298  and  A269 );
 a33932a <=( (not A267)  and  a33931a );
 a33936a <=( (not A302)  and  A301 );
 a33937a <=( A299  and  a33936a );
 a33938a <=( a33937a  and  a33932a );
 a33942a <=( A200  and  (not A166) );
 a33943a <=( (not A167)  and  a33942a );
 a33947a <=( A266  and  A265 );
 a33948a <=( A201  and  a33947a );
 a33949a <=( a33948a  and  a33943a );
 a33953a <=( A298  and  A269 );
 a33954a <=( (not A267)  and  a33953a );
 a33958a <=( A302  and  (not A301) );
 a33959a <=( (not A299)  and  a33958a );
 a33960a <=( a33959a  and  a33954a );
 a33964a <=( A200  and  (not A166) );
 a33965a <=( (not A167)  and  a33964a );
 a33969a <=( A266  and  A265 );
 a33970a <=( A201  and  a33969a );
 a33971a <=( a33970a  and  a33965a );
 a33975a <=( (not A298)  and  A269 );
 a33976a <=( (not A267)  and  a33975a );
 a33980a <=( A302  and  (not A301) );
 a33981a <=( A299  and  a33980a );
 a33982a <=( a33981a  and  a33976a );
 a33986a <=( A200  and  (not A166) );
 a33987a <=( (not A167)  and  a33986a );
 a33991a <=( A266  and  A265 );
 a33992a <=( A201  and  a33991a );
 a33993a <=( a33992a  and  a33987a );
 a33997a <=( (not A298)  and  A269 );
 a33998a <=( (not A267)  and  a33997a );
 a34002a <=( (not A302)  and  A301 );
 a34003a <=( (not A299)  and  a34002a );
 a34004a <=( a34003a  and  a33998a );
 a34008a <=( A200  and  (not A166) );
 a34009a <=( (not A167)  and  a34008a );
 a34013a <=( A266  and  (not A265) );
 a34014a <=( A201  and  a34013a );
 a34015a <=( a34014a  and  a34009a );
 a34019a <=( A298  and  A268 );
 a34020a <=( (not A267)  and  a34019a );
 a34024a <=( (not A302)  and  A301 );
 a34025a <=( A299  and  a34024a );
 a34026a <=( a34025a  and  a34020a );
 a34030a <=( A200  and  (not A166) );
 a34031a <=( (not A167)  and  a34030a );
 a34035a <=( A266  and  (not A265) );
 a34036a <=( A201  and  a34035a );
 a34037a <=( a34036a  and  a34031a );
 a34041a <=( A298  and  A268 );
 a34042a <=( (not A267)  and  a34041a );
 a34046a <=( A302  and  (not A301) );
 a34047a <=( (not A299)  and  a34046a );
 a34048a <=( a34047a  and  a34042a );
 a34052a <=( A200  and  (not A166) );
 a34053a <=( (not A167)  and  a34052a );
 a34057a <=( A266  and  (not A265) );
 a34058a <=( A201  and  a34057a );
 a34059a <=( a34058a  and  a34053a );
 a34063a <=( (not A298)  and  A268 );
 a34064a <=( (not A267)  and  a34063a );
 a34068a <=( A302  and  (not A301) );
 a34069a <=( A299  and  a34068a );
 a34070a <=( a34069a  and  a34064a );
 a34074a <=( A200  and  (not A166) );
 a34075a <=( (not A167)  and  a34074a );
 a34079a <=( A266  and  (not A265) );
 a34080a <=( A201  and  a34079a );
 a34081a <=( a34080a  and  a34075a );
 a34085a <=( (not A298)  and  A268 );
 a34086a <=( (not A267)  and  a34085a );
 a34090a <=( (not A302)  and  A301 );
 a34091a <=( (not A299)  and  a34090a );
 a34092a <=( a34091a  and  a34086a );
 a34096a <=( A200  and  (not A166) );
 a34097a <=( (not A167)  and  a34096a );
 a34101a <=( A266  and  (not A265) );
 a34102a <=( A201  and  a34101a );
 a34103a <=( a34102a  and  a34097a );
 a34107a <=( A298  and  (not A269) );
 a34108a <=( (not A267)  and  a34107a );
 a34112a <=( (not A302)  and  A301 );
 a34113a <=( A299  and  a34112a );
 a34114a <=( a34113a  and  a34108a );
 a34118a <=( A200  and  (not A166) );
 a34119a <=( (not A167)  and  a34118a );
 a34123a <=( A266  and  (not A265) );
 a34124a <=( A201  and  a34123a );
 a34125a <=( a34124a  and  a34119a );
 a34129a <=( A298  and  (not A269) );
 a34130a <=( (not A267)  and  a34129a );
 a34134a <=( A302  and  (not A301) );
 a34135a <=( (not A299)  and  a34134a );
 a34136a <=( a34135a  and  a34130a );
 a34140a <=( A200  and  (not A166) );
 a34141a <=( (not A167)  and  a34140a );
 a34145a <=( A266  and  (not A265) );
 a34146a <=( A201  and  a34145a );
 a34147a <=( a34146a  and  a34141a );
 a34151a <=( (not A298)  and  (not A269) );
 a34152a <=( (not A267)  and  a34151a );
 a34156a <=( A302  and  (not A301) );
 a34157a <=( A299  and  a34156a );
 a34158a <=( a34157a  and  a34152a );
 a34162a <=( A200  and  (not A166) );
 a34163a <=( (not A167)  and  a34162a );
 a34167a <=( A266  and  (not A265) );
 a34168a <=( A201  and  a34167a );
 a34169a <=( a34168a  and  a34163a );
 a34173a <=( (not A298)  and  (not A269) );
 a34174a <=( (not A267)  and  a34173a );
 a34178a <=( (not A302)  and  A301 );
 a34179a <=( (not A299)  and  a34178a );
 a34180a <=( a34179a  and  a34174a );
 a34184a <=( A200  and  (not A166) );
 a34185a <=( (not A167)  and  a34184a );
 a34189a <=( (not A266)  and  A265 );
 a34190a <=( A201  and  a34189a );
 a34191a <=( a34190a  and  a34185a );
 a34195a <=( A298  and  A268 );
 a34196a <=( (not A267)  and  a34195a );
 a34200a <=( (not A302)  and  A301 );
 a34201a <=( A299  and  a34200a );
 a34202a <=( a34201a  and  a34196a );
 a34206a <=( A200  and  (not A166) );
 a34207a <=( (not A167)  and  a34206a );
 a34211a <=( (not A266)  and  A265 );
 a34212a <=( A201  and  a34211a );
 a34213a <=( a34212a  and  a34207a );
 a34217a <=( A298  and  A268 );
 a34218a <=( (not A267)  and  a34217a );
 a34222a <=( A302  and  (not A301) );
 a34223a <=( (not A299)  and  a34222a );
 a34224a <=( a34223a  and  a34218a );
 a34228a <=( A200  and  (not A166) );
 a34229a <=( (not A167)  and  a34228a );
 a34233a <=( (not A266)  and  A265 );
 a34234a <=( A201  and  a34233a );
 a34235a <=( a34234a  and  a34229a );
 a34239a <=( (not A298)  and  A268 );
 a34240a <=( (not A267)  and  a34239a );
 a34244a <=( A302  and  (not A301) );
 a34245a <=( A299  and  a34244a );
 a34246a <=( a34245a  and  a34240a );
 a34250a <=( A200  and  (not A166) );
 a34251a <=( (not A167)  and  a34250a );
 a34255a <=( (not A266)  and  A265 );
 a34256a <=( A201  and  a34255a );
 a34257a <=( a34256a  and  a34251a );
 a34261a <=( (not A298)  and  A268 );
 a34262a <=( (not A267)  and  a34261a );
 a34266a <=( (not A302)  and  A301 );
 a34267a <=( (not A299)  and  a34266a );
 a34268a <=( a34267a  and  a34262a );
 a34272a <=( A200  and  (not A166) );
 a34273a <=( (not A167)  and  a34272a );
 a34277a <=( (not A266)  and  A265 );
 a34278a <=( A201  and  a34277a );
 a34279a <=( a34278a  and  a34273a );
 a34283a <=( A298  and  (not A269) );
 a34284a <=( (not A267)  and  a34283a );
 a34288a <=( (not A302)  and  A301 );
 a34289a <=( A299  and  a34288a );
 a34290a <=( a34289a  and  a34284a );
 a34294a <=( A200  and  (not A166) );
 a34295a <=( (not A167)  and  a34294a );
 a34299a <=( (not A266)  and  A265 );
 a34300a <=( A201  and  a34299a );
 a34301a <=( a34300a  and  a34295a );
 a34305a <=( A298  and  (not A269) );
 a34306a <=( (not A267)  and  a34305a );
 a34310a <=( A302  and  (not A301) );
 a34311a <=( (not A299)  and  a34310a );
 a34312a <=( a34311a  and  a34306a );
 a34316a <=( A200  and  (not A166) );
 a34317a <=( (not A167)  and  a34316a );
 a34321a <=( (not A266)  and  A265 );
 a34322a <=( A201  and  a34321a );
 a34323a <=( a34322a  and  a34317a );
 a34327a <=( (not A298)  and  (not A269) );
 a34328a <=( (not A267)  and  a34327a );
 a34332a <=( A302  and  (not A301) );
 a34333a <=( A299  and  a34332a );
 a34334a <=( a34333a  and  a34328a );
 a34338a <=( A200  and  (not A166) );
 a34339a <=( (not A167)  and  a34338a );
 a34343a <=( (not A266)  and  A265 );
 a34344a <=( A201  and  a34343a );
 a34345a <=( a34344a  and  a34339a );
 a34349a <=( (not A298)  and  (not A269) );
 a34350a <=( (not A267)  and  a34349a );
 a34354a <=( (not A302)  and  A301 );
 a34355a <=( (not A299)  and  a34354a );
 a34356a <=( a34355a  and  a34350a );
 a34360a <=( A199  and  (not A166) );
 a34361a <=( (not A167)  and  a34360a );
 a34365a <=( (not A203)  and  A202 );
 a34366a <=( A200  and  a34365a );
 a34367a <=( a34366a  and  a34361a );
 a34371a <=( (not A267)  and  A266 );
 a34372a <=( A265  and  a34371a );
 a34376a <=( A300  and  A299 );
 a34377a <=( (not A268)  and  a34376a );
 a34378a <=( a34377a  and  a34372a );
 a34382a <=( A199  and  (not A166) );
 a34383a <=( (not A167)  and  a34382a );
 a34387a <=( (not A203)  and  A202 );
 a34388a <=( A200  and  a34387a );
 a34389a <=( a34388a  and  a34383a );
 a34393a <=( (not A267)  and  A266 );
 a34394a <=( A265  and  a34393a );
 a34398a <=( A300  and  A298 );
 a34399a <=( (not A268)  and  a34398a );
 a34400a <=( a34399a  and  a34394a );
 a34404a <=( A199  and  (not A166) );
 a34405a <=( (not A167)  and  a34404a );
 a34409a <=( (not A203)  and  A202 );
 a34410a <=( A200  and  a34409a );
 a34411a <=( a34410a  and  a34405a );
 a34415a <=( (not A267)  and  A266 );
 a34416a <=( A265  and  a34415a );
 a34420a <=( A300  and  A299 );
 a34421a <=( A269  and  a34420a );
 a34422a <=( a34421a  and  a34416a );
 a34426a <=( A199  and  (not A166) );
 a34427a <=( (not A167)  and  a34426a );
 a34431a <=( (not A203)  and  A202 );
 a34432a <=( A200  and  a34431a );
 a34433a <=( a34432a  and  a34427a );
 a34437a <=( (not A267)  and  A266 );
 a34438a <=( A265  and  a34437a );
 a34442a <=( A300  and  A298 );
 a34443a <=( A269  and  a34442a );
 a34444a <=( a34443a  and  a34438a );
 a34448a <=( A199  and  (not A166) );
 a34449a <=( (not A167)  and  a34448a );
 a34453a <=( (not A203)  and  A202 );
 a34454a <=( A200  and  a34453a );
 a34455a <=( a34454a  and  a34449a );
 a34459a <=( (not A267)  and  A266 );
 a34460a <=( (not A265)  and  a34459a );
 a34464a <=( A300  and  A299 );
 a34465a <=( A268  and  a34464a );
 a34466a <=( a34465a  and  a34460a );
 a34470a <=( A199  and  (not A166) );
 a34471a <=( (not A167)  and  a34470a );
 a34475a <=( (not A203)  and  A202 );
 a34476a <=( A200  and  a34475a );
 a34477a <=( a34476a  and  a34471a );
 a34481a <=( (not A267)  and  A266 );
 a34482a <=( (not A265)  and  a34481a );
 a34486a <=( A300  and  A298 );
 a34487a <=( A268  and  a34486a );
 a34488a <=( a34487a  and  a34482a );
 a34492a <=( A199  and  (not A166) );
 a34493a <=( (not A167)  and  a34492a );
 a34497a <=( (not A203)  and  A202 );
 a34498a <=( A200  and  a34497a );
 a34499a <=( a34498a  and  a34493a );
 a34503a <=( (not A267)  and  A266 );
 a34504a <=( (not A265)  and  a34503a );
 a34508a <=( A300  and  A299 );
 a34509a <=( (not A269)  and  a34508a );
 a34510a <=( a34509a  and  a34504a );
 a34514a <=( A199  and  (not A166) );
 a34515a <=( (not A167)  and  a34514a );
 a34519a <=( (not A203)  and  A202 );
 a34520a <=( A200  and  a34519a );
 a34521a <=( a34520a  and  a34515a );
 a34525a <=( (not A267)  and  A266 );
 a34526a <=( (not A265)  and  a34525a );
 a34530a <=( A300  and  A298 );
 a34531a <=( (not A269)  and  a34530a );
 a34532a <=( a34531a  and  a34526a );
 a34536a <=( A199  and  (not A166) );
 a34537a <=( (not A167)  and  a34536a );
 a34541a <=( (not A203)  and  A202 );
 a34542a <=( A200  and  a34541a );
 a34543a <=( a34542a  and  a34537a );
 a34547a <=( (not A267)  and  (not A266) );
 a34548a <=( A265  and  a34547a );
 a34552a <=( A300  and  A299 );
 a34553a <=( A268  and  a34552a );
 a34554a <=( a34553a  and  a34548a );
 a34558a <=( A199  and  (not A166) );
 a34559a <=( (not A167)  and  a34558a );
 a34563a <=( (not A203)  and  A202 );
 a34564a <=( A200  and  a34563a );
 a34565a <=( a34564a  and  a34559a );
 a34569a <=( (not A267)  and  (not A266) );
 a34570a <=( A265  and  a34569a );
 a34574a <=( A300  and  A298 );
 a34575a <=( A268  and  a34574a );
 a34576a <=( a34575a  and  a34570a );
 a34580a <=( A199  and  (not A166) );
 a34581a <=( (not A167)  and  a34580a );
 a34585a <=( (not A203)  and  A202 );
 a34586a <=( A200  and  a34585a );
 a34587a <=( a34586a  and  a34581a );
 a34591a <=( (not A267)  and  (not A266) );
 a34592a <=( A265  and  a34591a );
 a34596a <=( A300  and  A299 );
 a34597a <=( (not A269)  and  a34596a );
 a34598a <=( a34597a  and  a34592a );
 a34602a <=( A199  and  (not A166) );
 a34603a <=( (not A167)  and  a34602a );
 a34607a <=( (not A203)  and  A202 );
 a34608a <=( A200  and  a34607a );
 a34609a <=( a34608a  and  a34603a );
 a34613a <=( (not A267)  and  (not A266) );
 a34614a <=( A265  and  a34613a );
 a34618a <=( A300  and  A298 );
 a34619a <=( (not A269)  and  a34618a );
 a34620a <=( a34619a  and  a34614a );
 a34624a <=( A199  and  (not A166) );
 a34625a <=( (not A167)  and  a34624a );
 a34629a <=( (not A202)  and  (not A201) );
 a34630a <=( A200  and  a34629a );
 a34631a <=( a34630a  and  a34625a );
 a34635a <=( A298  and  A267 );
 a34636a <=( A265  and  a34635a );
 a34640a <=( (not A301)  and  (not A300) );
 a34641a <=( A299  and  a34640a );
 a34642a <=( a34641a  and  a34636a );
 a34646a <=( A199  and  (not A166) );
 a34647a <=( (not A167)  and  a34646a );
 a34651a <=( (not A202)  and  (not A201) );
 a34652a <=( A200  and  a34651a );
 a34653a <=( a34652a  and  a34647a );
 a34657a <=( A298  and  A267 );
 a34658a <=( A265  and  a34657a );
 a34662a <=( A302  and  (not A300) );
 a34663a <=( A299  and  a34662a );
 a34664a <=( a34663a  and  a34658a );
 a34668a <=( A199  and  (not A166) );
 a34669a <=( (not A167)  and  a34668a );
 a34673a <=( (not A202)  and  (not A201) );
 a34674a <=( A200  and  a34673a );
 a34675a <=( a34674a  and  a34669a );
 a34679a <=( A298  and  A267 );
 a34680a <=( A265  and  a34679a );
 a34684a <=( A301  and  (not A300) );
 a34685a <=( (not A299)  and  a34684a );
 a34686a <=( a34685a  and  a34680a );
 a34690a <=( A199  and  (not A166) );
 a34691a <=( (not A167)  and  a34690a );
 a34695a <=( (not A202)  and  (not A201) );
 a34696a <=( A200  and  a34695a );
 a34697a <=( a34696a  and  a34691a );
 a34701a <=( A298  and  A267 );
 a34702a <=( A265  and  a34701a );
 a34706a <=( (not A302)  and  (not A300) );
 a34707a <=( (not A299)  and  a34706a );
 a34708a <=( a34707a  and  a34702a );
 a34712a <=( A199  and  (not A166) );
 a34713a <=( (not A167)  and  a34712a );
 a34717a <=( (not A202)  and  (not A201) );
 a34718a <=( A200  and  a34717a );
 a34719a <=( a34718a  and  a34713a );
 a34723a <=( (not A298)  and  A267 );
 a34724a <=( A265  and  a34723a );
 a34728a <=( A301  and  (not A300) );
 a34729a <=( A299  and  a34728a );
 a34730a <=( a34729a  and  a34724a );
 a34734a <=( A199  and  (not A166) );
 a34735a <=( (not A167)  and  a34734a );
 a34739a <=( (not A202)  and  (not A201) );
 a34740a <=( A200  and  a34739a );
 a34741a <=( a34740a  and  a34735a );
 a34745a <=( (not A298)  and  A267 );
 a34746a <=( A265  and  a34745a );
 a34750a <=( (not A302)  and  (not A300) );
 a34751a <=( A299  and  a34750a );
 a34752a <=( a34751a  and  a34746a );
 a34756a <=( A199  and  (not A166) );
 a34757a <=( (not A167)  and  a34756a );
 a34761a <=( (not A202)  and  (not A201) );
 a34762a <=( A200  and  a34761a );
 a34763a <=( a34762a  and  a34757a );
 a34767a <=( A298  and  A267 );
 a34768a <=( A266  and  a34767a );
 a34772a <=( (not A301)  and  (not A300) );
 a34773a <=( A299  and  a34772a );
 a34774a <=( a34773a  and  a34768a );
 a34778a <=( A199  and  (not A166) );
 a34779a <=( (not A167)  and  a34778a );
 a34783a <=( (not A202)  and  (not A201) );
 a34784a <=( A200  and  a34783a );
 a34785a <=( a34784a  and  a34779a );
 a34789a <=( A298  and  A267 );
 a34790a <=( A266  and  a34789a );
 a34794a <=( A302  and  (not A300) );
 a34795a <=( A299  and  a34794a );
 a34796a <=( a34795a  and  a34790a );
 a34800a <=( A199  and  (not A166) );
 a34801a <=( (not A167)  and  a34800a );
 a34805a <=( (not A202)  and  (not A201) );
 a34806a <=( A200  and  a34805a );
 a34807a <=( a34806a  and  a34801a );
 a34811a <=( A298  and  A267 );
 a34812a <=( A266  and  a34811a );
 a34816a <=( A301  and  (not A300) );
 a34817a <=( (not A299)  and  a34816a );
 a34818a <=( a34817a  and  a34812a );
 a34822a <=( A199  and  (not A166) );
 a34823a <=( (not A167)  and  a34822a );
 a34827a <=( (not A202)  and  (not A201) );
 a34828a <=( A200  and  a34827a );
 a34829a <=( a34828a  and  a34823a );
 a34833a <=( A298  and  A267 );
 a34834a <=( A266  and  a34833a );
 a34838a <=( (not A302)  and  (not A300) );
 a34839a <=( (not A299)  and  a34838a );
 a34840a <=( a34839a  and  a34834a );
 a34844a <=( A199  and  (not A166) );
 a34845a <=( (not A167)  and  a34844a );
 a34849a <=( (not A202)  and  (not A201) );
 a34850a <=( A200  and  a34849a );
 a34851a <=( a34850a  and  a34845a );
 a34855a <=( (not A298)  and  A267 );
 a34856a <=( A266  and  a34855a );
 a34860a <=( A301  and  (not A300) );
 a34861a <=( A299  and  a34860a );
 a34862a <=( a34861a  and  a34856a );
 a34866a <=( A199  and  (not A166) );
 a34867a <=( (not A167)  and  a34866a );
 a34871a <=( (not A202)  and  (not A201) );
 a34872a <=( A200  and  a34871a );
 a34873a <=( a34872a  and  a34867a );
 a34877a <=( (not A298)  and  A267 );
 a34878a <=( A266  and  a34877a );
 a34882a <=( (not A302)  and  (not A300) );
 a34883a <=( A299  and  a34882a );
 a34884a <=( a34883a  and  a34878a );
 a34888a <=( A199  and  (not A166) );
 a34889a <=( (not A167)  and  a34888a );
 a34893a <=( A203  and  (not A201) );
 a34894a <=( A200  and  a34893a );
 a34895a <=( a34894a  and  a34889a );
 a34899a <=( A298  and  A267 );
 a34900a <=( A265  and  a34899a );
 a34904a <=( (not A301)  and  (not A300) );
 a34905a <=( A299  and  a34904a );
 a34906a <=( a34905a  and  a34900a );
 a34910a <=( A199  and  (not A166) );
 a34911a <=( (not A167)  and  a34910a );
 a34915a <=( A203  and  (not A201) );
 a34916a <=( A200  and  a34915a );
 a34917a <=( a34916a  and  a34911a );
 a34921a <=( A298  and  A267 );
 a34922a <=( A265  and  a34921a );
 a34926a <=( A302  and  (not A300) );
 a34927a <=( A299  and  a34926a );
 a34928a <=( a34927a  and  a34922a );
 a34932a <=( A199  and  (not A166) );
 a34933a <=( (not A167)  and  a34932a );
 a34937a <=( A203  and  (not A201) );
 a34938a <=( A200  and  a34937a );
 a34939a <=( a34938a  and  a34933a );
 a34943a <=( A298  and  A267 );
 a34944a <=( A265  and  a34943a );
 a34948a <=( A301  and  (not A300) );
 a34949a <=( (not A299)  and  a34948a );
 a34950a <=( a34949a  and  a34944a );
 a34954a <=( A199  and  (not A166) );
 a34955a <=( (not A167)  and  a34954a );
 a34959a <=( A203  and  (not A201) );
 a34960a <=( A200  and  a34959a );
 a34961a <=( a34960a  and  a34955a );
 a34965a <=( A298  and  A267 );
 a34966a <=( A265  and  a34965a );
 a34970a <=( (not A302)  and  (not A300) );
 a34971a <=( (not A299)  and  a34970a );
 a34972a <=( a34971a  and  a34966a );
 a34976a <=( A199  and  (not A166) );
 a34977a <=( (not A167)  and  a34976a );
 a34981a <=( A203  and  (not A201) );
 a34982a <=( A200  and  a34981a );
 a34983a <=( a34982a  and  a34977a );
 a34987a <=( (not A298)  and  A267 );
 a34988a <=( A265  and  a34987a );
 a34992a <=( A301  and  (not A300) );
 a34993a <=( A299  and  a34992a );
 a34994a <=( a34993a  and  a34988a );
 a34998a <=( A199  and  (not A166) );
 a34999a <=( (not A167)  and  a34998a );
 a35003a <=( A203  and  (not A201) );
 a35004a <=( A200  and  a35003a );
 a35005a <=( a35004a  and  a34999a );
 a35009a <=( (not A298)  and  A267 );
 a35010a <=( A265  and  a35009a );
 a35014a <=( (not A302)  and  (not A300) );
 a35015a <=( A299  and  a35014a );
 a35016a <=( a35015a  and  a35010a );
 a35020a <=( A199  and  (not A166) );
 a35021a <=( (not A167)  and  a35020a );
 a35025a <=( A203  and  (not A201) );
 a35026a <=( A200  and  a35025a );
 a35027a <=( a35026a  and  a35021a );
 a35031a <=( A298  and  A267 );
 a35032a <=( A266  and  a35031a );
 a35036a <=( (not A301)  and  (not A300) );
 a35037a <=( A299  and  a35036a );
 a35038a <=( a35037a  and  a35032a );
 a35042a <=( A199  and  (not A166) );
 a35043a <=( (not A167)  and  a35042a );
 a35047a <=( A203  and  (not A201) );
 a35048a <=( A200  and  a35047a );
 a35049a <=( a35048a  and  a35043a );
 a35053a <=( A298  and  A267 );
 a35054a <=( A266  and  a35053a );
 a35058a <=( A302  and  (not A300) );
 a35059a <=( A299  and  a35058a );
 a35060a <=( a35059a  and  a35054a );
 a35064a <=( A199  and  (not A166) );
 a35065a <=( (not A167)  and  a35064a );
 a35069a <=( A203  and  (not A201) );
 a35070a <=( A200  and  a35069a );
 a35071a <=( a35070a  and  a35065a );
 a35075a <=( A298  and  A267 );
 a35076a <=( A266  and  a35075a );
 a35080a <=( A301  and  (not A300) );
 a35081a <=( (not A299)  and  a35080a );
 a35082a <=( a35081a  and  a35076a );
 a35086a <=( A199  and  (not A166) );
 a35087a <=( (not A167)  and  a35086a );
 a35091a <=( A203  and  (not A201) );
 a35092a <=( A200  and  a35091a );
 a35093a <=( a35092a  and  a35087a );
 a35097a <=( A298  and  A267 );
 a35098a <=( A266  and  a35097a );
 a35102a <=( (not A302)  and  (not A300) );
 a35103a <=( (not A299)  and  a35102a );
 a35104a <=( a35103a  and  a35098a );
 a35108a <=( A199  and  (not A166) );
 a35109a <=( (not A167)  and  a35108a );
 a35113a <=( A203  and  (not A201) );
 a35114a <=( A200  and  a35113a );
 a35115a <=( a35114a  and  a35109a );
 a35119a <=( (not A298)  and  A267 );
 a35120a <=( A266  and  a35119a );
 a35124a <=( A301  and  (not A300) );
 a35125a <=( A299  and  a35124a );
 a35126a <=( a35125a  and  a35120a );
 a35130a <=( A199  and  (not A166) );
 a35131a <=( (not A167)  and  a35130a );
 a35135a <=( A203  and  (not A201) );
 a35136a <=( A200  and  a35135a );
 a35137a <=( a35136a  and  a35131a );
 a35141a <=( (not A298)  and  A267 );
 a35142a <=( A266  and  a35141a );
 a35146a <=( (not A302)  and  (not A300) );
 a35147a <=( A299  and  a35146a );
 a35148a <=( a35147a  and  a35142a );
 a35152a <=( (not A199)  and  (not A166) );
 a35153a <=( (not A167)  and  a35152a );
 a35157a <=( A203  and  (not A202) );
 a35158a <=( A200  and  a35157a );
 a35159a <=( a35158a  and  a35153a );
 a35163a <=( (not A267)  and  A266 );
 a35164a <=( A265  and  a35163a );
 a35168a <=( A300  and  A299 );
 a35169a <=( (not A268)  and  a35168a );
 a35170a <=( a35169a  and  a35164a );
 a35174a <=( (not A199)  and  (not A166) );
 a35175a <=( (not A167)  and  a35174a );
 a35179a <=( A203  and  (not A202) );
 a35180a <=( A200  and  a35179a );
 a35181a <=( a35180a  and  a35175a );
 a35185a <=( (not A267)  and  A266 );
 a35186a <=( A265  and  a35185a );
 a35190a <=( A300  and  A298 );
 a35191a <=( (not A268)  and  a35190a );
 a35192a <=( a35191a  and  a35186a );
 a35196a <=( (not A199)  and  (not A166) );
 a35197a <=( (not A167)  and  a35196a );
 a35201a <=( A203  and  (not A202) );
 a35202a <=( A200  and  a35201a );
 a35203a <=( a35202a  and  a35197a );
 a35207a <=( (not A267)  and  A266 );
 a35208a <=( A265  and  a35207a );
 a35212a <=( A300  and  A299 );
 a35213a <=( A269  and  a35212a );
 a35214a <=( a35213a  and  a35208a );
 a35218a <=( (not A199)  and  (not A166) );
 a35219a <=( (not A167)  and  a35218a );
 a35223a <=( A203  and  (not A202) );
 a35224a <=( A200  and  a35223a );
 a35225a <=( a35224a  and  a35219a );
 a35229a <=( (not A267)  and  A266 );
 a35230a <=( A265  and  a35229a );
 a35234a <=( A300  and  A298 );
 a35235a <=( A269  and  a35234a );
 a35236a <=( a35235a  and  a35230a );
 a35240a <=( (not A199)  and  (not A166) );
 a35241a <=( (not A167)  and  a35240a );
 a35245a <=( A203  and  (not A202) );
 a35246a <=( A200  and  a35245a );
 a35247a <=( a35246a  and  a35241a );
 a35251a <=( (not A267)  and  A266 );
 a35252a <=( (not A265)  and  a35251a );
 a35256a <=( A300  and  A299 );
 a35257a <=( A268  and  a35256a );
 a35258a <=( a35257a  and  a35252a );
 a35262a <=( (not A199)  and  (not A166) );
 a35263a <=( (not A167)  and  a35262a );
 a35267a <=( A203  and  (not A202) );
 a35268a <=( A200  and  a35267a );
 a35269a <=( a35268a  and  a35263a );
 a35273a <=( (not A267)  and  A266 );
 a35274a <=( (not A265)  and  a35273a );
 a35278a <=( A300  and  A298 );
 a35279a <=( A268  and  a35278a );
 a35280a <=( a35279a  and  a35274a );
 a35284a <=( (not A199)  and  (not A166) );
 a35285a <=( (not A167)  and  a35284a );
 a35289a <=( A203  and  (not A202) );
 a35290a <=( A200  and  a35289a );
 a35291a <=( a35290a  and  a35285a );
 a35295a <=( (not A267)  and  A266 );
 a35296a <=( (not A265)  and  a35295a );
 a35300a <=( A300  and  A299 );
 a35301a <=( (not A269)  and  a35300a );
 a35302a <=( a35301a  and  a35296a );
 a35306a <=( (not A199)  and  (not A166) );
 a35307a <=( (not A167)  and  a35306a );
 a35311a <=( A203  and  (not A202) );
 a35312a <=( A200  and  a35311a );
 a35313a <=( a35312a  and  a35307a );
 a35317a <=( (not A267)  and  A266 );
 a35318a <=( (not A265)  and  a35317a );
 a35322a <=( A300  and  A298 );
 a35323a <=( (not A269)  and  a35322a );
 a35324a <=( a35323a  and  a35318a );
 a35328a <=( (not A199)  and  (not A166) );
 a35329a <=( (not A167)  and  a35328a );
 a35333a <=( A203  and  (not A202) );
 a35334a <=( A200  and  a35333a );
 a35335a <=( a35334a  and  a35329a );
 a35339a <=( (not A267)  and  (not A266) );
 a35340a <=( A265  and  a35339a );
 a35344a <=( A300  and  A299 );
 a35345a <=( A268  and  a35344a );
 a35346a <=( a35345a  and  a35340a );
 a35350a <=( (not A199)  and  (not A166) );
 a35351a <=( (not A167)  and  a35350a );
 a35355a <=( A203  and  (not A202) );
 a35356a <=( A200  and  a35355a );
 a35357a <=( a35356a  and  a35351a );
 a35361a <=( (not A267)  and  (not A266) );
 a35362a <=( A265  and  a35361a );
 a35366a <=( A300  and  A298 );
 a35367a <=( A268  and  a35366a );
 a35368a <=( a35367a  and  a35362a );
 a35372a <=( (not A199)  and  (not A166) );
 a35373a <=( (not A167)  and  a35372a );
 a35377a <=( A203  and  (not A202) );
 a35378a <=( A200  and  a35377a );
 a35379a <=( a35378a  and  a35373a );
 a35383a <=( (not A267)  and  (not A266) );
 a35384a <=( A265  and  a35383a );
 a35388a <=( A300  and  A299 );
 a35389a <=( (not A269)  and  a35388a );
 a35390a <=( a35389a  and  a35384a );
 a35394a <=( (not A199)  and  (not A166) );
 a35395a <=( (not A167)  and  a35394a );
 a35399a <=( A203  and  (not A202) );
 a35400a <=( A200  and  a35399a );
 a35401a <=( a35400a  and  a35395a );
 a35405a <=( (not A267)  and  (not A266) );
 a35406a <=( A265  and  a35405a );
 a35410a <=( A300  and  A298 );
 a35411a <=( (not A269)  and  a35410a );
 a35412a <=( a35411a  and  a35406a );
 a35416a <=( (not A199)  and  (not A166) );
 a35417a <=( (not A167)  and  a35416a );
 a35421a <=( A202  and  (not A201) );
 a35422a <=( A200  and  a35421a );
 a35423a <=( a35422a  and  a35417a );
 a35427a <=( A298  and  A267 );
 a35428a <=( A265  and  a35427a );
 a35432a <=( (not A301)  and  (not A300) );
 a35433a <=( A299  and  a35432a );
 a35434a <=( a35433a  and  a35428a );
 a35438a <=( (not A199)  and  (not A166) );
 a35439a <=( (not A167)  and  a35438a );
 a35443a <=( A202  and  (not A201) );
 a35444a <=( A200  and  a35443a );
 a35445a <=( a35444a  and  a35439a );
 a35449a <=( A298  and  A267 );
 a35450a <=( A265  and  a35449a );
 a35454a <=( A302  and  (not A300) );
 a35455a <=( A299  and  a35454a );
 a35456a <=( a35455a  and  a35450a );
 a35460a <=( (not A199)  and  (not A166) );
 a35461a <=( (not A167)  and  a35460a );
 a35465a <=( A202  and  (not A201) );
 a35466a <=( A200  and  a35465a );
 a35467a <=( a35466a  and  a35461a );
 a35471a <=( A298  and  A267 );
 a35472a <=( A265  and  a35471a );
 a35476a <=( A301  and  (not A300) );
 a35477a <=( (not A299)  and  a35476a );
 a35478a <=( a35477a  and  a35472a );
 a35482a <=( (not A199)  and  (not A166) );
 a35483a <=( (not A167)  and  a35482a );
 a35487a <=( A202  and  (not A201) );
 a35488a <=( A200  and  a35487a );
 a35489a <=( a35488a  and  a35483a );
 a35493a <=( A298  and  A267 );
 a35494a <=( A265  and  a35493a );
 a35498a <=( (not A302)  and  (not A300) );
 a35499a <=( (not A299)  and  a35498a );
 a35500a <=( a35499a  and  a35494a );
 a35504a <=( (not A199)  and  (not A166) );
 a35505a <=( (not A167)  and  a35504a );
 a35509a <=( A202  and  (not A201) );
 a35510a <=( A200  and  a35509a );
 a35511a <=( a35510a  and  a35505a );
 a35515a <=( (not A298)  and  A267 );
 a35516a <=( A265  and  a35515a );
 a35520a <=( A301  and  (not A300) );
 a35521a <=( A299  and  a35520a );
 a35522a <=( a35521a  and  a35516a );
 a35526a <=( (not A199)  and  (not A166) );
 a35527a <=( (not A167)  and  a35526a );
 a35531a <=( A202  and  (not A201) );
 a35532a <=( A200  and  a35531a );
 a35533a <=( a35532a  and  a35527a );
 a35537a <=( (not A298)  and  A267 );
 a35538a <=( A265  and  a35537a );
 a35542a <=( (not A302)  and  (not A300) );
 a35543a <=( A299  and  a35542a );
 a35544a <=( a35543a  and  a35538a );
 a35548a <=( (not A199)  and  (not A166) );
 a35549a <=( (not A167)  and  a35548a );
 a35553a <=( A202  and  (not A201) );
 a35554a <=( A200  and  a35553a );
 a35555a <=( a35554a  and  a35549a );
 a35559a <=( A298  and  A267 );
 a35560a <=( A266  and  a35559a );
 a35564a <=( (not A301)  and  (not A300) );
 a35565a <=( A299  and  a35564a );
 a35566a <=( a35565a  and  a35560a );
 a35570a <=( (not A199)  and  (not A166) );
 a35571a <=( (not A167)  and  a35570a );
 a35575a <=( A202  and  (not A201) );
 a35576a <=( A200  and  a35575a );
 a35577a <=( a35576a  and  a35571a );
 a35581a <=( A298  and  A267 );
 a35582a <=( A266  and  a35581a );
 a35586a <=( A302  and  (not A300) );
 a35587a <=( A299  and  a35586a );
 a35588a <=( a35587a  and  a35582a );
 a35592a <=( (not A199)  and  (not A166) );
 a35593a <=( (not A167)  and  a35592a );
 a35597a <=( A202  and  (not A201) );
 a35598a <=( A200  and  a35597a );
 a35599a <=( a35598a  and  a35593a );
 a35603a <=( A298  and  A267 );
 a35604a <=( A266  and  a35603a );
 a35608a <=( A301  and  (not A300) );
 a35609a <=( (not A299)  and  a35608a );
 a35610a <=( a35609a  and  a35604a );
 a35614a <=( (not A199)  and  (not A166) );
 a35615a <=( (not A167)  and  a35614a );
 a35619a <=( A202  and  (not A201) );
 a35620a <=( A200  and  a35619a );
 a35621a <=( a35620a  and  a35615a );
 a35625a <=( A298  and  A267 );
 a35626a <=( A266  and  a35625a );
 a35630a <=( (not A302)  and  (not A300) );
 a35631a <=( (not A299)  and  a35630a );
 a35632a <=( a35631a  and  a35626a );
 a35636a <=( (not A199)  and  (not A166) );
 a35637a <=( (not A167)  and  a35636a );
 a35641a <=( A202  and  (not A201) );
 a35642a <=( A200  and  a35641a );
 a35643a <=( a35642a  and  a35637a );
 a35647a <=( (not A298)  and  A267 );
 a35648a <=( A266  and  a35647a );
 a35652a <=( A301  and  (not A300) );
 a35653a <=( A299  and  a35652a );
 a35654a <=( a35653a  and  a35648a );
 a35658a <=( (not A199)  and  (not A166) );
 a35659a <=( (not A167)  and  a35658a );
 a35663a <=( A202  and  (not A201) );
 a35664a <=( A200  and  a35663a );
 a35665a <=( a35664a  and  a35659a );
 a35669a <=( (not A298)  and  A267 );
 a35670a <=( A266  and  a35669a );
 a35674a <=( (not A302)  and  (not A300) );
 a35675a <=( A299  and  a35674a );
 a35676a <=( a35675a  and  a35670a );
 a35680a <=( (not A199)  and  (not A166) );
 a35681a <=( (not A167)  and  a35680a );
 a35685a <=( (not A203)  and  (not A201) );
 a35686a <=( A200  and  a35685a );
 a35687a <=( a35686a  and  a35681a );
 a35691a <=( A298  and  A267 );
 a35692a <=( A265  and  a35691a );
 a35696a <=( (not A301)  and  (not A300) );
 a35697a <=( A299  and  a35696a );
 a35698a <=( a35697a  and  a35692a );
 a35702a <=( (not A199)  and  (not A166) );
 a35703a <=( (not A167)  and  a35702a );
 a35707a <=( (not A203)  and  (not A201) );
 a35708a <=( A200  and  a35707a );
 a35709a <=( a35708a  and  a35703a );
 a35713a <=( A298  and  A267 );
 a35714a <=( A265  and  a35713a );
 a35718a <=( A302  and  (not A300) );
 a35719a <=( A299  and  a35718a );
 a35720a <=( a35719a  and  a35714a );
 a35724a <=( (not A199)  and  (not A166) );
 a35725a <=( (not A167)  and  a35724a );
 a35729a <=( (not A203)  and  (not A201) );
 a35730a <=( A200  and  a35729a );
 a35731a <=( a35730a  and  a35725a );
 a35735a <=( A298  and  A267 );
 a35736a <=( A265  and  a35735a );
 a35740a <=( A301  and  (not A300) );
 a35741a <=( (not A299)  and  a35740a );
 a35742a <=( a35741a  and  a35736a );
 a35746a <=( (not A199)  and  (not A166) );
 a35747a <=( (not A167)  and  a35746a );
 a35751a <=( (not A203)  and  (not A201) );
 a35752a <=( A200  and  a35751a );
 a35753a <=( a35752a  and  a35747a );
 a35757a <=( A298  and  A267 );
 a35758a <=( A265  and  a35757a );
 a35762a <=( (not A302)  and  (not A300) );
 a35763a <=( (not A299)  and  a35762a );
 a35764a <=( a35763a  and  a35758a );
 a35768a <=( (not A199)  and  (not A166) );
 a35769a <=( (not A167)  and  a35768a );
 a35773a <=( (not A203)  and  (not A201) );
 a35774a <=( A200  and  a35773a );
 a35775a <=( a35774a  and  a35769a );
 a35779a <=( (not A298)  and  A267 );
 a35780a <=( A265  and  a35779a );
 a35784a <=( A301  and  (not A300) );
 a35785a <=( A299  and  a35784a );
 a35786a <=( a35785a  and  a35780a );
 a35790a <=( (not A199)  and  (not A166) );
 a35791a <=( (not A167)  and  a35790a );
 a35795a <=( (not A203)  and  (not A201) );
 a35796a <=( A200  and  a35795a );
 a35797a <=( a35796a  and  a35791a );
 a35801a <=( (not A298)  and  A267 );
 a35802a <=( A265  and  a35801a );
 a35806a <=( (not A302)  and  (not A300) );
 a35807a <=( A299  and  a35806a );
 a35808a <=( a35807a  and  a35802a );
 a35812a <=( (not A199)  and  (not A166) );
 a35813a <=( (not A167)  and  a35812a );
 a35817a <=( (not A203)  and  (not A201) );
 a35818a <=( A200  and  a35817a );
 a35819a <=( a35818a  and  a35813a );
 a35823a <=( A298  and  A267 );
 a35824a <=( A266  and  a35823a );
 a35828a <=( (not A301)  and  (not A300) );
 a35829a <=( A299  and  a35828a );
 a35830a <=( a35829a  and  a35824a );
 a35834a <=( (not A199)  and  (not A166) );
 a35835a <=( (not A167)  and  a35834a );
 a35839a <=( (not A203)  and  (not A201) );
 a35840a <=( A200  and  a35839a );
 a35841a <=( a35840a  and  a35835a );
 a35845a <=( A298  and  A267 );
 a35846a <=( A266  and  a35845a );
 a35850a <=( A302  and  (not A300) );
 a35851a <=( A299  and  a35850a );
 a35852a <=( a35851a  and  a35846a );
 a35856a <=( (not A199)  and  (not A166) );
 a35857a <=( (not A167)  and  a35856a );
 a35861a <=( (not A203)  and  (not A201) );
 a35862a <=( A200  and  a35861a );
 a35863a <=( a35862a  and  a35857a );
 a35867a <=( A298  and  A267 );
 a35868a <=( A266  and  a35867a );
 a35872a <=( A301  and  (not A300) );
 a35873a <=( (not A299)  and  a35872a );
 a35874a <=( a35873a  and  a35868a );
 a35878a <=( (not A199)  and  (not A166) );
 a35879a <=( (not A167)  and  a35878a );
 a35883a <=( (not A203)  and  (not A201) );
 a35884a <=( A200  and  a35883a );
 a35885a <=( a35884a  and  a35879a );
 a35889a <=( A298  and  A267 );
 a35890a <=( A266  and  a35889a );
 a35894a <=( (not A302)  and  (not A300) );
 a35895a <=( (not A299)  and  a35894a );
 a35896a <=( a35895a  and  a35890a );
 a35900a <=( (not A199)  and  (not A166) );
 a35901a <=( (not A167)  and  a35900a );
 a35905a <=( (not A203)  and  (not A201) );
 a35906a <=( A200  and  a35905a );
 a35907a <=( a35906a  and  a35901a );
 a35911a <=( (not A298)  and  A267 );
 a35912a <=( A266  and  a35911a );
 a35916a <=( A301  and  (not A300) );
 a35917a <=( A299  and  a35916a );
 a35918a <=( a35917a  and  a35912a );
 a35922a <=( (not A199)  and  (not A166) );
 a35923a <=( (not A167)  and  a35922a );
 a35927a <=( (not A203)  and  (not A201) );
 a35928a <=( A200  and  a35927a );
 a35929a <=( a35928a  and  a35923a );
 a35933a <=( (not A298)  and  A267 );
 a35934a <=( A266  and  a35933a );
 a35938a <=( (not A302)  and  (not A300) );
 a35939a <=( A299  and  a35938a );
 a35940a <=( a35939a  and  a35934a );
 a35944a <=( A199  and  (not A166) );
 a35945a <=( (not A167)  and  a35944a );
 a35949a <=( A203  and  (not A202) );
 a35950a <=( (not A200)  and  a35949a );
 a35951a <=( a35950a  and  a35945a );
 a35955a <=( (not A267)  and  A266 );
 a35956a <=( A265  and  a35955a );
 a35960a <=( A300  and  A299 );
 a35961a <=( (not A268)  and  a35960a );
 a35962a <=( a35961a  and  a35956a );
 a35966a <=( A199  and  (not A166) );
 a35967a <=( (not A167)  and  a35966a );
 a35971a <=( A203  and  (not A202) );
 a35972a <=( (not A200)  and  a35971a );
 a35973a <=( a35972a  and  a35967a );
 a35977a <=( (not A267)  and  A266 );
 a35978a <=( A265  and  a35977a );
 a35982a <=( A300  and  A298 );
 a35983a <=( (not A268)  and  a35982a );
 a35984a <=( a35983a  and  a35978a );
 a35988a <=( A199  and  (not A166) );
 a35989a <=( (not A167)  and  a35988a );
 a35993a <=( A203  and  (not A202) );
 a35994a <=( (not A200)  and  a35993a );
 a35995a <=( a35994a  and  a35989a );
 a35999a <=( (not A267)  and  A266 );
 a36000a <=( A265  and  a35999a );
 a36004a <=( A300  and  A299 );
 a36005a <=( A269  and  a36004a );
 a36006a <=( a36005a  and  a36000a );
 a36010a <=( A199  and  (not A166) );
 a36011a <=( (not A167)  and  a36010a );
 a36015a <=( A203  and  (not A202) );
 a36016a <=( (not A200)  and  a36015a );
 a36017a <=( a36016a  and  a36011a );
 a36021a <=( (not A267)  and  A266 );
 a36022a <=( A265  and  a36021a );
 a36026a <=( A300  and  A298 );
 a36027a <=( A269  and  a36026a );
 a36028a <=( a36027a  and  a36022a );
 a36032a <=( A199  and  (not A166) );
 a36033a <=( (not A167)  and  a36032a );
 a36037a <=( A203  and  (not A202) );
 a36038a <=( (not A200)  and  a36037a );
 a36039a <=( a36038a  and  a36033a );
 a36043a <=( (not A267)  and  A266 );
 a36044a <=( (not A265)  and  a36043a );
 a36048a <=( A300  and  A299 );
 a36049a <=( A268  and  a36048a );
 a36050a <=( a36049a  and  a36044a );
 a36054a <=( A199  and  (not A166) );
 a36055a <=( (not A167)  and  a36054a );
 a36059a <=( A203  and  (not A202) );
 a36060a <=( (not A200)  and  a36059a );
 a36061a <=( a36060a  and  a36055a );
 a36065a <=( (not A267)  and  A266 );
 a36066a <=( (not A265)  and  a36065a );
 a36070a <=( A300  and  A298 );
 a36071a <=( A268  and  a36070a );
 a36072a <=( a36071a  and  a36066a );
 a36076a <=( A199  and  (not A166) );
 a36077a <=( (not A167)  and  a36076a );
 a36081a <=( A203  and  (not A202) );
 a36082a <=( (not A200)  and  a36081a );
 a36083a <=( a36082a  and  a36077a );
 a36087a <=( (not A267)  and  A266 );
 a36088a <=( (not A265)  and  a36087a );
 a36092a <=( A300  and  A299 );
 a36093a <=( (not A269)  and  a36092a );
 a36094a <=( a36093a  and  a36088a );
 a36098a <=( A199  and  (not A166) );
 a36099a <=( (not A167)  and  a36098a );
 a36103a <=( A203  and  (not A202) );
 a36104a <=( (not A200)  and  a36103a );
 a36105a <=( a36104a  and  a36099a );
 a36109a <=( (not A267)  and  A266 );
 a36110a <=( (not A265)  and  a36109a );
 a36114a <=( A300  and  A298 );
 a36115a <=( (not A269)  and  a36114a );
 a36116a <=( a36115a  and  a36110a );
 a36120a <=( A199  and  (not A166) );
 a36121a <=( (not A167)  and  a36120a );
 a36125a <=( A203  and  (not A202) );
 a36126a <=( (not A200)  and  a36125a );
 a36127a <=( a36126a  and  a36121a );
 a36131a <=( (not A267)  and  (not A266) );
 a36132a <=( A265  and  a36131a );
 a36136a <=( A300  and  A299 );
 a36137a <=( A268  and  a36136a );
 a36138a <=( a36137a  and  a36132a );
 a36142a <=( A199  and  (not A166) );
 a36143a <=( (not A167)  and  a36142a );
 a36147a <=( A203  and  (not A202) );
 a36148a <=( (not A200)  and  a36147a );
 a36149a <=( a36148a  and  a36143a );
 a36153a <=( (not A267)  and  (not A266) );
 a36154a <=( A265  and  a36153a );
 a36158a <=( A300  and  A298 );
 a36159a <=( A268  and  a36158a );
 a36160a <=( a36159a  and  a36154a );
 a36164a <=( A199  and  (not A166) );
 a36165a <=( (not A167)  and  a36164a );
 a36169a <=( A203  and  (not A202) );
 a36170a <=( (not A200)  and  a36169a );
 a36171a <=( a36170a  and  a36165a );
 a36175a <=( (not A267)  and  (not A266) );
 a36176a <=( A265  and  a36175a );
 a36180a <=( A300  and  A299 );
 a36181a <=( (not A269)  and  a36180a );
 a36182a <=( a36181a  and  a36176a );
 a36186a <=( A199  and  (not A166) );
 a36187a <=( (not A167)  and  a36186a );
 a36191a <=( A203  and  (not A202) );
 a36192a <=( (not A200)  and  a36191a );
 a36193a <=( a36192a  and  a36187a );
 a36197a <=( (not A267)  and  (not A266) );
 a36198a <=( A265  and  a36197a );
 a36202a <=( A300  and  A298 );
 a36203a <=( (not A269)  and  a36202a );
 a36204a <=( a36203a  and  a36198a );
 a36208a <=( A199  and  (not A166) );
 a36209a <=( (not A167)  and  a36208a );
 a36213a <=( A202  and  (not A201) );
 a36214a <=( (not A200)  and  a36213a );
 a36215a <=( a36214a  and  a36209a );
 a36219a <=( A298  and  A267 );
 a36220a <=( A265  and  a36219a );
 a36224a <=( (not A301)  and  (not A300) );
 a36225a <=( A299  and  a36224a );
 a36226a <=( a36225a  and  a36220a );
 a36230a <=( A199  and  (not A166) );
 a36231a <=( (not A167)  and  a36230a );
 a36235a <=( A202  and  (not A201) );
 a36236a <=( (not A200)  and  a36235a );
 a36237a <=( a36236a  and  a36231a );
 a36241a <=( A298  and  A267 );
 a36242a <=( A265  and  a36241a );
 a36246a <=( A302  and  (not A300) );
 a36247a <=( A299  and  a36246a );
 a36248a <=( a36247a  and  a36242a );
 a36252a <=( A199  and  (not A166) );
 a36253a <=( (not A167)  and  a36252a );
 a36257a <=( A202  and  (not A201) );
 a36258a <=( (not A200)  and  a36257a );
 a36259a <=( a36258a  and  a36253a );
 a36263a <=( A298  and  A267 );
 a36264a <=( A265  and  a36263a );
 a36268a <=( A301  and  (not A300) );
 a36269a <=( (not A299)  and  a36268a );
 a36270a <=( a36269a  and  a36264a );
 a36274a <=( A199  and  (not A166) );
 a36275a <=( (not A167)  and  a36274a );
 a36279a <=( A202  and  (not A201) );
 a36280a <=( (not A200)  and  a36279a );
 a36281a <=( a36280a  and  a36275a );
 a36285a <=( A298  and  A267 );
 a36286a <=( A265  and  a36285a );
 a36290a <=( (not A302)  and  (not A300) );
 a36291a <=( (not A299)  and  a36290a );
 a36292a <=( a36291a  and  a36286a );
 a36296a <=( A199  and  (not A166) );
 a36297a <=( (not A167)  and  a36296a );
 a36301a <=( A202  and  (not A201) );
 a36302a <=( (not A200)  and  a36301a );
 a36303a <=( a36302a  and  a36297a );
 a36307a <=( (not A298)  and  A267 );
 a36308a <=( A265  and  a36307a );
 a36312a <=( A301  and  (not A300) );
 a36313a <=( A299  and  a36312a );
 a36314a <=( a36313a  and  a36308a );
 a36318a <=( A199  and  (not A166) );
 a36319a <=( (not A167)  and  a36318a );
 a36323a <=( A202  and  (not A201) );
 a36324a <=( (not A200)  and  a36323a );
 a36325a <=( a36324a  and  a36319a );
 a36329a <=( (not A298)  and  A267 );
 a36330a <=( A265  and  a36329a );
 a36334a <=( (not A302)  and  (not A300) );
 a36335a <=( A299  and  a36334a );
 a36336a <=( a36335a  and  a36330a );
 a36340a <=( A199  and  (not A166) );
 a36341a <=( (not A167)  and  a36340a );
 a36345a <=( A202  and  (not A201) );
 a36346a <=( (not A200)  and  a36345a );
 a36347a <=( a36346a  and  a36341a );
 a36351a <=( A298  and  A267 );
 a36352a <=( A266  and  a36351a );
 a36356a <=( (not A301)  and  (not A300) );
 a36357a <=( A299  and  a36356a );
 a36358a <=( a36357a  and  a36352a );
 a36362a <=( A199  and  (not A166) );
 a36363a <=( (not A167)  and  a36362a );
 a36367a <=( A202  and  (not A201) );
 a36368a <=( (not A200)  and  a36367a );
 a36369a <=( a36368a  and  a36363a );
 a36373a <=( A298  and  A267 );
 a36374a <=( A266  and  a36373a );
 a36378a <=( A302  and  (not A300) );
 a36379a <=( A299  and  a36378a );
 a36380a <=( a36379a  and  a36374a );
 a36384a <=( A199  and  (not A166) );
 a36385a <=( (not A167)  and  a36384a );
 a36389a <=( A202  and  (not A201) );
 a36390a <=( (not A200)  and  a36389a );
 a36391a <=( a36390a  and  a36385a );
 a36395a <=( A298  and  A267 );
 a36396a <=( A266  and  a36395a );
 a36400a <=( A301  and  (not A300) );
 a36401a <=( (not A299)  and  a36400a );
 a36402a <=( a36401a  and  a36396a );
 a36406a <=( A199  and  (not A166) );
 a36407a <=( (not A167)  and  a36406a );
 a36411a <=( A202  and  (not A201) );
 a36412a <=( (not A200)  and  a36411a );
 a36413a <=( a36412a  and  a36407a );
 a36417a <=( A298  and  A267 );
 a36418a <=( A266  and  a36417a );
 a36422a <=( (not A302)  and  (not A300) );
 a36423a <=( (not A299)  and  a36422a );
 a36424a <=( a36423a  and  a36418a );
 a36428a <=( A199  and  (not A166) );
 a36429a <=( (not A167)  and  a36428a );
 a36433a <=( A202  and  (not A201) );
 a36434a <=( (not A200)  and  a36433a );
 a36435a <=( a36434a  and  a36429a );
 a36439a <=( (not A298)  and  A267 );
 a36440a <=( A266  and  a36439a );
 a36444a <=( A301  and  (not A300) );
 a36445a <=( A299  and  a36444a );
 a36446a <=( a36445a  and  a36440a );
 a36450a <=( A199  and  (not A166) );
 a36451a <=( (not A167)  and  a36450a );
 a36455a <=( A202  and  (not A201) );
 a36456a <=( (not A200)  and  a36455a );
 a36457a <=( a36456a  and  a36451a );
 a36461a <=( (not A298)  and  A267 );
 a36462a <=( A266  and  a36461a );
 a36466a <=( (not A302)  and  (not A300) );
 a36467a <=( A299  and  a36466a );
 a36468a <=( a36467a  and  a36462a );
 a36472a <=( A199  and  (not A166) );
 a36473a <=( (not A167)  and  a36472a );
 a36477a <=( (not A203)  and  (not A201) );
 a36478a <=( (not A200)  and  a36477a );
 a36479a <=( a36478a  and  a36473a );
 a36483a <=( A298  and  A267 );
 a36484a <=( A265  and  a36483a );
 a36488a <=( (not A301)  and  (not A300) );
 a36489a <=( A299  and  a36488a );
 a36490a <=( a36489a  and  a36484a );
 a36494a <=( A199  and  (not A166) );
 a36495a <=( (not A167)  and  a36494a );
 a36499a <=( (not A203)  and  (not A201) );
 a36500a <=( (not A200)  and  a36499a );
 a36501a <=( a36500a  and  a36495a );
 a36505a <=( A298  and  A267 );
 a36506a <=( A265  and  a36505a );
 a36510a <=( A302  and  (not A300) );
 a36511a <=( A299  and  a36510a );
 a36512a <=( a36511a  and  a36506a );
 a36516a <=( A199  and  (not A166) );
 a36517a <=( (not A167)  and  a36516a );
 a36521a <=( (not A203)  and  (not A201) );
 a36522a <=( (not A200)  and  a36521a );
 a36523a <=( a36522a  and  a36517a );
 a36527a <=( A298  and  A267 );
 a36528a <=( A265  and  a36527a );
 a36532a <=( A301  and  (not A300) );
 a36533a <=( (not A299)  and  a36532a );
 a36534a <=( a36533a  and  a36528a );
 a36538a <=( A199  and  (not A166) );
 a36539a <=( (not A167)  and  a36538a );
 a36543a <=( (not A203)  and  (not A201) );
 a36544a <=( (not A200)  and  a36543a );
 a36545a <=( a36544a  and  a36539a );
 a36549a <=( A298  and  A267 );
 a36550a <=( A265  and  a36549a );
 a36554a <=( (not A302)  and  (not A300) );
 a36555a <=( (not A299)  and  a36554a );
 a36556a <=( a36555a  and  a36550a );
 a36560a <=( A199  and  (not A166) );
 a36561a <=( (not A167)  and  a36560a );
 a36565a <=( (not A203)  and  (not A201) );
 a36566a <=( (not A200)  and  a36565a );
 a36567a <=( a36566a  and  a36561a );
 a36571a <=( (not A298)  and  A267 );
 a36572a <=( A265  and  a36571a );
 a36576a <=( A301  and  (not A300) );
 a36577a <=( A299  and  a36576a );
 a36578a <=( a36577a  and  a36572a );
 a36582a <=( A199  and  (not A166) );
 a36583a <=( (not A167)  and  a36582a );
 a36587a <=( (not A203)  and  (not A201) );
 a36588a <=( (not A200)  and  a36587a );
 a36589a <=( a36588a  and  a36583a );
 a36593a <=( (not A298)  and  A267 );
 a36594a <=( A265  and  a36593a );
 a36598a <=( (not A302)  and  (not A300) );
 a36599a <=( A299  and  a36598a );
 a36600a <=( a36599a  and  a36594a );
 a36604a <=( A199  and  (not A166) );
 a36605a <=( (not A167)  and  a36604a );
 a36609a <=( (not A203)  and  (not A201) );
 a36610a <=( (not A200)  and  a36609a );
 a36611a <=( a36610a  and  a36605a );
 a36615a <=( A298  and  A267 );
 a36616a <=( A266  and  a36615a );
 a36620a <=( (not A301)  and  (not A300) );
 a36621a <=( A299  and  a36620a );
 a36622a <=( a36621a  and  a36616a );
 a36626a <=( A199  and  (not A166) );
 a36627a <=( (not A167)  and  a36626a );
 a36631a <=( (not A203)  and  (not A201) );
 a36632a <=( (not A200)  and  a36631a );
 a36633a <=( a36632a  and  a36627a );
 a36637a <=( A298  and  A267 );
 a36638a <=( A266  and  a36637a );
 a36642a <=( A302  and  (not A300) );
 a36643a <=( A299  and  a36642a );
 a36644a <=( a36643a  and  a36638a );
 a36648a <=( A199  and  (not A166) );
 a36649a <=( (not A167)  and  a36648a );
 a36653a <=( (not A203)  and  (not A201) );
 a36654a <=( (not A200)  and  a36653a );
 a36655a <=( a36654a  and  a36649a );
 a36659a <=( A298  and  A267 );
 a36660a <=( A266  and  a36659a );
 a36664a <=( A301  and  (not A300) );
 a36665a <=( (not A299)  and  a36664a );
 a36666a <=( a36665a  and  a36660a );
 a36670a <=( A199  and  (not A166) );
 a36671a <=( (not A167)  and  a36670a );
 a36675a <=( (not A203)  and  (not A201) );
 a36676a <=( (not A200)  and  a36675a );
 a36677a <=( a36676a  and  a36671a );
 a36681a <=( A298  and  A267 );
 a36682a <=( A266  and  a36681a );
 a36686a <=( (not A302)  and  (not A300) );
 a36687a <=( (not A299)  and  a36686a );
 a36688a <=( a36687a  and  a36682a );
 a36692a <=( A199  and  (not A166) );
 a36693a <=( (not A167)  and  a36692a );
 a36697a <=( (not A203)  and  (not A201) );
 a36698a <=( (not A200)  and  a36697a );
 a36699a <=( a36698a  and  a36693a );
 a36703a <=( (not A298)  and  A267 );
 a36704a <=( A266  and  a36703a );
 a36708a <=( A301  and  (not A300) );
 a36709a <=( A299  and  a36708a );
 a36710a <=( a36709a  and  a36704a );
 a36714a <=( A199  and  (not A166) );
 a36715a <=( (not A167)  and  a36714a );
 a36719a <=( (not A203)  and  (not A201) );
 a36720a <=( (not A200)  and  a36719a );
 a36721a <=( a36720a  and  a36715a );
 a36725a <=( (not A298)  and  A267 );
 a36726a <=( A266  and  a36725a );
 a36730a <=( (not A302)  and  (not A300) );
 a36731a <=( A299  and  a36730a );
 a36732a <=( a36731a  and  a36726a );
 a36736a <=( (not A199)  and  (not A166) );
 a36737a <=( (not A167)  and  a36736a );
 a36741a <=( A265  and  (not A202) );
 a36742a <=( (not A200)  and  a36741a );
 a36743a <=( a36742a  and  a36737a );
 a36747a <=( (not A269)  and  A268 );
 a36748a <=( A266  and  a36747a );
 a36752a <=( (not A301)  and  (not A299) );
 a36753a <=( (not A298)  and  a36752a );
 a36754a <=( a36753a  and  a36748a );
 a36758a <=( (not A199)  and  (not A166) );
 a36759a <=( (not A167)  and  a36758a );
 a36763a <=( A265  and  (not A202) );
 a36764a <=( (not A200)  and  a36763a );
 a36765a <=( a36764a  and  a36759a );
 a36769a <=( (not A269)  and  A268 );
 a36770a <=( A266  and  a36769a );
 a36774a <=( A302  and  (not A299) );
 a36775a <=( (not A298)  and  a36774a );
 a36776a <=( a36775a  and  a36770a );
 a36780a <=( (not A199)  and  (not A166) );
 a36781a <=( (not A167)  and  a36780a );
 a36785a <=( (not A265)  and  (not A202) );
 a36786a <=( (not A200)  and  a36785a );
 a36787a <=( a36786a  and  a36781a );
 a36791a <=( A269  and  (not A268) );
 a36792a <=( A266  and  a36791a );
 a36796a <=( (not A301)  and  (not A299) );
 a36797a <=( (not A298)  and  a36796a );
 a36798a <=( a36797a  and  a36792a );
 a36802a <=( (not A199)  and  (not A166) );
 a36803a <=( (not A167)  and  a36802a );
 a36807a <=( (not A265)  and  (not A202) );
 a36808a <=( (not A200)  and  a36807a );
 a36809a <=( a36808a  and  a36803a );
 a36813a <=( A269  and  (not A268) );
 a36814a <=( A266  and  a36813a );
 a36818a <=( A302  and  (not A299) );
 a36819a <=( (not A298)  and  a36818a );
 a36820a <=( a36819a  and  a36814a );
 a36824a <=( (not A199)  and  (not A166) );
 a36825a <=( (not A167)  and  a36824a );
 a36829a <=( A265  and  (not A202) );
 a36830a <=( (not A200)  and  a36829a );
 a36831a <=( a36830a  and  a36825a );
 a36835a <=( A269  and  (not A268) );
 a36836a <=( (not A266)  and  a36835a );
 a36840a <=( (not A301)  and  (not A299) );
 a36841a <=( (not A298)  and  a36840a );
 a36842a <=( a36841a  and  a36836a );
 a36846a <=( (not A199)  and  (not A166) );
 a36847a <=( (not A167)  and  a36846a );
 a36851a <=( A265  and  (not A202) );
 a36852a <=( (not A200)  and  a36851a );
 a36853a <=( a36852a  and  a36847a );
 a36857a <=( A269  and  (not A268) );
 a36858a <=( (not A266)  and  a36857a );
 a36862a <=( A302  and  (not A299) );
 a36863a <=( (not A298)  and  a36862a );
 a36864a <=( a36863a  and  a36858a );
 a36868a <=( (not A199)  and  (not A166) );
 a36869a <=( (not A167)  and  a36868a );
 a36873a <=( (not A265)  and  (not A202) );
 a36874a <=( (not A200)  and  a36873a );
 a36875a <=( a36874a  and  a36869a );
 a36879a <=( (not A269)  and  A268 );
 a36880a <=( (not A266)  and  a36879a );
 a36884a <=( (not A301)  and  (not A299) );
 a36885a <=( (not A298)  and  a36884a );
 a36886a <=( a36885a  and  a36880a );
 a36890a <=( (not A199)  and  (not A166) );
 a36891a <=( (not A167)  and  a36890a );
 a36895a <=( (not A265)  and  (not A202) );
 a36896a <=( (not A200)  and  a36895a );
 a36897a <=( a36896a  and  a36891a );
 a36901a <=( (not A269)  and  A268 );
 a36902a <=( (not A266)  and  a36901a );
 a36906a <=( A302  and  (not A299) );
 a36907a <=( (not A298)  and  a36906a );
 a36908a <=( a36907a  and  a36902a );
 a36912a <=( (not A199)  and  (not A166) );
 a36913a <=( (not A167)  and  a36912a );
 a36917a <=( A265  and  A203 );
 a36918a <=( (not A200)  and  a36917a );
 a36919a <=( a36918a  and  a36913a );
 a36923a <=( (not A269)  and  A268 );
 a36924a <=( A266  and  a36923a );
 a36928a <=( (not A301)  and  (not A299) );
 a36929a <=( (not A298)  and  a36928a );
 a36930a <=( a36929a  and  a36924a );
 a36934a <=( (not A199)  and  (not A166) );
 a36935a <=( (not A167)  and  a36934a );
 a36939a <=( A265  and  A203 );
 a36940a <=( (not A200)  and  a36939a );
 a36941a <=( a36940a  and  a36935a );
 a36945a <=( (not A269)  and  A268 );
 a36946a <=( A266  and  a36945a );
 a36950a <=( A302  and  (not A299) );
 a36951a <=( (not A298)  and  a36950a );
 a36952a <=( a36951a  and  a36946a );
 a36956a <=( (not A199)  and  (not A166) );
 a36957a <=( (not A167)  and  a36956a );
 a36961a <=( (not A265)  and  A203 );
 a36962a <=( (not A200)  and  a36961a );
 a36963a <=( a36962a  and  a36957a );
 a36967a <=( A269  and  (not A268) );
 a36968a <=( A266  and  a36967a );
 a36972a <=( (not A301)  and  (not A299) );
 a36973a <=( (not A298)  and  a36972a );
 a36974a <=( a36973a  and  a36968a );
 a36978a <=( (not A199)  and  (not A166) );
 a36979a <=( (not A167)  and  a36978a );
 a36983a <=( (not A265)  and  A203 );
 a36984a <=( (not A200)  and  a36983a );
 a36985a <=( a36984a  and  a36979a );
 a36989a <=( A269  and  (not A268) );
 a36990a <=( A266  and  a36989a );
 a36994a <=( A302  and  (not A299) );
 a36995a <=( (not A298)  and  a36994a );
 a36996a <=( a36995a  and  a36990a );
 a37000a <=( (not A199)  and  (not A166) );
 a37001a <=( (not A167)  and  a37000a );
 a37005a <=( A265  and  A203 );
 a37006a <=( (not A200)  and  a37005a );
 a37007a <=( a37006a  and  a37001a );
 a37011a <=( A269  and  (not A268) );
 a37012a <=( (not A266)  and  a37011a );
 a37016a <=( (not A301)  and  (not A299) );
 a37017a <=( (not A298)  and  a37016a );
 a37018a <=( a37017a  and  a37012a );
 a37022a <=( (not A199)  and  (not A166) );
 a37023a <=( (not A167)  and  a37022a );
 a37027a <=( A265  and  A203 );
 a37028a <=( (not A200)  and  a37027a );
 a37029a <=( a37028a  and  a37023a );
 a37033a <=( A269  and  (not A268) );
 a37034a <=( (not A266)  and  a37033a );
 a37038a <=( A302  and  (not A299) );
 a37039a <=( (not A298)  and  a37038a );
 a37040a <=( a37039a  and  a37034a );
 a37044a <=( (not A199)  and  (not A166) );
 a37045a <=( (not A167)  and  a37044a );
 a37049a <=( (not A265)  and  A203 );
 a37050a <=( (not A200)  and  a37049a );
 a37051a <=( a37050a  and  a37045a );
 a37055a <=( (not A269)  and  A268 );
 a37056a <=( (not A266)  and  a37055a );
 a37060a <=( (not A301)  and  (not A299) );
 a37061a <=( (not A298)  and  a37060a );
 a37062a <=( a37061a  and  a37056a );
 a37066a <=( (not A199)  and  (not A166) );
 a37067a <=( (not A167)  and  a37066a );
 a37071a <=( (not A265)  and  A203 );
 a37072a <=( (not A200)  and  a37071a );
 a37073a <=( a37072a  and  a37067a );
 a37077a <=( (not A269)  and  A268 );
 a37078a <=( (not A266)  and  a37077a );
 a37082a <=( A302  and  (not A299) );
 a37083a <=( (not A298)  and  a37082a );
 a37084a <=( a37083a  and  a37078a );
 a37088a <=( (not A199)  and  (not A166) );
 a37089a <=( (not A167)  and  a37088a );
 a37093a <=( (not A203)  and  A202 );
 a37094a <=( (not A200)  and  a37093a );
 a37095a <=( a37094a  and  a37089a );
 a37099a <=( (not A267)  and  A266 );
 a37100a <=( A265  and  a37099a );
 a37104a <=( A300  and  A299 );
 a37105a <=( (not A268)  and  a37104a );
 a37106a <=( a37105a  and  a37100a );
 a37110a <=( (not A199)  and  (not A166) );
 a37111a <=( (not A167)  and  a37110a );
 a37115a <=( (not A203)  and  A202 );
 a37116a <=( (not A200)  and  a37115a );
 a37117a <=( a37116a  and  a37111a );
 a37121a <=( (not A267)  and  A266 );
 a37122a <=( A265  and  a37121a );
 a37126a <=( A300  and  A298 );
 a37127a <=( (not A268)  and  a37126a );
 a37128a <=( a37127a  and  a37122a );
 a37132a <=( (not A199)  and  (not A166) );
 a37133a <=( (not A167)  and  a37132a );
 a37137a <=( (not A203)  and  A202 );
 a37138a <=( (not A200)  and  a37137a );
 a37139a <=( a37138a  and  a37133a );
 a37143a <=( (not A267)  and  A266 );
 a37144a <=( A265  and  a37143a );
 a37148a <=( A300  and  A299 );
 a37149a <=( A269  and  a37148a );
 a37150a <=( a37149a  and  a37144a );
 a37154a <=( (not A199)  and  (not A166) );
 a37155a <=( (not A167)  and  a37154a );
 a37159a <=( (not A203)  and  A202 );
 a37160a <=( (not A200)  and  a37159a );
 a37161a <=( a37160a  and  a37155a );
 a37165a <=( (not A267)  and  A266 );
 a37166a <=( A265  and  a37165a );
 a37170a <=( A300  and  A298 );
 a37171a <=( A269  and  a37170a );
 a37172a <=( a37171a  and  a37166a );
 a37176a <=( (not A199)  and  (not A166) );
 a37177a <=( (not A167)  and  a37176a );
 a37181a <=( (not A203)  and  A202 );
 a37182a <=( (not A200)  and  a37181a );
 a37183a <=( a37182a  and  a37177a );
 a37187a <=( (not A267)  and  A266 );
 a37188a <=( (not A265)  and  a37187a );
 a37192a <=( A300  and  A299 );
 a37193a <=( A268  and  a37192a );
 a37194a <=( a37193a  and  a37188a );
 a37198a <=( (not A199)  and  (not A166) );
 a37199a <=( (not A167)  and  a37198a );
 a37203a <=( (not A203)  and  A202 );
 a37204a <=( (not A200)  and  a37203a );
 a37205a <=( a37204a  and  a37199a );
 a37209a <=( (not A267)  and  A266 );
 a37210a <=( (not A265)  and  a37209a );
 a37214a <=( A300  and  A298 );
 a37215a <=( A268  and  a37214a );
 a37216a <=( a37215a  and  a37210a );
 a37220a <=( (not A199)  and  (not A166) );
 a37221a <=( (not A167)  and  a37220a );
 a37225a <=( (not A203)  and  A202 );
 a37226a <=( (not A200)  and  a37225a );
 a37227a <=( a37226a  and  a37221a );
 a37231a <=( (not A267)  and  A266 );
 a37232a <=( (not A265)  and  a37231a );
 a37236a <=( A300  and  A299 );
 a37237a <=( (not A269)  and  a37236a );
 a37238a <=( a37237a  and  a37232a );
 a37242a <=( (not A199)  and  (not A166) );
 a37243a <=( (not A167)  and  a37242a );
 a37247a <=( (not A203)  and  A202 );
 a37248a <=( (not A200)  and  a37247a );
 a37249a <=( a37248a  and  a37243a );
 a37253a <=( (not A267)  and  A266 );
 a37254a <=( (not A265)  and  a37253a );
 a37258a <=( A300  and  A298 );
 a37259a <=( (not A269)  and  a37258a );
 a37260a <=( a37259a  and  a37254a );
 a37264a <=( (not A199)  and  (not A166) );
 a37265a <=( (not A167)  and  a37264a );
 a37269a <=( (not A203)  and  A202 );
 a37270a <=( (not A200)  and  a37269a );
 a37271a <=( a37270a  and  a37265a );
 a37275a <=( (not A267)  and  (not A266) );
 a37276a <=( A265  and  a37275a );
 a37280a <=( A300  and  A299 );
 a37281a <=( A268  and  a37280a );
 a37282a <=( a37281a  and  a37276a );
 a37286a <=( (not A199)  and  (not A166) );
 a37287a <=( (not A167)  and  a37286a );
 a37291a <=( (not A203)  and  A202 );
 a37292a <=( (not A200)  and  a37291a );
 a37293a <=( a37292a  and  a37287a );
 a37297a <=( (not A267)  and  (not A266) );
 a37298a <=( A265  and  a37297a );
 a37302a <=( A300  and  A298 );
 a37303a <=( A268  and  a37302a );
 a37304a <=( a37303a  and  a37298a );
 a37308a <=( (not A199)  and  (not A166) );
 a37309a <=( (not A167)  and  a37308a );
 a37313a <=( (not A203)  and  A202 );
 a37314a <=( (not A200)  and  a37313a );
 a37315a <=( a37314a  and  a37309a );
 a37319a <=( (not A267)  and  (not A266) );
 a37320a <=( A265  and  a37319a );
 a37324a <=( A300  and  A299 );
 a37325a <=( (not A269)  and  a37324a );
 a37326a <=( a37325a  and  a37320a );
 a37330a <=( (not A199)  and  (not A166) );
 a37331a <=( (not A167)  and  a37330a );
 a37335a <=( (not A203)  and  A202 );
 a37336a <=( (not A200)  and  a37335a );
 a37337a <=( a37336a  and  a37331a );
 a37341a <=( (not A267)  and  (not A266) );
 a37342a <=( A265  and  a37341a );
 a37346a <=( A300  and  A298 );
 a37347a <=( (not A269)  and  a37346a );
 a37348a <=( a37347a  and  a37342a );
 a37352a <=( A199  and  (not A167) );
 a37353a <=( (not A168)  and  a37352a );
 a37357a <=( A266  and  A265 );
 a37358a <=( A201  and  a37357a );
 a37359a <=( a37358a  and  a37353a );
 a37363a <=( A298  and  (not A268) );
 a37364a <=( (not A267)  and  a37363a );
 a37368a <=( (not A302)  and  A301 );
 a37369a <=( A299  and  a37368a );
 a37370a <=( a37369a  and  a37364a );
 a37374a <=( A199  and  (not A167) );
 a37375a <=( (not A168)  and  a37374a );
 a37379a <=( A266  and  A265 );
 a37380a <=( A201  and  a37379a );
 a37381a <=( a37380a  and  a37375a );
 a37385a <=( A298  and  (not A268) );
 a37386a <=( (not A267)  and  a37385a );
 a37390a <=( A302  and  (not A301) );
 a37391a <=( (not A299)  and  a37390a );
 a37392a <=( a37391a  and  a37386a );
 a37396a <=( A199  and  (not A167) );
 a37397a <=( (not A168)  and  a37396a );
 a37401a <=( A266  and  A265 );
 a37402a <=( A201  and  a37401a );
 a37403a <=( a37402a  and  a37397a );
 a37407a <=( (not A298)  and  (not A268) );
 a37408a <=( (not A267)  and  a37407a );
 a37412a <=( A302  and  (not A301) );
 a37413a <=( A299  and  a37412a );
 a37414a <=( a37413a  and  a37408a );
 a37418a <=( A199  and  (not A167) );
 a37419a <=( (not A168)  and  a37418a );
 a37423a <=( A266  and  A265 );
 a37424a <=( A201  and  a37423a );
 a37425a <=( a37424a  and  a37419a );
 a37429a <=( (not A298)  and  (not A268) );
 a37430a <=( (not A267)  and  a37429a );
 a37434a <=( (not A302)  and  A301 );
 a37435a <=( (not A299)  and  a37434a );
 a37436a <=( a37435a  and  a37430a );
 a37440a <=( A199  and  (not A167) );
 a37441a <=( (not A168)  and  a37440a );
 a37445a <=( A266  and  A265 );
 a37446a <=( A201  and  a37445a );
 a37447a <=( a37446a  and  a37441a );
 a37451a <=( A298  and  A269 );
 a37452a <=( (not A267)  and  a37451a );
 a37456a <=( (not A302)  and  A301 );
 a37457a <=( A299  and  a37456a );
 a37458a <=( a37457a  and  a37452a );
 a37462a <=( A199  and  (not A167) );
 a37463a <=( (not A168)  and  a37462a );
 a37467a <=( A266  and  A265 );
 a37468a <=( A201  and  a37467a );
 a37469a <=( a37468a  and  a37463a );
 a37473a <=( A298  and  A269 );
 a37474a <=( (not A267)  and  a37473a );
 a37478a <=( A302  and  (not A301) );
 a37479a <=( (not A299)  and  a37478a );
 a37480a <=( a37479a  and  a37474a );
 a37484a <=( A199  and  (not A167) );
 a37485a <=( (not A168)  and  a37484a );
 a37489a <=( A266  and  A265 );
 a37490a <=( A201  and  a37489a );
 a37491a <=( a37490a  and  a37485a );
 a37495a <=( (not A298)  and  A269 );
 a37496a <=( (not A267)  and  a37495a );
 a37500a <=( A302  and  (not A301) );
 a37501a <=( A299  and  a37500a );
 a37502a <=( a37501a  and  a37496a );
 a37506a <=( A199  and  (not A167) );
 a37507a <=( (not A168)  and  a37506a );
 a37511a <=( A266  and  A265 );
 a37512a <=( A201  and  a37511a );
 a37513a <=( a37512a  and  a37507a );
 a37517a <=( (not A298)  and  A269 );
 a37518a <=( (not A267)  and  a37517a );
 a37522a <=( (not A302)  and  A301 );
 a37523a <=( (not A299)  and  a37522a );
 a37524a <=( a37523a  and  a37518a );
 a37528a <=( A199  and  (not A167) );
 a37529a <=( (not A168)  and  a37528a );
 a37533a <=( A266  and  (not A265) );
 a37534a <=( A201  and  a37533a );
 a37535a <=( a37534a  and  a37529a );
 a37539a <=( A298  and  A268 );
 a37540a <=( (not A267)  and  a37539a );
 a37544a <=( (not A302)  and  A301 );
 a37545a <=( A299  and  a37544a );
 a37546a <=( a37545a  and  a37540a );
 a37550a <=( A199  and  (not A167) );
 a37551a <=( (not A168)  and  a37550a );
 a37555a <=( A266  and  (not A265) );
 a37556a <=( A201  and  a37555a );
 a37557a <=( a37556a  and  a37551a );
 a37561a <=( A298  and  A268 );
 a37562a <=( (not A267)  and  a37561a );
 a37566a <=( A302  and  (not A301) );
 a37567a <=( (not A299)  and  a37566a );
 a37568a <=( a37567a  and  a37562a );
 a37572a <=( A199  and  (not A167) );
 a37573a <=( (not A168)  and  a37572a );
 a37577a <=( A266  and  (not A265) );
 a37578a <=( A201  and  a37577a );
 a37579a <=( a37578a  and  a37573a );
 a37583a <=( (not A298)  and  A268 );
 a37584a <=( (not A267)  and  a37583a );
 a37588a <=( A302  and  (not A301) );
 a37589a <=( A299  and  a37588a );
 a37590a <=( a37589a  and  a37584a );
 a37594a <=( A199  and  (not A167) );
 a37595a <=( (not A168)  and  a37594a );
 a37599a <=( A266  and  (not A265) );
 a37600a <=( A201  and  a37599a );
 a37601a <=( a37600a  and  a37595a );
 a37605a <=( (not A298)  and  A268 );
 a37606a <=( (not A267)  and  a37605a );
 a37610a <=( (not A302)  and  A301 );
 a37611a <=( (not A299)  and  a37610a );
 a37612a <=( a37611a  and  a37606a );
 a37616a <=( A199  and  (not A167) );
 a37617a <=( (not A168)  and  a37616a );
 a37621a <=( A266  and  (not A265) );
 a37622a <=( A201  and  a37621a );
 a37623a <=( a37622a  and  a37617a );
 a37627a <=( A298  and  (not A269) );
 a37628a <=( (not A267)  and  a37627a );
 a37632a <=( (not A302)  and  A301 );
 a37633a <=( A299  and  a37632a );
 a37634a <=( a37633a  and  a37628a );
 a37638a <=( A199  and  (not A167) );
 a37639a <=( (not A168)  and  a37638a );
 a37643a <=( A266  and  (not A265) );
 a37644a <=( A201  and  a37643a );
 a37645a <=( a37644a  and  a37639a );
 a37649a <=( A298  and  (not A269) );
 a37650a <=( (not A267)  and  a37649a );
 a37654a <=( A302  and  (not A301) );
 a37655a <=( (not A299)  and  a37654a );
 a37656a <=( a37655a  and  a37650a );
 a37660a <=( A199  and  (not A167) );
 a37661a <=( (not A168)  and  a37660a );
 a37665a <=( A266  and  (not A265) );
 a37666a <=( A201  and  a37665a );
 a37667a <=( a37666a  and  a37661a );
 a37671a <=( (not A298)  and  (not A269) );
 a37672a <=( (not A267)  and  a37671a );
 a37676a <=( A302  and  (not A301) );
 a37677a <=( A299  and  a37676a );
 a37678a <=( a37677a  and  a37672a );
 a37682a <=( A199  and  (not A167) );
 a37683a <=( (not A168)  and  a37682a );
 a37687a <=( A266  and  (not A265) );
 a37688a <=( A201  and  a37687a );
 a37689a <=( a37688a  and  a37683a );
 a37693a <=( (not A298)  and  (not A269) );
 a37694a <=( (not A267)  and  a37693a );
 a37698a <=( (not A302)  and  A301 );
 a37699a <=( (not A299)  and  a37698a );
 a37700a <=( a37699a  and  a37694a );
 a37704a <=( A199  and  (not A167) );
 a37705a <=( (not A168)  and  a37704a );
 a37709a <=( (not A266)  and  A265 );
 a37710a <=( A201  and  a37709a );
 a37711a <=( a37710a  and  a37705a );
 a37715a <=( A298  and  A268 );
 a37716a <=( (not A267)  and  a37715a );
 a37720a <=( (not A302)  and  A301 );
 a37721a <=( A299  and  a37720a );
 a37722a <=( a37721a  and  a37716a );
 a37726a <=( A199  and  (not A167) );
 a37727a <=( (not A168)  and  a37726a );
 a37731a <=( (not A266)  and  A265 );
 a37732a <=( A201  and  a37731a );
 a37733a <=( a37732a  and  a37727a );
 a37737a <=( A298  and  A268 );
 a37738a <=( (not A267)  and  a37737a );
 a37742a <=( A302  and  (not A301) );
 a37743a <=( (not A299)  and  a37742a );
 a37744a <=( a37743a  and  a37738a );
 a37748a <=( A199  and  (not A167) );
 a37749a <=( (not A168)  and  a37748a );
 a37753a <=( (not A266)  and  A265 );
 a37754a <=( A201  and  a37753a );
 a37755a <=( a37754a  and  a37749a );
 a37759a <=( (not A298)  and  A268 );
 a37760a <=( (not A267)  and  a37759a );
 a37764a <=( A302  and  (not A301) );
 a37765a <=( A299  and  a37764a );
 a37766a <=( a37765a  and  a37760a );
 a37770a <=( A199  and  (not A167) );
 a37771a <=( (not A168)  and  a37770a );
 a37775a <=( (not A266)  and  A265 );
 a37776a <=( A201  and  a37775a );
 a37777a <=( a37776a  and  a37771a );
 a37781a <=( (not A298)  and  A268 );
 a37782a <=( (not A267)  and  a37781a );
 a37786a <=( (not A302)  and  A301 );
 a37787a <=( (not A299)  and  a37786a );
 a37788a <=( a37787a  and  a37782a );
 a37792a <=( A199  and  (not A167) );
 a37793a <=( (not A168)  and  a37792a );
 a37797a <=( (not A266)  and  A265 );
 a37798a <=( A201  and  a37797a );
 a37799a <=( a37798a  and  a37793a );
 a37803a <=( A298  and  (not A269) );
 a37804a <=( (not A267)  and  a37803a );
 a37808a <=( (not A302)  and  A301 );
 a37809a <=( A299  and  a37808a );
 a37810a <=( a37809a  and  a37804a );
 a37814a <=( A199  and  (not A167) );
 a37815a <=( (not A168)  and  a37814a );
 a37819a <=( (not A266)  and  A265 );
 a37820a <=( A201  and  a37819a );
 a37821a <=( a37820a  and  a37815a );
 a37825a <=( A298  and  (not A269) );
 a37826a <=( (not A267)  and  a37825a );
 a37830a <=( A302  and  (not A301) );
 a37831a <=( (not A299)  and  a37830a );
 a37832a <=( a37831a  and  a37826a );
 a37836a <=( A199  and  (not A167) );
 a37837a <=( (not A168)  and  a37836a );
 a37841a <=( (not A266)  and  A265 );
 a37842a <=( A201  and  a37841a );
 a37843a <=( a37842a  and  a37837a );
 a37847a <=( (not A298)  and  (not A269) );
 a37848a <=( (not A267)  and  a37847a );
 a37852a <=( A302  and  (not A301) );
 a37853a <=( A299  and  a37852a );
 a37854a <=( a37853a  and  a37848a );
 a37858a <=( A199  and  (not A167) );
 a37859a <=( (not A168)  and  a37858a );
 a37863a <=( (not A266)  and  A265 );
 a37864a <=( A201  and  a37863a );
 a37865a <=( a37864a  and  a37859a );
 a37869a <=( (not A298)  and  (not A269) );
 a37870a <=( (not A267)  and  a37869a );
 a37874a <=( (not A302)  and  A301 );
 a37875a <=( (not A299)  and  a37874a );
 a37876a <=( a37875a  and  a37870a );
 a37880a <=( A200  and  (not A167) );
 a37881a <=( (not A168)  and  a37880a );
 a37885a <=( A266  and  A265 );
 a37886a <=( A201  and  a37885a );
 a37887a <=( a37886a  and  a37881a );
 a37891a <=( A298  and  (not A268) );
 a37892a <=( (not A267)  and  a37891a );
 a37896a <=( (not A302)  and  A301 );
 a37897a <=( A299  and  a37896a );
 a37898a <=( a37897a  and  a37892a );
 a37902a <=( A200  and  (not A167) );
 a37903a <=( (not A168)  and  a37902a );
 a37907a <=( A266  and  A265 );
 a37908a <=( A201  and  a37907a );
 a37909a <=( a37908a  and  a37903a );
 a37913a <=( A298  and  (not A268) );
 a37914a <=( (not A267)  and  a37913a );
 a37918a <=( A302  and  (not A301) );
 a37919a <=( (not A299)  and  a37918a );
 a37920a <=( a37919a  and  a37914a );
 a37924a <=( A200  and  (not A167) );
 a37925a <=( (not A168)  and  a37924a );
 a37929a <=( A266  and  A265 );
 a37930a <=( A201  and  a37929a );
 a37931a <=( a37930a  and  a37925a );
 a37935a <=( (not A298)  and  (not A268) );
 a37936a <=( (not A267)  and  a37935a );
 a37940a <=( A302  and  (not A301) );
 a37941a <=( A299  and  a37940a );
 a37942a <=( a37941a  and  a37936a );
 a37946a <=( A200  and  (not A167) );
 a37947a <=( (not A168)  and  a37946a );
 a37951a <=( A266  and  A265 );
 a37952a <=( A201  and  a37951a );
 a37953a <=( a37952a  and  a37947a );
 a37957a <=( (not A298)  and  (not A268) );
 a37958a <=( (not A267)  and  a37957a );
 a37962a <=( (not A302)  and  A301 );
 a37963a <=( (not A299)  and  a37962a );
 a37964a <=( a37963a  and  a37958a );
 a37968a <=( A200  and  (not A167) );
 a37969a <=( (not A168)  and  a37968a );
 a37973a <=( A266  and  A265 );
 a37974a <=( A201  and  a37973a );
 a37975a <=( a37974a  and  a37969a );
 a37979a <=( A298  and  A269 );
 a37980a <=( (not A267)  and  a37979a );
 a37984a <=( (not A302)  and  A301 );
 a37985a <=( A299  and  a37984a );
 a37986a <=( a37985a  and  a37980a );
 a37990a <=( A200  and  (not A167) );
 a37991a <=( (not A168)  and  a37990a );
 a37995a <=( A266  and  A265 );
 a37996a <=( A201  and  a37995a );
 a37997a <=( a37996a  and  a37991a );
 a38001a <=( A298  and  A269 );
 a38002a <=( (not A267)  and  a38001a );
 a38006a <=( A302  and  (not A301) );
 a38007a <=( (not A299)  and  a38006a );
 a38008a <=( a38007a  and  a38002a );
 a38012a <=( A200  and  (not A167) );
 a38013a <=( (not A168)  and  a38012a );
 a38017a <=( A266  and  A265 );
 a38018a <=( A201  and  a38017a );
 a38019a <=( a38018a  and  a38013a );
 a38023a <=( (not A298)  and  A269 );
 a38024a <=( (not A267)  and  a38023a );
 a38028a <=( A302  and  (not A301) );
 a38029a <=( A299  and  a38028a );
 a38030a <=( a38029a  and  a38024a );
 a38034a <=( A200  and  (not A167) );
 a38035a <=( (not A168)  and  a38034a );
 a38039a <=( A266  and  A265 );
 a38040a <=( A201  and  a38039a );
 a38041a <=( a38040a  and  a38035a );
 a38045a <=( (not A298)  and  A269 );
 a38046a <=( (not A267)  and  a38045a );
 a38050a <=( (not A302)  and  A301 );
 a38051a <=( (not A299)  and  a38050a );
 a38052a <=( a38051a  and  a38046a );
 a38056a <=( A200  and  (not A167) );
 a38057a <=( (not A168)  and  a38056a );
 a38061a <=( A266  and  (not A265) );
 a38062a <=( A201  and  a38061a );
 a38063a <=( a38062a  and  a38057a );
 a38067a <=( A298  and  A268 );
 a38068a <=( (not A267)  and  a38067a );
 a38072a <=( (not A302)  and  A301 );
 a38073a <=( A299  and  a38072a );
 a38074a <=( a38073a  and  a38068a );
 a38078a <=( A200  and  (not A167) );
 a38079a <=( (not A168)  and  a38078a );
 a38083a <=( A266  and  (not A265) );
 a38084a <=( A201  and  a38083a );
 a38085a <=( a38084a  and  a38079a );
 a38089a <=( A298  and  A268 );
 a38090a <=( (not A267)  and  a38089a );
 a38094a <=( A302  and  (not A301) );
 a38095a <=( (not A299)  and  a38094a );
 a38096a <=( a38095a  and  a38090a );
 a38100a <=( A200  and  (not A167) );
 a38101a <=( (not A168)  and  a38100a );
 a38105a <=( A266  and  (not A265) );
 a38106a <=( A201  and  a38105a );
 a38107a <=( a38106a  and  a38101a );
 a38111a <=( (not A298)  and  A268 );
 a38112a <=( (not A267)  and  a38111a );
 a38116a <=( A302  and  (not A301) );
 a38117a <=( A299  and  a38116a );
 a38118a <=( a38117a  and  a38112a );
 a38122a <=( A200  and  (not A167) );
 a38123a <=( (not A168)  and  a38122a );
 a38127a <=( A266  and  (not A265) );
 a38128a <=( A201  and  a38127a );
 a38129a <=( a38128a  and  a38123a );
 a38133a <=( (not A298)  and  A268 );
 a38134a <=( (not A267)  and  a38133a );
 a38138a <=( (not A302)  and  A301 );
 a38139a <=( (not A299)  and  a38138a );
 a38140a <=( a38139a  and  a38134a );
 a38144a <=( A200  and  (not A167) );
 a38145a <=( (not A168)  and  a38144a );
 a38149a <=( A266  and  (not A265) );
 a38150a <=( A201  and  a38149a );
 a38151a <=( a38150a  and  a38145a );
 a38155a <=( A298  and  (not A269) );
 a38156a <=( (not A267)  and  a38155a );
 a38160a <=( (not A302)  and  A301 );
 a38161a <=( A299  and  a38160a );
 a38162a <=( a38161a  and  a38156a );
 a38166a <=( A200  and  (not A167) );
 a38167a <=( (not A168)  and  a38166a );
 a38171a <=( A266  and  (not A265) );
 a38172a <=( A201  and  a38171a );
 a38173a <=( a38172a  and  a38167a );
 a38177a <=( A298  and  (not A269) );
 a38178a <=( (not A267)  and  a38177a );
 a38182a <=( A302  and  (not A301) );
 a38183a <=( (not A299)  and  a38182a );
 a38184a <=( a38183a  and  a38178a );
 a38188a <=( A200  and  (not A167) );
 a38189a <=( (not A168)  and  a38188a );
 a38193a <=( A266  and  (not A265) );
 a38194a <=( A201  and  a38193a );
 a38195a <=( a38194a  and  a38189a );
 a38199a <=( (not A298)  and  (not A269) );
 a38200a <=( (not A267)  and  a38199a );
 a38204a <=( A302  and  (not A301) );
 a38205a <=( A299  and  a38204a );
 a38206a <=( a38205a  and  a38200a );
 a38210a <=( A200  and  (not A167) );
 a38211a <=( (not A168)  and  a38210a );
 a38215a <=( A266  and  (not A265) );
 a38216a <=( A201  and  a38215a );
 a38217a <=( a38216a  and  a38211a );
 a38221a <=( (not A298)  and  (not A269) );
 a38222a <=( (not A267)  and  a38221a );
 a38226a <=( (not A302)  and  A301 );
 a38227a <=( (not A299)  and  a38226a );
 a38228a <=( a38227a  and  a38222a );
 a38232a <=( A200  and  (not A167) );
 a38233a <=( (not A168)  and  a38232a );
 a38237a <=( (not A266)  and  A265 );
 a38238a <=( A201  and  a38237a );
 a38239a <=( a38238a  and  a38233a );
 a38243a <=( A298  and  A268 );
 a38244a <=( (not A267)  and  a38243a );
 a38248a <=( (not A302)  and  A301 );
 a38249a <=( A299  and  a38248a );
 a38250a <=( a38249a  and  a38244a );
 a38254a <=( A200  and  (not A167) );
 a38255a <=( (not A168)  and  a38254a );
 a38259a <=( (not A266)  and  A265 );
 a38260a <=( A201  and  a38259a );
 a38261a <=( a38260a  and  a38255a );
 a38265a <=( A298  and  A268 );
 a38266a <=( (not A267)  and  a38265a );
 a38270a <=( A302  and  (not A301) );
 a38271a <=( (not A299)  and  a38270a );
 a38272a <=( a38271a  and  a38266a );
 a38276a <=( A200  and  (not A167) );
 a38277a <=( (not A168)  and  a38276a );
 a38281a <=( (not A266)  and  A265 );
 a38282a <=( A201  and  a38281a );
 a38283a <=( a38282a  and  a38277a );
 a38287a <=( (not A298)  and  A268 );
 a38288a <=( (not A267)  and  a38287a );
 a38292a <=( A302  and  (not A301) );
 a38293a <=( A299  and  a38292a );
 a38294a <=( a38293a  and  a38288a );
 a38298a <=( A200  and  (not A167) );
 a38299a <=( (not A168)  and  a38298a );
 a38303a <=( (not A266)  and  A265 );
 a38304a <=( A201  and  a38303a );
 a38305a <=( a38304a  and  a38299a );
 a38309a <=( (not A298)  and  A268 );
 a38310a <=( (not A267)  and  a38309a );
 a38314a <=( (not A302)  and  A301 );
 a38315a <=( (not A299)  and  a38314a );
 a38316a <=( a38315a  and  a38310a );
 a38320a <=( A200  and  (not A167) );
 a38321a <=( (not A168)  and  a38320a );
 a38325a <=( (not A266)  and  A265 );
 a38326a <=( A201  and  a38325a );
 a38327a <=( a38326a  and  a38321a );
 a38331a <=( A298  and  (not A269) );
 a38332a <=( (not A267)  and  a38331a );
 a38336a <=( (not A302)  and  A301 );
 a38337a <=( A299  and  a38336a );
 a38338a <=( a38337a  and  a38332a );
 a38342a <=( A200  and  (not A167) );
 a38343a <=( (not A168)  and  a38342a );
 a38347a <=( (not A266)  and  A265 );
 a38348a <=( A201  and  a38347a );
 a38349a <=( a38348a  and  a38343a );
 a38353a <=( A298  and  (not A269) );
 a38354a <=( (not A267)  and  a38353a );
 a38358a <=( A302  and  (not A301) );
 a38359a <=( (not A299)  and  a38358a );
 a38360a <=( a38359a  and  a38354a );
 a38364a <=( A200  and  (not A167) );
 a38365a <=( (not A168)  and  a38364a );
 a38369a <=( (not A266)  and  A265 );
 a38370a <=( A201  and  a38369a );
 a38371a <=( a38370a  and  a38365a );
 a38375a <=( (not A298)  and  (not A269) );
 a38376a <=( (not A267)  and  a38375a );
 a38380a <=( A302  and  (not A301) );
 a38381a <=( A299  and  a38380a );
 a38382a <=( a38381a  and  a38376a );
 a38386a <=( A200  and  (not A167) );
 a38387a <=( (not A168)  and  a38386a );
 a38391a <=( (not A266)  and  A265 );
 a38392a <=( A201  and  a38391a );
 a38393a <=( a38392a  and  a38387a );
 a38397a <=( (not A298)  and  (not A269) );
 a38398a <=( (not A267)  and  a38397a );
 a38402a <=( (not A302)  and  A301 );
 a38403a <=( (not A299)  and  a38402a );
 a38404a <=( a38403a  and  a38398a );
 a38408a <=( A199  and  (not A167) );
 a38409a <=( (not A168)  and  a38408a );
 a38413a <=( (not A203)  and  A202 );
 a38414a <=( A200  and  a38413a );
 a38415a <=( a38414a  and  a38409a );
 a38419a <=( (not A267)  and  A266 );
 a38420a <=( A265  and  a38419a );
 a38424a <=( A300  and  A299 );
 a38425a <=( (not A268)  and  a38424a );
 a38426a <=( a38425a  and  a38420a );
 a38430a <=( A199  and  (not A167) );
 a38431a <=( (not A168)  and  a38430a );
 a38435a <=( (not A203)  and  A202 );
 a38436a <=( A200  and  a38435a );
 a38437a <=( a38436a  and  a38431a );
 a38441a <=( (not A267)  and  A266 );
 a38442a <=( A265  and  a38441a );
 a38446a <=( A300  and  A298 );
 a38447a <=( (not A268)  and  a38446a );
 a38448a <=( a38447a  and  a38442a );
 a38452a <=( A199  and  (not A167) );
 a38453a <=( (not A168)  and  a38452a );
 a38457a <=( (not A203)  and  A202 );
 a38458a <=( A200  and  a38457a );
 a38459a <=( a38458a  and  a38453a );
 a38463a <=( (not A267)  and  A266 );
 a38464a <=( A265  and  a38463a );
 a38468a <=( A300  and  A299 );
 a38469a <=( A269  and  a38468a );
 a38470a <=( a38469a  and  a38464a );
 a38474a <=( A199  and  (not A167) );
 a38475a <=( (not A168)  and  a38474a );
 a38479a <=( (not A203)  and  A202 );
 a38480a <=( A200  and  a38479a );
 a38481a <=( a38480a  and  a38475a );
 a38485a <=( (not A267)  and  A266 );
 a38486a <=( A265  and  a38485a );
 a38490a <=( A300  and  A298 );
 a38491a <=( A269  and  a38490a );
 a38492a <=( a38491a  and  a38486a );
 a38496a <=( A199  and  (not A167) );
 a38497a <=( (not A168)  and  a38496a );
 a38501a <=( (not A203)  and  A202 );
 a38502a <=( A200  and  a38501a );
 a38503a <=( a38502a  and  a38497a );
 a38507a <=( (not A267)  and  A266 );
 a38508a <=( (not A265)  and  a38507a );
 a38512a <=( A300  and  A299 );
 a38513a <=( A268  and  a38512a );
 a38514a <=( a38513a  and  a38508a );
 a38518a <=( A199  and  (not A167) );
 a38519a <=( (not A168)  and  a38518a );
 a38523a <=( (not A203)  and  A202 );
 a38524a <=( A200  and  a38523a );
 a38525a <=( a38524a  and  a38519a );
 a38529a <=( (not A267)  and  A266 );
 a38530a <=( (not A265)  and  a38529a );
 a38534a <=( A300  and  A298 );
 a38535a <=( A268  and  a38534a );
 a38536a <=( a38535a  and  a38530a );
 a38540a <=( A199  and  (not A167) );
 a38541a <=( (not A168)  and  a38540a );
 a38545a <=( (not A203)  and  A202 );
 a38546a <=( A200  and  a38545a );
 a38547a <=( a38546a  and  a38541a );
 a38551a <=( (not A267)  and  A266 );
 a38552a <=( (not A265)  and  a38551a );
 a38556a <=( A300  and  A299 );
 a38557a <=( (not A269)  and  a38556a );
 a38558a <=( a38557a  and  a38552a );
 a38562a <=( A199  and  (not A167) );
 a38563a <=( (not A168)  and  a38562a );
 a38567a <=( (not A203)  and  A202 );
 a38568a <=( A200  and  a38567a );
 a38569a <=( a38568a  and  a38563a );
 a38573a <=( (not A267)  and  A266 );
 a38574a <=( (not A265)  and  a38573a );
 a38578a <=( A300  and  A298 );
 a38579a <=( (not A269)  and  a38578a );
 a38580a <=( a38579a  and  a38574a );
 a38584a <=( A199  and  (not A167) );
 a38585a <=( (not A168)  and  a38584a );
 a38589a <=( (not A203)  and  A202 );
 a38590a <=( A200  and  a38589a );
 a38591a <=( a38590a  and  a38585a );
 a38595a <=( (not A267)  and  (not A266) );
 a38596a <=( A265  and  a38595a );
 a38600a <=( A300  and  A299 );
 a38601a <=( A268  and  a38600a );
 a38602a <=( a38601a  and  a38596a );
 a38606a <=( A199  and  (not A167) );
 a38607a <=( (not A168)  and  a38606a );
 a38611a <=( (not A203)  and  A202 );
 a38612a <=( A200  and  a38611a );
 a38613a <=( a38612a  and  a38607a );
 a38617a <=( (not A267)  and  (not A266) );
 a38618a <=( A265  and  a38617a );
 a38622a <=( A300  and  A298 );
 a38623a <=( A268  and  a38622a );
 a38624a <=( a38623a  and  a38618a );
 a38628a <=( A199  and  (not A167) );
 a38629a <=( (not A168)  and  a38628a );
 a38633a <=( (not A203)  and  A202 );
 a38634a <=( A200  and  a38633a );
 a38635a <=( a38634a  and  a38629a );
 a38639a <=( (not A267)  and  (not A266) );
 a38640a <=( A265  and  a38639a );
 a38644a <=( A300  and  A299 );
 a38645a <=( (not A269)  and  a38644a );
 a38646a <=( a38645a  and  a38640a );
 a38650a <=( A199  and  (not A167) );
 a38651a <=( (not A168)  and  a38650a );
 a38655a <=( (not A203)  and  A202 );
 a38656a <=( A200  and  a38655a );
 a38657a <=( a38656a  and  a38651a );
 a38661a <=( (not A267)  and  (not A266) );
 a38662a <=( A265  and  a38661a );
 a38666a <=( A300  and  A298 );
 a38667a <=( (not A269)  and  a38666a );
 a38668a <=( a38667a  and  a38662a );
 a38672a <=( A199  and  (not A167) );
 a38673a <=( (not A168)  and  a38672a );
 a38677a <=( (not A202)  and  (not A201) );
 a38678a <=( A200  and  a38677a );
 a38679a <=( a38678a  and  a38673a );
 a38683a <=( A298  and  A267 );
 a38684a <=( A265  and  a38683a );
 a38688a <=( (not A301)  and  (not A300) );
 a38689a <=( A299  and  a38688a );
 a38690a <=( a38689a  and  a38684a );
 a38694a <=( A199  and  (not A167) );
 a38695a <=( (not A168)  and  a38694a );
 a38699a <=( (not A202)  and  (not A201) );
 a38700a <=( A200  and  a38699a );
 a38701a <=( a38700a  and  a38695a );
 a38705a <=( A298  and  A267 );
 a38706a <=( A265  and  a38705a );
 a38710a <=( A302  and  (not A300) );
 a38711a <=( A299  and  a38710a );
 a38712a <=( a38711a  and  a38706a );
 a38716a <=( A199  and  (not A167) );
 a38717a <=( (not A168)  and  a38716a );
 a38721a <=( (not A202)  and  (not A201) );
 a38722a <=( A200  and  a38721a );
 a38723a <=( a38722a  and  a38717a );
 a38727a <=( A298  and  A267 );
 a38728a <=( A265  and  a38727a );
 a38732a <=( A301  and  (not A300) );
 a38733a <=( (not A299)  and  a38732a );
 a38734a <=( a38733a  and  a38728a );
 a38738a <=( A199  and  (not A167) );
 a38739a <=( (not A168)  and  a38738a );
 a38743a <=( (not A202)  and  (not A201) );
 a38744a <=( A200  and  a38743a );
 a38745a <=( a38744a  and  a38739a );
 a38749a <=( A298  and  A267 );
 a38750a <=( A265  and  a38749a );
 a38754a <=( (not A302)  and  (not A300) );
 a38755a <=( (not A299)  and  a38754a );
 a38756a <=( a38755a  and  a38750a );
 a38760a <=( A199  and  (not A167) );
 a38761a <=( (not A168)  and  a38760a );
 a38765a <=( (not A202)  and  (not A201) );
 a38766a <=( A200  and  a38765a );
 a38767a <=( a38766a  and  a38761a );
 a38771a <=( (not A298)  and  A267 );
 a38772a <=( A265  and  a38771a );
 a38776a <=( A301  and  (not A300) );
 a38777a <=( A299  and  a38776a );
 a38778a <=( a38777a  and  a38772a );
 a38782a <=( A199  and  (not A167) );
 a38783a <=( (not A168)  and  a38782a );
 a38787a <=( (not A202)  and  (not A201) );
 a38788a <=( A200  and  a38787a );
 a38789a <=( a38788a  and  a38783a );
 a38793a <=( (not A298)  and  A267 );
 a38794a <=( A265  and  a38793a );
 a38798a <=( (not A302)  and  (not A300) );
 a38799a <=( A299  and  a38798a );
 a38800a <=( a38799a  and  a38794a );
 a38804a <=( A199  and  (not A167) );
 a38805a <=( (not A168)  and  a38804a );
 a38809a <=( (not A202)  and  (not A201) );
 a38810a <=( A200  and  a38809a );
 a38811a <=( a38810a  and  a38805a );
 a38815a <=( A298  and  A267 );
 a38816a <=( A266  and  a38815a );
 a38820a <=( (not A301)  and  (not A300) );
 a38821a <=( A299  and  a38820a );
 a38822a <=( a38821a  and  a38816a );
 a38826a <=( A199  and  (not A167) );
 a38827a <=( (not A168)  and  a38826a );
 a38831a <=( (not A202)  and  (not A201) );
 a38832a <=( A200  and  a38831a );
 a38833a <=( a38832a  and  a38827a );
 a38837a <=( A298  and  A267 );
 a38838a <=( A266  and  a38837a );
 a38842a <=( A302  and  (not A300) );
 a38843a <=( A299  and  a38842a );
 a38844a <=( a38843a  and  a38838a );
 a38848a <=( A199  and  (not A167) );
 a38849a <=( (not A168)  and  a38848a );
 a38853a <=( (not A202)  and  (not A201) );
 a38854a <=( A200  and  a38853a );
 a38855a <=( a38854a  and  a38849a );
 a38859a <=( A298  and  A267 );
 a38860a <=( A266  and  a38859a );
 a38864a <=( A301  and  (not A300) );
 a38865a <=( (not A299)  and  a38864a );
 a38866a <=( a38865a  and  a38860a );
 a38870a <=( A199  and  (not A167) );
 a38871a <=( (not A168)  and  a38870a );
 a38875a <=( (not A202)  and  (not A201) );
 a38876a <=( A200  and  a38875a );
 a38877a <=( a38876a  and  a38871a );
 a38881a <=( A298  and  A267 );
 a38882a <=( A266  and  a38881a );
 a38886a <=( (not A302)  and  (not A300) );
 a38887a <=( (not A299)  and  a38886a );
 a38888a <=( a38887a  and  a38882a );
 a38892a <=( A199  and  (not A167) );
 a38893a <=( (not A168)  and  a38892a );
 a38897a <=( (not A202)  and  (not A201) );
 a38898a <=( A200  and  a38897a );
 a38899a <=( a38898a  and  a38893a );
 a38903a <=( (not A298)  and  A267 );
 a38904a <=( A266  and  a38903a );
 a38908a <=( A301  and  (not A300) );
 a38909a <=( A299  and  a38908a );
 a38910a <=( a38909a  and  a38904a );
 a38914a <=( A199  and  (not A167) );
 a38915a <=( (not A168)  and  a38914a );
 a38919a <=( (not A202)  and  (not A201) );
 a38920a <=( A200  and  a38919a );
 a38921a <=( a38920a  and  a38915a );
 a38925a <=( (not A298)  and  A267 );
 a38926a <=( A266  and  a38925a );
 a38930a <=( (not A302)  and  (not A300) );
 a38931a <=( A299  and  a38930a );
 a38932a <=( a38931a  and  a38926a );
 a38936a <=( A199  and  (not A167) );
 a38937a <=( (not A168)  and  a38936a );
 a38941a <=( A203  and  (not A201) );
 a38942a <=( A200  and  a38941a );
 a38943a <=( a38942a  and  a38937a );
 a38947a <=( A298  and  A267 );
 a38948a <=( A265  and  a38947a );
 a38952a <=( (not A301)  and  (not A300) );
 a38953a <=( A299  and  a38952a );
 a38954a <=( a38953a  and  a38948a );
 a38958a <=( A199  and  (not A167) );
 a38959a <=( (not A168)  and  a38958a );
 a38963a <=( A203  and  (not A201) );
 a38964a <=( A200  and  a38963a );
 a38965a <=( a38964a  and  a38959a );
 a38969a <=( A298  and  A267 );
 a38970a <=( A265  and  a38969a );
 a38974a <=( A302  and  (not A300) );
 a38975a <=( A299  and  a38974a );
 a38976a <=( a38975a  and  a38970a );
 a38980a <=( A199  and  (not A167) );
 a38981a <=( (not A168)  and  a38980a );
 a38985a <=( A203  and  (not A201) );
 a38986a <=( A200  and  a38985a );
 a38987a <=( a38986a  and  a38981a );
 a38991a <=( A298  and  A267 );
 a38992a <=( A265  and  a38991a );
 a38996a <=( A301  and  (not A300) );
 a38997a <=( (not A299)  and  a38996a );
 a38998a <=( a38997a  and  a38992a );
 a39002a <=( A199  and  (not A167) );
 a39003a <=( (not A168)  and  a39002a );
 a39007a <=( A203  and  (not A201) );
 a39008a <=( A200  and  a39007a );
 a39009a <=( a39008a  and  a39003a );
 a39013a <=( A298  and  A267 );
 a39014a <=( A265  and  a39013a );
 a39018a <=( (not A302)  and  (not A300) );
 a39019a <=( (not A299)  and  a39018a );
 a39020a <=( a39019a  and  a39014a );
 a39024a <=( A199  and  (not A167) );
 a39025a <=( (not A168)  and  a39024a );
 a39029a <=( A203  and  (not A201) );
 a39030a <=( A200  and  a39029a );
 a39031a <=( a39030a  and  a39025a );
 a39035a <=( (not A298)  and  A267 );
 a39036a <=( A265  and  a39035a );
 a39040a <=( A301  and  (not A300) );
 a39041a <=( A299  and  a39040a );
 a39042a <=( a39041a  and  a39036a );
 a39046a <=( A199  and  (not A167) );
 a39047a <=( (not A168)  and  a39046a );
 a39051a <=( A203  and  (not A201) );
 a39052a <=( A200  and  a39051a );
 a39053a <=( a39052a  and  a39047a );
 a39057a <=( (not A298)  and  A267 );
 a39058a <=( A265  and  a39057a );
 a39062a <=( (not A302)  and  (not A300) );
 a39063a <=( A299  and  a39062a );
 a39064a <=( a39063a  and  a39058a );
 a39068a <=( A199  and  (not A167) );
 a39069a <=( (not A168)  and  a39068a );
 a39073a <=( A203  and  (not A201) );
 a39074a <=( A200  and  a39073a );
 a39075a <=( a39074a  and  a39069a );
 a39079a <=( A298  and  A267 );
 a39080a <=( A266  and  a39079a );
 a39084a <=( (not A301)  and  (not A300) );
 a39085a <=( A299  and  a39084a );
 a39086a <=( a39085a  and  a39080a );
 a39090a <=( A199  and  (not A167) );
 a39091a <=( (not A168)  and  a39090a );
 a39095a <=( A203  and  (not A201) );
 a39096a <=( A200  and  a39095a );
 a39097a <=( a39096a  and  a39091a );
 a39101a <=( A298  and  A267 );
 a39102a <=( A266  and  a39101a );
 a39106a <=( A302  and  (not A300) );
 a39107a <=( A299  and  a39106a );
 a39108a <=( a39107a  and  a39102a );
 a39112a <=( A199  and  (not A167) );
 a39113a <=( (not A168)  and  a39112a );
 a39117a <=( A203  and  (not A201) );
 a39118a <=( A200  and  a39117a );
 a39119a <=( a39118a  and  a39113a );
 a39123a <=( A298  and  A267 );
 a39124a <=( A266  and  a39123a );
 a39128a <=( A301  and  (not A300) );
 a39129a <=( (not A299)  and  a39128a );
 a39130a <=( a39129a  and  a39124a );
 a39134a <=( A199  and  (not A167) );
 a39135a <=( (not A168)  and  a39134a );
 a39139a <=( A203  and  (not A201) );
 a39140a <=( A200  and  a39139a );
 a39141a <=( a39140a  and  a39135a );
 a39145a <=( A298  and  A267 );
 a39146a <=( A266  and  a39145a );
 a39150a <=( (not A302)  and  (not A300) );
 a39151a <=( (not A299)  and  a39150a );
 a39152a <=( a39151a  and  a39146a );
 a39156a <=( A199  and  (not A167) );
 a39157a <=( (not A168)  and  a39156a );
 a39161a <=( A203  and  (not A201) );
 a39162a <=( A200  and  a39161a );
 a39163a <=( a39162a  and  a39157a );
 a39167a <=( (not A298)  and  A267 );
 a39168a <=( A266  and  a39167a );
 a39172a <=( A301  and  (not A300) );
 a39173a <=( A299  and  a39172a );
 a39174a <=( a39173a  and  a39168a );
 a39178a <=( A199  and  (not A167) );
 a39179a <=( (not A168)  and  a39178a );
 a39183a <=( A203  and  (not A201) );
 a39184a <=( A200  and  a39183a );
 a39185a <=( a39184a  and  a39179a );
 a39189a <=( (not A298)  and  A267 );
 a39190a <=( A266  and  a39189a );
 a39194a <=( (not A302)  and  (not A300) );
 a39195a <=( A299  and  a39194a );
 a39196a <=( a39195a  and  a39190a );
 a39200a <=( (not A199)  and  (not A167) );
 a39201a <=( (not A168)  and  a39200a );
 a39205a <=( A203  and  (not A202) );
 a39206a <=( A200  and  a39205a );
 a39207a <=( a39206a  and  a39201a );
 a39211a <=( (not A267)  and  A266 );
 a39212a <=( A265  and  a39211a );
 a39216a <=( A300  and  A299 );
 a39217a <=( (not A268)  and  a39216a );
 a39218a <=( a39217a  and  a39212a );
 a39222a <=( (not A199)  and  (not A167) );
 a39223a <=( (not A168)  and  a39222a );
 a39227a <=( A203  and  (not A202) );
 a39228a <=( A200  and  a39227a );
 a39229a <=( a39228a  and  a39223a );
 a39233a <=( (not A267)  and  A266 );
 a39234a <=( A265  and  a39233a );
 a39238a <=( A300  and  A298 );
 a39239a <=( (not A268)  and  a39238a );
 a39240a <=( a39239a  and  a39234a );
 a39244a <=( (not A199)  and  (not A167) );
 a39245a <=( (not A168)  and  a39244a );
 a39249a <=( A203  and  (not A202) );
 a39250a <=( A200  and  a39249a );
 a39251a <=( a39250a  and  a39245a );
 a39255a <=( (not A267)  and  A266 );
 a39256a <=( A265  and  a39255a );
 a39260a <=( A300  and  A299 );
 a39261a <=( A269  and  a39260a );
 a39262a <=( a39261a  and  a39256a );
 a39266a <=( (not A199)  and  (not A167) );
 a39267a <=( (not A168)  and  a39266a );
 a39271a <=( A203  and  (not A202) );
 a39272a <=( A200  and  a39271a );
 a39273a <=( a39272a  and  a39267a );
 a39277a <=( (not A267)  and  A266 );
 a39278a <=( A265  and  a39277a );
 a39282a <=( A300  and  A298 );
 a39283a <=( A269  and  a39282a );
 a39284a <=( a39283a  and  a39278a );
 a39288a <=( (not A199)  and  (not A167) );
 a39289a <=( (not A168)  and  a39288a );
 a39293a <=( A203  and  (not A202) );
 a39294a <=( A200  and  a39293a );
 a39295a <=( a39294a  and  a39289a );
 a39299a <=( (not A267)  and  A266 );
 a39300a <=( (not A265)  and  a39299a );
 a39304a <=( A300  and  A299 );
 a39305a <=( A268  and  a39304a );
 a39306a <=( a39305a  and  a39300a );
 a39310a <=( (not A199)  and  (not A167) );
 a39311a <=( (not A168)  and  a39310a );
 a39315a <=( A203  and  (not A202) );
 a39316a <=( A200  and  a39315a );
 a39317a <=( a39316a  and  a39311a );
 a39321a <=( (not A267)  and  A266 );
 a39322a <=( (not A265)  and  a39321a );
 a39326a <=( A300  and  A298 );
 a39327a <=( A268  and  a39326a );
 a39328a <=( a39327a  and  a39322a );
 a39332a <=( (not A199)  and  (not A167) );
 a39333a <=( (not A168)  and  a39332a );
 a39337a <=( A203  and  (not A202) );
 a39338a <=( A200  and  a39337a );
 a39339a <=( a39338a  and  a39333a );
 a39343a <=( (not A267)  and  A266 );
 a39344a <=( (not A265)  and  a39343a );
 a39348a <=( A300  and  A299 );
 a39349a <=( (not A269)  and  a39348a );
 a39350a <=( a39349a  and  a39344a );
 a39354a <=( (not A199)  and  (not A167) );
 a39355a <=( (not A168)  and  a39354a );
 a39359a <=( A203  and  (not A202) );
 a39360a <=( A200  and  a39359a );
 a39361a <=( a39360a  and  a39355a );
 a39365a <=( (not A267)  and  A266 );
 a39366a <=( (not A265)  and  a39365a );
 a39370a <=( A300  and  A298 );
 a39371a <=( (not A269)  and  a39370a );
 a39372a <=( a39371a  and  a39366a );
 a39376a <=( (not A199)  and  (not A167) );
 a39377a <=( (not A168)  and  a39376a );
 a39381a <=( A203  and  (not A202) );
 a39382a <=( A200  and  a39381a );
 a39383a <=( a39382a  and  a39377a );
 a39387a <=( (not A267)  and  (not A266) );
 a39388a <=( A265  and  a39387a );
 a39392a <=( A300  and  A299 );
 a39393a <=( A268  and  a39392a );
 a39394a <=( a39393a  and  a39388a );
 a39398a <=( (not A199)  and  (not A167) );
 a39399a <=( (not A168)  and  a39398a );
 a39403a <=( A203  and  (not A202) );
 a39404a <=( A200  and  a39403a );
 a39405a <=( a39404a  and  a39399a );
 a39409a <=( (not A267)  and  (not A266) );
 a39410a <=( A265  and  a39409a );
 a39414a <=( A300  and  A298 );
 a39415a <=( A268  and  a39414a );
 a39416a <=( a39415a  and  a39410a );
 a39420a <=( (not A199)  and  (not A167) );
 a39421a <=( (not A168)  and  a39420a );
 a39425a <=( A203  and  (not A202) );
 a39426a <=( A200  and  a39425a );
 a39427a <=( a39426a  and  a39421a );
 a39431a <=( (not A267)  and  (not A266) );
 a39432a <=( A265  and  a39431a );
 a39436a <=( A300  and  A299 );
 a39437a <=( (not A269)  and  a39436a );
 a39438a <=( a39437a  and  a39432a );
 a39442a <=( (not A199)  and  (not A167) );
 a39443a <=( (not A168)  and  a39442a );
 a39447a <=( A203  and  (not A202) );
 a39448a <=( A200  and  a39447a );
 a39449a <=( a39448a  and  a39443a );
 a39453a <=( (not A267)  and  (not A266) );
 a39454a <=( A265  and  a39453a );
 a39458a <=( A300  and  A298 );
 a39459a <=( (not A269)  and  a39458a );
 a39460a <=( a39459a  and  a39454a );
 a39464a <=( (not A199)  and  (not A167) );
 a39465a <=( (not A168)  and  a39464a );
 a39469a <=( A202  and  (not A201) );
 a39470a <=( A200  and  a39469a );
 a39471a <=( a39470a  and  a39465a );
 a39475a <=( A298  and  A267 );
 a39476a <=( A265  and  a39475a );
 a39480a <=( (not A301)  and  (not A300) );
 a39481a <=( A299  and  a39480a );
 a39482a <=( a39481a  and  a39476a );
 a39486a <=( (not A199)  and  (not A167) );
 a39487a <=( (not A168)  and  a39486a );
 a39491a <=( A202  and  (not A201) );
 a39492a <=( A200  and  a39491a );
 a39493a <=( a39492a  and  a39487a );
 a39497a <=( A298  and  A267 );
 a39498a <=( A265  and  a39497a );
 a39502a <=( A302  and  (not A300) );
 a39503a <=( A299  and  a39502a );
 a39504a <=( a39503a  and  a39498a );
 a39508a <=( (not A199)  and  (not A167) );
 a39509a <=( (not A168)  and  a39508a );
 a39513a <=( A202  and  (not A201) );
 a39514a <=( A200  and  a39513a );
 a39515a <=( a39514a  and  a39509a );
 a39519a <=( A298  and  A267 );
 a39520a <=( A265  and  a39519a );
 a39524a <=( A301  and  (not A300) );
 a39525a <=( (not A299)  and  a39524a );
 a39526a <=( a39525a  and  a39520a );
 a39530a <=( (not A199)  and  (not A167) );
 a39531a <=( (not A168)  and  a39530a );
 a39535a <=( A202  and  (not A201) );
 a39536a <=( A200  and  a39535a );
 a39537a <=( a39536a  and  a39531a );
 a39541a <=( A298  and  A267 );
 a39542a <=( A265  and  a39541a );
 a39546a <=( (not A302)  and  (not A300) );
 a39547a <=( (not A299)  and  a39546a );
 a39548a <=( a39547a  and  a39542a );
 a39552a <=( (not A199)  and  (not A167) );
 a39553a <=( (not A168)  and  a39552a );
 a39557a <=( A202  and  (not A201) );
 a39558a <=( A200  and  a39557a );
 a39559a <=( a39558a  and  a39553a );
 a39563a <=( (not A298)  and  A267 );
 a39564a <=( A265  and  a39563a );
 a39568a <=( A301  and  (not A300) );
 a39569a <=( A299  and  a39568a );
 a39570a <=( a39569a  and  a39564a );
 a39574a <=( (not A199)  and  (not A167) );
 a39575a <=( (not A168)  and  a39574a );
 a39579a <=( A202  and  (not A201) );
 a39580a <=( A200  and  a39579a );
 a39581a <=( a39580a  and  a39575a );
 a39585a <=( (not A298)  and  A267 );
 a39586a <=( A265  and  a39585a );
 a39590a <=( (not A302)  and  (not A300) );
 a39591a <=( A299  and  a39590a );
 a39592a <=( a39591a  and  a39586a );
 a39596a <=( (not A199)  and  (not A167) );
 a39597a <=( (not A168)  and  a39596a );
 a39601a <=( A202  and  (not A201) );
 a39602a <=( A200  and  a39601a );
 a39603a <=( a39602a  and  a39597a );
 a39607a <=( A298  and  A267 );
 a39608a <=( A266  and  a39607a );
 a39612a <=( (not A301)  and  (not A300) );
 a39613a <=( A299  and  a39612a );
 a39614a <=( a39613a  and  a39608a );
 a39618a <=( (not A199)  and  (not A167) );
 a39619a <=( (not A168)  and  a39618a );
 a39623a <=( A202  and  (not A201) );
 a39624a <=( A200  and  a39623a );
 a39625a <=( a39624a  and  a39619a );
 a39629a <=( A298  and  A267 );
 a39630a <=( A266  and  a39629a );
 a39634a <=( A302  and  (not A300) );
 a39635a <=( A299  and  a39634a );
 a39636a <=( a39635a  and  a39630a );
 a39640a <=( (not A199)  and  (not A167) );
 a39641a <=( (not A168)  and  a39640a );
 a39645a <=( A202  and  (not A201) );
 a39646a <=( A200  and  a39645a );
 a39647a <=( a39646a  and  a39641a );
 a39651a <=( A298  and  A267 );
 a39652a <=( A266  and  a39651a );
 a39656a <=( A301  and  (not A300) );
 a39657a <=( (not A299)  and  a39656a );
 a39658a <=( a39657a  and  a39652a );
 a39662a <=( (not A199)  and  (not A167) );
 a39663a <=( (not A168)  and  a39662a );
 a39667a <=( A202  and  (not A201) );
 a39668a <=( A200  and  a39667a );
 a39669a <=( a39668a  and  a39663a );
 a39673a <=( A298  and  A267 );
 a39674a <=( A266  and  a39673a );
 a39678a <=( (not A302)  and  (not A300) );
 a39679a <=( (not A299)  and  a39678a );
 a39680a <=( a39679a  and  a39674a );
 a39684a <=( (not A199)  and  (not A167) );
 a39685a <=( (not A168)  and  a39684a );
 a39689a <=( A202  and  (not A201) );
 a39690a <=( A200  and  a39689a );
 a39691a <=( a39690a  and  a39685a );
 a39695a <=( (not A298)  and  A267 );
 a39696a <=( A266  and  a39695a );
 a39700a <=( A301  and  (not A300) );
 a39701a <=( A299  and  a39700a );
 a39702a <=( a39701a  and  a39696a );
 a39706a <=( (not A199)  and  (not A167) );
 a39707a <=( (not A168)  and  a39706a );
 a39711a <=( A202  and  (not A201) );
 a39712a <=( A200  and  a39711a );
 a39713a <=( a39712a  and  a39707a );
 a39717a <=( (not A298)  and  A267 );
 a39718a <=( A266  and  a39717a );
 a39722a <=( (not A302)  and  (not A300) );
 a39723a <=( A299  and  a39722a );
 a39724a <=( a39723a  and  a39718a );
 a39728a <=( (not A199)  and  (not A167) );
 a39729a <=( (not A168)  and  a39728a );
 a39733a <=( (not A203)  and  (not A201) );
 a39734a <=( A200  and  a39733a );
 a39735a <=( a39734a  and  a39729a );
 a39739a <=( A298  and  A267 );
 a39740a <=( A265  and  a39739a );
 a39744a <=( (not A301)  and  (not A300) );
 a39745a <=( A299  and  a39744a );
 a39746a <=( a39745a  and  a39740a );
 a39750a <=( (not A199)  and  (not A167) );
 a39751a <=( (not A168)  and  a39750a );
 a39755a <=( (not A203)  and  (not A201) );
 a39756a <=( A200  and  a39755a );
 a39757a <=( a39756a  and  a39751a );
 a39761a <=( A298  and  A267 );
 a39762a <=( A265  and  a39761a );
 a39766a <=( A302  and  (not A300) );
 a39767a <=( A299  and  a39766a );
 a39768a <=( a39767a  and  a39762a );
 a39772a <=( (not A199)  and  (not A167) );
 a39773a <=( (not A168)  and  a39772a );
 a39777a <=( (not A203)  and  (not A201) );
 a39778a <=( A200  and  a39777a );
 a39779a <=( a39778a  and  a39773a );
 a39783a <=( A298  and  A267 );
 a39784a <=( A265  and  a39783a );
 a39788a <=( A301  and  (not A300) );
 a39789a <=( (not A299)  and  a39788a );
 a39790a <=( a39789a  and  a39784a );
 a39794a <=( (not A199)  and  (not A167) );
 a39795a <=( (not A168)  and  a39794a );
 a39799a <=( (not A203)  and  (not A201) );
 a39800a <=( A200  and  a39799a );
 a39801a <=( a39800a  and  a39795a );
 a39805a <=( A298  and  A267 );
 a39806a <=( A265  and  a39805a );
 a39810a <=( (not A302)  and  (not A300) );
 a39811a <=( (not A299)  and  a39810a );
 a39812a <=( a39811a  and  a39806a );
 a39816a <=( (not A199)  and  (not A167) );
 a39817a <=( (not A168)  and  a39816a );
 a39821a <=( (not A203)  and  (not A201) );
 a39822a <=( A200  and  a39821a );
 a39823a <=( a39822a  and  a39817a );
 a39827a <=( (not A298)  and  A267 );
 a39828a <=( A265  and  a39827a );
 a39832a <=( A301  and  (not A300) );
 a39833a <=( A299  and  a39832a );
 a39834a <=( a39833a  and  a39828a );
 a39838a <=( (not A199)  and  (not A167) );
 a39839a <=( (not A168)  and  a39838a );
 a39843a <=( (not A203)  and  (not A201) );
 a39844a <=( A200  and  a39843a );
 a39845a <=( a39844a  and  a39839a );
 a39849a <=( (not A298)  and  A267 );
 a39850a <=( A265  and  a39849a );
 a39854a <=( (not A302)  and  (not A300) );
 a39855a <=( A299  and  a39854a );
 a39856a <=( a39855a  and  a39850a );
 a39860a <=( (not A199)  and  (not A167) );
 a39861a <=( (not A168)  and  a39860a );
 a39865a <=( (not A203)  and  (not A201) );
 a39866a <=( A200  and  a39865a );
 a39867a <=( a39866a  and  a39861a );
 a39871a <=( A298  and  A267 );
 a39872a <=( A266  and  a39871a );
 a39876a <=( (not A301)  and  (not A300) );
 a39877a <=( A299  and  a39876a );
 a39878a <=( a39877a  and  a39872a );
 a39882a <=( (not A199)  and  (not A167) );
 a39883a <=( (not A168)  and  a39882a );
 a39887a <=( (not A203)  and  (not A201) );
 a39888a <=( A200  and  a39887a );
 a39889a <=( a39888a  and  a39883a );
 a39893a <=( A298  and  A267 );
 a39894a <=( A266  and  a39893a );
 a39898a <=( A302  and  (not A300) );
 a39899a <=( A299  and  a39898a );
 a39900a <=( a39899a  and  a39894a );
 a39904a <=( (not A199)  and  (not A167) );
 a39905a <=( (not A168)  and  a39904a );
 a39909a <=( (not A203)  and  (not A201) );
 a39910a <=( A200  and  a39909a );
 a39911a <=( a39910a  and  a39905a );
 a39915a <=( A298  and  A267 );
 a39916a <=( A266  and  a39915a );
 a39920a <=( A301  and  (not A300) );
 a39921a <=( (not A299)  and  a39920a );
 a39922a <=( a39921a  and  a39916a );
 a39926a <=( (not A199)  and  (not A167) );
 a39927a <=( (not A168)  and  a39926a );
 a39931a <=( (not A203)  and  (not A201) );
 a39932a <=( A200  and  a39931a );
 a39933a <=( a39932a  and  a39927a );
 a39937a <=( A298  and  A267 );
 a39938a <=( A266  and  a39937a );
 a39942a <=( (not A302)  and  (not A300) );
 a39943a <=( (not A299)  and  a39942a );
 a39944a <=( a39943a  and  a39938a );
 a39948a <=( (not A199)  and  (not A167) );
 a39949a <=( (not A168)  and  a39948a );
 a39953a <=( (not A203)  and  (not A201) );
 a39954a <=( A200  and  a39953a );
 a39955a <=( a39954a  and  a39949a );
 a39959a <=( (not A298)  and  A267 );
 a39960a <=( A266  and  a39959a );
 a39964a <=( A301  and  (not A300) );
 a39965a <=( A299  and  a39964a );
 a39966a <=( a39965a  and  a39960a );
 a39970a <=( (not A199)  and  (not A167) );
 a39971a <=( (not A168)  and  a39970a );
 a39975a <=( (not A203)  and  (not A201) );
 a39976a <=( A200  and  a39975a );
 a39977a <=( a39976a  and  a39971a );
 a39981a <=( (not A298)  and  A267 );
 a39982a <=( A266  and  a39981a );
 a39986a <=( (not A302)  and  (not A300) );
 a39987a <=( A299  and  a39986a );
 a39988a <=( a39987a  and  a39982a );
 a39992a <=( A199  and  (not A167) );
 a39993a <=( (not A168)  and  a39992a );
 a39997a <=( A203  and  (not A202) );
 a39998a <=( (not A200)  and  a39997a );
 a39999a <=( a39998a  and  a39993a );
 a40003a <=( (not A267)  and  A266 );
 a40004a <=( A265  and  a40003a );
 a40008a <=( A300  and  A299 );
 a40009a <=( (not A268)  and  a40008a );
 a40010a <=( a40009a  and  a40004a );
 a40014a <=( A199  and  (not A167) );
 a40015a <=( (not A168)  and  a40014a );
 a40019a <=( A203  and  (not A202) );
 a40020a <=( (not A200)  and  a40019a );
 a40021a <=( a40020a  and  a40015a );
 a40025a <=( (not A267)  and  A266 );
 a40026a <=( A265  and  a40025a );
 a40030a <=( A300  and  A298 );
 a40031a <=( (not A268)  and  a40030a );
 a40032a <=( a40031a  and  a40026a );
 a40036a <=( A199  and  (not A167) );
 a40037a <=( (not A168)  and  a40036a );
 a40041a <=( A203  and  (not A202) );
 a40042a <=( (not A200)  and  a40041a );
 a40043a <=( a40042a  and  a40037a );
 a40047a <=( (not A267)  and  A266 );
 a40048a <=( A265  and  a40047a );
 a40052a <=( A300  and  A299 );
 a40053a <=( A269  and  a40052a );
 a40054a <=( a40053a  and  a40048a );
 a40058a <=( A199  and  (not A167) );
 a40059a <=( (not A168)  and  a40058a );
 a40063a <=( A203  and  (not A202) );
 a40064a <=( (not A200)  and  a40063a );
 a40065a <=( a40064a  and  a40059a );
 a40069a <=( (not A267)  and  A266 );
 a40070a <=( A265  and  a40069a );
 a40074a <=( A300  and  A298 );
 a40075a <=( A269  and  a40074a );
 a40076a <=( a40075a  and  a40070a );
 a40080a <=( A199  and  (not A167) );
 a40081a <=( (not A168)  and  a40080a );
 a40085a <=( A203  and  (not A202) );
 a40086a <=( (not A200)  and  a40085a );
 a40087a <=( a40086a  and  a40081a );
 a40091a <=( (not A267)  and  A266 );
 a40092a <=( (not A265)  and  a40091a );
 a40096a <=( A300  and  A299 );
 a40097a <=( A268  and  a40096a );
 a40098a <=( a40097a  and  a40092a );
 a40102a <=( A199  and  (not A167) );
 a40103a <=( (not A168)  and  a40102a );
 a40107a <=( A203  and  (not A202) );
 a40108a <=( (not A200)  and  a40107a );
 a40109a <=( a40108a  and  a40103a );
 a40113a <=( (not A267)  and  A266 );
 a40114a <=( (not A265)  and  a40113a );
 a40118a <=( A300  and  A298 );
 a40119a <=( A268  and  a40118a );
 a40120a <=( a40119a  and  a40114a );
 a40124a <=( A199  and  (not A167) );
 a40125a <=( (not A168)  and  a40124a );
 a40129a <=( A203  and  (not A202) );
 a40130a <=( (not A200)  and  a40129a );
 a40131a <=( a40130a  and  a40125a );
 a40135a <=( (not A267)  and  A266 );
 a40136a <=( (not A265)  and  a40135a );
 a40140a <=( A300  and  A299 );
 a40141a <=( (not A269)  and  a40140a );
 a40142a <=( a40141a  and  a40136a );
 a40146a <=( A199  and  (not A167) );
 a40147a <=( (not A168)  and  a40146a );
 a40151a <=( A203  and  (not A202) );
 a40152a <=( (not A200)  and  a40151a );
 a40153a <=( a40152a  and  a40147a );
 a40157a <=( (not A267)  and  A266 );
 a40158a <=( (not A265)  and  a40157a );
 a40162a <=( A300  and  A298 );
 a40163a <=( (not A269)  and  a40162a );
 a40164a <=( a40163a  and  a40158a );
 a40168a <=( A199  and  (not A167) );
 a40169a <=( (not A168)  and  a40168a );
 a40173a <=( A203  and  (not A202) );
 a40174a <=( (not A200)  and  a40173a );
 a40175a <=( a40174a  and  a40169a );
 a40179a <=( (not A267)  and  (not A266) );
 a40180a <=( A265  and  a40179a );
 a40184a <=( A300  and  A299 );
 a40185a <=( A268  and  a40184a );
 a40186a <=( a40185a  and  a40180a );
 a40190a <=( A199  and  (not A167) );
 a40191a <=( (not A168)  and  a40190a );
 a40195a <=( A203  and  (not A202) );
 a40196a <=( (not A200)  and  a40195a );
 a40197a <=( a40196a  and  a40191a );
 a40201a <=( (not A267)  and  (not A266) );
 a40202a <=( A265  and  a40201a );
 a40206a <=( A300  and  A298 );
 a40207a <=( A268  and  a40206a );
 a40208a <=( a40207a  and  a40202a );
 a40212a <=( A199  and  (not A167) );
 a40213a <=( (not A168)  and  a40212a );
 a40217a <=( A203  and  (not A202) );
 a40218a <=( (not A200)  and  a40217a );
 a40219a <=( a40218a  and  a40213a );
 a40223a <=( (not A267)  and  (not A266) );
 a40224a <=( A265  and  a40223a );
 a40228a <=( A300  and  A299 );
 a40229a <=( (not A269)  and  a40228a );
 a40230a <=( a40229a  and  a40224a );
 a40234a <=( A199  and  (not A167) );
 a40235a <=( (not A168)  and  a40234a );
 a40239a <=( A203  and  (not A202) );
 a40240a <=( (not A200)  and  a40239a );
 a40241a <=( a40240a  and  a40235a );
 a40245a <=( (not A267)  and  (not A266) );
 a40246a <=( A265  and  a40245a );
 a40250a <=( A300  and  A298 );
 a40251a <=( (not A269)  and  a40250a );
 a40252a <=( a40251a  and  a40246a );
 a40256a <=( A199  and  (not A167) );
 a40257a <=( (not A168)  and  a40256a );
 a40261a <=( A202  and  (not A201) );
 a40262a <=( (not A200)  and  a40261a );
 a40263a <=( a40262a  and  a40257a );
 a40267a <=( A298  and  A267 );
 a40268a <=( A265  and  a40267a );
 a40272a <=( (not A301)  and  (not A300) );
 a40273a <=( A299  and  a40272a );
 a40274a <=( a40273a  and  a40268a );
 a40278a <=( A199  and  (not A167) );
 a40279a <=( (not A168)  and  a40278a );
 a40283a <=( A202  and  (not A201) );
 a40284a <=( (not A200)  and  a40283a );
 a40285a <=( a40284a  and  a40279a );
 a40289a <=( A298  and  A267 );
 a40290a <=( A265  and  a40289a );
 a40294a <=( A302  and  (not A300) );
 a40295a <=( A299  and  a40294a );
 a40296a <=( a40295a  and  a40290a );
 a40300a <=( A199  and  (not A167) );
 a40301a <=( (not A168)  and  a40300a );
 a40305a <=( A202  and  (not A201) );
 a40306a <=( (not A200)  and  a40305a );
 a40307a <=( a40306a  and  a40301a );
 a40311a <=( A298  and  A267 );
 a40312a <=( A265  and  a40311a );
 a40316a <=( A301  and  (not A300) );
 a40317a <=( (not A299)  and  a40316a );
 a40318a <=( a40317a  and  a40312a );
 a40322a <=( A199  and  (not A167) );
 a40323a <=( (not A168)  and  a40322a );
 a40327a <=( A202  and  (not A201) );
 a40328a <=( (not A200)  and  a40327a );
 a40329a <=( a40328a  and  a40323a );
 a40333a <=( A298  and  A267 );
 a40334a <=( A265  and  a40333a );
 a40338a <=( (not A302)  and  (not A300) );
 a40339a <=( (not A299)  and  a40338a );
 a40340a <=( a40339a  and  a40334a );
 a40344a <=( A199  and  (not A167) );
 a40345a <=( (not A168)  and  a40344a );
 a40349a <=( A202  and  (not A201) );
 a40350a <=( (not A200)  and  a40349a );
 a40351a <=( a40350a  and  a40345a );
 a40355a <=( (not A298)  and  A267 );
 a40356a <=( A265  and  a40355a );
 a40360a <=( A301  and  (not A300) );
 a40361a <=( A299  and  a40360a );
 a40362a <=( a40361a  and  a40356a );
 a40366a <=( A199  and  (not A167) );
 a40367a <=( (not A168)  and  a40366a );
 a40371a <=( A202  and  (not A201) );
 a40372a <=( (not A200)  and  a40371a );
 a40373a <=( a40372a  and  a40367a );
 a40377a <=( (not A298)  and  A267 );
 a40378a <=( A265  and  a40377a );
 a40382a <=( (not A302)  and  (not A300) );
 a40383a <=( A299  and  a40382a );
 a40384a <=( a40383a  and  a40378a );
 a40388a <=( A199  and  (not A167) );
 a40389a <=( (not A168)  and  a40388a );
 a40393a <=( A202  and  (not A201) );
 a40394a <=( (not A200)  and  a40393a );
 a40395a <=( a40394a  and  a40389a );
 a40399a <=( A298  and  A267 );
 a40400a <=( A266  and  a40399a );
 a40404a <=( (not A301)  and  (not A300) );
 a40405a <=( A299  and  a40404a );
 a40406a <=( a40405a  and  a40400a );
 a40410a <=( A199  and  (not A167) );
 a40411a <=( (not A168)  and  a40410a );
 a40415a <=( A202  and  (not A201) );
 a40416a <=( (not A200)  and  a40415a );
 a40417a <=( a40416a  and  a40411a );
 a40421a <=( A298  and  A267 );
 a40422a <=( A266  and  a40421a );
 a40426a <=( A302  and  (not A300) );
 a40427a <=( A299  and  a40426a );
 a40428a <=( a40427a  and  a40422a );
 a40432a <=( A199  and  (not A167) );
 a40433a <=( (not A168)  and  a40432a );
 a40437a <=( A202  and  (not A201) );
 a40438a <=( (not A200)  and  a40437a );
 a40439a <=( a40438a  and  a40433a );
 a40443a <=( A298  and  A267 );
 a40444a <=( A266  and  a40443a );
 a40448a <=( A301  and  (not A300) );
 a40449a <=( (not A299)  and  a40448a );
 a40450a <=( a40449a  and  a40444a );
 a40454a <=( A199  and  (not A167) );
 a40455a <=( (not A168)  and  a40454a );
 a40459a <=( A202  and  (not A201) );
 a40460a <=( (not A200)  and  a40459a );
 a40461a <=( a40460a  and  a40455a );
 a40465a <=( A298  and  A267 );
 a40466a <=( A266  and  a40465a );
 a40470a <=( (not A302)  and  (not A300) );
 a40471a <=( (not A299)  and  a40470a );
 a40472a <=( a40471a  and  a40466a );
 a40476a <=( A199  and  (not A167) );
 a40477a <=( (not A168)  and  a40476a );
 a40481a <=( A202  and  (not A201) );
 a40482a <=( (not A200)  and  a40481a );
 a40483a <=( a40482a  and  a40477a );
 a40487a <=( (not A298)  and  A267 );
 a40488a <=( A266  and  a40487a );
 a40492a <=( A301  and  (not A300) );
 a40493a <=( A299  and  a40492a );
 a40494a <=( a40493a  and  a40488a );
 a40498a <=( A199  and  (not A167) );
 a40499a <=( (not A168)  and  a40498a );
 a40503a <=( A202  and  (not A201) );
 a40504a <=( (not A200)  and  a40503a );
 a40505a <=( a40504a  and  a40499a );
 a40509a <=( (not A298)  and  A267 );
 a40510a <=( A266  and  a40509a );
 a40514a <=( (not A302)  and  (not A300) );
 a40515a <=( A299  and  a40514a );
 a40516a <=( a40515a  and  a40510a );
 a40520a <=( A199  and  (not A167) );
 a40521a <=( (not A168)  and  a40520a );
 a40525a <=( (not A203)  and  (not A201) );
 a40526a <=( (not A200)  and  a40525a );
 a40527a <=( a40526a  and  a40521a );
 a40531a <=( A298  and  A267 );
 a40532a <=( A265  and  a40531a );
 a40536a <=( (not A301)  and  (not A300) );
 a40537a <=( A299  and  a40536a );
 a40538a <=( a40537a  and  a40532a );
 a40542a <=( A199  and  (not A167) );
 a40543a <=( (not A168)  and  a40542a );
 a40547a <=( (not A203)  and  (not A201) );
 a40548a <=( (not A200)  and  a40547a );
 a40549a <=( a40548a  and  a40543a );
 a40553a <=( A298  and  A267 );
 a40554a <=( A265  and  a40553a );
 a40558a <=( A302  and  (not A300) );
 a40559a <=( A299  and  a40558a );
 a40560a <=( a40559a  and  a40554a );
 a40564a <=( A199  and  (not A167) );
 a40565a <=( (not A168)  and  a40564a );
 a40569a <=( (not A203)  and  (not A201) );
 a40570a <=( (not A200)  and  a40569a );
 a40571a <=( a40570a  and  a40565a );
 a40575a <=( A298  and  A267 );
 a40576a <=( A265  and  a40575a );
 a40580a <=( A301  and  (not A300) );
 a40581a <=( (not A299)  and  a40580a );
 a40582a <=( a40581a  and  a40576a );
 a40586a <=( A199  and  (not A167) );
 a40587a <=( (not A168)  and  a40586a );
 a40591a <=( (not A203)  and  (not A201) );
 a40592a <=( (not A200)  and  a40591a );
 a40593a <=( a40592a  and  a40587a );
 a40597a <=( A298  and  A267 );
 a40598a <=( A265  and  a40597a );
 a40602a <=( (not A302)  and  (not A300) );
 a40603a <=( (not A299)  and  a40602a );
 a40604a <=( a40603a  and  a40598a );
 a40608a <=( A199  and  (not A167) );
 a40609a <=( (not A168)  and  a40608a );
 a40613a <=( (not A203)  and  (not A201) );
 a40614a <=( (not A200)  and  a40613a );
 a40615a <=( a40614a  and  a40609a );
 a40619a <=( (not A298)  and  A267 );
 a40620a <=( A265  and  a40619a );
 a40624a <=( A301  and  (not A300) );
 a40625a <=( A299  and  a40624a );
 a40626a <=( a40625a  and  a40620a );
 a40630a <=( A199  and  (not A167) );
 a40631a <=( (not A168)  and  a40630a );
 a40635a <=( (not A203)  and  (not A201) );
 a40636a <=( (not A200)  and  a40635a );
 a40637a <=( a40636a  and  a40631a );
 a40641a <=( (not A298)  and  A267 );
 a40642a <=( A265  and  a40641a );
 a40646a <=( (not A302)  and  (not A300) );
 a40647a <=( A299  and  a40646a );
 a40648a <=( a40647a  and  a40642a );
 a40652a <=( A199  and  (not A167) );
 a40653a <=( (not A168)  and  a40652a );
 a40657a <=( (not A203)  and  (not A201) );
 a40658a <=( (not A200)  and  a40657a );
 a40659a <=( a40658a  and  a40653a );
 a40663a <=( A298  and  A267 );
 a40664a <=( A266  and  a40663a );
 a40668a <=( (not A301)  and  (not A300) );
 a40669a <=( A299  and  a40668a );
 a40670a <=( a40669a  and  a40664a );
 a40674a <=( A199  and  (not A167) );
 a40675a <=( (not A168)  and  a40674a );
 a40679a <=( (not A203)  and  (not A201) );
 a40680a <=( (not A200)  and  a40679a );
 a40681a <=( a40680a  and  a40675a );
 a40685a <=( A298  and  A267 );
 a40686a <=( A266  and  a40685a );
 a40690a <=( A302  and  (not A300) );
 a40691a <=( A299  and  a40690a );
 a40692a <=( a40691a  and  a40686a );
 a40696a <=( A199  and  (not A167) );
 a40697a <=( (not A168)  and  a40696a );
 a40701a <=( (not A203)  and  (not A201) );
 a40702a <=( (not A200)  and  a40701a );
 a40703a <=( a40702a  and  a40697a );
 a40707a <=( A298  and  A267 );
 a40708a <=( A266  and  a40707a );
 a40712a <=( A301  and  (not A300) );
 a40713a <=( (not A299)  and  a40712a );
 a40714a <=( a40713a  and  a40708a );
 a40718a <=( A199  and  (not A167) );
 a40719a <=( (not A168)  and  a40718a );
 a40723a <=( (not A203)  and  (not A201) );
 a40724a <=( (not A200)  and  a40723a );
 a40725a <=( a40724a  and  a40719a );
 a40729a <=( A298  and  A267 );
 a40730a <=( A266  and  a40729a );
 a40734a <=( (not A302)  and  (not A300) );
 a40735a <=( (not A299)  and  a40734a );
 a40736a <=( a40735a  and  a40730a );
 a40740a <=( A199  and  (not A167) );
 a40741a <=( (not A168)  and  a40740a );
 a40745a <=( (not A203)  and  (not A201) );
 a40746a <=( (not A200)  and  a40745a );
 a40747a <=( a40746a  and  a40741a );
 a40751a <=( (not A298)  and  A267 );
 a40752a <=( A266  and  a40751a );
 a40756a <=( A301  and  (not A300) );
 a40757a <=( A299  and  a40756a );
 a40758a <=( a40757a  and  a40752a );
 a40762a <=( A199  and  (not A167) );
 a40763a <=( (not A168)  and  a40762a );
 a40767a <=( (not A203)  and  (not A201) );
 a40768a <=( (not A200)  and  a40767a );
 a40769a <=( a40768a  and  a40763a );
 a40773a <=( (not A298)  and  A267 );
 a40774a <=( A266  and  a40773a );
 a40778a <=( (not A302)  and  (not A300) );
 a40779a <=( A299  and  a40778a );
 a40780a <=( a40779a  and  a40774a );
 a40784a <=( (not A199)  and  (not A167) );
 a40785a <=( (not A168)  and  a40784a );
 a40789a <=( A265  and  (not A202) );
 a40790a <=( (not A200)  and  a40789a );
 a40791a <=( a40790a  and  a40785a );
 a40795a <=( (not A269)  and  A268 );
 a40796a <=( A266  and  a40795a );
 a40800a <=( (not A301)  and  (not A299) );
 a40801a <=( (not A298)  and  a40800a );
 a40802a <=( a40801a  and  a40796a );
 a40806a <=( (not A199)  and  (not A167) );
 a40807a <=( (not A168)  and  a40806a );
 a40811a <=( A265  and  (not A202) );
 a40812a <=( (not A200)  and  a40811a );
 a40813a <=( a40812a  and  a40807a );
 a40817a <=( (not A269)  and  A268 );
 a40818a <=( A266  and  a40817a );
 a40822a <=( A302  and  (not A299) );
 a40823a <=( (not A298)  and  a40822a );
 a40824a <=( a40823a  and  a40818a );
 a40828a <=( (not A199)  and  (not A167) );
 a40829a <=( (not A168)  and  a40828a );
 a40833a <=( (not A265)  and  (not A202) );
 a40834a <=( (not A200)  and  a40833a );
 a40835a <=( a40834a  and  a40829a );
 a40839a <=( A269  and  (not A268) );
 a40840a <=( A266  and  a40839a );
 a40844a <=( (not A301)  and  (not A299) );
 a40845a <=( (not A298)  and  a40844a );
 a40846a <=( a40845a  and  a40840a );
 a40850a <=( (not A199)  and  (not A167) );
 a40851a <=( (not A168)  and  a40850a );
 a40855a <=( (not A265)  and  (not A202) );
 a40856a <=( (not A200)  and  a40855a );
 a40857a <=( a40856a  and  a40851a );
 a40861a <=( A269  and  (not A268) );
 a40862a <=( A266  and  a40861a );
 a40866a <=( A302  and  (not A299) );
 a40867a <=( (not A298)  and  a40866a );
 a40868a <=( a40867a  and  a40862a );
 a40872a <=( (not A199)  and  (not A167) );
 a40873a <=( (not A168)  and  a40872a );
 a40877a <=( A265  and  (not A202) );
 a40878a <=( (not A200)  and  a40877a );
 a40879a <=( a40878a  and  a40873a );
 a40883a <=( A269  and  (not A268) );
 a40884a <=( (not A266)  and  a40883a );
 a40888a <=( (not A301)  and  (not A299) );
 a40889a <=( (not A298)  and  a40888a );
 a40890a <=( a40889a  and  a40884a );
 a40894a <=( (not A199)  and  (not A167) );
 a40895a <=( (not A168)  and  a40894a );
 a40899a <=( A265  and  (not A202) );
 a40900a <=( (not A200)  and  a40899a );
 a40901a <=( a40900a  and  a40895a );
 a40905a <=( A269  and  (not A268) );
 a40906a <=( (not A266)  and  a40905a );
 a40910a <=( A302  and  (not A299) );
 a40911a <=( (not A298)  and  a40910a );
 a40912a <=( a40911a  and  a40906a );
 a40916a <=( (not A199)  and  (not A167) );
 a40917a <=( (not A168)  and  a40916a );
 a40921a <=( (not A265)  and  (not A202) );
 a40922a <=( (not A200)  and  a40921a );
 a40923a <=( a40922a  and  a40917a );
 a40927a <=( (not A269)  and  A268 );
 a40928a <=( (not A266)  and  a40927a );
 a40932a <=( (not A301)  and  (not A299) );
 a40933a <=( (not A298)  and  a40932a );
 a40934a <=( a40933a  and  a40928a );
 a40938a <=( (not A199)  and  (not A167) );
 a40939a <=( (not A168)  and  a40938a );
 a40943a <=( (not A265)  and  (not A202) );
 a40944a <=( (not A200)  and  a40943a );
 a40945a <=( a40944a  and  a40939a );
 a40949a <=( (not A269)  and  A268 );
 a40950a <=( (not A266)  and  a40949a );
 a40954a <=( A302  and  (not A299) );
 a40955a <=( (not A298)  and  a40954a );
 a40956a <=( a40955a  and  a40950a );
 a40960a <=( (not A199)  and  (not A167) );
 a40961a <=( (not A168)  and  a40960a );
 a40965a <=( A265  and  A203 );
 a40966a <=( (not A200)  and  a40965a );
 a40967a <=( a40966a  and  a40961a );
 a40971a <=( (not A269)  and  A268 );
 a40972a <=( A266  and  a40971a );
 a40976a <=( (not A301)  and  (not A299) );
 a40977a <=( (not A298)  and  a40976a );
 a40978a <=( a40977a  and  a40972a );
 a40982a <=( (not A199)  and  (not A167) );
 a40983a <=( (not A168)  and  a40982a );
 a40987a <=( A265  and  A203 );
 a40988a <=( (not A200)  and  a40987a );
 a40989a <=( a40988a  and  a40983a );
 a40993a <=( (not A269)  and  A268 );
 a40994a <=( A266  and  a40993a );
 a40998a <=( A302  and  (not A299) );
 a40999a <=( (not A298)  and  a40998a );
 a41000a <=( a40999a  and  a40994a );
 a41004a <=( (not A199)  and  (not A167) );
 a41005a <=( (not A168)  and  a41004a );
 a41009a <=( (not A265)  and  A203 );
 a41010a <=( (not A200)  and  a41009a );
 a41011a <=( a41010a  and  a41005a );
 a41015a <=( A269  and  (not A268) );
 a41016a <=( A266  and  a41015a );
 a41020a <=( (not A301)  and  (not A299) );
 a41021a <=( (not A298)  and  a41020a );
 a41022a <=( a41021a  and  a41016a );
 a41026a <=( (not A199)  and  (not A167) );
 a41027a <=( (not A168)  and  a41026a );
 a41031a <=( (not A265)  and  A203 );
 a41032a <=( (not A200)  and  a41031a );
 a41033a <=( a41032a  and  a41027a );
 a41037a <=( A269  and  (not A268) );
 a41038a <=( A266  and  a41037a );
 a41042a <=( A302  and  (not A299) );
 a41043a <=( (not A298)  and  a41042a );
 a41044a <=( a41043a  and  a41038a );
 a41048a <=( (not A199)  and  (not A167) );
 a41049a <=( (not A168)  and  a41048a );
 a41053a <=( A265  and  A203 );
 a41054a <=( (not A200)  and  a41053a );
 a41055a <=( a41054a  and  a41049a );
 a41059a <=( A269  and  (not A268) );
 a41060a <=( (not A266)  and  a41059a );
 a41064a <=( (not A301)  and  (not A299) );
 a41065a <=( (not A298)  and  a41064a );
 a41066a <=( a41065a  and  a41060a );
 a41070a <=( (not A199)  and  (not A167) );
 a41071a <=( (not A168)  and  a41070a );
 a41075a <=( A265  and  A203 );
 a41076a <=( (not A200)  and  a41075a );
 a41077a <=( a41076a  and  a41071a );
 a41081a <=( A269  and  (not A268) );
 a41082a <=( (not A266)  and  a41081a );
 a41086a <=( A302  and  (not A299) );
 a41087a <=( (not A298)  and  a41086a );
 a41088a <=( a41087a  and  a41082a );
 a41092a <=( (not A199)  and  (not A167) );
 a41093a <=( (not A168)  and  a41092a );
 a41097a <=( (not A265)  and  A203 );
 a41098a <=( (not A200)  and  a41097a );
 a41099a <=( a41098a  and  a41093a );
 a41103a <=( (not A269)  and  A268 );
 a41104a <=( (not A266)  and  a41103a );
 a41108a <=( (not A301)  and  (not A299) );
 a41109a <=( (not A298)  and  a41108a );
 a41110a <=( a41109a  and  a41104a );
 a41114a <=( (not A199)  and  (not A167) );
 a41115a <=( (not A168)  and  a41114a );
 a41119a <=( (not A265)  and  A203 );
 a41120a <=( (not A200)  and  a41119a );
 a41121a <=( a41120a  and  a41115a );
 a41125a <=( (not A269)  and  A268 );
 a41126a <=( (not A266)  and  a41125a );
 a41130a <=( A302  and  (not A299) );
 a41131a <=( (not A298)  and  a41130a );
 a41132a <=( a41131a  and  a41126a );
 a41136a <=( (not A199)  and  (not A167) );
 a41137a <=( (not A168)  and  a41136a );
 a41141a <=( (not A203)  and  A202 );
 a41142a <=( (not A200)  and  a41141a );
 a41143a <=( a41142a  and  a41137a );
 a41147a <=( (not A267)  and  A266 );
 a41148a <=( A265  and  a41147a );
 a41152a <=( A300  and  A299 );
 a41153a <=( (not A268)  and  a41152a );
 a41154a <=( a41153a  and  a41148a );
 a41158a <=( (not A199)  and  (not A167) );
 a41159a <=( (not A168)  and  a41158a );
 a41163a <=( (not A203)  and  A202 );
 a41164a <=( (not A200)  and  a41163a );
 a41165a <=( a41164a  and  a41159a );
 a41169a <=( (not A267)  and  A266 );
 a41170a <=( A265  and  a41169a );
 a41174a <=( A300  and  A298 );
 a41175a <=( (not A268)  and  a41174a );
 a41176a <=( a41175a  and  a41170a );
 a41180a <=( (not A199)  and  (not A167) );
 a41181a <=( (not A168)  and  a41180a );
 a41185a <=( (not A203)  and  A202 );
 a41186a <=( (not A200)  and  a41185a );
 a41187a <=( a41186a  and  a41181a );
 a41191a <=( (not A267)  and  A266 );
 a41192a <=( A265  and  a41191a );
 a41196a <=( A300  and  A299 );
 a41197a <=( A269  and  a41196a );
 a41198a <=( a41197a  and  a41192a );
 a41202a <=( (not A199)  and  (not A167) );
 a41203a <=( (not A168)  and  a41202a );
 a41207a <=( (not A203)  and  A202 );
 a41208a <=( (not A200)  and  a41207a );
 a41209a <=( a41208a  and  a41203a );
 a41213a <=( (not A267)  and  A266 );
 a41214a <=( A265  and  a41213a );
 a41218a <=( A300  and  A298 );
 a41219a <=( A269  and  a41218a );
 a41220a <=( a41219a  and  a41214a );
 a41224a <=( (not A199)  and  (not A167) );
 a41225a <=( (not A168)  and  a41224a );
 a41229a <=( (not A203)  and  A202 );
 a41230a <=( (not A200)  and  a41229a );
 a41231a <=( a41230a  and  a41225a );
 a41235a <=( (not A267)  and  A266 );
 a41236a <=( (not A265)  and  a41235a );
 a41240a <=( A300  and  A299 );
 a41241a <=( A268  and  a41240a );
 a41242a <=( a41241a  and  a41236a );
 a41246a <=( (not A199)  and  (not A167) );
 a41247a <=( (not A168)  and  a41246a );
 a41251a <=( (not A203)  and  A202 );
 a41252a <=( (not A200)  and  a41251a );
 a41253a <=( a41252a  and  a41247a );
 a41257a <=( (not A267)  and  A266 );
 a41258a <=( (not A265)  and  a41257a );
 a41262a <=( A300  and  A298 );
 a41263a <=( A268  and  a41262a );
 a41264a <=( a41263a  and  a41258a );
 a41268a <=( (not A199)  and  (not A167) );
 a41269a <=( (not A168)  and  a41268a );
 a41273a <=( (not A203)  and  A202 );
 a41274a <=( (not A200)  and  a41273a );
 a41275a <=( a41274a  and  a41269a );
 a41279a <=( (not A267)  and  A266 );
 a41280a <=( (not A265)  and  a41279a );
 a41284a <=( A300  and  A299 );
 a41285a <=( (not A269)  and  a41284a );
 a41286a <=( a41285a  and  a41280a );
 a41290a <=( (not A199)  and  (not A167) );
 a41291a <=( (not A168)  and  a41290a );
 a41295a <=( (not A203)  and  A202 );
 a41296a <=( (not A200)  and  a41295a );
 a41297a <=( a41296a  and  a41291a );
 a41301a <=( (not A267)  and  A266 );
 a41302a <=( (not A265)  and  a41301a );
 a41306a <=( A300  and  A298 );
 a41307a <=( (not A269)  and  a41306a );
 a41308a <=( a41307a  and  a41302a );
 a41312a <=( (not A199)  and  (not A167) );
 a41313a <=( (not A168)  and  a41312a );
 a41317a <=( (not A203)  and  A202 );
 a41318a <=( (not A200)  and  a41317a );
 a41319a <=( a41318a  and  a41313a );
 a41323a <=( (not A267)  and  (not A266) );
 a41324a <=( A265  and  a41323a );
 a41328a <=( A300  and  A299 );
 a41329a <=( A268  and  a41328a );
 a41330a <=( a41329a  and  a41324a );
 a41334a <=( (not A199)  and  (not A167) );
 a41335a <=( (not A168)  and  a41334a );
 a41339a <=( (not A203)  and  A202 );
 a41340a <=( (not A200)  and  a41339a );
 a41341a <=( a41340a  and  a41335a );
 a41345a <=( (not A267)  and  (not A266) );
 a41346a <=( A265  and  a41345a );
 a41350a <=( A300  and  A298 );
 a41351a <=( A268  and  a41350a );
 a41352a <=( a41351a  and  a41346a );
 a41356a <=( (not A199)  and  (not A167) );
 a41357a <=( (not A168)  and  a41356a );
 a41361a <=( (not A203)  and  A202 );
 a41362a <=( (not A200)  and  a41361a );
 a41363a <=( a41362a  and  a41357a );
 a41367a <=( (not A267)  and  (not A266) );
 a41368a <=( A265  and  a41367a );
 a41372a <=( A300  and  A299 );
 a41373a <=( (not A269)  and  a41372a );
 a41374a <=( a41373a  and  a41368a );
 a41378a <=( (not A199)  and  (not A167) );
 a41379a <=( (not A168)  and  a41378a );
 a41383a <=( (not A203)  and  A202 );
 a41384a <=( (not A200)  and  a41383a );
 a41385a <=( a41384a  and  a41379a );
 a41389a <=( (not A267)  and  (not A266) );
 a41390a <=( A265  and  a41389a );
 a41394a <=( A300  and  A298 );
 a41395a <=( (not A269)  and  a41394a );
 a41396a <=( a41395a  and  a41390a );
 a41400a <=( (not A167)  and  A168 );
 a41401a <=( A170  and  a41400a );
 a41405a <=( A201  and  A199 );
 a41406a <=( A166  and  a41405a );
 a41407a <=( a41406a  and  a41401a );
 a41411a <=( A298  and  A267 );
 a41412a <=( A265  and  a41411a );
 a41416a <=( (not A301)  and  (not A300) );
 a41417a <=( A299  and  a41416a );
 a41418a <=( a41417a  and  a41412a );
 a41422a <=( (not A167)  and  A168 );
 a41423a <=( A170  and  a41422a );
 a41427a <=( A201  and  A199 );
 a41428a <=( A166  and  a41427a );
 a41429a <=( a41428a  and  a41423a );
 a41433a <=( A298  and  A267 );
 a41434a <=( A265  and  a41433a );
 a41438a <=( A302  and  (not A300) );
 a41439a <=( A299  and  a41438a );
 a41440a <=( a41439a  and  a41434a );
 a41444a <=( (not A167)  and  A168 );
 a41445a <=( A170  and  a41444a );
 a41449a <=( A201  and  A199 );
 a41450a <=( A166  and  a41449a );
 a41451a <=( a41450a  and  a41445a );
 a41455a <=( A298  and  A267 );
 a41456a <=( A265  and  a41455a );
 a41460a <=( A301  and  (not A300) );
 a41461a <=( (not A299)  and  a41460a );
 a41462a <=( a41461a  and  a41456a );
 a41466a <=( (not A167)  and  A168 );
 a41467a <=( A170  and  a41466a );
 a41471a <=( A201  and  A199 );
 a41472a <=( A166  and  a41471a );
 a41473a <=( a41472a  and  a41467a );
 a41477a <=( A298  and  A267 );
 a41478a <=( A265  and  a41477a );
 a41482a <=( (not A302)  and  (not A300) );
 a41483a <=( (not A299)  and  a41482a );
 a41484a <=( a41483a  and  a41478a );
 a41488a <=( (not A167)  and  A168 );
 a41489a <=( A170  and  a41488a );
 a41493a <=( A201  and  A199 );
 a41494a <=( A166  and  a41493a );
 a41495a <=( a41494a  and  a41489a );
 a41499a <=( (not A298)  and  A267 );
 a41500a <=( A265  and  a41499a );
 a41504a <=( A301  and  (not A300) );
 a41505a <=( A299  and  a41504a );
 a41506a <=( a41505a  and  a41500a );
 a41510a <=( (not A167)  and  A168 );
 a41511a <=( A170  and  a41510a );
 a41515a <=( A201  and  A199 );
 a41516a <=( A166  and  a41515a );
 a41517a <=( a41516a  and  a41511a );
 a41521a <=( (not A298)  and  A267 );
 a41522a <=( A265  and  a41521a );
 a41526a <=( (not A302)  and  (not A300) );
 a41527a <=( A299  and  a41526a );
 a41528a <=( a41527a  and  a41522a );
 a41532a <=( (not A167)  and  A168 );
 a41533a <=( A170  and  a41532a );
 a41537a <=( A201  and  A199 );
 a41538a <=( A166  and  a41537a );
 a41539a <=( a41538a  and  a41533a );
 a41543a <=( A298  and  A267 );
 a41544a <=( A266  and  a41543a );
 a41548a <=( (not A301)  and  (not A300) );
 a41549a <=( A299  and  a41548a );
 a41550a <=( a41549a  and  a41544a );
 a41554a <=( (not A167)  and  A168 );
 a41555a <=( A170  and  a41554a );
 a41559a <=( A201  and  A199 );
 a41560a <=( A166  and  a41559a );
 a41561a <=( a41560a  and  a41555a );
 a41565a <=( A298  and  A267 );
 a41566a <=( A266  and  a41565a );
 a41570a <=( A302  and  (not A300) );
 a41571a <=( A299  and  a41570a );
 a41572a <=( a41571a  and  a41566a );
 a41576a <=( (not A167)  and  A168 );
 a41577a <=( A170  and  a41576a );
 a41581a <=( A201  and  A199 );
 a41582a <=( A166  and  a41581a );
 a41583a <=( a41582a  and  a41577a );
 a41587a <=( A298  and  A267 );
 a41588a <=( A266  and  a41587a );
 a41592a <=( A301  and  (not A300) );
 a41593a <=( (not A299)  and  a41592a );
 a41594a <=( a41593a  and  a41588a );
 a41598a <=( (not A167)  and  A168 );
 a41599a <=( A170  and  a41598a );
 a41603a <=( A201  and  A199 );
 a41604a <=( A166  and  a41603a );
 a41605a <=( a41604a  and  a41599a );
 a41609a <=( A298  and  A267 );
 a41610a <=( A266  and  a41609a );
 a41614a <=( (not A302)  and  (not A300) );
 a41615a <=( (not A299)  and  a41614a );
 a41616a <=( a41615a  and  a41610a );
 a41620a <=( (not A167)  and  A168 );
 a41621a <=( A170  and  a41620a );
 a41625a <=( A201  and  A199 );
 a41626a <=( A166  and  a41625a );
 a41627a <=( a41626a  and  a41621a );
 a41631a <=( (not A298)  and  A267 );
 a41632a <=( A266  and  a41631a );
 a41636a <=( A301  and  (not A300) );
 a41637a <=( A299  and  a41636a );
 a41638a <=( a41637a  and  a41632a );
 a41642a <=( (not A167)  and  A168 );
 a41643a <=( A170  and  a41642a );
 a41647a <=( A201  and  A199 );
 a41648a <=( A166  and  a41647a );
 a41649a <=( a41648a  and  a41643a );
 a41653a <=( (not A298)  and  A267 );
 a41654a <=( A266  and  a41653a );
 a41658a <=( (not A302)  and  (not A300) );
 a41659a <=( A299  and  a41658a );
 a41660a <=( a41659a  and  a41654a );
 a41664a <=( (not A167)  and  A168 );
 a41665a <=( A170  and  a41664a );
 a41669a <=( A201  and  A200 );
 a41670a <=( A166  and  a41669a );
 a41671a <=( a41670a  and  a41665a );
 a41675a <=( A298  and  A267 );
 a41676a <=( A265  and  a41675a );
 a41680a <=( (not A301)  and  (not A300) );
 a41681a <=( A299  and  a41680a );
 a41682a <=( a41681a  and  a41676a );
 a41686a <=( (not A167)  and  A168 );
 a41687a <=( A170  and  a41686a );
 a41691a <=( A201  and  A200 );
 a41692a <=( A166  and  a41691a );
 a41693a <=( a41692a  and  a41687a );
 a41697a <=( A298  and  A267 );
 a41698a <=( A265  and  a41697a );
 a41702a <=( A302  and  (not A300) );
 a41703a <=( A299  and  a41702a );
 a41704a <=( a41703a  and  a41698a );
 a41708a <=( (not A167)  and  A168 );
 a41709a <=( A170  and  a41708a );
 a41713a <=( A201  and  A200 );
 a41714a <=( A166  and  a41713a );
 a41715a <=( a41714a  and  a41709a );
 a41719a <=( A298  and  A267 );
 a41720a <=( A265  and  a41719a );
 a41724a <=( A301  and  (not A300) );
 a41725a <=( (not A299)  and  a41724a );
 a41726a <=( a41725a  and  a41720a );
 a41730a <=( (not A167)  and  A168 );
 a41731a <=( A170  and  a41730a );
 a41735a <=( A201  and  A200 );
 a41736a <=( A166  and  a41735a );
 a41737a <=( a41736a  and  a41731a );
 a41741a <=( A298  and  A267 );
 a41742a <=( A265  and  a41741a );
 a41746a <=( (not A302)  and  (not A300) );
 a41747a <=( (not A299)  and  a41746a );
 a41748a <=( a41747a  and  a41742a );
 a41752a <=( (not A167)  and  A168 );
 a41753a <=( A170  and  a41752a );
 a41757a <=( A201  and  A200 );
 a41758a <=( A166  and  a41757a );
 a41759a <=( a41758a  and  a41753a );
 a41763a <=( (not A298)  and  A267 );
 a41764a <=( A265  and  a41763a );
 a41768a <=( A301  and  (not A300) );
 a41769a <=( A299  and  a41768a );
 a41770a <=( a41769a  and  a41764a );
 a41774a <=( (not A167)  and  A168 );
 a41775a <=( A170  and  a41774a );
 a41779a <=( A201  and  A200 );
 a41780a <=( A166  and  a41779a );
 a41781a <=( a41780a  and  a41775a );
 a41785a <=( (not A298)  and  A267 );
 a41786a <=( A265  and  a41785a );
 a41790a <=( (not A302)  and  (not A300) );
 a41791a <=( A299  and  a41790a );
 a41792a <=( a41791a  and  a41786a );
 a41796a <=( (not A167)  and  A168 );
 a41797a <=( A170  and  a41796a );
 a41801a <=( A201  and  A200 );
 a41802a <=( A166  and  a41801a );
 a41803a <=( a41802a  and  a41797a );
 a41807a <=( A298  and  A267 );
 a41808a <=( A266  and  a41807a );
 a41812a <=( (not A301)  and  (not A300) );
 a41813a <=( A299  and  a41812a );
 a41814a <=( a41813a  and  a41808a );
 a41818a <=( (not A167)  and  A168 );
 a41819a <=( A170  and  a41818a );
 a41823a <=( A201  and  A200 );
 a41824a <=( A166  and  a41823a );
 a41825a <=( a41824a  and  a41819a );
 a41829a <=( A298  and  A267 );
 a41830a <=( A266  and  a41829a );
 a41834a <=( A302  and  (not A300) );
 a41835a <=( A299  and  a41834a );
 a41836a <=( a41835a  and  a41830a );
 a41840a <=( (not A167)  and  A168 );
 a41841a <=( A170  and  a41840a );
 a41845a <=( A201  and  A200 );
 a41846a <=( A166  and  a41845a );
 a41847a <=( a41846a  and  a41841a );
 a41851a <=( A298  and  A267 );
 a41852a <=( A266  and  a41851a );
 a41856a <=( A301  and  (not A300) );
 a41857a <=( (not A299)  and  a41856a );
 a41858a <=( a41857a  and  a41852a );
 a41862a <=( (not A167)  and  A168 );
 a41863a <=( A170  and  a41862a );
 a41867a <=( A201  and  A200 );
 a41868a <=( A166  and  a41867a );
 a41869a <=( a41868a  and  a41863a );
 a41873a <=( A298  and  A267 );
 a41874a <=( A266  and  a41873a );
 a41878a <=( (not A302)  and  (not A300) );
 a41879a <=( (not A299)  and  a41878a );
 a41880a <=( a41879a  and  a41874a );
 a41884a <=( (not A167)  and  A168 );
 a41885a <=( A170  and  a41884a );
 a41889a <=( A201  and  A200 );
 a41890a <=( A166  and  a41889a );
 a41891a <=( a41890a  and  a41885a );
 a41895a <=( (not A298)  and  A267 );
 a41896a <=( A266  and  a41895a );
 a41900a <=( A301  and  (not A300) );
 a41901a <=( A299  and  a41900a );
 a41902a <=( a41901a  and  a41896a );
 a41906a <=( (not A167)  and  A168 );
 a41907a <=( A170  and  a41906a );
 a41911a <=( A201  and  A200 );
 a41912a <=( A166  and  a41911a );
 a41913a <=( a41912a  and  a41907a );
 a41917a <=( (not A298)  and  A267 );
 a41918a <=( A266  and  a41917a );
 a41922a <=( (not A302)  and  (not A300) );
 a41923a <=( A299  and  a41922a );
 a41924a <=( a41923a  and  a41918a );
 a41928a <=( (not A167)  and  A168 );
 a41929a <=( A170  and  a41928a );
 a41933a <=( (not A200)  and  (not A199) );
 a41934a <=( A166  and  a41933a );
 a41935a <=( a41934a  and  a41929a );
 a41939a <=( (not A266)  and  (not A265) );
 a41940a <=( (not A202)  and  a41939a );
 a41944a <=( A300  and  A299 );
 a41945a <=( (not A268)  and  a41944a );
 a41946a <=( a41945a  and  a41940a );
 a41950a <=( (not A167)  and  A168 );
 a41951a <=( A170  and  a41950a );
 a41955a <=( (not A200)  and  (not A199) );
 a41956a <=( A166  and  a41955a );
 a41957a <=( a41956a  and  a41951a );
 a41961a <=( (not A266)  and  (not A265) );
 a41962a <=( (not A202)  and  a41961a );
 a41966a <=( A300  and  A298 );
 a41967a <=( (not A268)  and  a41966a );
 a41968a <=( a41967a  and  a41962a );
 a41972a <=( (not A167)  and  A168 );
 a41973a <=( A170  and  a41972a );
 a41977a <=( (not A200)  and  (not A199) );
 a41978a <=( A166  and  a41977a );
 a41979a <=( a41978a  and  a41973a );
 a41983a <=( (not A266)  and  (not A265) );
 a41984a <=( (not A202)  and  a41983a );
 a41988a <=( A300  and  A299 );
 a41989a <=( A269  and  a41988a );
 a41990a <=( a41989a  and  a41984a );
 a41994a <=( (not A167)  and  A168 );
 a41995a <=( A170  and  a41994a );
 a41999a <=( (not A200)  and  (not A199) );
 a42000a <=( A166  and  a41999a );
 a42001a <=( a42000a  and  a41995a );
 a42005a <=( (not A266)  and  (not A265) );
 a42006a <=( (not A202)  and  a42005a );
 a42010a <=( A300  and  A298 );
 a42011a <=( A269  and  a42010a );
 a42012a <=( a42011a  and  a42006a );
 a42016a <=( (not A167)  and  A168 );
 a42017a <=( A170  and  a42016a );
 a42021a <=( (not A200)  and  (not A199) );
 a42022a <=( A166  and  a42021a );
 a42023a <=( a42022a  and  a42017a );
 a42027a <=( (not A266)  and  (not A265) );
 a42028a <=( A203  and  a42027a );
 a42032a <=( A300  and  A299 );
 a42033a <=( (not A268)  and  a42032a );
 a42034a <=( a42033a  and  a42028a );
 a42038a <=( (not A167)  and  A168 );
 a42039a <=( A170  and  a42038a );
 a42043a <=( (not A200)  and  (not A199) );
 a42044a <=( A166  and  a42043a );
 a42045a <=( a42044a  and  a42039a );
 a42049a <=( (not A266)  and  (not A265) );
 a42050a <=( A203  and  a42049a );
 a42054a <=( A300  and  A298 );
 a42055a <=( (not A268)  and  a42054a );
 a42056a <=( a42055a  and  a42050a );
 a42060a <=( (not A167)  and  A168 );
 a42061a <=( A170  and  a42060a );
 a42065a <=( (not A200)  and  (not A199) );
 a42066a <=( A166  and  a42065a );
 a42067a <=( a42066a  and  a42061a );
 a42071a <=( (not A266)  and  (not A265) );
 a42072a <=( A203  and  a42071a );
 a42076a <=( A300  and  A299 );
 a42077a <=( A269  and  a42076a );
 a42078a <=( a42077a  and  a42072a );
 a42082a <=( (not A167)  and  A168 );
 a42083a <=( A170  and  a42082a );
 a42087a <=( (not A200)  and  (not A199) );
 a42088a <=( A166  and  a42087a );
 a42089a <=( a42088a  and  a42083a );
 a42093a <=( (not A266)  and  (not A265) );
 a42094a <=( A203  and  a42093a );
 a42098a <=( A300  and  A298 );
 a42099a <=( A269  and  a42098a );
 a42100a <=( a42099a  and  a42094a );
 a42104a <=( (not A167)  and  A168 );
 a42105a <=( A169  and  a42104a );
 a42109a <=( A201  and  A199 );
 a42110a <=( A166  and  a42109a );
 a42111a <=( a42110a  and  a42105a );
 a42115a <=( A298  and  A267 );
 a42116a <=( A265  and  a42115a );
 a42120a <=( (not A301)  and  (not A300) );
 a42121a <=( A299  and  a42120a );
 a42122a <=( a42121a  and  a42116a );
 a42126a <=( (not A167)  and  A168 );
 a42127a <=( A169  and  a42126a );
 a42131a <=( A201  and  A199 );
 a42132a <=( A166  and  a42131a );
 a42133a <=( a42132a  and  a42127a );
 a42137a <=( A298  and  A267 );
 a42138a <=( A265  and  a42137a );
 a42142a <=( A302  and  (not A300) );
 a42143a <=( A299  and  a42142a );
 a42144a <=( a42143a  and  a42138a );
 a42148a <=( (not A167)  and  A168 );
 a42149a <=( A169  and  a42148a );
 a42153a <=( A201  and  A199 );
 a42154a <=( A166  and  a42153a );
 a42155a <=( a42154a  and  a42149a );
 a42159a <=( A298  and  A267 );
 a42160a <=( A265  and  a42159a );
 a42164a <=( A301  and  (not A300) );
 a42165a <=( (not A299)  and  a42164a );
 a42166a <=( a42165a  and  a42160a );
 a42170a <=( (not A167)  and  A168 );
 a42171a <=( A169  and  a42170a );
 a42175a <=( A201  and  A199 );
 a42176a <=( A166  and  a42175a );
 a42177a <=( a42176a  and  a42171a );
 a42181a <=( A298  and  A267 );
 a42182a <=( A265  and  a42181a );
 a42186a <=( (not A302)  and  (not A300) );
 a42187a <=( (not A299)  and  a42186a );
 a42188a <=( a42187a  and  a42182a );
 a42192a <=( (not A167)  and  A168 );
 a42193a <=( A169  and  a42192a );
 a42197a <=( A201  and  A199 );
 a42198a <=( A166  and  a42197a );
 a42199a <=( a42198a  and  a42193a );
 a42203a <=( (not A298)  and  A267 );
 a42204a <=( A265  and  a42203a );
 a42208a <=( A301  and  (not A300) );
 a42209a <=( A299  and  a42208a );
 a42210a <=( a42209a  and  a42204a );
 a42214a <=( (not A167)  and  A168 );
 a42215a <=( A169  and  a42214a );
 a42219a <=( A201  and  A199 );
 a42220a <=( A166  and  a42219a );
 a42221a <=( a42220a  and  a42215a );
 a42225a <=( (not A298)  and  A267 );
 a42226a <=( A265  and  a42225a );
 a42230a <=( (not A302)  and  (not A300) );
 a42231a <=( A299  and  a42230a );
 a42232a <=( a42231a  and  a42226a );
 a42236a <=( (not A167)  and  A168 );
 a42237a <=( A169  and  a42236a );
 a42241a <=( A201  and  A199 );
 a42242a <=( A166  and  a42241a );
 a42243a <=( a42242a  and  a42237a );
 a42247a <=( A298  and  A267 );
 a42248a <=( A266  and  a42247a );
 a42252a <=( (not A301)  and  (not A300) );
 a42253a <=( A299  and  a42252a );
 a42254a <=( a42253a  and  a42248a );
 a42258a <=( (not A167)  and  A168 );
 a42259a <=( A169  and  a42258a );
 a42263a <=( A201  and  A199 );
 a42264a <=( A166  and  a42263a );
 a42265a <=( a42264a  and  a42259a );
 a42269a <=( A298  and  A267 );
 a42270a <=( A266  and  a42269a );
 a42274a <=( A302  and  (not A300) );
 a42275a <=( A299  and  a42274a );
 a42276a <=( a42275a  and  a42270a );
 a42280a <=( (not A167)  and  A168 );
 a42281a <=( A169  and  a42280a );
 a42285a <=( A201  and  A199 );
 a42286a <=( A166  and  a42285a );
 a42287a <=( a42286a  and  a42281a );
 a42291a <=( A298  and  A267 );
 a42292a <=( A266  and  a42291a );
 a42296a <=( A301  and  (not A300) );
 a42297a <=( (not A299)  and  a42296a );
 a42298a <=( a42297a  and  a42292a );
 a42302a <=( (not A167)  and  A168 );
 a42303a <=( A169  and  a42302a );
 a42307a <=( A201  and  A199 );
 a42308a <=( A166  and  a42307a );
 a42309a <=( a42308a  and  a42303a );
 a42313a <=( A298  and  A267 );
 a42314a <=( A266  and  a42313a );
 a42318a <=( (not A302)  and  (not A300) );
 a42319a <=( (not A299)  and  a42318a );
 a42320a <=( a42319a  and  a42314a );
 a42324a <=( (not A167)  and  A168 );
 a42325a <=( A169  and  a42324a );
 a42329a <=( A201  and  A199 );
 a42330a <=( A166  and  a42329a );
 a42331a <=( a42330a  and  a42325a );
 a42335a <=( (not A298)  and  A267 );
 a42336a <=( A266  and  a42335a );
 a42340a <=( A301  and  (not A300) );
 a42341a <=( A299  and  a42340a );
 a42342a <=( a42341a  and  a42336a );
 a42346a <=( (not A167)  and  A168 );
 a42347a <=( A169  and  a42346a );
 a42351a <=( A201  and  A199 );
 a42352a <=( A166  and  a42351a );
 a42353a <=( a42352a  and  a42347a );
 a42357a <=( (not A298)  and  A267 );
 a42358a <=( A266  and  a42357a );
 a42362a <=( (not A302)  and  (not A300) );
 a42363a <=( A299  and  a42362a );
 a42364a <=( a42363a  and  a42358a );
 a42368a <=( (not A167)  and  A168 );
 a42369a <=( A169  and  a42368a );
 a42373a <=( A201  and  A200 );
 a42374a <=( A166  and  a42373a );
 a42375a <=( a42374a  and  a42369a );
 a42379a <=( A298  and  A267 );
 a42380a <=( A265  and  a42379a );
 a42384a <=( (not A301)  and  (not A300) );
 a42385a <=( A299  and  a42384a );
 a42386a <=( a42385a  and  a42380a );
 a42390a <=( (not A167)  and  A168 );
 a42391a <=( A169  and  a42390a );
 a42395a <=( A201  and  A200 );
 a42396a <=( A166  and  a42395a );
 a42397a <=( a42396a  and  a42391a );
 a42401a <=( A298  and  A267 );
 a42402a <=( A265  and  a42401a );
 a42406a <=( A302  and  (not A300) );
 a42407a <=( A299  and  a42406a );
 a42408a <=( a42407a  and  a42402a );
 a42412a <=( (not A167)  and  A168 );
 a42413a <=( A169  and  a42412a );
 a42417a <=( A201  and  A200 );
 a42418a <=( A166  and  a42417a );
 a42419a <=( a42418a  and  a42413a );
 a42423a <=( A298  and  A267 );
 a42424a <=( A265  and  a42423a );
 a42428a <=( A301  and  (not A300) );
 a42429a <=( (not A299)  and  a42428a );
 a42430a <=( a42429a  and  a42424a );
 a42434a <=( (not A167)  and  A168 );
 a42435a <=( A169  and  a42434a );
 a42439a <=( A201  and  A200 );
 a42440a <=( A166  and  a42439a );
 a42441a <=( a42440a  and  a42435a );
 a42445a <=( A298  and  A267 );
 a42446a <=( A265  and  a42445a );
 a42450a <=( (not A302)  and  (not A300) );
 a42451a <=( (not A299)  and  a42450a );
 a42452a <=( a42451a  and  a42446a );
 a42456a <=( (not A167)  and  A168 );
 a42457a <=( A169  and  a42456a );
 a42461a <=( A201  and  A200 );
 a42462a <=( A166  and  a42461a );
 a42463a <=( a42462a  and  a42457a );
 a42467a <=( (not A298)  and  A267 );
 a42468a <=( A265  and  a42467a );
 a42472a <=( A301  and  (not A300) );
 a42473a <=( A299  and  a42472a );
 a42474a <=( a42473a  and  a42468a );
 a42478a <=( (not A167)  and  A168 );
 a42479a <=( A169  and  a42478a );
 a42483a <=( A201  and  A200 );
 a42484a <=( A166  and  a42483a );
 a42485a <=( a42484a  and  a42479a );
 a42489a <=( (not A298)  and  A267 );
 a42490a <=( A265  and  a42489a );
 a42494a <=( (not A302)  and  (not A300) );
 a42495a <=( A299  and  a42494a );
 a42496a <=( a42495a  and  a42490a );
 a42500a <=( (not A167)  and  A168 );
 a42501a <=( A169  and  a42500a );
 a42505a <=( A201  and  A200 );
 a42506a <=( A166  and  a42505a );
 a42507a <=( a42506a  and  a42501a );
 a42511a <=( A298  and  A267 );
 a42512a <=( A266  and  a42511a );
 a42516a <=( (not A301)  and  (not A300) );
 a42517a <=( A299  and  a42516a );
 a42518a <=( a42517a  and  a42512a );
 a42522a <=( (not A167)  and  A168 );
 a42523a <=( A169  and  a42522a );
 a42527a <=( A201  and  A200 );
 a42528a <=( A166  and  a42527a );
 a42529a <=( a42528a  and  a42523a );
 a42533a <=( A298  and  A267 );
 a42534a <=( A266  and  a42533a );
 a42538a <=( A302  and  (not A300) );
 a42539a <=( A299  and  a42538a );
 a42540a <=( a42539a  and  a42534a );
 a42544a <=( (not A167)  and  A168 );
 a42545a <=( A169  and  a42544a );
 a42549a <=( A201  and  A200 );
 a42550a <=( A166  and  a42549a );
 a42551a <=( a42550a  and  a42545a );
 a42555a <=( A298  and  A267 );
 a42556a <=( A266  and  a42555a );
 a42560a <=( A301  and  (not A300) );
 a42561a <=( (not A299)  and  a42560a );
 a42562a <=( a42561a  and  a42556a );
 a42566a <=( (not A167)  and  A168 );
 a42567a <=( A169  and  a42566a );
 a42571a <=( A201  and  A200 );
 a42572a <=( A166  and  a42571a );
 a42573a <=( a42572a  and  a42567a );
 a42577a <=( A298  and  A267 );
 a42578a <=( A266  and  a42577a );
 a42582a <=( (not A302)  and  (not A300) );
 a42583a <=( (not A299)  and  a42582a );
 a42584a <=( a42583a  and  a42578a );
 a42588a <=( (not A167)  and  A168 );
 a42589a <=( A169  and  a42588a );
 a42593a <=( A201  and  A200 );
 a42594a <=( A166  and  a42593a );
 a42595a <=( a42594a  and  a42589a );
 a42599a <=( (not A298)  and  A267 );
 a42600a <=( A266  and  a42599a );
 a42604a <=( A301  and  (not A300) );
 a42605a <=( A299  and  a42604a );
 a42606a <=( a42605a  and  a42600a );
 a42610a <=( (not A167)  and  A168 );
 a42611a <=( A169  and  a42610a );
 a42615a <=( A201  and  A200 );
 a42616a <=( A166  and  a42615a );
 a42617a <=( a42616a  and  a42611a );
 a42621a <=( (not A298)  and  A267 );
 a42622a <=( A266  and  a42621a );
 a42626a <=( (not A302)  and  (not A300) );
 a42627a <=( A299  and  a42626a );
 a42628a <=( a42627a  and  a42622a );
 a42632a <=( (not A167)  and  A168 );
 a42633a <=( A169  and  a42632a );
 a42637a <=( (not A200)  and  (not A199) );
 a42638a <=( A166  and  a42637a );
 a42639a <=( a42638a  and  a42633a );
 a42643a <=( (not A266)  and  (not A265) );
 a42644a <=( (not A202)  and  a42643a );
 a42648a <=( A300  and  A299 );
 a42649a <=( (not A268)  and  a42648a );
 a42650a <=( a42649a  and  a42644a );
 a42654a <=( (not A167)  and  A168 );
 a42655a <=( A169  and  a42654a );
 a42659a <=( (not A200)  and  (not A199) );
 a42660a <=( A166  and  a42659a );
 a42661a <=( a42660a  and  a42655a );
 a42665a <=( (not A266)  and  (not A265) );
 a42666a <=( (not A202)  and  a42665a );
 a42670a <=( A300  and  A298 );
 a42671a <=( (not A268)  and  a42670a );
 a42672a <=( a42671a  and  a42666a );
 a42676a <=( (not A167)  and  A168 );
 a42677a <=( A169  and  a42676a );
 a42681a <=( (not A200)  and  (not A199) );
 a42682a <=( A166  and  a42681a );
 a42683a <=( a42682a  and  a42677a );
 a42687a <=( (not A266)  and  (not A265) );
 a42688a <=( (not A202)  and  a42687a );
 a42692a <=( A300  and  A299 );
 a42693a <=( A269  and  a42692a );
 a42694a <=( a42693a  and  a42688a );
 a42698a <=( (not A167)  and  A168 );
 a42699a <=( A169  and  a42698a );
 a42703a <=( (not A200)  and  (not A199) );
 a42704a <=( A166  and  a42703a );
 a42705a <=( a42704a  and  a42699a );
 a42709a <=( (not A266)  and  (not A265) );
 a42710a <=( (not A202)  and  a42709a );
 a42714a <=( A300  and  A298 );
 a42715a <=( A269  and  a42714a );
 a42716a <=( a42715a  and  a42710a );
 a42720a <=( (not A167)  and  A168 );
 a42721a <=( A169  and  a42720a );
 a42725a <=( (not A200)  and  (not A199) );
 a42726a <=( A166  and  a42725a );
 a42727a <=( a42726a  and  a42721a );
 a42731a <=( (not A266)  and  (not A265) );
 a42732a <=( A203  and  a42731a );
 a42736a <=( A300  and  A299 );
 a42737a <=( (not A268)  and  a42736a );
 a42738a <=( a42737a  and  a42732a );
 a42742a <=( (not A167)  and  A168 );
 a42743a <=( A169  and  a42742a );
 a42747a <=( (not A200)  and  (not A199) );
 a42748a <=( A166  and  a42747a );
 a42749a <=( a42748a  and  a42743a );
 a42753a <=( (not A266)  and  (not A265) );
 a42754a <=( A203  and  a42753a );
 a42758a <=( A300  and  A298 );
 a42759a <=( (not A268)  and  a42758a );
 a42760a <=( a42759a  and  a42754a );
 a42764a <=( (not A167)  and  A168 );
 a42765a <=( A169  and  a42764a );
 a42769a <=( (not A200)  and  (not A199) );
 a42770a <=( A166  and  a42769a );
 a42771a <=( a42770a  and  a42765a );
 a42775a <=( (not A266)  and  (not A265) );
 a42776a <=( A203  and  a42775a );
 a42780a <=( A300  and  A299 );
 a42781a <=( A269  and  a42780a );
 a42782a <=( a42781a  and  a42776a );
 a42786a <=( (not A167)  and  A168 );
 a42787a <=( A169  and  a42786a );
 a42791a <=( (not A200)  and  (not A199) );
 a42792a <=( A166  and  a42791a );
 a42793a <=( a42792a  and  a42787a );
 a42797a <=( (not A266)  and  (not A265) );
 a42798a <=( A203  and  a42797a );
 a42802a <=( A300  and  A298 );
 a42803a <=( A269  and  a42802a );
 a42804a <=( a42803a  and  a42798a );
 a42808a <=( (not A167)  and  (not A169) );
 a42809a <=( (not A170)  and  a42808a );
 a42813a <=( (not A265)  and  A201 );
 a42814a <=( A199  and  a42813a );
 a42815a <=( a42814a  and  a42809a );
 a42819a <=( A298  and  (not A268) );
 a42820a <=( (not A266)  and  a42819a );
 a42824a <=( (not A302)  and  A301 );
 a42825a <=( A299  and  a42824a );
 a42826a <=( a42825a  and  a42820a );
 a42830a <=( (not A167)  and  (not A169) );
 a42831a <=( (not A170)  and  a42830a );
 a42835a <=( (not A265)  and  A201 );
 a42836a <=( A199  and  a42835a );
 a42837a <=( a42836a  and  a42831a );
 a42841a <=( A298  and  (not A268) );
 a42842a <=( (not A266)  and  a42841a );
 a42846a <=( A302  and  (not A301) );
 a42847a <=( (not A299)  and  a42846a );
 a42848a <=( a42847a  and  a42842a );
 a42852a <=( (not A167)  and  (not A169) );
 a42853a <=( (not A170)  and  a42852a );
 a42857a <=( (not A265)  and  A201 );
 a42858a <=( A199  and  a42857a );
 a42859a <=( a42858a  and  a42853a );
 a42863a <=( (not A298)  and  (not A268) );
 a42864a <=( (not A266)  and  a42863a );
 a42868a <=( A302  and  (not A301) );
 a42869a <=( A299  and  a42868a );
 a42870a <=( a42869a  and  a42864a );
 a42874a <=( (not A167)  and  (not A169) );
 a42875a <=( (not A170)  and  a42874a );
 a42879a <=( (not A265)  and  A201 );
 a42880a <=( A199  and  a42879a );
 a42881a <=( a42880a  and  a42875a );
 a42885a <=( (not A298)  and  (not A268) );
 a42886a <=( (not A266)  and  a42885a );
 a42890a <=( (not A302)  and  A301 );
 a42891a <=( (not A299)  and  a42890a );
 a42892a <=( a42891a  and  a42886a );
 a42896a <=( (not A167)  and  (not A169) );
 a42897a <=( (not A170)  and  a42896a );
 a42901a <=( (not A265)  and  A201 );
 a42902a <=( A199  and  a42901a );
 a42903a <=( a42902a  and  a42897a );
 a42907a <=( A298  and  A269 );
 a42908a <=( (not A266)  and  a42907a );
 a42912a <=( (not A302)  and  A301 );
 a42913a <=( A299  and  a42912a );
 a42914a <=( a42913a  and  a42908a );
 a42918a <=( (not A167)  and  (not A169) );
 a42919a <=( (not A170)  and  a42918a );
 a42923a <=( (not A265)  and  A201 );
 a42924a <=( A199  and  a42923a );
 a42925a <=( a42924a  and  a42919a );
 a42929a <=( A298  and  A269 );
 a42930a <=( (not A266)  and  a42929a );
 a42934a <=( A302  and  (not A301) );
 a42935a <=( (not A299)  and  a42934a );
 a42936a <=( a42935a  and  a42930a );
 a42940a <=( (not A167)  and  (not A169) );
 a42941a <=( (not A170)  and  a42940a );
 a42945a <=( (not A265)  and  A201 );
 a42946a <=( A199  and  a42945a );
 a42947a <=( a42946a  and  a42941a );
 a42951a <=( (not A298)  and  A269 );
 a42952a <=( (not A266)  and  a42951a );
 a42956a <=( A302  and  (not A301) );
 a42957a <=( A299  and  a42956a );
 a42958a <=( a42957a  and  a42952a );
 a42962a <=( (not A167)  and  (not A169) );
 a42963a <=( (not A170)  and  a42962a );
 a42967a <=( (not A265)  and  A201 );
 a42968a <=( A199  and  a42967a );
 a42969a <=( a42968a  and  a42963a );
 a42973a <=( (not A298)  and  A269 );
 a42974a <=( (not A266)  and  a42973a );
 a42978a <=( (not A302)  and  A301 );
 a42979a <=( (not A299)  and  a42978a );
 a42980a <=( a42979a  and  a42974a );
 a42984a <=( (not A167)  and  (not A169) );
 a42985a <=( (not A170)  and  a42984a );
 a42989a <=( (not A265)  and  A201 );
 a42990a <=( A200  and  a42989a );
 a42991a <=( a42990a  and  a42985a );
 a42995a <=( A298  and  (not A268) );
 a42996a <=( (not A266)  and  a42995a );
 a43000a <=( (not A302)  and  A301 );
 a43001a <=( A299  and  a43000a );
 a43002a <=( a43001a  and  a42996a );
 a43006a <=( (not A167)  and  (not A169) );
 a43007a <=( (not A170)  and  a43006a );
 a43011a <=( (not A265)  and  A201 );
 a43012a <=( A200  and  a43011a );
 a43013a <=( a43012a  and  a43007a );
 a43017a <=( A298  and  (not A268) );
 a43018a <=( (not A266)  and  a43017a );
 a43022a <=( A302  and  (not A301) );
 a43023a <=( (not A299)  and  a43022a );
 a43024a <=( a43023a  and  a43018a );
 a43028a <=( (not A167)  and  (not A169) );
 a43029a <=( (not A170)  and  a43028a );
 a43033a <=( (not A265)  and  A201 );
 a43034a <=( A200  and  a43033a );
 a43035a <=( a43034a  and  a43029a );
 a43039a <=( (not A298)  and  (not A268) );
 a43040a <=( (not A266)  and  a43039a );
 a43044a <=( A302  and  (not A301) );
 a43045a <=( A299  and  a43044a );
 a43046a <=( a43045a  and  a43040a );
 a43050a <=( (not A167)  and  (not A169) );
 a43051a <=( (not A170)  and  a43050a );
 a43055a <=( (not A265)  and  A201 );
 a43056a <=( A200  and  a43055a );
 a43057a <=( a43056a  and  a43051a );
 a43061a <=( (not A298)  and  (not A268) );
 a43062a <=( (not A266)  and  a43061a );
 a43066a <=( (not A302)  and  A301 );
 a43067a <=( (not A299)  and  a43066a );
 a43068a <=( a43067a  and  a43062a );
 a43072a <=( (not A167)  and  (not A169) );
 a43073a <=( (not A170)  and  a43072a );
 a43077a <=( (not A265)  and  A201 );
 a43078a <=( A200  and  a43077a );
 a43079a <=( a43078a  and  a43073a );
 a43083a <=( A298  and  A269 );
 a43084a <=( (not A266)  and  a43083a );
 a43088a <=( (not A302)  and  A301 );
 a43089a <=( A299  and  a43088a );
 a43090a <=( a43089a  and  a43084a );
 a43094a <=( (not A167)  and  (not A169) );
 a43095a <=( (not A170)  and  a43094a );
 a43099a <=( (not A265)  and  A201 );
 a43100a <=( A200  and  a43099a );
 a43101a <=( a43100a  and  a43095a );
 a43105a <=( A298  and  A269 );
 a43106a <=( (not A266)  and  a43105a );
 a43110a <=( A302  and  (not A301) );
 a43111a <=( (not A299)  and  a43110a );
 a43112a <=( a43111a  and  a43106a );
 a43116a <=( (not A167)  and  (not A169) );
 a43117a <=( (not A170)  and  a43116a );
 a43121a <=( (not A265)  and  A201 );
 a43122a <=( A200  and  a43121a );
 a43123a <=( a43122a  and  a43117a );
 a43127a <=( (not A298)  and  A269 );
 a43128a <=( (not A266)  and  a43127a );
 a43132a <=( A302  and  (not A301) );
 a43133a <=( A299  and  a43132a );
 a43134a <=( a43133a  and  a43128a );
 a43138a <=( (not A167)  and  (not A169) );
 a43139a <=( (not A170)  and  a43138a );
 a43143a <=( (not A265)  and  A201 );
 a43144a <=( A200  and  a43143a );
 a43145a <=( a43144a  and  a43139a );
 a43149a <=( (not A298)  and  A269 );
 a43150a <=( (not A266)  and  a43149a );
 a43154a <=( (not A302)  and  A301 );
 a43155a <=( (not A299)  and  a43154a );
 a43156a <=( a43155a  and  a43150a );
 a43160a <=( (not A167)  and  (not A169) );
 a43161a <=( (not A170)  and  a43160a );
 a43165a <=( A202  and  A200 );
 a43166a <=( A199  and  a43165a );
 a43167a <=( a43166a  and  a43161a );
 a43171a <=( (not A266)  and  (not A265) );
 a43172a <=( (not A203)  and  a43171a );
 a43176a <=( A300  and  A299 );
 a43177a <=( (not A268)  and  a43176a );
 a43178a <=( a43177a  and  a43172a );
 a43182a <=( (not A167)  and  (not A169) );
 a43183a <=( (not A170)  and  a43182a );
 a43187a <=( A202  and  A200 );
 a43188a <=( A199  and  a43187a );
 a43189a <=( a43188a  and  a43183a );
 a43193a <=( (not A266)  and  (not A265) );
 a43194a <=( (not A203)  and  a43193a );
 a43198a <=( A300  and  A298 );
 a43199a <=( (not A268)  and  a43198a );
 a43200a <=( a43199a  and  a43194a );
 a43204a <=( (not A167)  and  (not A169) );
 a43205a <=( (not A170)  and  a43204a );
 a43209a <=( A202  and  A200 );
 a43210a <=( A199  and  a43209a );
 a43211a <=( a43210a  and  a43205a );
 a43215a <=( (not A266)  and  (not A265) );
 a43216a <=( (not A203)  and  a43215a );
 a43220a <=( A300  and  A299 );
 a43221a <=( A269  and  a43220a );
 a43222a <=( a43221a  and  a43216a );
 a43226a <=( (not A167)  and  (not A169) );
 a43227a <=( (not A170)  and  a43226a );
 a43231a <=( A202  and  A200 );
 a43232a <=( A199  and  a43231a );
 a43233a <=( a43232a  and  a43227a );
 a43237a <=( (not A266)  and  (not A265) );
 a43238a <=( (not A203)  and  a43237a );
 a43242a <=( A300  and  A298 );
 a43243a <=( A269  and  a43242a );
 a43244a <=( a43243a  and  a43238a );
 a43248a <=( (not A167)  and  (not A169) );
 a43249a <=( (not A170)  and  a43248a );
 a43253a <=( (not A201)  and  A200 );
 a43254a <=( A199  and  a43253a );
 a43255a <=( a43254a  and  a43249a );
 a43259a <=( A267  and  A265 );
 a43260a <=( (not A202)  and  a43259a );
 a43264a <=( (not A301)  and  (not A299) );
 a43265a <=( (not A298)  and  a43264a );
 a43266a <=( a43265a  and  a43260a );
 a43270a <=( (not A167)  and  (not A169) );
 a43271a <=( (not A170)  and  a43270a );
 a43275a <=( (not A201)  and  A200 );
 a43276a <=( A199  and  a43275a );
 a43277a <=( a43276a  and  a43271a );
 a43281a <=( A267  and  A265 );
 a43282a <=( (not A202)  and  a43281a );
 a43286a <=( A302  and  (not A299) );
 a43287a <=( (not A298)  and  a43286a );
 a43288a <=( a43287a  and  a43282a );
 a43292a <=( (not A167)  and  (not A169) );
 a43293a <=( (not A170)  and  a43292a );
 a43297a <=( (not A201)  and  A200 );
 a43298a <=( A199  and  a43297a );
 a43299a <=( a43298a  and  a43293a );
 a43303a <=( A267  and  A266 );
 a43304a <=( (not A202)  and  a43303a );
 a43308a <=( (not A301)  and  (not A299) );
 a43309a <=( (not A298)  and  a43308a );
 a43310a <=( a43309a  and  a43304a );
 a43314a <=( (not A167)  and  (not A169) );
 a43315a <=( (not A170)  and  a43314a );
 a43319a <=( (not A201)  and  A200 );
 a43320a <=( A199  and  a43319a );
 a43321a <=( a43320a  and  a43315a );
 a43325a <=( A267  and  A266 );
 a43326a <=( (not A202)  and  a43325a );
 a43330a <=( A302  and  (not A299) );
 a43331a <=( (not A298)  and  a43330a );
 a43332a <=( a43331a  and  a43326a );
 a43336a <=( (not A167)  and  (not A169) );
 a43337a <=( (not A170)  and  a43336a );
 a43341a <=( (not A201)  and  A200 );
 a43342a <=( A199  and  a43341a );
 a43343a <=( a43342a  and  a43337a );
 a43347a <=( A267  and  A265 );
 a43348a <=( A203  and  a43347a );
 a43352a <=( (not A301)  and  (not A299) );
 a43353a <=( (not A298)  and  a43352a );
 a43354a <=( a43353a  and  a43348a );
 a43358a <=( (not A167)  and  (not A169) );
 a43359a <=( (not A170)  and  a43358a );
 a43363a <=( (not A201)  and  A200 );
 a43364a <=( A199  and  a43363a );
 a43365a <=( a43364a  and  a43359a );
 a43369a <=( A267  and  A265 );
 a43370a <=( A203  and  a43369a );
 a43374a <=( A302  and  (not A299) );
 a43375a <=( (not A298)  and  a43374a );
 a43376a <=( a43375a  and  a43370a );
 a43380a <=( (not A167)  and  (not A169) );
 a43381a <=( (not A170)  and  a43380a );
 a43385a <=( (not A201)  and  A200 );
 a43386a <=( A199  and  a43385a );
 a43387a <=( a43386a  and  a43381a );
 a43391a <=( A267  and  A266 );
 a43392a <=( A203  and  a43391a );
 a43396a <=( (not A301)  and  (not A299) );
 a43397a <=( (not A298)  and  a43396a );
 a43398a <=( a43397a  and  a43392a );
 a43402a <=( (not A167)  and  (not A169) );
 a43403a <=( (not A170)  and  a43402a );
 a43407a <=( (not A201)  and  A200 );
 a43408a <=( A199  and  a43407a );
 a43409a <=( a43408a  and  a43403a );
 a43413a <=( A267  and  A266 );
 a43414a <=( A203  and  a43413a );
 a43418a <=( A302  and  (not A299) );
 a43419a <=( (not A298)  and  a43418a );
 a43420a <=( a43419a  and  a43414a );
 a43424a <=( (not A167)  and  (not A169) );
 a43425a <=( (not A170)  and  a43424a );
 a43429a <=( (not A202)  and  A200 );
 a43430a <=( (not A199)  and  a43429a );
 a43431a <=( a43430a  and  a43425a );
 a43435a <=( (not A266)  and  (not A265) );
 a43436a <=( A203  and  a43435a );
 a43440a <=( A300  and  A299 );
 a43441a <=( (not A268)  and  a43440a );
 a43442a <=( a43441a  and  a43436a );
 a43446a <=( (not A167)  and  (not A169) );
 a43447a <=( (not A170)  and  a43446a );
 a43451a <=( (not A202)  and  A200 );
 a43452a <=( (not A199)  and  a43451a );
 a43453a <=( a43452a  and  a43447a );
 a43457a <=( (not A266)  and  (not A265) );
 a43458a <=( A203  and  a43457a );
 a43462a <=( A300  and  A298 );
 a43463a <=( (not A268)  and  a43462a );
 a43464a <=( a43463a  and  a43458a );
 a43468a <=( (not A167)  and  (not A169) );
 a43469a <=( (not A170)  and  a43468a );
 a43473a <=( (not A202)  and  A200 );
 a43474a <=( (not A199)  and  a43473a );
 a43475a <=( a43474a  and  a43469a );
 a43479a <=( (not A266)  and  (not A265) );
 a43480a <=( A203  and  a43479a );
 a43484a <=( A300  and  A299 );
 a43485a <=( A269  and  a43484a );
 a43486a <=( a43485a  and  a43480a );
 a43490a <=( (not A167)  and  (not A169) );
 a43491a <=( (not A170)  and  a43490a );
 a43495a <=( (not A202)  and  A200 );
 a43496a <=( (not A199)  and  a43495a );
 a43497a <=( a43496a  and  a43491a );
 a43501a <=( (not A266)  and  (not A265) );
 a43502a <=( A203  and  a43501a );
 a43506a <=( A300  and  A298 );
 a43507a <=( A269  and  a43506a );
 a43508a <=( a43507a  and  a43502a );
 a43512a <=( (not A167)  and  (not A169) );
 a43513a <=( (not A170)  and  a43512a );
 a43517a <=( (not A201)  and  A200 );
 a43518a <=( (not A199)  and  a43517a );
 a43519a <=( a43518a  and  a43513a );
 a43523a <=( A267  and  A265 );
 a43524a <=( A202  and  a43523a );
 a43528a <=( (not A301)  and  (not A299) );
 a43529a <=( (not A298)  and  a43528a );
 a43530a <=( a43529a  and  a43524a );
 a43534a <=( (not A167)  and  (not A169) );
 a43535a <=( (not A170)  and  a43534a );
 a43539a <=( (not A201)  and  A200 );
 a43540a <=( (not A199)  and  a43539a );
 a43541a <=( a43540a  and  a43535a );
 a43545a <=( A267  and  A265 );
 a43546a <=( A202  and  a43545a );
 a43550a <=( A302  and  (not A299) );
 a43551a <=( (not A298)  and  a43550a );
 a43552a <=( a43551a  and  a43546a );
 a43556a <=( (not A167)  and  (not A169) );
 a43557a <=( (not A170)  and  a43556a );
 a43561a <=( (not A201)  and  A200 );
 a43562a <=( (not A199)  and  a43561a );
 a43563a <=( a43562a  and  a43557a );
 a43567a <=( A267  and  A266 );
 a43568a <=( A202  and  a43567a );
 a43572a <=( (not A301)  and  (not A299) );
 a43573a <=( (not A298)  and  a43572a );
 a43574a <=( a43573a  and  a43568a );
 a43578a <=( (not A167)  and  (not A169) );
 a43579a <=( (not A170)  and  a43578a );
 a43583a <=( (not A201)  and  A200 );
 a43584a <=( (not A199)  and  a43583a );
 a43585a <=( a43584a  and  a43579a );
 a43589a <=( A267  and  A266 );
 a43590a <=( A202  and  a43589a );
 a43594a <=( A302  and  (not A299) );
 a43595a <=( (not A298)  and  a43594a );
 a43596a <=( a43595a  and  a43590a );
 a43600a <=( (not A167)  and  (not A169) );
 a43601a <=( (not A170)  and  a43600a );
 a43605a <=( (not A201)  and  A200 );
 a43606a <=( (not A199)  and  a43605a );
 a43607a <=( a43606a  and  a43601a );
 a43611a <=( A267  and  A265 );
 a43612a <=( (not A203)  and  a43611a );
 a43616a <=( (not A301)  and  (not A299) );
 a43617a <=( (not A298)  and  a43616a );
 a43618a <=( a43617a  and  a43612a );
 a43622a <=( (not A167)  and  (not A169) );
 a43623a <=( (not A170)  and  a43622a );
 a43627a <=( (not A201)  and  A200 );
 a43628a <=( (not A199)  and  a43627a );
 a43629a <=( a43628a  and  a43623a );
 a43633a <=( A267  and  A265 );
 a43634a <=( (not A203)  and  a43633a );
 a43638a <=( A302  and  (not A299) );
 a43639a <=( (not A298)  and  a43638a );
 a43640a <=( a43639a  and  a43634a );
 a43644a <=( (not A167)  and  (not A169) );
 a43645a <=( (not A170)  and  a43644a );
 a43649a <=( (not A201)  and  A200 );
 a43650a <=( (not A199)  and  a43649a );
 a43651a <=( a43650a  and  a43645a );
 a43655a <=( A267  and  A266 );
 a43656a <=( (not A203)  and  a43655a );
 a43660a <=( (not A301)  and  (not A299) );
 a43661a <=( (not A298)  and  a43660a );
 a43662a <=( a43661a  and  a43656a );
 a43666a <=( (not A167)  and  (not A169) );
 a43667a <=( (not A170)  and  a43666a );
 a43671a <=( (not A201)  and  A200 );
 a43672a <=( (not A199)  and  a43671a );
 a43673a <=( a43672a  and  a43667a );
 a43677a <=( A267  and  A266 );
 a43678a <=( (not A203)  and  a43677a );
 a43682a <=( A302  and  (not A299) );
 a43683a <=( (not A298)  and  a43682a );
 a43684a <=( a43683a  and  a43678a );
 a43688a <=( (not A167)  and  (not A169) );
 a43689a <=( (not A170)  and  a43688a );
 a43693a <=( (not A202)  and  (not A200) );
 a43694a <=( A199  and  a43693a );
 a43695a <=( a43694a  and  a43689a );
 a43699a <=( (not A266)  and  (not A265) );
 a43700a <=( A203  and  a43699a );
 a43704a <=( A300  and  A299 );
 a43705a <=( (not A268)  and  a43704a );
 a43706a <=( a43705a  and  a43700a );
 a43710a <=( (not A167)  and  (not A169) );
 a43711a <=( (not A170)  and  a43710a );
 a43715a <=( (not A202)  and  (not A200) );
 a43716a <=( A199  and  a43715a );
 a43717a <=( a43716a  and  a43711a );
 a43721a <=( (not A266)  and  (not A265) );
 a43722a <=( A203  and  a43721a );
 a43726a <=( A300  and  A298 );
 a43727a <=( (not A268)  and  a43726a );
 a43728a <=( a43727a  and  a43722a );
 a43732a <=( (not A167)  and  (not A169) );
 a43733a <=( (not A170)  and  a43732a );
 a43737a <=( (not A202)  and  (not A200) );
 a43738a <=( A199  and  a43737a );
 a43739a <=( a43738a  and  a43733a );
 a43743a <=( (not A266)  and  (not A265) );
 a43744a <=( A203  and  a43743a );
 a43748a <=( A300  and  A299 );
 a43749a <=( A269  and  a43748a );
 a43750a <=( a43749a  and  a43744a );
 a43754a <=( (not A167)  and  (not A169) );
 a43755a <=( (not A170)  and  a43754a );
 a43759a <=( (not A202)  and  (not A200) );
 a43760a <=( A199  and  a43759a );
 a43761a <=( a43760a  and  a43755a );
 a43765a <=( (not A266)  and  (not A265) );
 a43766a <=( A203  and  a43765a );
 a43770a <=( A300  and  A298 );
 a43771a <=( A269  and  a43770a );
 a43772a <=( a43771a  and  a43766a );
 a43776a <=( (not A167)  and  (not A169) );
 a43777a <=( (not A170)  and  a43776a );
 a43781a <=( (not A201)  and  (not A200) );
 a43782a <=( A199  and  a43781a );
 a43783a <=( a43782a  and  a43777a );
 a43787a <=( A267  and  A265 );
 a43788a <=( A202  and  a43787a );
 a43792a <=( (not A301)  and  (not A299) );
 a43793a <=( (not A298)  and  a43792a );
 a43794a <=( a43793a  and  a43788a );
 a43798a <=( (not A167)  and  (not A169) );
 a43799a <=( (not A170)  and  a43798a );
 a43803a <=( (not A201)  and  (not A200) );
 a43804a <=( A199  and  a43803a );
 a43805a <=( a43804a  and  a43799a );
 a43809a <=( A267  and  A265 );
 a43810a <=( A202  and  a43809a );
 a43814a <=( A302  and  (not A299) );
 a43815a <=( (not A298)  and  a43814a );
 a43816a <=( a43815a  and  a43810a );
 a43820a <=( (not A167)  and  (not A169) );
 a43821a <=( (not A170)  and  a43820a );
 a43825a <=( (not A201)  and  (not A200) );
 a43826a <=( A199  and  a43825a );
 a43827a <=( a43826a  and  a43821a );
 a43831a <=( A267  and  A266 );
 a43832a <=( A202  and  a43831a );
 a43836a <=( (not A301)  and  (not A299) );
 a43837a <=( (not A298)  and  a43836a );
 a43838a <=( a43837a  and  a43832a );
 a43842a <=( (not A167)  and  (not A169) );
 a43843a <=( (not A170)  and  a43842a );
 a43847a <=( (not A201)  and  (not A200) );
 a43848a <=( A199  and  a43847a );
 a43849a <=( a43848a  and  a43843a );
 a43853a <=( A267  and  A266 );
 a43854a <=( A202  and  a43853a );
 a43858a <=( A302  and  (not A299) );
 a43859a <=( (not A298)  and  a43858a );
 a43860a <=( a43859a  and  a43854a );
 a43864a <=( (not A167)  and  (not A169) );
 a43865a <=( (not A170)  and  a43864a );
 a43869a <=( (not A201)  and  (not A200) );
 a43870a <=( A199  and  a43869a );
 a43871a <=( a43870a  and  a43865a );
 a43875a <=( A267  and  A265 );
 a43876a <=( (not A203)  and  a43875a );
 a43880a <=( (not A301)  and  (not A299) );
 a43881a <=( (not A298)  and  a43880a );
 a43882a <=( a43881a  and  a43876a );
 a43886a <=( (not A167)  and  (not A169) );
 a43887a <=( (not A170)  and  a43886a );
 a43891a <=( (not A201)  and  (not A200) );
 a43892a <=( A199  and  a43891a );
 a43893a <=( a43892a  and  a43887a );
 a43897a <=( A267  and  A265 );
 a43898a <=( (not A203)  and  a43897a );
 a43902a <=( A302  and  (not A299) );
 a43903a <=( (not A298)  and  a43902a );
 a43904a <=( a43903a  and  a43898a );
 a43908a <=( (not A167)  and  (not A169) );
 a43909a <=( (not A170)  and  a43908a );
 a43913a <=( (not A201)  and  (not A200) );
 a43914a <=( A199  and  a43913a );
 a43915a <=( a43914a  and  a43909a );
 a43919a <=( A267  and  A266 );
 a43920a <=( (not A203)  and  a43919a );
 a43924a <=( (not A301)  and  (not A299) );
 a43925a <=( (not A298)  and  a43924a );
 a43926a <=( a43925a  and  a43920a );
 a43930a <=( (not A167)  and  (not A169) );
 a43931a <=( (not A170)  and  a43930a );
 a43935a <=( (not A201)  and  (not A200) );
 a43936a <=( A199  and  a43935a );
 a43937a <=( a43936a  and  a43931a );
 a43941a <=( A267  and  A266 );
 a43942a <=( (not A203)  and  a43941a );
 a43946a <=( A302  and  (not A299) );
 a43947a <=( (not A298)  and  a43946a );
 a43948a <=( a43947a  and  a43942a );
 a43952a <=( (not A167)  and  (not A169) );
 a43953a <=( (not A170)  and  a43952a );
 a43957a <=( (not A202)  and  (not A200) );
 a43958a <=( (not A199)  and  a43957a );
 a43959a <=( a43958a  and  a43953a );
 a43963a <=( A298  and  A267 );
 a43964a <=( A265  and  a43963a );
 a43968a <=( (not A301)  and  (not A300) );
 a43969a <=( A299  and  a43968a );
 a43970a <=( a43969a  and  a43964a );
 a43974a <=( (not A167)  and  (not A169) );
 a43975a <=( (not A170)  and  a43974a );
 a43979a <=( (not A202)  and  (not A200) );
 a43980a <=( (not A199)  and  a43979a );
 a43981a <=( a43980a  and  a43975a );
 a43985a <=( A298  and  A267 );
 a43986a <=( A265  and  a43985a );
 a43990a <=( A302  and  (not A300) );
 a43991a <=( A299  and  a43990a );
 a43992a <=( a43991a  and  a43986a );
 a43996a <=( (not A167)  and  (not A169) );
 a43997a <=( (not A170)  and  a43996a );
 a44001a <=( (not A202)  and  (not A200) );
 a44002a <=( (not A199)  and  a44001a );
 a44003a <=( a44002a  and  a43997a );
 a44007a <=( A298  and  A267 );
 a44008a <=( A265  and  a44007a );
 a44012a <=( A301  and  (not A300) );
 a44013a <=( (not A299)  and  a44012a );
 a44014a <=( a44013a  and  a44008a );
 a44018a <=( (not A167)  and  (not A169) );
 a44019a <=( (not A170)  and  a44018a );
 a44023a <=( (not A202)  and  (not A200) );
 a44024a <=( (not A199)  and  a44023a );
 a44025a <=( a44024a  and  a44019a );
 a44029a <=( A298  and  A267 );
 a44030a <=( A265  and  a44029a );
 a44034a <=( (not A302)  and  (not A300) );
 a44035a <=( (not A299)  and  a44034a );
 a44036a <=( a44035a  and  a44030a );
 a44040a <=( (not A167)  and  (not A169) );
 a44041a <=( (not A170)  and  a44040a );
 a44045a <=( (not A202)  and  (not A200) );
 a44046a <=( (not A199)  and  a44045a );
 a44047a <=( a44046a  and  a44041a );
 a44051a <=( (not A298)  and  A267 );
 a44052a <=( A265  and  a44051a );
 a44056a <=( A301  and  (not A300) );
 a44057a <=( A299  and  a44056a );
 a44058a <=( a44057a  and  a44052a );
 a44062a <=( (not A167)  and  (not A169) );
 a44063a <=( (not A170)  and  a44062a );
 a44067a <=( (not A202)  and  (not A200) );
 a44068a <=( (not A199)  and  a44067a );
 a44069a <=( a44068a  and  a44063a );
 a44073a <=( (not A298)  and  A267 );
 a44074a <=( A265  and  a44073a );
 a44078a <=( (not A302)  and  (not A300) );
 a44079a <=( A299  and  a44078a );
 a44080a <=( a44079a  and  a44074a );
 a44084a <=( (not A167)  and  (not A169) );
 a44085a <=( (not A170)  and  a44084a );
 a44089a <=( (not A202)  and  (not A200) );
 a44090a <=( (not A199)  and  a44089a );
 a44091a <=( a44090a  and  a44085a );
 a44095a <=( A298  and  A267 );
 a44096a <=( A266  and  a44095a );
 a44100a <=( (not A301)  and  (not A300) );
 a44101a <=( A299  and  a44100a );
 a44102a <=( a44101a  and  a44096a );
 a44106a <=( (not A167)  and  (not A169) );
 a44107a <=( (not A170)  and  a44106a );
 a44111a <=( (not A202)  and  (not A200) );
 a44112a <=( (not A199)  and  a44111a );
 a44113a <=( a44112a  and  a44107a );
 a44117a <=( A298  and  A267 );
 a44118a <=( A266  and  a44117a );
 a44122a <=( A302  and  (not A300) );
 a44123a <=( A299  and  a44122a );
 a44124a <=( a44123a  and  a44118a );
 a44128a <=( (not A167)  and  (not A169) );
 a44129a <=( (not A170)  and  a44128a );
 a44133a <=( (not A202)  and  (not A200) );
 a44134a <=( (not A199)  and  a44133a );
 a44135a <=( a44134a  and  a44129a );
 a44139a <=( A298  and  A267 );
 a44140a <=( A266  and  a44139a );
 a44144a <=( A301  and  (not A300) );
 a44145a <=( (not A299)  and  a44144a );
 a44146a <=( a44145a  and  a44140a );
 a44150a <=( (not A167)  and  (not A169) );
 a44151a <=( (not A170)  and  a44150a );
 a44155a <=( (not A202)  and  (not A200) );
 a44156a <=( (not A199)  and  a44155a );
 a44157a <=( a44156a  and  a44151a );
 a44161a <=( A298  and  A267 );
 a44162a <=( A266  and  a44161a );
 a44166a <=( (not A302)  and  (not A300) );
 a44167a <=( (not A299)  and  a44166a );
 a44168a <=( a44167a  and  a44162a );
 a44172a <=( (not A167)  and  (not A169) );
 a44173a <=( (not A170)  and  a44172a );
 a44177a <=( (not A202)  and  (not A200) );
 a44178a <=( (not A199)  and  a44177a );
 a44179a <=( a44178a  and  a44173a );
 a44183a <=( (not A298)  and  A267 );
 a44184a <=( A266  and  a44183a );
 a44188a <=( A301  and  (not A300) );
 a44189a <=( A299  and  a44188a );
 a44190a <=( a44189a  and  a44184a );
 a44194a <=( (not A167)  and  (not A169) );
 a44195a <=( (not A170)  and  a44194a );
 a44199a <=( (not A202)  and  (not A200) );
 a44200a <=( (not A199)  and  a44199a );
 a44201a <=( a44200a  and  a44195a );
 a44205a <=( (not A298)  and  A267 );
 a44206a <=( A266  and  a44205a );
 a44210a <=( (not A302)  and  (not A300) );
 a44211a <=( A299  and  a44210a );
 a44212a <=( a44211a  and  a44206a );
 a44216a <=( (not A167)  and  (not A169) );
 a44217a <=( (not A170)  and  a44216a );
 a44221a <=( A203  and  (not A200) );
 a44222a <=( (not A199)  and  a44221a );
 a44223a <=( a44222a  and  a44217a );
 a44227a <=( A298  and  A267 );
 a44228a <=( A265  and  a44227a );
 a44232a <=( (not A301)  and  (not A300) );
 a44233a <=( A299  and  a44232a );
 a44234a <=( a44233a  and  a44228a );
 a44238a <=( (not A167)  and  (not A169) );
 a44239a <=( (not A170)  and  a44238a );
 a44243a <=( A203  and  (not A200) );
 a44244a <=( (not A199)  and  a44243a );
 a44245a <=( a44244a  and  a44239a );
 a44249a <=( A298  and  A267 );
 a44250a <=( A265  and  a44249a );
 a44254a <=( A302  and  (not A300) );
 a44255a <=( A299  and  a44254a );
 a44256a <=( a44255a  and  a44250a );
 a44260a <=( (not A167)  and  (not A169) );
 a44261a <=( (not A170)  and  a44260a );
 a44265a <=( A203  and  (not A200) );
 a44266a <=( (not A199)  and  a44265a );
 a44267a <=( a44266a  and  a44261a );
 a44271a <=( A298  and  A267 );
 a44272a <=( A265  and  a44271a );
 a44276a <=( A301  and  (not A300) );
 a44277a <=( (not A299)  and  a44276a );
 a44278a <=( a44277a  and  a44272a );
 a44282a <=( (not A167)  and  (not A169) );
 a44283a <=( (not A170)  and  a44282a );
 a44287a <=( A203  and  (not A200) );
 a44288a <=( (not A199)  and  a44287a );
 a44289a <=( a44288a  and  a44283a );
 a44293a <=( A298  and  A267 );
 a44294a <=( A265  and  a44293a );
 a44298a <=( (not A302)  and  (not A300) );
 a44299a <=( (not A299)  and  a44298a );
 a44300a <=( a44299a  and  a44294a );
 a44304a <=( (not A167)  and  (not A169) );
 a44305a <=( (not A170)  and  a44304a );
 a44309a <=( A203  and  (not A200) );
 a44310a <=( (not A199)  and  a44309a );
 a44311a <=( a44310a  and  a44305a );
 a44315a <=( (not A298)  and  A267 );
 a44316a <=( A265  and  a44315a );
 a44320a <=( A301  and  (not A300) );
 a44321a <=( A299  and  a44320a );
 a44322a <=( a44321a  and  a44316a );
 a44326a <=( (not A167)  and  (not A169) );
 a44327a <=( (not A170)  and  a44326a );
 a44331a <=( A203  and  (not A200) );
 a44332a <=( (not A199)  and  a44331a );
 a44333a <=( a44332a  and  a44327a );
 a44337a <=( (not A298)  and  A267 );
 a44338a <=( A265  and  a44337a );
 a44342a <=( (not A302)  and  (not A300) );
 a44343a <=( A299  and  a44342a );
 a44344a <=( a44343a  and  a44338a );
 a44348a <=( (not A167)  and  (not A169) );
 a44349a <=( (not A170)  and  a44348a );
 a44353a <=( A203  and  (not A200) );
 a44354a <=( (not A199)  and  a44353a );
 a44355a <=( a44354a  and  a44349a );
 a44359a <=( A298  and  A267 );
 a44360a <=( A266  and  a44359a );
 a44364a <=( (not A301)  and  (not A300) );
 a44365a <=( A299  and  a44364a );
 a44366a <=( a44365a  and  a44360a );
 a44370a <=( (not A167)  and  (not A169) );
 a44371a <=( (not A170)  and  a44370a );
 a44375a <=( A203  and  (not A200) );
 a44376a <=( (not A199)  and  a44375a );
 a44377a <=( a44376a  and  a44371a );
 a44381a <=( A298  and  A267 );
 a44382a <=( A266  and  a44381a );
 a44386a <=( A302  and  (not A300) );
 a44387a <=( A299  and  a44386a );
 a44388a <=( a44387a  and  a44382a );
 a44392a <=( (not A167)  and  (not A169) );
 a44393a <=( (not A170)  and  a44392a );
 a44397a <=( A203  and  (not A200) );
 a44398a <=( (not A199)  and  a44397a );
 a44399a <=( a44398a  and  a44393a );
 a44403a <=( A298  and  A267 );
 a44404a <=( A266  and  a44403a );
 a44408a <=( A301  and  (not A300) );
 a44409a <=( (not A299)  and  a44408a );
 a44410a <=( a44409a  and  a44404a );
 a44414a <=( (not A167)  and  (not A169) );
 a44415a <=( (not A170)  and  a44414a );
 a44419a <=( A203  and  (not A200) );
 a44420a <=( (not A199)  and  a44419a );
 a44421a <=( a44420a  and  a44415a );
 a44425a <=( A298  and  A267 );
 a44426a <=( A266  and  a44425a );
 a44430a <=( (not A302)  and  (not A300) );
 a44431a <=( (not A299)  and  a44430a );
 a44432a <=( a44431a  and  a44426a );
 a44436a <=( (not A167)  and  (not A169) );
 a44437a <=( (not A170)  and  a44436a );
 a44441a <=( A203  and  (not A200) );
 a44442a <=( (not A199)  and  a44441a );
 a44443a <=( a44442a  and  a44437a );
 a44447a <=( (not A298)  and  A267 );
 a44448a <=( A266  and  a44447a );
 a44452a <=( A301  and  (not A300) );
 a44453a <=( A299  and  a44452a );
 a44454a <=( a44453a  and  a44448a );
 a44458a <=( (not A167)  and  (not A169) );
 a44459a <=( (not A170)  and  a44458a );
 a44463a <=( A203  and  (not A200) );
 a44464a <=( (not A199)  and  a44463a );
 a44465a <=( a44464a  and  a44459a );
 a44469a <=( (not A298)  and  A267 );
 a44470a <=( A266  and  a44469a );
 a44474a <=( (not A302)  and  (not A300) );
 a44475a <=( A299  and  a44474a );
 a44476a <=( a44475a  and  a44470a );
 a44480a <=( (not A167)  and  (not A169) );
 a44481a <=( (not A170)  and  a44480a );
 a44485a <=( A202  and  (not A200) );
 a44486a <=( (not A199)  and  a44485a );
 a44487a <=( a44486a  and  a44481a );
 a44491a <=( (not A266)  and  (not A265) );
 a44492a <=( (not A203)  and  a44491a );
 a44496a <=( A300  and  A299 );
 a44497a <=( (not A268)  and  a44496a );
 a44498a <=( a44497a  and  a44492a );
 a44502a <=( (not A167)  and  (not A169) );
 a44503a <=( (not A170)  and  a44502a );
 a44507a <=( A202  and  (not A200) );
 a44508a <=( (not A199)  and  a44507a );
 a44509a <=( a44508a  and  a44503a );
 a44513a <=( (not A266)  and  (not A265) );
 a44514a <=( (not A203)  and  a44513a );
 a44518a <=( A300  and  A298 );
 a44519a <=( (not A268)  and  a44518a );
 a44520a <=( a44519a  and  a44514a );
 a44524a <=( (not A167)  and  (not A169) );
 a44525a <=( (not A170)  and  a44524a );
 a44529a <=( A202  and  (not A200) );
 a44530a <=( (not A199)  and  a44529a );
 a44531a <=( a44530a  and  a44525a );
 a44535a <=( (not A266)  and  (not A265) );
 a44536a <=( (not A203)  and  a44535a );
 a44540a <=( A300  and  A299 );
 a44541a <=( A269  and  a44540a );
 a44542a <=( a44541a  and  a44536a );
 a44546a <=( (not A167)  and  (not A169) );
 a44547a <=( (not A170)  and  a44546a );
 a44551a <=( A202  and  (not A200) );
 a44552a <=( (not A199)  and  a44551a );
 a44553a <=( a44552a  and  a44547a );
 a44557a <=( (not A266)  and  (not A265) );
 a44558a <=( (not A203)  and  a44557a );
 a44562a <=( A300  and  A298 );
 a44563a <=( A269  and  a44562a );
 a44564a <=( a44563a  and  a44558a );
 a44568a <=( A199  and  A166 );
 a44569a <=( A167  and  a44568a );
 a44573a <=( (not A203)  and  A202 );
 a44574a <=( A200  and  a44573a );
 a44575a <=( a44574a  and  a44569a );
 a44579a <=( (not A268)  and  (not A266) );
 a44580a <=( (not A265)  and  a44579a );
 a44583a <=( A299  and  A298 );
 a44586a <=( (not A302)  and  A301 );
 a44587a <=( a44586a  and  a44583a );
 a44588a <=( a44587a  and  a44580a );
 a44592a <=( A199  and  A166 );
 a44593a <=( A167  and  a44592a );
 a44597a <=( (not A203)  and  A202 );
 a44598a <=( A200  and  a44597a );
 a44599a <=( a44598a  and  a44593a );
 a44603a <=( (not A268)  and  (not A266) );
 a44604a <=( (not A265)  and  a44603a );
 a44607a <=( (not A299)  and  A298 );
 a44610a <=( A302  and  (not A301) );
 a44611a <=( a44610a  and  a44607a );
 a44612a <=( a44611a  and  a44604a );
 a44616a <=( A199  and  A166 );
 a44617a <=( A167  and  a44616a );
 a44621a <=( (not A203)  and  A202 );
 a44622a <=( A200  and  a44621a );
 a44623a <=( a44622a  and  a44617a );
 a44627a <=( (not A268)  and  (not A266) );
 a44628a <=( (not A265)  and  a44627a );
 a44631a <=( A299  and  (not A298) );
 a44634a <=( A302  and  (not A301) );
 a44635a <=( a44634a  and  a44631a );
 a44636a <=( a44635a  and  a44628a );
 a44640a <=( A199  and  A166 );
 a44641a <=( A167  and  a44640a );
 a44645a <=( (not A203)  and  A202 );
 a44646a <=( A200  and  a44645a );
 a44647a <=( a44646a  and  a44641a );
 a44651a <=( (not A268)  and  (not A266) );
 a44652a <=( (not A265)  and  a44651a );
 a44655a <=( (not A299)  and  (not A298) );
 a44658a <=( (not A302)  and  A301 );
 a44659a <=( a44658a  and  a44655a );
 a44660a <=( a44659a  and  a44652a );
 a44664a <=( A199  and  A166 );
 a44665a <=( A167  and  a44664a );
 a44669a <=( (not A203)  and  A202 );
 a44670a <=( A200  and  a44669a );
 a44671a <=( a44670a  and  a44665a );
 a44675a <=( A269  and  (not A266) );
 a44676a <=( (not A265)  and  a44675a );
 a44679a <=( A299  and  A298 );
 a44682a <=( (not A302)  and  A301 );
 a44683a <=( a44682a  and  a44679a );
 a44684a <=( a44683a  and  a44676a );
 a44688a <=( A199  and  A166 );
 a44689a <=( A167  and  a44688a );
 a44693a <=( (not A203)  and  A202 );
 a44694a <=( A200  and  a44693a );
 a44695a <=( a44694a  and  a44689a );
 a44699a <=( A269  and  (not A266) );
 a44700a <=( (not A265)  and  a44699a );
 a44703a <=( (not A299)  and  A298 );
 a44706a <=( A302  and  (not A301) );
 a44707a <=( a44706a  and  a44703a );
 a44708a <=( a44707a  and  a44700a );
 a44712a <=( A199  and  A166 );
 a44713a <=( A167  and  a44712a );
 a44717a <=( (not A203)  and  A202 );
 a44718a <=( A200  and  a44717a );
 a44719a <=( a44718a  and  a44713a );
 a44723a <=( A269  and  (not A266) );
 a44724a <=( (not A265)  and  a44723a );
 a44727a <=( A299  and  (not A298) );
 a44730a <=( A302  and  (not A301) );
 a44731a <=( a44730a  and  a44727a );
 a44732a <=( a44731a  and  a44724a );
 a44736a <=( A199  and  A166 );
 a44737a <=( A167  and  a44736a );
 a44741a <=( (not A203)  and  A202 );
 a44742a <=( A200  and  a44741a );
 a44743a <=( a44742a  and  a44737a );
 a44747a <=( A269  and  (not A266) );
 a44748a <=( (not A265)  and  a44747a );
 a44751a <=( (not A299)  and  (not A298) );
 a44754a <=( (not A302)  and  A301 );
 a44755a <=( a44754a  and  a44751a );
 a44756a <=( a44755a  and  a44748a );
 a44760a <=( A199  and  A166 );
 a44761a <=( A167  and  a44760a );
 a44765a <=( (not A202)  and  (not A201) );
 a44766a <=( A200  and  a44765a );
 a44767a <=( a44766a  and  a44761a );
 a44771a <=( A268  and  A266 );
 a44772a <=( A265  and  a44771a );
 a44775a <=( (not A298)  and  (not A269) );
 a44778a <=( (not A301)  and  (not A299) );
 a44779a <=( a44778a  and  a44775a );
 a44780a <=( a44779a  and  a44772a );
 a44784a <=( A199  and  A166 );
 a44785a <=( A167  and  a44784a );
 a44789a <=( (not A202)  and  (not A201) );
 a44790a <=( A200  and  a44789a );
 a44791a <=( a44790a  and  a44785a );
 a44795a <=( A268  and  A266 );
 a44796a <=( A265  and  a44795a );
 a44799a <=( (not A298)  and  (not A269) );
 a44802a <=( A302  and  (not A299) );
 a44803a <=( a44802a  and  a44799a );
 a44804a <=( a44803a  and  a44796a );
 a44808a <=( A199  and  A166 );
 a44809a <=( A167  and  a44808a );
 a44813a <=( (not A202)  and  (not A201) );
 a44814a <=( A200  and  a44813a );
 a44815a <=( a44814a  and  a44809a );
 a44819a <=( (not A268)  and  A266 );
 a44820a <=( (not A265)  and  a44819a );
 a44823a <=( (not A298)  and  A269 );
 a44826a <=( (not A301)  and  (not A299) );
 a44827a <=( a44826a  and  a44823a );
 a44828a <=( a44827a  and  a44820a );
 a44832a <=( A199  and  A166 );
 a44833a <=( A167  and  a44832a );
 a44837a <=( (not A202)  and  (not A201) );
 a44838a <=( A200  and  a44837a );
 a44839a <=( a44838a  and  a44833a );
 a44843a <=( (not A268)  and  A266 );
 a44844a <=( (not A265)  and  a44843a );
 a44847a <=( (not A298)  and  A269 );
 a44850a <=( A302  and  (not A299) );
 a44851a <=( a44850a  and  a44847a );
 a44852a <=( a44851a  and  a44844a );
 a44856a <=( A199  and  A166 );
 a44857a <=( A167  and  a44856a );
 a44861a <=( (not A202)  and  (not A201) );
 a44862a <=( A200  and  a44861a );
 a44863a <=( a44862a  and  a44857a );
 a44867a <=( (not A268)  and  (not A266) );
 a44868a <=( A265  and  a44867a );
 a44871a <=( (not A298)  and  A269 );
 a44874a <=( (not A301)  and  (not A299) );
 a44875a <=( a44874a  and  a44871a );
 a44876a <=( a44875a  and  a44868a );
 a44880a <=( A199  and  A166 );
 a44881a <=( A167  and  a44880a );
 a44885a <=( (not A202)  and  (not A201) );
 a44886a <=( A200  and  a44885a );
 a44887a <=( a44886a  and  a44881a );
 a44891a <=( (not A268)  and  (not A266) );
 a44892a <=( A265  and  a44891a );
 a44895a <=( (not A298)  and  A269 );
 a44898a <=( A302  and  (not A299) );
 a44899a <=( a44898a  and  a44895a );
 a44900a <=( a44899a  and  a44892a );
 a44904a <=( A199  and  A166 );
 a44905a <=( A167  and  a44904a );
 a44909a <=( (not A202)  and  (not A201) );
 a44910a <=( A200  and  a44909a );
 a44911a <=( a44910a  and  a44905a );
 a44915a <=( A268  and  (not A266) );
 a44916a <=( (not A265)  and  a44915a );
 a44919a <=( (not A298)  and  (not A269) );
 a44922a <=( (not A301)  and  (not A299) );
 a44923a <=( a44922a  and  a44919a );
 a44924a <=( a44923a  and  a44916a );
 a44928a <=( A199  and  A166 );
 a44929a <=( A167  and  a44928a );
 a44933a <=( (not A202)  and  (not A201) );
 a44934a <=( A200  and  a44933a );
 a44935a <=( a44934a  and  a44929a );
 a44939a <=( A268  and  (not A266) );
 a44940a <=( (not A265)  and  a44939a );
 a44943a <=( (not A298)  and  (not A269) );
 a44946a <=( A302  and  (not A299) );
 a44947a <=( a44946a  and  a44943a );
 a44948a <=( a44947a  and  a44940a );
 a44952a <=( A199  and  A166 );
 a44953a <=( A167  and  a44952a );
 a44957a <=( A203  and  (not A201) );
 a44958a <=( A200  and  a44957a );
 a44959a <=( a44958a  and  a44953a );
 a44963a <=( A268  and  A266 );
 a44964a <=( A265  and  a44963a );
 a44967a <=( (not A298)  and  (not A269) );
 a44970a <=( (not A301)  and  (not A299) );
 a44971a <=( a44970a  and  a44967a );
 a44972a <=( a44971a  and  a44964a );
 a44976a <=( A199  and  A166 );
 a44977a <=( A167  and  a44976a );
 a44981a <=( A203  and  (not A201) );
 a44982a <=( A200  and  a44981a );
 a44983a <=( a44982a  and  a44977a );
 a44987a <=( A268  and  A266 );
 a44988a <=( A265  and  a44987a );
 a44991a <=( (not A298)  and  (not A269) );
 a44994a <=( A302  and  (not A299) );
 a44995a <=( a44994a  and  a44991a );
 a44996a <=( a44995a  and  a44988a );
 a45000a <=( A199  and  A166 );
 a45001a <=( A167  and  a45000a );
 a45005a <=( A203  and  (not A201) );
 a45006a <=( A200  and  a45005a );
 a45007a <=( a45006a  and  a45001a );
 a45011a <=( (not A268)  and  A266 );
 a45012a <=( (not A265)  and  a45011a );
 a45015a <=( (not A298)  and  A269 );
 a45018a <=( (not A301)  and  (not A299) );
 a45019a <=( a45018a  and  a45015a );
 a45020a <=( a45019a  and  a45012a );
 a45024a <=( A199  and  A166 );
 a45025a <=( A167  and  a45024a );
 a45029a <=( A203  and  (not A201) );
 a45030a <=( A200  and  a45029a );
 a45031a <=( a45030a  and  a45025a );
 a45035a <=( (not A268)  and  A266 );
 a45036a <=( (not A265)  and  a45035a );
 a45039a <=( (not A298)  and  A269 );
 a45042a <=( A302  and  (not A299) );
 a45043a <=( a45042a  and  a45039a );
 a45044a <=( a45043a  and  a45036a );
 a45048a <=( A199  and  A166 );
 a45049a <=( A167  and  a45048a );
 a45053a <=( A203  and  (not A201) );
 a45054a <=( A200  and  a45053a );
 a45055a <=( a45054a  and  a45049a );
 a45059a <=( (not A268)  and  (not A266) );
 a45060a <=( A265  and  a45059a );
 a45063a <=( (not A298)  and  A269 );
 a45066a <=( (not A301)  and  (not A299) );
 a45067a <=( a45066a  and  a45063a );
 a45068a <=( a45067a  and  a45060a );
 a45072a <=( A199  and  A166 );
 a45073a <=( A167  and  a45072a );
 a45077a <=( A203  and  (not A201) );
 a45078a <=( A200  and  a45077a );
 a45079a <=( a45078a  and  a45073a );
 a45083a <=( (not A268)  and  (not A266) );
 a45084a <=( A265  and  a45083a );
 a45087a <=( (not A298)  and  A269 );
 a45090a <=( A302  and  (not A299) );
 a45091a <=( a45090a  and  a45087a );
 a45092a <=( a45091a  and  a45084a );
 a45096a <=( A199  and  A166 );
 a45097a <=( A167  and  a45096a );
 a45101a <=( A203  and  (not A201) );
 a45102a <=( A200  and  a45101a );
 a45103a <=( a45102a  and  a45097a );
 a45107a <=( A268  and  (not A266) );
 a45108a <=( (not A265)  and  a45107a );
 a45111a <=( (not A298)  and  (not A269) );
 a45114a <=( (not A301)  and  (not A299) );
 a45115a <=( a45114a  and  a45111a );
 a45116a <=( a45115a  and  a45108a );
 a45120a <=( A199  and  A166 );
 a45121a <=( A167  and  a45120a );
 a45125a <=( A203  and  (not A201) );
 a45126a <=( A200  and  a45125a );
 a45127a <=( a45126a  and  a45121a );
 a45131a <=( A268  and  (not A266) );
 a45132a <=( (not A265)  and  a45131a );
 a45135a <=( (not A298)  and  (not A269) );
 a45138a <=( A302  and  (not A299) );
 a45139a <=( a45138a  and  a45135a );
 a45140a <=( a45139a  and  a45132a );
 a45144a <=( (not A199)  and  A166 );
 a45145a <=( A167  and  a45144a );
 a45149a <=( A203  and  (not A202) );
 a45150a <=( A200  and  a45149a );
 a45151a <=( a45150a  and  a45145a );
 a45155a <=( (not A268)  and  (not A266) );
 a45156a <=( (not A265)  and  a45155a );
 a45159a <=( A299  and  A298 );
 a45162a <=( (not A302)  and  A301 );
 a45163a <=( a45162a  and  a45159a );
 a45164a <=( a45163a  and  a45156a );
 a45168a <=( (not A199)  and  A166 );
 a45169a <=( A167  and  a45168a );
 a45173a <=( A203  and  (not A202) );
 a45174a <=( A200  and  a45173a );
 a45175a <=( a45174a  and  a45169a );
 a45179a <=( (not A268)  and  (not A266) );
 a45180a <=( (not A265)  and  a45179a );
 a45183a <=( (not A299)  and  A298 );
 a45186a <=( A302  and  (not A301) );
 a45187a <=( a45186a  and  a45183a );
 a45188a <=( a45187a  and  a45180a );
 a45192a <=( (not A199)  and  A166 );
 a45193a <=( A167  and  a45192a );
 a45197a <=( A203  and  (not A202) );
 a45198a <=( A200  and  a45197a );
 a45199a <=( a45198a  and  a45193a );
 a45203a <=( (not A268)  and  (not A266) );
 a45204a <=( (not A265)  and  a45203a );
 a45207a <=( A299  and  (not A298) );
 a45210a <=( A302  and  (not A301) );
 a45211a <=( a45210a  and  a45207a );
 a45212a <=( a45211a  and  a45204a );
 a45216a <=( (not A199)  and  A166 );
 a45217a <=( A167  and  a45216a );
 a45221a <=( A203  and  (not A202) );
 a45222a <=( A200  and  a45221a );
 a45223a <=( a45222a  and  a45217a );
 a45227a <=( (not A268)  and  (not A266) );
 a45228a <=( (not A265)  and  a45227a );
 a45231a <=( (not A299)  and  (not A298) );
 a45234a <=( (not A302)  and  A301 );
 a45235a <=( a45234a  and  a45231a );
 a45236a <=( a45235a  and  a45228a );
 a45240a <=( (not A199)  and  A166 );
 a45241a <=( A167  and  a45240a );
 a45245a <=( A203  and  (not A202) );
 a45246a <=( A200  and  a45245a );
 a45247a <=( a45246a  and  a45241a );
 a45251a <=( A269  and  (not A266) );
 a45252a <=( (not A265)  and  a45251a );
 a45255a <=( A299  and  A298 );
 a45258a <=( (not A302)  and  A301 );
 a45259a <=( a45258a  and  a45255a );
 a45260a <=( a45259a  and  a45252a );
 a45264a <=( (not A199)  and  A166 );
 a45265a <=( A167  and  a45264a );
 a45269a <=( A203  and  (not A202) );
 a45270a <=( A200  and  a45269a );
 a45271a <=( a45270a  and  a45265a );
 a45275a <=( A269  and  (not A266) );
 a45276a <=( (not A265)  and  a45275a );
 a45279a <=( (not A299)  and  A298 );
 a45282a <=( A302  and  (not A301) );
 a45283a <=( a45282a  and  a45279a );
 a45284a <=( a45283a  and  a45276a );
 a45288a <=( (not A199)  and  A166 );
 a45289a <=( A167  and  a45288a );
 a45293a <=( A203  and  (not A202) );
 a45294a <=( A200  and  a45293a );
 a45295a <=( a45294a  and  a45289a );
 a45299a <=( A269  and  (not A266) );
 a45300a <=( (not A265)  and  a45299a );
 a45303a <=( A299  and  (not A298) );
 a45306a <=( A302  and  (not A301) );
 a45307a <=( a45306a  and  a45303a );
 a45308a <=( a45307a  and  a45300a );
 a45312a <=( (not A199)  and  A166 );
 a45313a <=( A167  and  a45312a );
 a45317a <=( A203  and  (not A202) );
 a45318a <=( A200  and  a45317a );
 a45319a <=( a45318a  and  a45313a );
 a45323a <=( A269  and  (not A266) );
 a45324a <=( (not A265)  and  a45323a );
 a45327a <=( (not A299)  and  (not A298) );
 a45330a <=( (not A302)  and  A301 );
 a45331a <=( a45330a  and  a45327a );
 a45332a <=( a45331a  and  a45324a );
 a45336a <=( (not A199)  and  A166 );
 a45337a <=( A167  and  a45336a );
 a45341a <=( A202  and  (not A201) );
 a45342a <=( A200  and  a45341a );
 a45343a <=( a45342a  and  a45337a );
 a45347a <=( A268  and  A266 );
 a45348a <=( A265  and  a45347a );
 a45351a <=( (not A298)  and  (not A269) );
 a45354a <=( (not A301)  and  (not A299) );
 a45355a <=( a45354a  and  a45351a );
 a45356a <=( a45355a  and  a45348a );
 a45360a <=( (not A199)  and  A166 );
 a45361a <=( A167  and  a45360a );
 a45365a <=( A202  and  (not A201) );
 a45366a <=( A200  and  a45365a );
 a45367a <=( a45366a  and  a45361a );
 a45371a <=( A268  and  A266 );
 a45372a <=( A265  and  a45371a );
 a45375a <=( (not A298)  and  (not A269) );
 a45378a <=( A302  and  (not A299) );
 a45379a <=( a45378a  and  a45375a );
 a45380a <=( a45379a  and  a45372a );
 a45384a <=( (not A199)  and  A166 );
 a45385a <=( A167  and  a45384a );
 a45389a <=( A202  and  (not A201) );
 a45390a <=( A200  and  a45389a );
 a45391a <=( a45390a  and  a45385a );
 a45395a <=( (not A268)  and  A266 );
 a45396a <=( (not A265)  and  a45395a );
 a45399a <=( (not A298)  and  A269 );
 a45402a <=( (not A301)  and  (not A299) );
 a45403a <=( a45402a  and  a45399a );
 a45404a <=( a45403a  and  a45396a );
 a45408a <=( (not A199)  and  A166 );
 a45409a <=( A167  and  a45408a );
 a45413a <=( A202  and  (not A201) );
 a45414a <=( A200  and  a45413a );
 a45415a <=( a45414a  and  a45409a );
 a45419a <=( (not A268)  and  A266 );
 a45420a <=( (not A265)  and  a45419a );
 a45423a <=( (not A298)  and  A269 );
 a45426a <=( A302  and  (not A299) );
 a45427a <=( a45426a  and  a45423a );
 a45428a <=( a45427a  and  a45420a );
 a45432a <=( (not A199)  and  A166 );
 a45433a <=( A167  and  a45432a );
 a45437a <=( A202  and  (not A201) );
 a45438a <=( A200  and  a45437a );
 a45439a <=( a45438a  and  a45433a );
 a45443a <=( (not A268)  and  (not A266) );
 a45444a <=( A265  and  a45443a );
 a45447a <=( (not A298)  and  A269 );
 a45450a <=( (not A301)  and  (not A299) );
 a45451a <=( a45450a  and  a45447a );
 a45452a <=( a45451a  and  a45444a );
 a45456a <=( (not A199)  and  A166 );
 a45457a <=( A167  and  a45456a );
 a45461a <=( A202  and  (not A201) );
 a45462a <=( A200  and  a45461a );
 a45463a <=( a45462a  and  a45457a );
 a45467a <=( (not A268)  and  (not A266) );
 a45468a <=( A265  and  a45467a );
 a45471a <=( (not A298)  and  A269 );
 a45474a <=( A302  and  (not A299) );
 a45475a <=( a45474a  and  a45471a );
 a45476a <=( a45475a  and  a45468a );
 a45480a <=( (not A199)  and  A166 );
 a45481a <=( A167  and  a45480a );
 a45485a <=( A202  and  (not A201) );
 a45486a <=( A200  and  a45485a );
 a45487a <=( a45486a  and  a45481a );
 a45491a <=( A268  and  (not A266) );
 a45492a <=( (not A265)  and  a45491a );
 a45495a <=( (not A298)  and  (not A269) );
 a45498a <=( (not A301)  and  (not A299) );
 a45499a <=( a45498a  and  a45495a );
 a45500a <=( a45499a  and  a45492a );
 a45504a <=( (not A199)  and  A166 );
 a45505a <=( A167  and  a45504a );
 a45509a <=( A202  and  (not A201) );
 a45510a <=( A200  and  a45509a );
 a45511a <=( a45510a  and  a45505a );
 a45515a <=( A268  and  (not A266) );
 a45516a <=( (not A265)  and  a45515a );
 a45519a <=( (not A298)  and  (not A269) );
 a45522a <=( A302  and  (not A299) );
 a45523a <=( a45522a  and  a45519a );
 a45524a <=( a45523a  and  a45516a );
 a45528a <=( (not A199)  and  A166 );
 a45529a <=( A167  and  a45528a );
 a45533a <=( (not A203)  and  (not A201) );
 a45534a <=( A200  and  a45533a );
 a45535a <=( a45534a  and  a45529a );
 a45539a <=( A268  and  A266 );
 a45540a <=( A265  and  a45539a );
 a45543a <=( (not A298)  and  (not A269) );
 a45546a <=( (not A301)  and  (not A299) );
 a45547a <=( a45546a  and  a45543a );
 a45548a <=( a45547a  and  a45540a );
 a45552a <=( (not A199)  and  A166 );
 a45553a <=( A167  and  a45552a );
 a45557a <=( (not A203)  and  (not A201) );
 a45558a <=( A200  and  a45557a );
 a45559a <=( a45558a  and  a45553a );
 a45563a <=( A268  and  A266 );
 a45564a <=( A265  and  a45563a );
 a45567a <=( (not A298)  and  (not A269) );
 a45570a <=( A302  and  (not A299) );
 a45571a <=( a45570a  and  a45567a );
 a45572a <=( a45571a  and  a45564a );
 a45576a <=( (not A199)  and  A166 );
 a45577a <=( A167  and  a45576a );
 a45581a <=( (not A203)  and  (not A201) );
 a45582a <=( A200  and  a45581a );
 a45583a <=( a45582a  and  a45577a );
 a45587a <=( (not A268)  and  A266 );
 a45588a <=( (not A265)  and  a45587a );
 a45591a <=( (not A298)  and  A269 );
 a45594a <=( (not A301)  and  (not A299) );
 a45595a <=( a45594a  and  a45591a );
 a45596a <=( a45595a  and  a45588a );
 a45600a <=( (not A199)  and  A166 );
 a45601a <=( A167  and  a45600a );
 a45605a <=( (not A203)  and  (not A201) );
 a45606a <=( A200  and  a45605a );
 a45607a <=( a45606a  and  a45601a );
 a45611a <=( (not A268)  and  A266 );
 a45612a <=( (not A265)  and  a45611a );
 a45615a <=( (not A298)  and  A269 );
 a45618a <=( A302  and  (not A299) );
 a45619a <=( a45618a  and  a45615a );
 a45620a <=( a45619a  and  a45612a );
 a45624a <=( (not A199)  and  A166 );
 a45625a <=( A167  and  a45624a );
 a45629a <=( (not A203)  and  (not A201) );
 a45630a <=( A200  and  a45629a );
 a45631a <=( a45630a  and  a45625a );
 a45635a <=( (not A268)  and  (not A266) );
 a45636a <=( A265  and  a45635a );
 a45639a <=( (not A298)  and  A269 );
 a45642a <=( (not A301)  and  (not A299) );
 a45643a <=( a45642a  and  a45639a );
 a45644a <=( a45643a  and  a45636a );
 a45648a <=( (not A199)  and  A166 );
 a45649a <=( A167  and  a45648a );
 a45653a <=( (not A203)  and  (not A201) );
 a45654a <=( A200  and  a45653a );
 a45655a <=( a45654a  and  a45649a );
 a45659a <=( (not A268)  and  (not A266) );
 a45660a <=( A265  and  a45659a );
 a45663a <=( (not A298)  and  A269 );
 a45666a <=( A302  and  (not A299) );
 a45667a <=( a45666a  and  a45663a );
 a45668a <=( a45667a  and  a45660a );
 a45672a <=( (not A199)  and  A166 );
 a45673a <=( A167  and  a45672a );
 a45677a <=( (not A203)  and  (not A201) );
 a45678a <=( A200  and  a45677a );
 a45679a <=( a45678a  and  a45673a );
 a45683a <=( A268  and  (not A266) );
 a45684a <=( (not A265)  and  a45683a );
 a45687a <=( (not A298)  and  (not A269) );
 a45690a <=( (not A301)  and  (not A299) );
 a45691a <=( a45690a  and  a45687a );
 a45692a <=( a45691a  and  a45684a );
 a45696a <=( (not A199)  and  A166 );
 a45697a <=( A167  and  a45696a );
 a45701a <=( (not A203)  and  (not A201) );
 a45702a <=( A200  and  a45701a );
 a45703a <=( a45702a  and  a45697a );
 a45707a <=( A268  and  (not A266) );
 a45708a <=( (not A265)  and  a45707a );
 a45711a <=( (not A298)  and  (not A269) );
 a45714a <=( A302  and  (not A299) );
 a45715a <=( a45714a  and  a45711a );
 a45716a <=( a45715a  and  a45708a );
 a45720a <=( A199  and  A166 );
 a45721a <=( A167  and  a45720a );
 a45725a <=( A203  and  (not A202) );
 a45726a <=( (not A200)  and  a45725a );
 a45727a <=( a45726a  and  a45721a );
 a45731a <=( (not A268)  and  (not A266) );
 a45732a <=( (not A265)  and  a45731a );
 a45735a <=( A299  and  A298 );
 a45738a <=( (not A302)  and  A301 );
 a45739a <=( a45738a  and  a45735a );
 a45740a <=( a45739a  and  a45732a );
 a45744a <=( A199  and  A166 );
 a45745a <=( A167  and  a45744a );
 a45749a <=( A203  and  (not A202) );
 a45750a <=( (not A200)  and  a45749a );
 a45751a <=( a45750a  and  a45745a );
 a45755a <=( (not A268)  and  (not A266) );
 a45756a <=( (not A265)  and  a45755a );
 a45759a <=( (not A299)  and  A298 );
 a45762a <=( A302  and  (not A301) );
 a45763a <=( a45762a  and  a45759a );
 a45764a <=( a45763a  and  a45756a );
 a45768a <=( A199  and  A166 );
 a45769a <=( A167  and  a45768a );
 a45773a <=( A203  and  (not A202) );
 a45774a <=( (not A200)  and  a45773a );
 a45775a <=( a45774a  and  a45769a );
 a45779a <=( (not A268)  and  (not A266) );
 a45780a <=( (not A265)  and  a45779a );
 a45783a <=( A299  and  (not A298) );
 a45786a <=( A302  and  (not A301) );
 a45787a <=( a45786a  and  a45783a );
 a45788a <=( a45787a  and  a45780a );
 a45792a <=( A199  and  A166 );
 a45793a <=( A167  and  a45792a );
 a45797a <=( A203  and  (not A202) );
 a45798a <=( (not A200)  and  a45797a );
 a45799a <=( a45798a  and  a45793a );
 a45803a <=( (not A268)  and  (not A266) );
 a45804a <=( (not A265)  and  a45803a );
 a45807a <=( (not A299)  and  (not A298) );
 a45810a <=( (not A302)  and  A301 );
 a45811a <=( a45810a  and  a45807a );
 a45812a <=( a45811a  and  a45804a );
 a45816a <=( A199  and  A166 );
 a45817a <=( A167  and  a45816a );
 a45821a <=( A203  and  (not A202) );
 a45822a <=( (not A200)  and  a45821a );
 a45823a <=( a45822a  and  a45817a );
 a45827a <=( A269  and  (not A266) );
 a45828a <=( (not A265)  and  a45827a );
 a45831a <=( A299  and  A298 );
 a45834a <=( (not A302)  and  A301 );
 a45835a <=( a45834a  and  a45831a );
 a45836a <=( a45835a  and  a45828a );
 a45840a <=( A199  and  A166 );
 a45841a <=( A167  and  a45840a );
 a45845a <=( A203  and  (not A202) );
 a45846a <=( (not A200)  and  a45845a );
 a45847a <=( a45846a  and  a45841a );
 a45851a <=( A269  and  (not A266) );
 a45852a <=( (not A265)  and  a45851a );
 a45855a <=( (not A299)  and  A298 );
 a45858a <=( A302  and  (not A301) );
 a45859a <=( a45858a  and  a45855a );
 a45860a <=( a45859a  and  a45852a );
 a45864a <=( A199  and  A166 );
 a45865a <=( A167  and  a45864a );
 a45869a <=( A203  and  (not A202) );
 a45870a <=( (not A200)  and  a45869a );
 a45871a <=( a45870a  and  a45865a );
 a45875a <=( A269  and  (not A266) );
 a45876a <=( (not A265)  and  a45875a );
 a45879a <=( A299  and  (not A298) );
 a45882a <=( A302  and  (not A301) );
 a45883a <=( a45882a  and  a45879a );
 a45884a <=( a45883a  and  a45876a );
 a45888a <=( A199  and  A166 );
 a45889a <=( A167  and  a45888a );
 a45893a <=( A203  and  (not A202) );
 a45894a <=( (not A200)  and  a45893a );
 a45895a <=( a45894a  and  a45889a );
 a45899a <=( A269  and  (not A266) );
 a45900a <=( (not A265)  and  a45899a );
 a45903a <=( (not A299)  and  (not A298) );
 a45906a <=( (not A302)  and  A301 );
 a45907a <=( a45906a  and  a45903a );
 a45908a <=( a45907a  and  a45900a );
 a45912a <=( A199  and  A166 );
 a45913a <=( A167  and  a45912a );
 a45917a <=( A202  and  (not A201) );
 a45918a <=( (not A200)  and  a45917a );
 a45919a <=( a45918a  and  a45913a );
 a45923a <=( A268  and  A266 );
 a45924a <=( A265  and  a45923a );
 a45927a <=( (not A298)  and  (not A269) );
 a45930a <=( (not A301)  and  (not A299) );
 a45931a <=( a45930a  and  a45927a );
 a45932a <=( a45931a  and  a45924a );
 a45936a <=( A199  and  A166 );
 a45937a <=( A167  and  a45936a );
 a45941a <=( A202  and  (not A201) );
 a45942a <=( (not A200)  and  a45941a );
 a45943a <=( a45942a  and  a45937a );
 a45947a <=( A268  and  A266 );
 a45948a <=( A265  and  a45947a );
 a45951a <=( (not A298)  and  (not A269) );
 a45954a <=( A302  and  (not A299) );
 a45955a <=( a45954a  and  a45951a );
 a45956a <=( a45955a  and  a45948a );
 a45960a <=( A199  and  A166 );
 a45961a <=( A167  and  a45960a );
 a45965a <=( A202  and  (not A201) );
 a45966a <=( (not A200)  and  a45965a );
 a45967a <=( a45966a  and  a45961a );
 a45971a <=( (not A268)  and  A266 );
 a45972a <=( (not A265)  and  a45971a );
 a45975a <=( (not A298)  and  A269 );
 a45978a <=( (not A301)  and  (not A299) );
 a45979a <=( a45978a  and  a45975a );
 a45980a <=( a45979a  and  a45972a );
 a45984a <=( A199  and  A166 );
 a45985a <=( A167  and  a45984a );
 a45989a <=( A202  and  (not A201) );
 a45990a <=( (not A200)  and  a45989a );
 a45991a <=( a45990a  and  a45985a );
 a45995a <=( (not A268)  and  A266 );
 a45996a <=( (not A265)  and  a45995a );
 a45999a <=( (not A298)  and  A269 );
 a46002a <=( A302  and  (not A299) );
 a46003a <=( a46002a  and  a45999a );
 a46004a <=( a46003a  and  a45996a );
 a46008a <=( A199  and  A166 );
 a46009a <=( A167  and  a46008a );
 a46013a <=( A202  and  (not A201) );
 a46014a <=( (not A200)  and  a46013a );
 a46015a <=( a46014a  and  a46009a );
 a46019a <=( (not A268)  and  (not A266) );
 a46020a <=( A265  and  a46019a );
 a46023a <=( (not A298)  and  A269 );
 a46026a <=( (not A301)  and  (not A299) );
 a46027a <=( a46026a  and  a46023a );
 a46028a <=( a46027a  and  a46020a );
 a46032a <=( A199  and  A166 );
 a46033a <=( A167  and  a46032a );
 a46037a <=( A202  and  (not A201) );
 a46038a <=( (not A200)  and  a46037a );
 a46039a <=( a46038a  and  a46033a );
 a46043a <=( (not A268)  and  (not A266) );
 a46044a <=( A265  and  a46043a );
 a46047a <=( (not A298)  and  A269 );
 a46050a <=( A302  and  (not A299) );
 a46051a <=( a46050a  and  a46047a );
 a46052a <=( a46051a  and  a46044a );
 a46056a <=( A199  and  A166 );
 a46057a <=( A167  and  a46056a );
 a46061a <=( A202  and  (not A201) );
 a46062a <=( (not A200)  and  a46061a );
 a46063a <=( a46062a  and  a46057a );
 a46067a <=( A268  and  (not A266) );
 a46068a <=( (not A265)  and  a46067a );
 a46071a <=( (not A298)  and  (not A269) );
 a46074a <=( (not A301)  and  (not A299) );
 a46075a <=( a46074a  and  a46071a );
 a46076a <=( a46075a  and  a46068a );
 a46080a <=( A199  and  A166 );
 a46081a <=( A167  and  a46080a );
 a46085a <=( A202  and  (not A201) );
 a46086a <=( (not A200)  and  a46085a );
 a46087a <=( a46086a  and  a46081a );
 a46091a <=( A268  and  (not A266) );
 a46092a <=( (not A265)  and  a46091a );
 a46095a <=( (not A298)  and  (not A269) );
 a46098a <=( A302  and  (not A299) );
 a46099a <=( a46098a  and  a46095a );
 a46100a <=( a46099a  and  a46092a );
 a46104a <=( A199  and  A166 );
 a46105a <=( A167  and  a46104a );
 a46109a <=( (not A203)  and  (not A201) );
 a46110a <=( (not A200)  and  a46109a );
 a46111a <=( a46110a  and  a46105a );
 a46115a <=( A268  and  A266 );
 a46116a <=( A265  and  a46115a );
 a46119a <=( (not A298)  and  (not A269) );
 a46122a <=( (not A301)  and  (not A299) );
 a46123a <=( a46122a  and  a46119a );
 a46124a <=( a46123a  and  a46116a );
 a46128a <=( A199  and  A166 );
 a46129a <=( A167  and  a46128a );
 a46133a <=( (not A203)  and  (not A201) );
 a46134a <=( (not A200)  and  a46133a );
 a46135a <=( a46134a  and  a46129a );
 a46139a <=( A268  and  A266 );
 a46140a <=( A265  and  a46139a );
 a46143a <=( (not A298)  and  (not A269) );
 a46146a <=( A302  and  (not A299) );
 a46147a <=( a46146a  and  a46143a );
 a46148a <=( a46147a  and  a46140a );
 a46152a <=( A199  and  A166 );
 a46153a <=( A167  and  a46152a );
 a46157a <=( (not A203)  and  (not A201) );
 a46158a <=( (not A200)  and  a46157a );
 a46159a <=( a46158a  and  a46153a );
 a46163a <=( (not A268)  and  A266 );
 a46164a <=( (not A265)  and  a46163a );
 a46167a <=( (not A298)  and  A269 );
 a46170a <=( (not A301)  and  (not A299) );
 a46171a <=( a46170a  and  a46167a );
 a46172a <=( a46171a  and  a46164a );
 a46176a <=( A199  and  A166 );
 a46177a <=( A167  and  a46176a );
 a46181a <=( (not A203)  and  (not A201) );
 a46182a <=( (not A200)  and  a46181a );
 a46183a <=( a46182a  and  a46177a );
 a46187a <=( (not A268)  and  A266 );
 a46188a <=( (not A265)  and  a46187a );
 a46191a <=( (not A298)  and  A269 );
 a46194a <=( A302  and  (not A299) );
 a46195a <=( a46194a  and  a46191a );
 a46196a <=( a46195a  and  a46188a );
 a46200a <=( A199  and  A166 );
 a46201a <=( A167  and  a46200a );
 a46205a <=( (not A203)  and  (not A201) );
 a46206a <=( (not A200)  and  a46205a );
 a46207a <=( a46206a  and  a46201a );
 a46211a <=( (not A268)  and  (not A266) );
 a46212a <=( A265  and  a46211a );
 a46215a <=( (not A298)  and  A269 );
 a46218a <=( (not A301)  and  (not A299) );
 a46219a <=( a46218a  and  a46215a );
 a46220a <=( a46219a  and  a46212a );
 a46224a <=( A199  and  A166 );
 a46225a <=( A167  and  a46224a );
 a46229a <=( (not A203)  and  (not A201) );
 a46230a <=( (not A200)  and  a46229a );
 a46231a <=( a46230a  and  a46225a );
 a46235a <=( (not A268)  and  (not A266) );
 a46236a <=( A265  and  a46235a );
 a46239a <=( (not A298)  and  A269 );
 a46242a <=( A302  and  (not A299) );
 a46243a <=( a46242a  and  a46239a );
 a46244a <=( a46243a  and  a46236a );
 a46248a <=( A199  and  A166 );
 a46249a <=( A167  and  a46248a );
 a46253a <=( (not A203)  and  (not A201) );
 a46254a <=( (not A200)  and  a46253a );
 a46255a <=( a46254a  and  a46249a );
 a46259a <=( A268  and  (not A266) );
 a46260a <=( (not A265)  and  a46259a );
 a46263a <=( (not A298)  and  (not A269) );
 a46266a <=( (not A301)  and  (not A299) );
 a46267a <=( a46266a  and  a46263a );
 a46268a <=( a46267a  and  a46260a );
 a46272a <=( A199  and  A166 );
 a46273a <=( A167  and  a46272a );
 a46277a <=( (not A203)  and  (not A201) );
 a46278a <=( (not A200)  and  a46277a );
 a46279a <=( a46278a  and  a46273a );
 a46283a <=( A268  and  (not A266) );
 a46284a <=( (not A265)  and  a46283a );
 a46287a <=( (not A298)  and  (not A269) );
 a46290a <=( A302  and  (not A299) );
 a46291a <=( a46290a  and  a46287a );
 a46292a <=( a46291a  and  a46284a );
 a46296a <=( (not A199)  and  A166 );
 a46297a <=( A167  and  a46296a );
 a46301a <=( A265  and  (not A202) );
 a46302a <=( (not A200)  and  a46301a );
 a46303a <=( a46302a  and  a46297a );
 a46307a <=( (not A269)  and  A268 );
 a46308a <=( A266  and  a46307a );
 a46311a <=( A299  and  A298 );
 a46314a <=( (not A301)  and  (not A300) );
 a46315a <=( a46314a  and  a46311a );
 a46316a <=( a46315a  and  a46308a );
 a46320a <=( (not A199)  and  A166 );
 a46321a <=( A167  and  a46320a );
 a46325a <=( A265  and  (not A202) );
 a46326a <=( (not A200)  and  a46325a );
 a46327a <=( a46326a  and  a46321a );
 a46331a <=( (not A269)  and  A268 );
 a46332a <=( A266  and  a46331a );
 a46335a <=( A299  and  A298 );
 a46338a <=( A302  and  (not A300) );
 a46339a <=( a46338a  and  a46335a );
 a46340a <=( a46339a  and  a46332a );
 a46344a <=( (not A199)  and  A166 );
 a46345a <=( A167  and  a46344a );
 a46349a <=( A265  and  (not A202) );
 a46350a <=( (not A200)  and  a46349a );
 a46351a <=( a46350a  and  a46345a );
 a46355a <=( (not A269)  and  A268 );
 a46356a <=( A266  and  a46355a );
 a46359a <=( (not A299)  and  A298 );
 a46362a <=( A301  and  (not A300) );
 a46363a <=( a46362a  and  a46359a );
 a46364a <=( a46363a  and  a46356a );
 a46368a <=( (not A199)  and  A166 );
 a46369a <=( A167  and  a46368a );
 a46373a <=( A265  and  (not A202) );
 a46374a <=( (not A200)  and  a46373a );
 a46375a <=( a46374a  and  a46369a );
 a46379a <=( (not A269)  and  A268 );
 a46380a <=( A266  and  a46379a );
 a46383a <=( (not A299)  and  A298 );
 a46386a <=( (not A302)  and  (not A300) );
 a46387a <=( a46386a  and  a46383a );
 a46388a <=( a46387a  and  a46380a );
 a46392a <=( (not A199)  and  A166 );
 a46393a <=( A167  and  a46392a );
 a46397a <=( A265  and  (not A202) );
 a46398a <=( (not A200)  and  a46397a );
 a46399a <=( a46398a  and  a46393a );
 a46403a <=( (not A269)  and  A268 );
 a46404a <=( A266  and  a46403a );
 a46407a <=( A299  and  (not A298) );
 a46410a <=( A301  and  (not A300) );
 a46411a <=( a46410a  and  a46407a );
 a46412a <=( a46411a  and  a46404a );
 a46416a <=( (not A199)  and  A166 );
 a46417a <=( A167  and  a46416a );
 a46421a <=( A265  and  (not A202) );
 a46422a <=( (not A200)  and  a46421a );
 a46423a <=( a46422a  and  a46417a );
 a46427a <=( (not A269)  and  A268 );
 a46428a <=( A266  and  a46427a );
 a46431a <=( A299  and  (not A298) );
 a46434a <=( (not A302)  and  (not A300) );
 a46435a <=( a46434a  and  a46431a );
 a46436a <=( a46435a  and  a46428a );
 a46440a <=( (not A199)  and  A166 );
 a46441a <=( A167  and  a46440a );
 a46445a <=( (not A265)  and  (not A202) );
 a46446a <=( (not A200)  and  a46445a );
 a46447a <=( a46446a  and  a46441a );
 a46451a <=( A269  and  (not A268) );
 a46452a <=( A266  and  a46451a );
 a46455a <=( A299  and  A298 );
 a46458a <=( (not A301)  and  (not A300) );
 a46459a <=( a46458a  and  a46455a );
 a46460a <=( a46459a  and  a46452a );
 a46464a <=( (not A199)  and  A166 );
 a46465a <=( A167  and  a46464a );
 a46469a <=( (not A265)  and  (not A202) );
 a46470a <=( (not A200)  and  a46469a );
 a46471a <=( a46470a  and  a46465a );
 a46475a <=( A269  and  (not A268) );
 a46476a <=( A266  and  a46475a );
 a46479a <=( A299  and  A298 );
 a46482a <=( A302  and  (not A300) );
 a46483a <=( a46482a  and  a46479a );
 a46484a <=( a46483a  and  a46476a );
 a46488a <=( (not A199)  and  A166 );
 a46489a <=( A167  and  a46488a );
 a46493a <=( (not A265)  and  (not A202) );
 a46494a <=( (not A200)  and  a46493a );
 a46495a <=( a46494a  and  a46489a );
 a46499a <=( A269  and  (not A268) );
 a46500a <=( A266  and  a46499a );
 a46503a <=( (not A299)  and  A298 );
 a46506a <=( A301  and  (not A300) );
 a46507a <=( a46506a  and  a46503a );
 a46508a <=( a46507a  and  a46500a );
 a46512a <=( (not A199)  and  A166 );
 a46513a <=( A167  and  a46512a );
 a46517a <=( (not A265)  and  (not A202) );
 a46518a <=( (not A200)  and  a46517a );
 a46519a <=( a46518a  and  a46513a );
 a46523a <=( A269  and  (not A268) );
 a46524a <=( A266  and  a46523a );
 a46527a <=( (not A299)  and  A298 );
 a46530a <=( (not A302)  and  (not A300) );
 a46531a <=( a46530a  and  a46527a );
 a46532a <=( a46531a  and  a46524a );
 a46536a <=( (not A199)  and  A166 );
 a46537a <=( A167  and  a46536a );
 a46541a <=( (not A265)  and  (not A202) );
 a46542a <=( (not A200)  and  a46541a );
 a46543a <=( a46542a  and  a46537a );
 a46547a <=( A269  and  (not A268) );
 a46548a <=( A266  and  a46547a );
 a46551a <=( A299  and  (not A298) );
 a46554a <=( A301  and  (not A300) );
 a46555a <=( a46554a  and  a46551a );
 a46556a <=( a46555a  and  a46548a );
 a46560a <=( (not A199)  and  A166 );
 a46561a <=( A167  and  a46560a );
 a46565a <=( (not A265)  and  (not A202) );
 a46566a <=( (not A200)  and  a46565a );
 a46567a <=( a46566a  and  a46561a );
 a46571a <=( A269  and  (not A268) );
 a46572a <=( A266  and  a46571a );
 a46575a <=( A299  and  (not A298) );
 a46578a <=( (not A302)  and  (not A300) );
 a46579a <=( a46578a  and  a46575a );
 a46580a <=( a46579a  and  a46572a );
 a46584a <=( (not A199)  and  A166 );
 a46585a <=( A167  and  a46584a );
 a46589a <=( A265  and  (not A202) );
 a46590a <=( (not A200)  and  a46589a );
 a46591a <=( a46590a  and  a46585a );
 a46595a <=( A269  and  (not A268) );
 a46596a <=( (not A266)  and  a46595a );
 a46599a <=( A299  and  A298 );
 a46602a <=( (not A301)  and  (not A300) );
 a46603a <=( a46602a  and  a46599a );
 a46604a <=( a46603a  and  a46596a );
 a46608a <=( (not A199)  and  A166 );
 a46609a <=( A167  and  a46608a );
 a46613a <=( A265  and  (not A202) );
 a46614a <=( (not A200)  and  a46613a );
 a46615a <=( a46614a  and  a46609a );
 a46619a <=( A269  and  (not A268) );
 a46620a <=( (not A266)  and  a46619a );
 a46623a <=( A299  and  A298 );
 a46626a <=( A302  and  (not A300) );
 a46627a <=( a46626a  and  a46623a );
 a46628a <=( a46627a  and  a46620a );
 a46632a <=( (not A199)  and  A166 );
 a46633a <=( A167  and  a46632a );
 a46637a <=( A265  and  (not A202) );
 a46638a <=( (not A200)  and  a46637a );
 a46639a <=( a46638a  and  a46633a );
 a46643a <=( A269  and  (not A268) );
 a46644a <=( (not A266)  and  a46643a );
 a46647a <=( (not A299)  and  A298 );
 a46650a <=( A301  and  (not A300) );
 a46651a <=( a46650a  and  a46647a );
 a46652a <=( a46651a  and  a46644a );
 a46656a <=( (not A199)  and  A166 );
 a46657a <=( A167  and  a46656a );
 a46661a <=( A265  and  (not A202) );
 a46662a <=( (not A200)  and  a46661a );
 a46663a <=( a46662a  and  a46657a );
 a46667a <=( A269  and  (not A268) );
 a46668a <=( (not A266)  and  a46667a );
 a46671a <=( (not A299)  and  A298 );
 a46674a <=( (not A302)  and  (not A300) );
 a46675a <=( a46674a  and  a46671a );
 a46676a <=( a46675a  and  a46668a );
 a46680a <=( (not A199)  and  A166 );
 a46681a <=( A167  and  a46680a );
 a46685a <=( A265  and  (not A202) );
 a46686a <=( (not A200)  and  a46685a );
 a46687a <=( a46686a  and  a46681a );
 a46691a <=( A269  and  (not A268) );
 a46692a <=( (not A266)  and  a46691a );
 a46695a <=( A299  and  (not A298) );
 a46698a <=( A301  and  (not A300) );
 a46699a <=( a46698a  and  a46695a );
 a46700a <=( a46699a  and  a46692a );
 a46704a <=( (not A199)  and  A166 );
 a46705a <=( A167  and  a46704a );
 a46709a <=( A265  and  (not A202) );
 a46710a <=( (not A200)  and  a46709a );
 a46711a <=( a46710a  and  a46705a );
 a46715a <=( A269  and  (not A268) );
 a46716a <=( (not A266)  and  a46715a );
 a46719a <=( A299  and  (not A298) );
 a46722a <=( (not A302)  and  (not A300) );
 a46723a <=( a46722a  and  a46719a );
 a46724a <=( a46723a  and  a46716a );
 a46728a <=( (not A199)  and  A166 );
 a46729a <=( A167  and  a46728a );
 a46733a <=( (not A265)  and  (not A202) );
 a46734a <=( (not A200)  and  a46733a );
 a46735a <=( a46734a  and  a46729a );
 a46739a <=( (not A269)  and  A268 );
 a46740a <=( (not A266)  and  a46739a );
 a46743a <=( A299  and  A298 );
 a46746a <=( (not A301)  and  (not A300) );
 a46747a <=( a46746a  and  a46743a );
 a46748a <=( a46747a  and  a46740a );
 a46752a <=( (not A199)  and  A166 );
 a46753a <=( A167  and  a46752a );
 a46757a <=( (not A265)  and  (not A202) );
 a46758a <=( (not A200)  and  a46757a );
 a46759a <=( a46758a  and  a46753a );
 a46763a <=( (not A269)  and  A268 );
 a46764a <=( (not A266)  and  a46763a );
 a46767a <=( A299  and  A298 );
 a46770a <=( A302  and  (not A300) );
 a46771a <=( a46770a  and  a46767a );
 a46772a <=( a46771a  and  a46764a );
 a46776a <=( (not A199)  and  A166 );
 a46777a <=( A167  and  a46776a );
 a46781a <=( (not A265)  and  (not A202) );
 a46782a <=( (not A200)  and  a46781a );
 a46783a <=( a46782a  and  a46777a );
 a46787a <=( (not A269)  and  A268 );
 a46788a <=( (not A266)  and  a46787a );
 a46791a <=( (not A299)  and  A298 );
 a46794a <=( A301  and  (not A300) );
 a46795a <=( a46794a  and  a46791a );
 a46796a <=( a46795a  and  a46788a );
 a46800a <=( (not A199)  and  A166 );
 a46801a <=( A167  and  a46800a );
 a46805a <=( (not A265)  and  (not A202) );
 a46806a <=( (not A200)  and  a46805a );
 a46807a <=( a46806a  and  a46801a );
 a46811a <=( (not A269)  and  A268 );
 a46812a <=( (not A266)  and  a46811a );
 a46815a <=( (not A299)  and  A298 );
 a46818a <=( (not A302)  and  (not A300) );
 a46819a <=( a46818a  and  a46815a );
 a46820a <=( a46819a  and  a46812a );
 a46824a <=( (not A199)  and  A166 );
 a46825a <=( A167  and  a46824a );
 a46829a <=( (not A265)  and  (not A202) );
 a46830a <=( (not A200)  and  a46829a );
 a46831a <=( a46830a  and  a46825a );
 a46835a <=( (not A269)  and  A268 );
 a46836a <=( (not A266)  and  a46835a );
 a46839a <=( A299  and  (not A298) );
 a46842a <=( A301  and  (not A300) );
 a46843a <=( a46842a  and  a46839a );
 a46844a <=( a46843a  and  a46836a );
 a46848a <=( (not A199)  and  A166 );
 a46849a <=( A167  and  a46848a );
 a46853a <=( (not A265)  and  (not A202) );
 a46854a <=( (not A200)  and  a46853a );
 a46855a <=( a46854a  and  a46849a );
 a46859a <=( (not A269)  and  A268 );
 a46860a <=( (not A266)  and  a46859a );
 a46863a <=( A299  and  (not A298) );
 a46866a <=( (not A302)  and  (not A300) );
 a46867a <=( a46866a  and  a46863a );
 a46868a <=( a46867a  and  a46860a );
 a46872a <=( (not A199)  and  A166 );
 a46873a <=( A167  and  a46872a );
 a46877a <=( A265  and  A203 );
 a46878a <=( (not A200)  and  a46877a );
 a46879a <=( a46878a  and  a46873a );
 a46883a <=( (not A269)  and  A268 );
 a46884a <=( A266  and  a46883a );
 a46887a <=( A299  and  A298 );
 a46890a <=( (not A301)  and  (not A300) );
 a46891a <=( a46890a  and  a46887a );
 a46892a <=( a46891a  and  a46884a );
 a46896a <=( (not A199)  and  A166 );
 a46897a <=( A167  and  a46896a );
 a46901a <=( A265  and  A203 );
 a46902a <=( (not A200)  and  a46901a );
 a46903a <=( a46902a  and  a46897a );
 a46907a <=( (not A269)  and  A268 );
 a46908a <=( A266  and  a46907a );
 a46911a <=( A299  and  A298 );
 a46914a <=( A302  and  (not A300) );
 a46915a <=( a46914a  and  a46911a );
 a46916a <=( a46915a  and  a46908a );
 a46920a <=( (not A199)  and  A166 );
 a46921a <=( A167  and  a46920a );
 a46925a <=( A265  and  A203 );
 a46926a <=( (not A200)  and  a46925a );
 a46927a <=( a46926a  and  a46921a );
 a46931a <=( (not A269)  and  A268 );
 a46932a <=( A266  and  a46931a );
 a46935a <=( (not A299)  and  A298 );
 a46938a <=( A301  and  (not A300) );
 a46939a <=( a46938a  and  a46935a );
 a46940a <=( a46939a  and  a46932a );
 a46944a <=( (not A199)  and  A166 );
 a46945a <=( A167  and  a46944a );
 a46949a <=( A265  and  A203 );
 a46950a <=( (not A200)  and  a46949a );
 a46951a <=( a46950a  and  a46945a );
 a46955a <=( (not A269)  and  A268 );
 a46956a <=( A266  and  a46955a );
 a46959a <=( (not A299)  and  A298 );
 a46962a <=( (not A302)  and  (not A300) );
 a46963a <=( a46962a  and  a46959a );
 a46964a <=( a46963a  and  a46956a );
 a46968a <=( (not A199)  and  A166 );
 a46969a <=( A167  and  a46968a );
 a46973a <=( A265  and  A203 );
 a46974a <=( (not A200)  and  a46973a );
 a46975a <=( a46974a  and  a46969a );
 a46979a <=( (not A269)  and  A268 );
 a46980a <=( A266  and  a46979a );
 a46983a <=( A299  and  (not A298) );
 a46986a <=( A301  and  (not A300) );
 a46987a <=( a46986a  and  a46983a );
 a46988a <=( a46987a  and  a46980a );
 a46992a <=( (not A199)  and  A166 );
 a46993a <=( A167  and  a46992a );
 a46997a <=( A265  and  A203 );
 a46998a <=( (not A200)  and  a46997a );
 a46999a <=( a46998a  and  a46993a );
 a47003a <=( (not A269)  and  A268 );
 a47004a <=( A266  and  a47003a );
 a47007a <=( A299  and  (not A298) );
 a47010a <=( (not A302)  and  (not A300) );
 a47011a <=( a47010a  and  a47007a );
 a47012a <=( a47011a  and  a47004a );
 a47016a <=( (not A199)  and  A166 );
 a47017a <=( A167  and  a47016a );
 a47021a <=( (not A265)  and  A203 );
 a47022a <=( (not A200)  and  a47021a );
 a47023a <=( a47022a  and  a47017a );
 a47027a <=( A269  and  (not A268) );
 a47028a <=( A266  and  a47027a );
 a47031a <=( A299  and  A298 );
 a47034a <=( (not A301)  and  (not A300) );
 a47035a <=( a47034a  and  a47031a );
 a47036a <=( a47035a  and  a47028a );
 a47040a <=( (not A199)  and  A166 );
 a47041a <=( A167  and  a47040a );
 a47045a <=( (not A265)  and  A203 );
 a47046a <=( (not A200)  and  a47045a );
 a47047a <=( a47046a  and  a47041a );
 a47051a <=( A269  and  (not A268) );
 a47052a <=( A266  and  a47051a );
 a47055a <=( A299  and  A298 );
 a47058a <=( A302  and  (not A300) );
 a47059a <=( a47058a  and  a47055a );
 a47060a <=( a47059a  and  a47052a );
 a47064a <=( (not A199)  and  A166 );
 a47065a <=( A167  and  a47064a );
 a47069a <=( (not A265)  and  A203 );
 a47070a <=( (not A200)  and  a47069a );
 a47071a <=( a47070a  and  a47065a );
 a47075a <=( A269  and  (not A268) );
 a47076a <=( A266  and  a47075a );
 a47079a <=( (not A299)  and  A298 );
 a47082a <=( A301  and  (not A300) );
 a47083a <=( a47082a  and  a47079a );
 a47084a <=( a47083a  and  a47076a );
 a47088a <=( (not A199)  and  A166 );
 a47089a <=( A167  and  a47088a );
 a47093a <=( (not A265)  and  A203 );
 a47094a <=( (not A200)  and  a47093a );
 a47095a <=( a47094a  and  a47089a );
 a47099a <=( A269  and  (not A268) );
 a47100a <=( A266  and  a47099a );
 a47103a <=( (not A299)  and  A298 );
 a47106a <=( (not A302)  and  (not A300) );
 a47107a <=( a47106a  and  a47103a );
 a47108a <=( a47107a  and  a47100a );
 a47112a <=( (not A199)  and  A166 );
 a47113a <=( A167  and  a47112a );
 a47117a <=( (not A265)  and  A203 );
 a47118a <=( (not A200)  and  a47117a );
 a47119a <=( a47118a  and  a47113a );
 a47123a <=( A269  and  (not A268) );
 a47124a <=( A266  and  a47123a );
 a47127a <=( A299  and  (not A298) );
 a47130a <=( A301  and  (not A300) );
 a47131a <=( a47130a  and  a47127a );
 a47132a <=( a47131a  and  a47124a );
 a47136a <=( (not A199)  and  A166 );
 a47137a <=( A167  and  a47136a );
 a47141a <=( (not A265)  and  A203 );
 a47142a <=( (not A200)  and  a47141a );
 a47143a <=( a47142a  and  a47137a );
 a47147a <=( A269  and  (not A268) );
 a47148a <=( A266  and  a47147a );
 a47151a <=( A299  and  (not A298) );
 a47154a <=( (not A302)  and  (not A300) );
 a47155a <=( a47154a  and  a47151a );
 a47156a <=( a47155a  and  a47148a );
 a47160a <=( (not A199)  and  A166 );
 a47161a <=( A167  and  a47160a );
 a47165a <=( A265  and  A203 );
 a47166a <=( (not A200)  and  a47165a );
 a47167a <=( a47166a  and  a47161a );
 a47171a <=( A269  and  (not A268) );
 a47172a <=( (not A266)  and  a47171a );
 a47175a <=( A299  and  A298 );
 a47178a <=( (not A301)  and  (not A300) );
 a47179a <=( a47178a  and  a47175a );
 a47180a <=( a47179a  and  a47172a );
 a47184a <=( (not A199)  and  A166 );
 a47185a <=( A167  and  a47184a );
 a47189a <=( A265  and  A203 );
 a47190a <=( (not A200)  and  a47189a );
 a47191a <=( a47190a  and  a47185a );
 a47195a <=( A269  and  (not A268) );
 a47196a <=( (not A266)  and  a47195a );
 a47199a <=( A299  and  A298 );
 a47202a <=( A302  and  (not A300) );
 a47203a <=( a47202a  and  a47199a );
 a47204a <=( a47203a  and  a47196a );
 a47208a <=( (not A199)  and  A166 );
 a47209a <=( A167  and  a47208a );
 a47213a <=( A265  and  A203 );
 a47214a <=( (not A200)  and  a47213a );
 a47215a <=( a47214a  and  a47209a );
 a47219a <=( A269  and  (not A268) );
 a47220a <=( (not A266)  and  a47219a );
 a47223a <=( (not A299)  and  A298 );
 a47226a <=( A301  and  (not A300) );
 a47227a <=( a47226a  and  a47223a );
 a47228a <=( a47227a  and  a47220a );
 a47232a <=( (not A199)  and  A166 );
 a47233a <=( A167  and  a47232a );
 a47237a <=( A265  and  A203 );
 a47238a <=( (not A200)  and  a47237a );
 a47239a <=( a47238a  and  a47233a );
 a47243a <=( A269  and  (not A268) );
 a47244a <=( (not A266)  and  a47243a );
 a47247a <=( (not A299)  and  A298 );
 a47250a <=( (not A302)  and  (not A300) );
 a47251a <=( a47250a  and  a47247a );
 a47252a <=( a47251a  and  a47244a );
 a47256a <=( (not A199)  and  A166 );
 a47257a <=( A167  and  a47256a );
 a47261a <=( A265  and  A203 );
 a47262a <=( (not A200)  and  a47261a );
 a47263a <=( a47262a  and  a47257a );
 a47267a <=( A269  and  (not A268) );
 a47268a <=( (not A266)  and  a47267a );
 a47271a <=( A299  and  (not A298) );
 a47274a <=( A301  and  (not A300) );
 a47275a <=( a47274a  and  a47271a );
 a47276a <=( a47275a  and  a47268a );
 a47280a <=( (not A199)  and  A166 );
 a47281a <=( A167  and  a47280a );
 a47285a <=( A265  and  A203 );
 a47286a <=( (not A200)  and  a47285a );
 a47287a <=( a47286a  and  a47281a );
 a47291a <=( A269  and  (not A268) );
 a47292a <=( (not A266)  and  a47291a );
 a47295a <=( A299  and  (not A298) );
 a47298a <=( (not A302)  and  (not A300) );
 a47299a <=( a47298a  and  a47295a );
 a47300a <=( a47299a  and  a47292a );
 a47304a <=( (not A199)  and  A166 );
 a47305a <=( A167  and  a47304a );
 a47309a <=( (not A265)  and  A203 );
 a47310a <=( (not A200)  and  a47309a );
 a47311a <=( a47310a  and  a47305a );
 a47315a <=( (not A269)  and  A268 );
 a47316a <=( (not A266)  and  a47315a );
 a47319a <=( A299  and  A298 );
 a47322a <=( (not A301)  and  (not A300) );
 a47323a <=( a47322a  and  a47319a );
 a47324a <=( a47323a  and  a47316a );
 a47328a <=( (not A199)  and  A166 );
 a47329a <=( A167  and  a47328a );
 a47333a <=( (not A265)  and  A203 );
 a47334a <=( (not A200)  and  a47333a );
 a47335a <=( a47334a  and  a47329a );
 a47339a <=( (not A269)  and  A268 );
 a47340a <=( (not A266)  and  a47339a );
 a47343a <=( A299  and  A298 );
 a47346a <=( A302  and  (not A300) );
 a47347a <=( a47346a  and  a47343a );
 a47348a <=( a47347a  and  a47340a );
 a47352a <=( (not A199)  and  A166 );
 a47353a <=( A167  and  a47352a );
 a47357a <=( (not A265)  and  A203 );
 a47358a <=( (not A200)  and  a47357a );
 a47359a <=( a47358a  and  a47353a );
 a47363a <=( (not A269)  and  A268 );
 a47364a <=( (not A266)  and  a47363a );
 a47367a <=( (not A299)  and  A298 );
 a47370a <=( A301  and  (not A300) );
 a47371a <=( a47370a  and  a47367a );
 a47372a <=( a47371a  and  a47364a );
 a47376a <=( (not A199)  and  A166 );
 a47377a <=( A167  and  a47376a );
 a47381a <=( (not A265)  and  A203 );
 a47382a <=( (not A200)  and  a47381a );
 a47383a <=( a47382a  and  a47377a );
 a47387a <=( (not A269)  and  A268 );
 a47388a <=( (not A266)  and  a47387a );
 a47391a <=( (not A299)  and  A298 );
 a47394a <=( (not A302)  and  (not A300) );
 a47395a <=( a47394a  and  a47391a );
 a47396a <=( a47395a  and  a47388a );
 a47400a <=( (not A199)  and  A166 );
 a47401a <=( A167  and  a47400a );
 a47405a <=( (not A265)  and  A203 );
 a47406a <=( (not A200)  and  a47405a );
 a47407a <=( a47406a  and  a47401a );
 a47411a <=( (not A269)  and  A268 );
 a47412a <=( (not A266)  and  a47411a );
 a47415a <=( A299  and  (not A298) );
 a47418a <=( A301  and  (not A300) );
 a47419a <=( a47418a  and  a47415a );
 a47420a <=( a47419a  and  a47412a );
 a47424a <=( (not A199)  and  A166 );
 a47425a <=( A167  and  a47424a );
 a47429a <=( (not A265)  and  A203 );
 a47430a <=( (not A200)  and  a47429a );
 a47431a <=( a47430a  and  a47425a );
 a47435a <=( (not A269)  and  A268 );
 a47436a <=( (not A266)  and  a47435a );
 a47439a <=( A299  and  (not A298) );
 a47442a <=( (not A302)  and  (not A300) );
 a47443a <=( a47442a  and  a47439a );
 a47444a <=( a47443a  and  a47436a );
 a47448a <=( (not A199)  and  A166 );
 a47449a <=( A167  and  a47448a );
 a47453a <=( (not A203)  and  A202 );
 a47454a <=( (not A200)  and  a47453a );
 a47455a <=( a47454a  and  a47449a );
 a47459a <=( (not A268)  and  (not A266) );
 a47460a <=( (not A265)  and  a47459a );
 a47463a <=( A299  and  A298 );
 a47466a <=( (not A302)  and  A301 );
 a47467a <=( a47466a  and  a47463a );
 a47468a <=( a47467a  and  a47460a );
 a47472a <=( (not A199)  and  A166 );
 a47473a <=( A167  and  a47472a );
 a47477a <=( (not A203)  and  A202 );
 a47478a <=( (not A200)  and  a47477a );
 a47479a <=( a47478a  and  a47473a );
 a47483a <=( (not A268)  and  (not A266) );
 a47484a <=( (not A265)  and  a47483a );
 a47487a <=( (not A299)  and  A298 );
 a47490a <=( A302  and  (not A301) );
 a47491a <=( a47490a  and  a47487a );
 a47492a <=( a47491a  and  a47484a );
 a47496a <=( (not A199)  and  A166 );
 a47497a <=( A167  and  a47496a );
 a47501a <=( (not A203)  and  A202 );
 a47502a <=( (not A200)  and  a47501a );
 a47503a <=( a47502a  and  a47497a );
 a47507a <=( (not A268)  and  (not A266) );
 a47508a <=( (not A265)  and  a47507a );
 a47511a <=( A299  and  (not A298) );
 a47514a <=( A302  and  (not A301) );
 a47515a <=( a47514a  and  a47511a );
 a47516a <=( a47515a  and  a47508a );
 a47520a <=( (not A199)  and  A166 );
 a47521a <=( A167  and  a47520a );
 a47525a <=( (not A203)  and  A202 );
 a47526a <=( (not A200)  and  a47525a );
 a47527a <=( a47526a  and  a47521a );
 a47531a <=( (not A268)  and  (not A266) );
 a47532a <=( (not A265)  and  a47531a );
 a47535a <=( (not A299)  and  (not A298) );
 a47538a <=( (not A302)  and  A301 );
 a47539a <=( a47538a  and  a47535a );
 a47540a <=( a47539a  and  a47532a );
 a47544a <=( (not A199)  and  A166 );
 a47545a <=( A167  and  a47544a );
 a47549a <=( (not A203)  and  A202 );
 a47550a <=( (not A200)  and  a47549a );
 a47551a <=( a47550a  and  a47545a );
 a47555a <=( A269  and  (not A266) );
 a47556a <=( (not A265)  and  a47555a );
 a47559a <=( A299  and  A298 );
 a47562a <=( (not A302)  and  A301 );
 a47563a <=( a47562a  and  a47559a );
 a47564a <=( a47563a  and  a47556a );
 a47568a <=( (not A199)  and  A166 );
 a47569a <=( A167  and  a47568a );
 a47573a <=( (not A203)  and  A202 );
 a47574a <=( (not A200)  and  a47573a );
 a47575a <=( a47574a  and  a47569a );
 a47579a <=( A269  and  (not A266) );
 a47580a <=( (not A265)  and  a47579a );
 a47583a <=( (not A299)  and  A298 );
 a47586a <=( A302  and  (not A301) );
 a47587a <=( a47586a  and  a47583a );
 a47588a <=( a47587a  and  a47580a );
 a47592a <=( (not A199)  and  A166 );
 a47593a <=( A167  and  a47592a );
 a47597a <=( (not A203)  and  A202 );
 a47598a <=( (not A200)  and  a47597a );
 a47599a <=( a47598a  and  a47593a );
 a47603a <=( A269  and  (not A266) );
 a47604a <=( (not A265)  and  a47603a );
 a47607a <=( A299  and  (not A298) );
 a47610a <=( A302  and  (not A301) );
 a47611a <=( a47610a  and  a47607a );
 a47612a <=( a47611a  and  a47604a );
 a47616a <=( (not A199)  and  A166 );
 a47617a <=( A167  and  a47616a );
 a47621a <=( (not A203)  and  A202 );
 a47622a <=( (not A200)  and  a47621a );
 a47623a <=( a47622a  and  a47617a );
 a47627a <=( A269  and  (not A266) );
 a47628a <=( (not A265)  and  a47627a );
 a47631a <=( (not A299)  and  (not A298) );
 a47634a <=( (not A302)  and  A301 );
 a47635a <=( a47634a  and  a47631a );
 a47636a <=( a47635a  and  a47628a );
 a47640a <=( A199  and  (not A166) );
 a47641a <=( A167  and  a47640a );
 a47645a <=( (not A203)  and  A202 );
 a47646a <=( A200  and  a47645a );
 a47647a <=( a47646a  and  a47641a );
 a47651a <=( A268  and  A266 );
 a47652a <=( A265  and  a47651a );
 a47655a <=( (not A298)  and  (not A269) );
 a47658a <=( (not A301)  and  (not A299) );
 a47659a <=( a47658a  and  a47655a );
 a47660a <=( a47659a  and  a47652a );
 a47664a <=( A199  and  (not A166) );
 a47665a <=( A167  and  a47664a );
 a47669a <=( (not A203)  and  A202 );
 a47670a <=( A200  and  a47669a );
 a47671a <=( a47670a  and  a47665a );
 a47675a <=( A268  and  A266 );
 a47676a <=( A265  and  a47675a );
 a47679a <=( (not A298)  and  (not A269) );
 a47682a <=( A302  and  (not A299) );
 a47683a <=( a47682a  and  a47679a );
 a47684a <=( a47683a  and  a47676a );
 a47688a <=( A199  and  (not A166) );
 a47689a <=( A167  and  a47688a );
 a47693a <=( (not A203)  and  A202 );
 a47694a <=( A200  and  a47693a );
 a47695a <=( a47694a  and  a47689a );
 a47699a <=( (not A268)  and  A266 );
 a47700a <=( (not A265)  and  a47699a );
 a47703a <=( (not A298)  and  A269 );
 a47706a <=( (not A301)  and  (not A299) );
 a47707a <=( a47706a  and  a47703a );
 a47708a <=( a47707a  and  a47700a );
 a47712a <=( A199  and  (not A166) );
 a47713a <=( A167  and  a47712a );
 a47717a <=( (not A203)  and  A202 );
 a47718a <=( A200  and  a47717a );
 a47719a <=( a47718a  and  a47713a );
 a47723a <=( (not A268)  and  A266 );
 a47724a <=( (not A265)  and  a47723a );
 a47727a <=( (not A298)  and  A269 );
 a47730a <=( A302  and  (not A299) );
 a47731a <=( a47730a  and  a47727a );
 a47732a <=( a47731a  and  a47724a );
 a47736a <=( A199  and  (not A166) );
 a47737a <=( A167  and  a47736a );
 a47741a <=( (not A203)  and  A202 );
 a47742a <=( A200  and  a47741a );
 a47743a <=( a47742a  and  a47737a );
 a47747a <=( (not A268)  and  (not A266) );
 a47748a <=( A265  and  a47747a );
 a47751a <=( (not A298)  and  A269 );
 a47754a <=( (not A301)  and  (not A299) );
 a47755a <=( a47754a  and  a47751a );
 a47756a <=( a47755a  and  a47748a );
 a47760a <=( A199  and  (not A166) );
 a47761a <=( A167  and  a47760a );
 a47765a <=( (not A203)  and  A202 );
 a47766a <=( A200  and  a47765a );
 a47767a <=( a47766a  and  a47761a );
 a47771a <=( (not A268)  and  (not A266) );
 a47772a <=( A265  and  a47771a );
 a47775a <=( (not A298)  and  A269 );
 a47778a <=( A302  and  (not A299) );
 a47779a <=( a47778a  and  a47775a );
 a47780a <=( a47779a  and  a47772a );
 a47784a <=( A199  and  (not A166) );
 a47785a <=( A167  and  a47784a );
 a47789a <=( (not A203)  and  A202 );
 a47790a <=( A200  and  a47789a );
 a47791a <=( a47790a  and  a47785a );
 a47795a <=( A268  and  (not A266) );
 a47796a <=( (not A265)  and  a47795a );
 a47799a <=( (not A298)  and  (not A269) );
 a47802a <=( (not A301)  and  (not A299) );
 a47803a <=( a47802a  and  a47799a );
 a47804a <=( a47803a  and  a47796a );
 a47808a <=( A199  and  (not A166) );
 a47809a <=( A167  and  a47808a );
 a47813a <=( (not A203)  and  A202 );
 a47814a <=( A200  and  a47813a );
 a47815a <=( a47814a  and  a47809a );
 a47819a <=( A268  and  (not A266) );
 a47820a <=( (not A265)  and  a47819a );
 a47823a <=( (not A298)  and  (not A269) );
 a47826a <=( A302  and  (not A299) );
 a47827a <=( a47826a  and  a47823a );
 a47828a <=( a47827a  and  a47820a );
 a47832a <=( A199  and  (not A166) );
 a47833a <=( A167  and  a47832a );
 a47837a <=( (not A202)  and  (not A201) );
 a47838a <=( A200  and  a47837a );
 a47839a <=( a47838a  and  a47833a );
 a47843a <=( (not A268)  and  (not A266) );
 a47844a <=( (not A265)  and  a47843a );
 a47847a <=( A299  and  A298 );
 a47850a <=( (not A302)  and  A301 );
 a47851a <=( a47850a  and  a47847a );
 a47852a <=( a47851a  and  a47844a );
 a47856a <=( A199  and  (not A166) );
 a47857a <=( A167  and  a47856a );
 a47861a <=( (not A202)  and  (not A201) );
 a47862a <=( A200  and  a47861a );
 a47863a <=( a47862a  and  a47857a );
 a47867a <=( (not A268)  and  (not A266) );
 a47868a <=( (not A265)  and  a47867a );
 a47871a <=( (not A299)  and  A298 );
 a47874a <=( A302  and  (not A301) );
 a47875a <=( a47874a  and  a47871a );
 a47876a <=( a47875a  and  a47868a );
 a47880a <=( A199  and  (not A166) );
 a47881a <=( A167  and  a47880a );
 a47885a <=( (not A202)  and  (not A201) );
 a47886a <=( A200  and  a47885a );
 a47887a <=( a47886a  and  a47881a );
 a47891a <=( (not A268)  and  (not A266) );
 a47892a <=( (not A265)  and  a47891a );
 a47895a <=( A299  and  (not A298) );
 a47898a <=( A302  and  (not A301) );
 a47899a <=( a47898a  and  a47895a );
 a47900a <=( a47899a  and  a47892a );
 a47904a <=( A199  and  (not A166) );
 a47905a <=( A167  and  a47904a );
 a47909a <=( (not A202)  and  (not A201) );
 a47910a <=( A200  and  a47909a );
 a47911a <=( a47910a  and  a47905a );
 a47915a <=( (not A268)  and  (not A266) );
 a47916a <=( (not A265)  and  a47915a );
 a47919a <=( (not A299)  and  (not A298) );
 a47922a <=( (not A302)  and  A301 );
 a47923a <=( a47922a  and  a47919a );
 a47924a <=( a47923a  and  a47916a );
 a47928a <=( A199  and  (not A166) );
 a47929a <=( A167  and  a47928a );
 a47933a <=( (not A202)  and  (not A201) );
 a47934a <=( A200  and  a47933a );
 a47935a <=( a47934a  and  a47929a );
 a47939a <=( A269  and  (not A266) );
 a47940a <=( (not A265)  and  a47939a );
 a47943a <=( A299  and  A298 );
 a47946a <=( (not A302)  and  A301 );
 a47947a <=( a47946a  and  a47943a );
 a47948a <=( a47947a  and  a47940a );
 a47952a <=( A199  and  (not A166) );
 a47953a <=( A167  and  a47952a );
 a47957a <=( (not A202)  and  (not A201) );
 a47958a <=( A200  and  a47957a );
 a47959a <=( a47958a  and  a47953a );
 a47963a <=( A269  and  (not A266) );
 a47964a <=( (not A265)  and  a47963a );
 a47967a <=( (not A299)  and  A298 );
 a47970a <=( A302  and  (not A301) );
 a47971a <=( a47970a  and  a47967a );
 a47972a <=( a47971a  and  a47964a );
 a47976a <=( A199  and  (not A166) );
 a47977a <=( A167  and  a47976a );
 a47981a <=( (not A202)  and  (not A201) );
 a47982a <=( A200  and  a47981a );
 a47983a <=( a47982a  and  a47977a );
 a47987a <=( A269  and  (not A266) );
 a47988a <=( (not A265)  and  a47987a );
 a47991a <=( A299  and  (not A298) );
 a47994a <=( A302  and  (not A301) );
 a47995a <=( a47994a  and  a47991a );
 a47996a <=( a47995a  and  a47988a );
 a48000a <=( A199  and  (not A166) );
 a48001a <=( A167  and  a48000a );
 a48005a <=( (not A202)  and  (not A201) );
 a48006a <=( A200  and  a48005a );
 a48007a <=( a48006a  and  a48001a );
 a48011a <=( A269  and  (not A266) );
 a48012a <=( (not A265)  and  a48011a );
 a48015a <=( (not A299)  and  (not A298) );
 a48018a <=( (not A302)  and  A301 );
 a48019a <=( a48018a  and  a48015a );
 a48020a <=( a48019a  and  a48012a );
 a48024a <=( A199  and  (not A166) );
 a48025a <=( A167  and  a48024a );
 a48029a <=( A203  and  (not A201) );
 a48030a <=( A200  and  a48029a );
 a48031a <=( a48030a  and  a48025a );
 a48035a <=( (not A268)  and  (not A266) );
 a48036a <=( (not A265)  and  a48035a );
 a48039a <=( A299  and  A298 );
 a48042a <=( (not A302)  and  A301 );
 a48043a <=( a48042a  and  a48039a );
 a48044a <=( a48043a  and  a48036a );
 a48048a <=( A199  and  (not A166) );
 a48049a <=( A167  and  a48048a );
 a48053a <=( A203  and  (not A201) );
 a48054a <=( A200  and  a48053a );
 a48055a <=( a48054a  and  a48049a );
 a48059a <=( (not A268)  and  (not A266) );
 a48060a <=( (not A265)  and  a48059a );
 a48063a <=( (not A299)  and  A298 );
 a48066a <=( A302  and  (not A301) );
 a48067a <=( a48066a  and  a48063a );
 a48068a <=( a48067a  and  a48060a );
 a48072a <=( A199  and  (not A166) );
 a48073a <=( A167  and  a48072a );
 a48077a <=( A203  and  (not A201) );
 a48078a <=( A200  and  a48077a );
 a48079a <=( a48078a  and  a48073a );
 a48083a <=( (not A268)  and  (not A266) );
 a48084a <=( (not A265)  and  a48083a );
 a48087a <=( A299  and  (not A298) );
 a48090a <=( A302  and  (not A301) );
 a48091a <=( a48090a  and  a48087a );
 a48092a <=( a48091a  and  a48084a );
 a48096a <=( A199  and  (not A166) );
 a48097a <=( A167  and  a48096a );
 a48101a <=( A203  and  (not A201) );
 a48102a <=( A200  and  a48101a );
 a48103a <=( a48102a  and  a48097a );
 a48107a <=( (not A268)  and  (not A266) );
 a48108a <=( (not A265)  and  a48107a );
 a48111a <=( (not A299)  and  (not A298) );
 a48114a <=( (not A302)  and  A301 );
 a48115a <=( a48114a  and  a48111a );
 a48116a <=( a48115a  and  a48108a );
 a48120a <=( A199  and  (not A166) );
 a48121a <=( A167  and  a48120a );
 a48125a <=( A203  and  (not A201) );
 a48126a <=( A200  and  a48125a );
 a48127a <=( a48126a  and  a48121a );
 a48131a <=( A269  and  (not A266) );
 a48132a <=( (not A265)  and  a48131a );
 a48135a <=( A299  and  A298 );
 a48138a <=( (not A302)  and  A301 );
 a48139a <=( a48138a  and  a48135a );
 a48140a <=( a48139a  and  a48132a );
 a48144a <=( A199  and  (not A166) );
 a48145a <=( A167  and  a48144a );
 a48149a <=( A203  and  (not A201) );
 a48150a <=( A200  and  a48149a );
 a48151a <=( a48150a  and  a48145a );
 a48155a <=( A269  and  (not A266) );
 a48156a <=( (not A265)  and  a48155a );
 a48159a <=( (not A299)  and  A298 );
 a48162a <=( A302  and  (not A301) );
 a48163a <=( a48162a  and  a48159a );
 a48164a <=( a48163a  and  a48156a );
 a48168a <=( A199  and  (not A166) );
 a48169a <=( A167  and  a48168a );
 a48173a <=( A203  and  (not A201) );
 a48174a <=( A200  and  a48173a );
 a48175a <=( a48174a  and  a48169a );
 a48179a <=( A269  and  (not A266) );
 a48180a <=( (not A265)  and  a48179a );
 a48183a <=( A299  and  (not A298) );
 a48186a <=( A302  and  (not A301) );
 a48187a <=( a48186a  and  a48183a );
 a48188a <=( a48187a  and  a48180a );
 a48192a <=( A199  and  (not A166) );
 a48193a <=( A167  and  a48192a );
 a48197a <=( A203  and  (not A201) );
 a48198a <=( A200  and  a48197a );
 a48199a <=( a48198a  and  a48193a );
 a48203a <=( A269  and  (not A266) );
 a48204a <=( (not A265)  and  a48203a );
 a48207a <=( (not A299)  and  (not A298) );
 a48210a <=( (not A302)  and  A301 );
 a48211a <=( a48210a  and  a48207a );
 a48212a <=( a48211a  and  a48204a );
 a48216a <=( (not A199)  and  (not A166) );
 a48217a <=( A167  and  a48216a );
 a48221a <=( A203  and  (not A202) );
 a48222a <=( A200  and  a48221a );
 a48223a <=( a48222a  and  a48217a );
 a48227a <=( A268  and  A266 );
 a48228a <=( A265  and  a48227a );
 a48231a <=( (not A298)  and  (not A269) );
 a48234a <=( (not A301)  and  (not A299) );
 a48235a <=( a48234a  and  a48231a );
 a48236a <=( a48235a  and  a48228a );
 a48240a <=( (not A199)  and  (not A166) );
 a48241a <=( A167  and  a48240a );
 a48245a <=( A203  and  (not A202) );
 a48246a <=( A200  and  a48245a );
 a48247a <=( a48246a  and  a48241a );
 a48251a <=( A268  and  A266 );
 a48252a <=( A265  and  a48251a );
 a48255a <=( (not A298)  and  (not A269) );
 a48258a <=( A302  and  (not A299) );
 a48259a <=( a48258a  and  a48255a );
 a48260a <=( a48259a  and  a48252a );
 a48264a <=( (not A199)  and  (not A166) );
 a48265a <=( A167  and  a48264a );
 a48269a <=( A203  and  (not A202) );
 a48270a <=( A200  and  a48269a );
 a48271a <=( a48270a  and  a48265a );
 a48275a <=( (not A268)  and  A266 );
 a48276a <=( (not A265)  and  a48275a );
 a48279a <=( (not A298)  and  A269 );
 a48282a <=( (not A301)  and  (not A299) );
 a48283a <=( a48282a  and  a48279a );
 a48284a <=( a48283a  and  a48276a );
 a48288a <=( (not A199)  and  (not A166) );
 a48289a <=( A167  and  a48288a );
 a48293a <=( A203  and  (not A202) );
 a48294a <=( A200  and  a48293a );
 a48295a <=( a48294a  and  a48289a );
 a48299a <=( (not A268)  and  A266 );
 a48300a <=( (not A265)  and  a48299a );
 a48303a <=( (not A298)  and  A269 );
 a48306a <=( A302  and  (not A299) );
 a48307a <=( a48306a  and  a48303a );
 a48308a <=( a48307a  and  a48300a );
 a48312a <=( (not A199)  and  (not A166) );
 a48313a <=( A167  and  a48312a );
 a48317a <=( A203  and  (not A202) );
 a48318a <=( A200  and  a48317a );
 a48319a <=( a48318a  and  a48313a );
 a48323a <=( (not A268)  and  (not A266) );
 a48324a <=( A265  and  a48323a );
 a48327a <=( (not A298)  and  A269 );
 a48330a <=( (not A301)  and  (not A299) );
 a48331a <=( a48330a  and  a48327a );
 a48332a <=( a48331a  and  a48324a );
 a48336a <=( (not A199)  and  (not A166) );
 a48337a <=( A167  and  a48336a );
 a48341a <=( A203  and  (not A202) );
 a48342a <=( A200  and  a48341a );
 a48343a <=( a48342a  and  a48337a );
 a48347a <=( (not A268)  and  (not A266) );
 a48348a <=( A265  and  a48347a );
 a48351a <=( (not A298)  and  A269 );
 a48354a <=( A302  and  (not A299) );
 a48355a <=( a48354a  and  a48351a );
 a48356a <=( a48355a  and  a48348a );
 a48360a <=( (not A199)  and  (not A166) );
 a48361a <=( A167  and  a48360a );
 a48365a <=( A203  and  (not A202) );
 a48366a <=( A200  and  a48365a );
 a48367a <=( a48366a  and  a48361a );
 a48371a <=( A268  and  (not A266) );
 a48372a <=( (not A265)  and  a48371a );
 a48375a <=( (not A298)  and  (not A269) );
 a48378a <=( (not A301)  and  (not A299) );
 a48379a <=( a48378a  and  a48375a );
 a48380a <=( a48379a  and  a48372a );
 a48384a <=( (not A199)  and  (not A166) );
 a48385a <=( A167  and  a48384a );
 a48389a <=( A203  and  (not A202) );
 a48390a <=( A200  and  a48389a );
 a48391a <=( a48390a  and  a48385a );
 a48395a <=( A268  and  (not A266) );
 a48396a <=( (not A265)  and  a48395a );
 a48399a <=( (not A298)  and  (not A269) );
 a48402a <=( A302  and  (not A299) );
 a48403a <=( a48402a  and  a48399a );
 a48404a <=( a48403a  and  a48396a );
 a48408a <=( (not A199)  and  (not A166) );
 a48409a <=( A167  and  a48408a );
 a48413a <=( A202  and  (not A201) );
 a48414a <=( A200  and  a48413a );
 a48415a <=( a48414a  and  a48409a );
 a48419a <=( (not A268)  and  (not A266) );
 a48420a <=( (not A265)  and  a48419a );
 a48423a <=( A299  and  A298 );
 a48426a <=( (not A302)  and  A301 );
 a48427a <=( a48426a  and  a48423a );
 a48428a <=( a48427a  and  a48420a );
 a48432a <=( (not A199)  and  (not A166) );
 a48433a <=( A167  and  a48432a );
 a48437a <=( A202  and  (not A201) );
 a48438a <=( A200  and  a48437a );
 a48439a <=( a48438a  and  a48433a );
 a48443a <=( (not A268)  and  (not A266) );
 a48444a <=( (not A265)  and  a48443a );
 a48447a <=( (not A299)  and  A298 );
 a48450a <=( A302  and  (not A301) );
 a48451a <=( a48450a  and  a48447a );
 a48452a <=( a48451a  and  a48444a );
 a48456a <=( (not A199)  and  (not A166) );
 a48457a <=( A167  and  a48456a );
 a48461a <=( A202  and  (not A201) );
 a48462a <=( A200  and  a48461a );
 a48463a <=( a48462a  and  a48457a );
 a48467a <=( (not A268)  and  (not A266) );
 a48468a <=( (not A265)  and  a48467a );
 a48471a <=( A299  and  (not A298) );
 a48474a <=( A302  and  (not A301) );
 a48475a <=( a48474a  and  a48471a );
 a48476a <=( a48475a  and  a48468a );
 a48480a <=( (not A199)  and  (not A166) );
 a48481a <=( A167  and  a48480a );
 a48485a <=( A202  and  (not A201) );
 a48486a <=( A200  and  a48485a );
 a48487a <=( a48486a  and  a48481a );
 a48491a <=( (not A268)  and  (not A266) );
 a48492a <=( (not A265)  and  a48491a );
 a48495a <=( (not A299)  and  (not A298) );
 a48498a <=( (not A302)  and  A301 );
 a48499a <=( a48498a  and  a48495a );
 a48500a <=( a48499a  and  a48492a );
 a48504a <=( (not A199)  and  (not A166) );
 a48505a <=( A167  and  a48504a );
 a48509a <=( A202  and  (not A201) );
 a48510a <=( A200  and  a48509a );
 a48511a <=( a48510a  and  a48505a );
 a48515a <=( A269  and  (not A266) );
 a48516a <=( (not A265)  and  a48515a );
 a48519a <=( A299  and  A298 );
 a48522a <=( (not A302)  and  A301 );
 a48523a <=( a48522a  and  a48519a );
 a48524a <=( a48523a  and  a48516a );
 a48528a <=( (not A199)  and  (not A166) );
 a48529a <=( A167  and  a48528a );
 a48533a <=( A202  and  (not A201) );
 a48534a <=( A200  and  a48533a );
 a48535a <=( a48534a  and  a48529a );
 a48539a <=( A269  and  (not A266) );
 a48540a <=( (not A265)  and  a48539a );
 a48543a <=( (not A299)  and  A298 );
 a48546a <=( A302  and  (not A301) );
 a48547a <=( a48546a  and  a48543a );
 a48548a <=( a48547a  and  a48540a );
 a48552a <=( (not A199)  and  (not A166) );
 a48553a <=( A167  and  a48552a );
 a48557a <=( A202  and  (not A201) );
 a48558a <=( A200  and  a48557a );
 a48559a <=( a48558a  and  a48553a );
 a48563a <=( A269  and  (not A266) );
 a48564a <=( (not A265)  and  a48563a );
 a48567a <=( A299  and  (not A298) );
 a48570a <=( A302  and  (not A301) );
 a48571a <=( a48570a  and  a48567a );
 a48572a <=( a48571a  and  a48564a );
 a48576a <=( (not A199)  and  (not A166) );
 a48577a <=( A167  and  a48576a );
 a48581a <=( A202  and  (not A201) );
 a48582a <=( A200  and  a48581a );
 a48583a <=( a48582a  and  a48577a );
 a48587a <=( A269  and  (not A266) );
 a48588a <=( (not A265)  and  a48587a );
 a48591a <=( (not A299)  and  (not A298) );
 a48594a <=( (not A302)  and  A301 );
 a48595a <=( a48594a  and  a48591a );
 a48596a <=( a48595a  and  a48588a );
 a48600a <=( (not A199)  and  (not A166) );
 a48601a <=( A167  and  a48600a );
 a48605a <=( (not A203)  and  (not A201) );
 a48606a <=( A200  and  a48605a );
 a48607a <=( a48606a  and  a48601a );
 a48611a <=( (not A268)  and  (not A266) );
 a48612a <=( (not A265)  and  a48611a );
 a48615a <=( A299  and  A298 );
 a48618a <=( (not A302)  and  A301 );
 a48619a <=( a48618a  and  a48615a );
 a48620a <=( a48619a  and  a48612a );
 a48624a <=( (not A199)  and  (not A166) );
 a48625a <=( A167  and  a48624a );
 a48629a <=( (not A203)  and  (not A201) );
 a48630a <=( A200  and  a48629a );
 a48631a <=( a48630a  and  a48625a );
 a48635a <=( (not A268)  and  (not A266) );
 a48636a <=( (not A265)  and  a48635a );
 a48639a <=( (not A299)  and  A298 );
 a48642a <=( A302  and  (not A301) );
 a48643a <=( a48642a  and  a48639a );
 a48644a <=( a48643a  and  a48636a );
 a48648a <=( (not A199)  and  (not A166) );
 a48649a <=( A167  and  a48648a );
 a48653a <=( (not A203)  and  (not A201) );
 a48654a <=( A200  and  a48653a );
 a48655a <=( a48654a  and  a48649a );
 a48659a <=( (not A268)  and  (not A266) );
 a48660a <=( (not A265)  and  a48659a );
 a48663a <=( A299  and  (not A298) );
 a48666a <=( A302  and  (not A301) );
 a48667a <=( a48666a  and  a48663a );
 a48668a <=( a48667a  and  a48660a );
 a48672a <=( (not A199)  and  (not A166) );
 a48673a <=( A167  and  a48672a );
 a48677a <=( (not A203)  and  (not A201) );
 a48678a <=( A200  and  a48677a );
 a48679a <=( a48678a  and  a48673a );
 a48683a <=( (not A268)  and  (not A266) );
 a48684a <=( (not A265)  and  a48683a );
 a48687a <=( (not A299)  and  (not A298) );
 a48690a <=( (not A302)  and  A301 );
 a48691a <=( a48690a  and  a48687a );
 a48692a <=( a48691a  and  a48684a );
 a48696a <=( (not A199)  and  (not A166) );
 a48697a <=( A167  and  a48696a );
 a48701a <=( (not A203)  and  (not A201) );
 a48702a <=( A200  and  a48701a );
 a48703a <=( a48702a  and  a48697a );
 a48707a <=( A269  and  (not A266) );
 a48708a <=( (not A265)  and  a48707a );
 a48711a <=( A299  and  A298 );
 a48714a <=( (not A302)  and  A301 );
 a48715a <=( a48714a  and  a48711a );
 a48716a <=( a48715a  and  a48708a );
 a48720a <=( (not A199)  and  (not A166) );
 a48721a <=( A167  and  a48720a );
 a48725a <=( (not A203)  and  (not A201) );
 a48726a <=( A200  and  a48725a );
 a48727a <=( a48726a  and  a48721a );
 a48731a <=( A269  and  (not A266) );
 a48732a <=( (not A265)  and  a48731a );
 a48735a <=( (not A299)  and  A298 );
 a48738a <=( A302  and  (not A301) );
 a48739a <=( a48738a  and  a48735a );
 a48740a <=( a48739a  and  a48732a );
 a48744a <=( (not A199)  and  (not A166) );
 a48745a <=( A167  and  a48744a );
 a48749a <=( (not A203)  and  (not A201) );
 a48750a <=( A200  and  a48749a );
 a48751a <=( a48750a  and  a48745a );
 a48755a <=( A269  and  (not A266) );
 a48756a <=( (not A265)  and  a48755a );
 a48759a <=( A299  and  (not A298) );
 a48762a <=( A302  and  (not A301) );
 a48763a <=( a48762a  and  a48759a );
 a48764a <=( a48763a  and  a48756a );
 a48768a <=( (not A199)  and  (not A166) );
 a48769a <=( A167  and  a48768a );
 a48773a <=( (not A203)  and  (not A201) );
 a48774a <=( A200  and  a48773a );
 a48775a <=( a48774a  and  a48769a );
 a48779a <=( A269  and  (not A266) );
 a48780a <=( (not A265)  and  a48779a );
 a48783a <=( (not A299)  and  (not A298) );
 a48786a <=( (not A302)  and  A301 );
 a48787a <=( a48786a  and  a48783a );
 a48788a <=( a48787a  and  a48780a );
 a48792a <=( A199  and  (not A166) );
 a48793a <=( A167  and  a48792a );
 a48797a <=( A203  and  (not A202) );
 a48798a <=( (not A200)  and  a48797a );
 a48799a <=( a48798a  and  a48793a );
 a48803a <=( A268  and  A266 );
 a48804a <=( A265  and  a48803a );
 a48807a <=( (not A298)  and  (not A269) );
 a48810a <=( (not A301)  and  (not A299) );
 a48811a <=( a48810a  and  a48807a );
 a48812a <=( a48811a  and  a48804a );
 a48816a <=( A199  and  (not A166) );
 a48817a <=( A167  and  a48816a );
 a48821a <=( A203  and  (not A202) );
 a48822a <=( (not A200)  and  a48821a );
 a48823a <=( a48822a  and  a48817a );
 a48827a <=( A268  and  A266 );
 a48828a <=( A265  and  a48827a );
 a48831a <=( (not A298)  and  (not A269) );
 a48834a <=( A302  and  (not A299) );
 a48835a <=( a48834a  and  a48831a );
 a48836a <=( a48835a  and  a48828a );
 a48840a <=( A199  and  (not A166) );
 a48841a <=( A167  and  a48840a );
 a48845a <=( A203  and  (not A202) );
 a48846a <=( (not A200)  and  a48845a );
 a48847a <=( a48846a  and  a48841a );
 a48851a <=( (not A268)  and  A266 );
 a48852a <=( (not A265)  and  a48851a );
 a48855a <=( (not A298)  and  A269 );
 a48858a <=( (not A301)  and  (not A299) );
 a48859a <=( a48858a  and  a48855a );
 a48860a <=( a48859a  and  a48852a );
 a48864a <=( A199  and  (not A166) );
 a48865a <=( A167  and  a48864a );
 a48869a <=( A203  and  (not A202) );
 a48870a <=( (not A200)  and  a48869a );
 a48871a <=( a48870a  and  a48865a );
 a48875a <=( (not A268)  and  A266 );
 a48876a <=( (not A265)  and  a48875a );
 a48879a <=( (not A298)  and  A269 );
 a48882a <=( A302  and  (not A299) );
 a48883a <=( a48882a  and  a48879a );
 a48884a <=( a48883a  and  a48876a );
 a48888a <=( A199  and  (not A166) );
 a48889a <=( A167  and  a48888a );
 a48893a <=( A203  and  (not A202) );
 a48894a <=( (not A200)  and  a48893a );
 a48895a <=( a48894a  and  a48889a );
 a48899a <=( (not A268)  and  (not A266) );
 a48900a <=( A265  and  a48899a );
 a48903a <=( (not A298)  and  A269 );
 a48906a <=( (not A301)  and  (not A299) );
 a48907a <=( a48906a  and  a48903a );
 a48908a <=( a48907a  and  a48900a );
 a48912a <=( A199  and  (not A166) );
 a48913a <=( A167  and  a48912a );
 a48917a <=( A203  and  (not A202) );
 a48918a <=( (not A200)  and  a48917a );
 a48919a <=( a48918a  and  a48913a );
 a48923a <=( (not A268)  and  (not A266) );
 a48924a <=( A265  and  a48923a );
 a48927a <=( (not A298)  and  A269 );
 a48930a <=( A302  and  (not A299) );
 a48931a <=( a48930a  and  a48927a );
 a48932a <=( a48931a  and  a48924a );
 a48936a <=( A199  and  (not A166) );
 a48937a <=( A167  and  a48936a );
 a48941a <=( A203  and  (not A202) );
 a48942a <=( (not A200)  and  a48941a );
 a48943a <=( a48942a  and  a48937a );
 a48947a <=( A268  and  (not A266) );
 a48948a <=( (not A265)  and  a48947a );
 a48951a <=( (not A298)  and  (not A269) );
 a48954a <=( (not A301)  and  (not A299) );
 a48955a <=( a48954a  and  a48951a );
 a48956a <=( a48955a  and  a48948a );
 a48960a <=( A199  and  (not A166) );
 a48961a <=( A167  and  a48960a );
 a48965a <=( A203  and  (not A202) );
 a48966a <=( (not A200)  and  a48965a );
 a48967a <=( a48966a  and  a48961a );
 a48971a <=( A268  and  (not A266) );
 a48972a <=( (not A265)  and  a48971a );
 a48975a <=( (not A298)  and  (not A269) );
 a48978a <=( A302  and  (not A299) );
 a48979a <=( a48978a  and  a48975a );
 a48980a <=( a48979a  and  a48972a );
 a48984a <=( A199  and  (not A166) );
 a48985a <=( A167  and  a48984a );
 a48989a <=( A202  and  (not A201) );
 a48990a <=( (not A200)  and  a48989a );
 a48991a <=( a48990a  and  a48985a );
 a48995a <=( (not A268)  and  (not A266) );
 a48996a <=( (not A265)  and  a48995a );
 a48999a <=( A299  and  A298 );
 a49002a <=( (not A302)  and  A301 );
 a49003a <=( a49002a  and  a48999a );
 a49004a <=( a49003a  and  a48996a );
 a49008a <=( A199  and  (not A166) );
 a49009a <=( A167  and  a49008a );
 a49013a <=( A202  and  (not A201) );
 a49014a <=( (not A200)  and  a49013a );
 a49015a <=( a49014a  and  a49009a );
 a49019a <=( (not A268)  and  (not A266) );
 a49020a <=( (not A265)  and  a49019a );
 a49023a <=( (not A299)  and  A298 );
 a49026a <=( A302  and  (not A301) );
 a49027a <=( a49026a  and  a49023a );
 a49028a <=( a49027a  and  a49020a );
 a49032a <=( A199  and  (not A166) );
 a49033a <=( A167  and  a49032a );
 a49037a <=( A202  and  (not A201) );
 a49038a <=( (not A200)  and  a49037a );
 a49039a <=( a49038a  and  a49033a );
 a49043a <=( (not A268)  and  (not A266) );
 a49044a <=( (not A265)  and  a49043a );
 a49047a <=( A299  and  (not A298) );
 a49050a <=( A302  and  (not A301) );
 a49051a <=( a49050a  and  a49047a );
 a49052a <=( a49051a  and  a49044a );
 a49056a <=( A199  and  (not A166) );
 a49057a <=( A167  and  a49056a );
 a49061a <=( A202  and  (not A201) );
 a49062a <=( (not A200)  and  a49061a );
 a49063a <=( a49062a  and  a49057a );
 a49067a <=( (not A268)  and  (not A266) );
 a49068a <=( (not A265)  and  a49067a );
 a49071a <=( (not A299)  and  (not A298) );
 a49074a <=( (not A302)  and  A301 );
 a49075a <=( a49074a  and  a49071a );
 a49076a <=( a49075a  and  a49068a );
 a49080a <=( A199  and  (not A166) );
 a49081a <=( A167  and  a49080a );
 a49085a <=( A202  and  (not A201) );
 a49086a <=( (not A200)  and  a49085a );
 a49087a <=( a49086a  and  a49081a );
 a49091a <=( A269  and  (not A266) );
 a49092a <=( (not A265)  and  a49091a );
 a49095a <=( A299  and  A298 );
 a49098a <=( (not A302)  and  A301 );
 a49099a <=( a49098a  and  a49095a );
 a49100a <=( a49099a  and  a49092a );
 a49104a <=( A199  and  (not A166) );
 a49105a <=( A167  and  a49104a );
 a49109a <=( A202  and  (not A201) );
 a49110a <=( (not A200)  and  a49109a );
 a49111a <=( a49110a  and  a49105a );
 a49115a <=( A269  and  (not A266) );
 a49116a <=( (not A265)  and  a49115a );
 a49119a <=( (not A299)  and  A298 );
 a49122a <=( A302  and  (not A301) );
 a49123a <=( a49122a  and  a49119a );
 a49124a <=( a49123a  and  a49116a );
 a49128a <=( A199  and  (not A166) );
 a49129a <=( A167  and  a49128a );
 a49133a <=( A202  and  (not A201) );
 a49134a <=( (not A200)  and  a49133a );
 a49135a <=( a49134a  and  a49129a );
 a49139a <=( A269  and  (not A266) );
 a49140a <=( (not A265)  and  a49139a );
 a49143a <=( A299  and  (not A298) );
 a49146a <=( A302  and  (not A301) );
 a49147a <=( a49146a  and  a49143a );
 a49148a <=( a49147a  and  a49140a );
 a49152a <=( A199  and  (not A166) );
 a49153a <=( A167  and  a49152a );
 a49157a <=( A202  and  (not A201) );
 a49158a <=( (not A200)  and  a49157a );
 a49159a <=( a49158a  and  a49153a );
 a49163a <=( A269  and  (not A266) );
 a49164a <=( (not A265)  and  a49163a );
 a49167a <=( (not A299)  and  (not A298) );
 a49170a <=( (not A302)  and  A301 );
 a49171a <=( a49170a  and  a49167a );
 a49172a <=( a49171a  and  a49164a );
 a49176a <=( A199  and  (not A166) );
 a49177a <=( A167  and  a49176a );
 a49181a <=( (not A203)  and  (not A201) );
 a49182a <=( (not A200)  and  a49181a );
 a49183a <=( a49182a  and  a49177a );
 a49187a <=( (not A268)  and  (not A266) );
 a49188a <=( (not A265)  and  a49187a );
 a49191a <=( A299  and  A298 );
 a49194a <=( (not A302)  and  A301 );
 a49195a <=( a49194a  and  a49191a );
 a49196a <=( a49195a  and  a49188a );
 a49200a <=( A199  and  (not A166) );
 a49201a <=( A167  and  a49200a );
 a49205a <=( (not A203)  and  (not A201) );
 a49206a <=( (not A200)  and  a49205a );
 a49207a <=( a49206a  and  a49201a );
 a49211a <=( (not A268)  and  (not A266) );
 a49212a <=( (not A265)  and  a49211a );
 a49215a <=( (not A299)  and  A298 );
 a49218a <=( A302  and  (not A301) );
 a49219a <=( a49218a  and  a49215a );
 a49220a <=( a49219a  and  a49212a );
 a49224a <=( A199  and  (not A166) );
 a49225a <=( A167  and  a49224a );
 a49229a <=( (not A203)  and  (not A201) );
 a49230a <=( (not A200)  and  a49229a );
 a49231a <=( a49230a  and  a49225a );
 a49235a <=( (not A268)  and  (not A266) );
 a49236a <=( (not A265)  and  a49235a );
 a49239a <=( A299  and  (not A298) );
 a49242a <=( A302  and  (not A301) );
 a49243a <=( a49242a  and  a49239a );
 a49244a <=( a49243a  and  a49236a );
 a49248a <=( A199  and  (not A166) );
 a49249a <=( A167  and  a49248a );
 a49253a <=( (not A203)  and  (not A201) );
 a49254a <=( (not A200)  and  a49253a );
 a49255a <=( a49254a  and  a49249a );
 a49259a <=( (not A268)  and  (not A266) );
 a49260a <=( (not A265)  and  a49259a );
 a49263a <=( (not A299)  and  (not A298) );
 a49266a <=( (not A302)  and  A301 );
 a49267a <=( a49266a  and  a49263a );
 a49268a <=( a49267a  and  a49260a );
 a49272a <=( A199  and  (not A166) );
 a49273a <=( A167  and  a49272a );
 a49277a <=( (not A203)  and  (not A201) );
 a49278a <=( (not A200)  and  a49277a );
 a49279a <=( a49278a  and  a49273a );
 a49283a <=( A269  and  (not A266) );
 a49284a <=( (not A265)  and  a49283a );
 a49287a <=( A299  and  A298 );
 a49290a <=( (not A302)  and  A301 );
 a49291a <=( a49290a  and  a49287a );
 a49292a <=( a49291a  and  a49284a );
 a49296a <=( A199  and  (not A166) );
 a49297a <=( A167  and  a49296a );
 a49301a <=( (not A203)  and  (not A201) );
 a49302a <=( (not A200)  and  a49301a );
 a49303a <=( a49302a  and  a49297a );
 a49307a <=( A269  and  (not A266) );
 a49308a <=( (not A265)  and  a49307a );
 a49311a <=( (not A299)  and  A298 );
 a49314a <=( A302  and  (not A301) );
 a49315a <=( a49314a  and  a49311a );
 a49316a <=( a49315a  and  a49308a );
 a49320a <=( A199  and  (not A166) );
 a49321a <=( A167  and  a49320a );
 a49325a <=( (not A203)  and  (not A201) );
 a49326a <=( (not A200)  and  a49325a );
 a49327a <=( a49326a  and  a49321a );
 a49331a <=( A269  and  (not A266) );
 a49332a <=( (not A265)  and  a49331a );
 a49335a <=( A299  and  (not A298) );
 a49338a <=( A302  and  (not A301) );
 a49339a <=( a49338a  and  a49335a );
 a49340a <=( a49339a  and  a49332a );
 a49344a <=( A199  and  (not A166) );
 a49345a <=( A167  and  a49344a );
 a49349a <=( (not A203)  and  (not A201) );
 a49350a <=( (not A200)  and  a49349a );
 a49351a <=( a49350a  and  a49345a );
 a49355a <=( A269  and  (not A266) );
 a49356a <=( (not A265)  and  a49355a );
 a49359a <=( (not A299)  and  (not A298) );
 a49362a <=( (not A302)  and  A301 );
 a49363a <=( a49362a  and  a49359a );
 a49364a <=( a49363a  and  a49356a );
 a49368a <=( (not A199)  and  (not A166) );
 a49369a <=( A167  and  a49368a );
 a49373a <=( A265  and  (not A202) );
 a49374a <=( (not A200)  and  a49373a );
 a49375a <=( a49374a  and  a49369a );
 a49379a <=( (not A268)  and  (not A267) );
 a49380a <=( A266  and  a49379a );
 a49383a <=( A299  and  A298 );
 a49386a <=( (not A302)  and  A301 );
 a49387a <=( a49386a  and  a49383a );
 a49388a <=( a49387a  and  a49380a );
 a49392a <=( (not A199)  and  (not A166) );
 a49393a <=( A167  and  a49392a );
 a49397a <=( A265  and  (not A202) );
 a49398a <=( (not A200)  and  a49397a );
 a49399a <=( a49398a  and  a49393a );
 a49403a <=( (not A268)  and  (not A267) );
 a49404a <=( A266  and  a49403a );
 a49407a <=( (not A299)  and  A298 );
 a49410a <=( A302  and  (not A301) );
 a49411a <=( a49410a  and  a49407a );
 a49412a <=( a49411a  and  a49404a );
 a49416a <=( (not A199)  and  (not A166) );
 a49417a <=( A167  and  a49416a );
 a49421a <=( A265  and  (not A202) );
 a49422a <=( (not A200)  and  a49421a );
 a49423a <=( a49422a  and  a49417a );
 a49427a <=( (not A268)  and  (not A267) );
 a49428a <=( A266  and  a49427a );
 a49431a <=( A299  and  (not A298) );
 a49434a <=( A302  and  (not A301) );
 a49435a <=( a49434a  and  a49431a );
 a49436a <=( a49435a  and  a49428a );
 a49440a <=( (not A199)  and  (not A166) );
 a49441a <=( A167  and  a49440a );
 a49445a <=( A265  and  (not A202) );
 a49446a <=( (not A200)  and  a49445a );
 a49447a <=( a49446a  and  a49441a );
 a49451a <=( (not A268)  and  (not A267) );
 a49452a <=( A266  and  a49451a );
 a49455a <=( (not A299)  and  (not A298) );
 a49458a <=( (not A302)  and  A301 );
 a49459a <=( a49458a  and  a49455a );
 a49460a <=( a49459a  and  a49452a );
 a49464a <=( (not A199)  and  (not A166) );
 a49465a <=( A167  and  a49464a );
 a49469a <=( A265  and  (not A202) );
 a49470a <=( (not A200)  and  a49469a );
 a49471a <=( a49470a  and  a49465a );
 a49475a <=( A269  and  (not A267) );
 a49476a <=( A266  and  a49475a );
 a49479a <=( A299  and  A298 );
 a49482a <=( (not A302)  and  A301 );
 a49483a <=( a49482a  and  a49479a );
 a49484a <=( a49483a  and  a49476a );
 a49488a <=( (not A199)  and  (not A166) );
 a49489a <=( A167  and  a49488a );
 a49493a <=( A265  and  (not A202) );
 a49494a <=( (not A200)  and  a49493a );
 a49495a <=( a49494a  and  a49489a );
 a49499a <=( A269  and  (not A267) );
 a49500a <=( A266  and  a49499a );
 a49503a <=( (not A299)  and  A298 );
 a49506a <=( A302  and  (not A301) );
 a49507a <=( a49506a  and  a49503a );
 a49508a <=( a49507a  and  a49500a );
 a49512a <=( (not A199)  and  (not A166) );
 a49513a <=( A167  and  a49512a );
 a49517a <=( A265  and  (not A202) );
 a49518a <=( (not A200)  and  a49517a );
 a49519a <=( a49518a  and  a49513a );
 a49523a <=( A269  and  (not A267) );
 a49524a <=( A266  and  a49523a );
 a49527a <=( A299  and  (not A298) );
 a49530a <=( A302  and  (not A301) );
 a49531a <=( a49530a  and  a49527a );
 a49532a <=( a49531a  and  a49524a );
 a49536a <=( (not A199)  and  (not A166) );
 a49537a <=( A167  and  a49536a );
 a49541a <=( A265  and  (not A202) );
 a49542a <=( (not A200)  and  a49541a );
 a49543a <=( a49542a  and  a49537a );
 a49547a <=( A269  and  (not A267) );
 a49548a <=( A266  and  a49547a );
 a49551a <=( (not A299)  and  (not A298) );
 a49554a <=( (not A302)  and  A301 );
 a49555a <=( a49554a  and  a49551a );
 a49556a <=( a49555a  and  a49548a );
 a49560a <=( (not A199)  and  (not A166) );
 a49561a <=( A167  and  a49560a );
 a49565a <=( (not A265)  and  (not A202) );
 a49566a <=( (not A200)  and  a49565a );
 a49567a <=( a49566a  and  a49561a );
 a49571a <=( A268  and  (not A267) );
 a49572a <=( A266  and  a49571a );
 a49575a <=( A299  and  A298 );
 a49578a <=( (not A302)  and  A301 );
 a49579a <=( a49578a  and  a49575a );
 a49580a <=( a49579a  and  a49572a );
 a49584a <=( (not A199)  and  (not A166) );
 a49585a <=( A167  and  a49584a );
 a49589a <=( (not A265)  and  (not A202) );
 a49590a <=( (not A200)  and  a49589a );
 a49591a <=( a49590a  and  a49585a );
 a49595a <=( A268  and  (not A267) );
 a49596a <=( A266  and  a49595a );
 a49599a <=( (not A299)  and  A298 );
 a49602a <=( A302  and  (not A301) );
 a49603a <=( a49602a  and  a49599a );
 a49604a <=( a49603a  and  a49596a );
 a49608a <=( (not A199)  and  (not A166) );
 a49609a <=( A167  and  a49608a );
 a49613a <=( (not A265)  and  (not A202) );
 a49614a <=( (not A200)  and  a49613a );
 a49615a <=( a49614a  and  a49609a );
 a49619a <=( A268  and  (not A267) );
 a49620a <=( A266  and  a49619a );
 a49623a <=( A299  and  (not A298) );
 a49626a <=( A302  and  (not A301) );
 a49627a <=( a49626a  and  a49623a );
 a49628a <=( a49627a  and  a49620a );
 a49632a <=( (not A199)  and  (not A166) );
 a49633a <=( A167  and  a49632a );
 a49637a <=( (not A265)  and  (not A202) );
 a49638a <=( (not A200)  and  a49637a );
 a49639a <=( a49638a  and  a49633a );
 a49643a <=( A268  and  (not A267) );
 a49644a <=( A266  and  a49643a );
 a49647a <=( (not A299)  and  (not A298) );
 a49650a <=( (not A302)  and  A301 );
 a49651a <=( a49650a  and  a49647a );
 a49652a <=( a49651a  and  a49644a );
 a49656a <=( (not A199)  and  (not A166) );
 a49657a <=( A167  and  a49656a );
 a49661a <=( (not A265)  and  (not A202) );
 a49662a <=( (not A200)  and  a49661a );
 a49663a <=( a49662a  and  a49657a );
 a49667a <=( (not A269)  and  (not A267) );
 a49668a <=( A266  and  a49667a );
 a49671a <=( A299  and  A298 );
 a49674a <=( (not A302)  and  A301 );
 a49675a <=( a49674a  and  a49671a );
 a49676a <=( a49675a  and  a49668a );
 a49680a <=( (not A199)  and  (not A166) );
 a49681a <=( A167  and  a49680a );
 a49685a <=( (not A265)  and  (not A202) );
 a49686a <=( (not A200)  and  a49685a );
 a49687a <=( a49686a  and  a49681a );
 a49691a <=( (not A269)  and  (not A267) );
 a49692a <=( A266  and  a49691a );
 a49695a <=( (not A299)  and  A298 );
 a49698a <=( A302  and  (not A301) );
 a49699a <=( a49698a  and  a49695a );
 a49700a <=( a49699a  and  a49692a );
 a49704a <=( (not A199)  and  (not A166) );
 a49705a <=( A167  and  a49704a );
 a49709a <=( (not A265)  and  (not A202) );
 a49710a <=( (not A200)  and  a49709a );
 a49711a <=( a49710a  and  a49705a );
 a49715a <=( (not A269)  and  (not A267) );
 a49716a <=( A266  and  a49715a );
 a49719a <=( A299  and  (not A298) );
 a49722a <=( A302  and  (not A301) );
 a49723a <=( a49722a  and  a49719a );
 a49724a <=( a49723a  and  a49716a );
 a49728a <=( (not A199)  and  (not A166) );
 a49729a <=( A167  and  a49728a );
 a49733a <=( (not A265)  and  (not A202) );
 a49734a <=( (not A200)  and  a49733a );
 a49735a <=( a49734a  and  a49729a );
 a49739a <=( (not A269)  and  (not A267) );
 a49740a <=( A266  and  a49739a );
 a49743a <=( (not A299)  and  (not A298) );
 a49746a <=( (not A302)  and  A301 );
 a49747a <=( a49746a  and  a49743a );
 a49748a <=( a49747a  and  a49740a );
 a49752a <=( (not A199)  and  (not A166) );
 a49753a <=( A167  and  a49752a );
 a49757a <=( A265  and  (not A202) );
 a49758a <=( (not A200)  and  a49757a );
 a49759a <=( a49758a  and  a49753a );
 a49763a <=( A268  and  (not A267) );
 a49764a <=( (not A266)  and  a49763a );
 a49767a <=( A299  and  A298 );
 a49770a <=( (not A302)  and  A301 );
 a49771a <=( a49770a  and  a49767a );
 a49772a <=( a49771a  and  a49764a );
 a49776a <=( (not A199)  and  (not A166) );
 a49777a <=( A167  and  a49776a );
 a49781a <=( A265  and  (not A202) );
 a49782a <=( (not A200)  and  a49781a );
 a49783a <=( a49782a  and  a49777a );
 a49787a <=( A268  and  (not A267) );
 a49788a <=( (not A266)  and  a49787a );
 a49791a <=( (not A299)  and  A298 );
 a49794a <=( A302  and  (not A301) );
 a49795a <=( a49794a  and  a49791a );
 a49796a <=( a49795a  and  a49788a );
 a49800a <=( (not A199)  and  (not A166) );
 a49801a <=( A167  and  a49800a );
 a49805a <=( A265  and  (not A202) );
 a49806a <=( (not A200)  and  a49805a );
 a49807a <=( a49806a  and  a49801a );
 a49811a <=( A268  and  (not A267) );
 a49812a <=( (not A266)  and  a49811a );
 a49815a <=( A299  and  (not A298) );
 a49818a <=( A302  and  (not A301) );
 a49819a <=( a49818a  and  a49815a );
 a49820a <=( a49819a  and  a49812a );
 a49824a <=( (not A199)  and  (not A166) );
 a49825a <=( A167  and  a49824a );
 a49829a <=( A265  and  (not A202) );
 a49830a <=( (not A200)  and  a49829a );
 a49831a <=( a49830a  and  a49825a );
 a49835a <=( A268  and  (not A267) );
 a49836a <=( (not A266)  and  a49835a );
 a49839a <=( (not A299)  and  (not A298) );
 a49842a <=( (not A302)  and  A301 );
 a49843a <=( a49842a  and  a49839a );
 a49844a <=( a49843a  and  a49836a );
 a49848a <=( (not A199)  and  (not A166) );
 a49849a <=( A167  and  a49848a );
 a49853a <=( A265  and  (not A202) );
 a49854a <=( (not A200)  and  a49853a );
 a49855a <=( a49854a  and  a49849a );
 a49859a <=( (not A269)  and  (not A267) );
 a49860a <=( (not A266)  and  a49859a );
 a49863a <=( A299  and  A298 );
 a49866a <=( (not A302)  and  A301 );
 a49867a <=( a49866a  and  a49863a );
 a49868a <=( a49867a  and  a49860a );
 a49872a <=( (not A199)  and  (not A166) );
 a49873a <=( A167  and  a49872a );
 a49877a <=( A265  and  (not A202) );
 a49878a <=( (not A200)  and  a49877a );
 a49879a <=( a49878a  and  a49873a );
 a49883a <=( (not A269)  and  (not A267) );
 a49884a <=( (not A266)  and  a49883a );
 a49887a <=( (not A299)  and  A298 );
 a49890a <=( A302  and  (not A301) );
 a49891a <=( a49890a  and  a49887a );
 a49892a <=( a49891a  and  a49884a );
 a49896a <=( (not A199)  and  (not A166) );
 a49897a <=( A167  and  a49896a );
 a49901a <=( A265  and  (not A202) );
 a49902a <=( (not A200)  and  a49901a );
 a49903a <=( a49902a  and  a49897a );
 a49907a <=( (not A269)  and  (not A267) );
 a49908a <=( (not A266)  and  a49907a );
 a49911a <=( A299  and  (not A298) );
 a49914a <=( A302  and  (not A301) );
 a49915a <=( a49914a  and  a49911a );
 a49916a <=( a49915a  and  a49908a );
 a49920a <=( (not A199)  and  (not A166) );
 a49921a <=( A167  and  a49920a );
 a49925a <=( A265  and  (not A202) );
 a49926a <=( (not A200)  and  a49925a );
 a49927a <=( a49926a  and  a49921a );
 a49931a <=( (not A269)  and  (not A267) );
 a49932a <=( (not A266)  and  a49931a );
 a49935a <=( (not A299)  and  (not A298) );
 a49938a <=( (not A302)  and  A301 );
 a49939a <=( a49938a  and  a49935a );
 a49940a <=( a49939a  and  a49932a );
 a49944a <=( (not A199)  and  (not A166) );
 a49945a <=( A167  and  a49944a );
 a49949a <=( A265  and  A203 );
 a49950a <=( (not A200)  and  a49949a );
 a49951a <=( a49950a  and  a49945a );
 a49955a <=( (not A268)  and  (not A267) );
 a49956a <=( A266  and  a49955a );
 a49959a <=( A299  and  A298 );
 a49962a <=( (not A302)  and  A301 );
 a49963a <=( a49962a  and  a49959a );
 a49964a <=( a49963a  and  a49956a );
 a49968a <=( (not A199)  and  (not A166) );
 a49969a <=( A167  and  a49968a );
 a49973a <=( A265  and  A203 );
 a49974a <=( (not A200)  and  a49973a );
 a49975a <=( a49974a  and  a49969a );
 a49979a <=( (not A268)  and  (not A267) );
 a49980a <=( A266  and  a49979a );
 a49983a <=( (not A299)  and  A298 );
 a49986a <=( A302  and  (not A301) );
 a49987a <=( a49986a  and  a49983a );
 a49988a <=( a49987a  and  a49980a );
 a49992a <=( (not A199)  and  (not A166) );
 a49993a <=( A167  and  a49992a );
 a49997a <=( A265  and  A203 );
 a49998a <=( (not A200)  and  a49997a );
 a49999a <=( a49998a  and  a49993a );
 a50003a <=( (not A268)  and  (not A267) );
 a50004a <=( A266  and  a50003a );
 a50007a <=( A299  and  (not A298) );
 a50010a <=( A302  and  (not A301) );
 a50011a <=( a50010a  and  a50007a );
 a50012a <=( a50011a  and  a50004a );
 a50016a <=( (not A199)  and  (not A166) );
 a50017a <=( A167  and  a50016a );
 a50021a <=( A265  and  A203 );
 a50022a <=( (not A200)  and  a50021a );
 a50023a <=( a50022a  and  a50017a );
 a50027a <=( (not A268)  and  (not A267) );
 a50028a <=( A266  and  a50027a );
 a50031a <=( (not A299)  and  (not A298) );
 a50034a <=( (not A302)  and  A301 );
 a50035a <=( a50034a  and  a50031a );
 a50036a <=( a50035a  and  a50028a );
 a50040a <=( (not A199)  and  (not A166) );
 a50041a <=( A167  and  a50040a );
 a50045a <=( A265  and  A203 );
 a50046a <=( (not A200)  and  a50045a );
 a50047a <=( a50046a  and  a50041a );
 a50051a <=( A269  and  (not A267) );
 a50052a <=( A266  and  a50051a );
 a50055a <=( A299  and  A298 );
 a50058a <=( (not A302)  and  A301 );
 a50059a <=( a50058a  and  a50055a );
 a50060a <=( a50059a  and  a50052a );
 a50064a <=( (not A199)  and  (not A166) );
 a50065a <=( A167  and  a50064a );
 a50069a <=( A265  and  A203 );
 a50070a <=( (not A200)  and  a50069a );
 a50071a <=( a50070a  and  a50065a );
 a50075a <=( A269  and  (not A267) );
 a50076a <=( A266  and  a50075a );
 a50079a <=( (not A299)  and  A298 );
 a50082a <=( A302  and  (not A301) );
 a50083a <=( a50082a  and  a50079a );
 a50084a <=( a50083a  and  a50076a );
 a50088a <=( (not A199)  and  (not A166) );
 a50089a <=( A167  and  a50088a );
 a50093a <=( A265  and  A203 );
 a50094a <=( (not A200)  and  a50093a );
 a50095a <=( a50094a  and  a50089a );
 a50099a <=( A269  and  (not A267) );
 a50100a <=( A266  and  a50099a );
 a50103a <=( A299  and  (not A298) );
 a50106a <=( A302  and  (not A301) );
 a50107a <=( a50106a  and  a50103a );
 a50108a <=( a50107a  and  a50100a );
 a50112a <=( (not A199)  and  (not A166) );
 a50113a <=( A167  and  a50112a );
 a50117a <=( A265  and  A203 );
 a50118a <=( (not A200)  and  a50117a );
 a50119a <=( a50118a  and  a50113a );
 a50123a <=( A269  and  (not A267) );
 a50124a <=( A266  and  a50123a );
 a50127a <=( (not A299)  and  (not A298) );
 a50130a <=( (not A302)  and  A301 );
 a50131a <=( a50130a  and  a50127a );
 a50132a <=( a50131a  and  a50124a );
 a50136a <=( (not A199)  and  (not A166) );
 a50137a <=( A167  and  a50136a );
 a50141a <=( (not A265)  and  A203 );
 a50142a <=( (not A200)  and  a50141a );
 a50143a <=( a50142a  and  a50137a );
 a50147a <=( A268  and  (not A267) );
 a50148a <=( A266  and  a50147a );
 a50151a <=( A299  and  A298 );
 a50154a <=( (not A302)  and  A301 );
 a50155a <=( a50154a  and  a50151a );
 a50156a <=( a50155a  and  a50148a );
 a50160a <=( (not A199)  and  (not A166) );
 a50161a <=( A167  and  a50160a );
 a50165a <=( (not A265)  and  A203 );
 a50166a <=( (not A200)  and  a50165a );
 a50167a <=( a50166a  and  a50161a );
 a50171a <=( A268  and  (not A267) );
 a50172a <=( A266  and  a50171a );
 a50175a <=( (not A299)  and  A298 );
 a50178a <=( A302  and  (not A301) );
 a50179a <=( a50178a  and  a50175a );
 a50180a <=( a50179a  and  a50172a );
 a50184a <=( (not A199)  and  (not A166) );
 a50185a <=( A167  and  a50184a );
 a50189a <=( (not A265)  and  A203 );
 a50190a <=( (not A200)  and  a50189a );
 a50191a <=( a50190a  and  a50185a );
 a50195a <=( A268  and  (not A267) );
 a50196a <=( A266  and  a50195a );
 a50199a <=( A299  and  (not A298) );
 a50202a <=( A302  and  (not A301) );
 a50203a <=( a50202a  and  a50199a );
 a50204a <=( a50203a  and  a50196a );
 a50208a <=( (not A199)  and  (not A166) );
 a50209a <=( A167  and  a50208a );
 a50213a <=( (not A265)  and  A203 );
 a50214a <=( (not A200)  and  a50213a );
 a50215a <=( a50214a  and  a50209a );
 a50219a <=( A268  and  (not A267) );
 a50220a <=( A266  and  a50219a );
 a50223a <=( (not A299)  and  (not A298) );
 a50226a <=( (not A302)  and  A301 );
 a50227a <=( a50226a  and  a50223a );
 a50228a <=( a50227a  and  a50220a );
 a50232a <=( (not A199)  and  (not A166) );
 a50233a <=( A167  and  a50232a );
 a50237a <=( (not A265)  and  A203 );
 a50238a <=( (not A200)  and  a50237a );
 a50239a <=( a50238a  and  a50233a );
 a50243a <=( (not A269)  and  (not A267) );
 a50244a <=( A266  and  a50243a );
 a50247a <=( A299  and  A298 );
 a50250a <=( (not A302)  and  A301 );
 a50251a <=( a50250a  and  a50247a );
 a50252a <=( a50251a  and  a50244a );
 a50256a <=( (not A199)  and  (not A166) );
 a50257a <=( A167  and  a50256a );
 a50261a <=( (not A265)  and  A203 );
 a50262a <=( (not A200)  and  a50261a );
 a50263a <=( a50262a  and  a50257a );
 a50267a <=( (not A269)  and  (not A267) );
 a50268a <=( A266  and  a50267a );
 a50271a <=( (not A299)  and  A298 );
 a50274a <=( A302  and  (not A301) );
 a50275a <=( a50274a  and  a50271a );
 a50276a <=( a50275a  and  a50268a );
 a50280a <=( (not A199)  and  (not A166) );
 a50281a <=( A167  and  a50280a );
 a50285a <=( (not A265)  and  A203 );
 a50286a <=( (not A200)  and  a50285a );
 a50287a <=( a50286a  and  a50281a );
 a50291a <=( (not A269)  and  (not A267) );
 a50292a <=( A266  and  a50291a );
 a50295a <=( A299  and  (not A298) );
 a50298a <=( A302  and  (not A301) );
 a50299a <=( a50298a  and  a50295a );
 a50300a <=( a50299a  and  a50292a );
 a50304a <=( (not A199)  and  (not A166) );
 a50305a <=( A167  and  a50304a );
 a50309a <=( (not A265)  and  A203 );
 a50310a <=( (not A200)  and  a50309a );
 a50311a <=( a50310a  and  a50305a );
 a50315a <=( (not A269)  and  (not A267) );
 a50316a <=( A266  and  a50315a );
 a50319a <=( (not A299)  and  (not A298) );
 a50322a <=( (not A302)  and  A301 );
 a50323a <=( a50322a  and  a50319a );
 a50324a <=( a50323a  and  a50316a );
 a50328a <=( (not A199)  and  (not A166) );
 a50329a <=( A167  and  a50328a );
 a50333a <=( A265  and  A203 );
 a50334a <=( (not A200)  and  a50333a );
 a50335a <=( a50334a  and  a50329a );
 a50339a <=( A268  and  (not A267) );
 a50340a <=( (not A266)  and  a50339a );
 a50343a <=( A299  and  A298 );
 a50346a <=( (not A302)  and  A301 );
 a50347a <=( a50346a  and  a50343a );
 a50348a <=( a50347a  and  a50340a );
 a50352a <=( (not A199)  and  (not A166) );
 a50353a <=( A167  and  a50352a );
 a50357a <=( A265  and  A203 );
 a50358a <=( (not A200)  and  a50357a );
 a50359a <=( a50358a  and  a50353a );
 a50363a <=( A268  and  (not A267) );
 a50364a <=( (not A266)  and  a50363a );
 a50367a <=( (not A299)  and  A298 );
 a50370a <=( A302  and  (not A301) );
 a50371a <=( a50370a  and  a50367a );
 a50372a <=( a50371a  and  a50364a );
 a50376a <=( (not A199)  and  (not A166) );
 a50377a <=( A167  and  a50376a );
 a50381a <=( A265  and  A203 );
 a50382a <=( (not A200)  and  a50381a );
 a50383a <=( a50382a  and  a50377a );
 a50387a <=( A268  and  (not A267) );
 a50388a <=( (not A266)  and  a50387a );
 a50391a <=( A299  and  (not A298) );
 a50394a <=( A302  and  (not A301) );
 a50395a <=( a50394a  and  a50391a );
 a50396a <=( a50395a  and  a50388a );
 a50400a <=( (not A199)  and  (not A166) );
 a50401a <=( A167  and  a50400a );
 a50405a <=( A265  and  A203 );
 a50406a <=( (not A200)  and  a50405a );
 a50407a <=( a50406a  and  a50401a );
 a50411a <=( A268  and  (not A267) );
 a50412a <=( (not A266)  and  a50411a );
 a50415a <=( (not A299)  and  (not A298) );
 a50418a <=( (not A302)  and  A301 );
 a50419a <=( a50418a  and  a50415a );
 a50420a <=( a50419a  and  a50412a );
 a50424a <=( (not A199)  and  (not A166) );
 a50425a <=( A167  and  a50424a );
 a50429a <=( A265  and  A203 );
 a50430a <=( (not A200)  and  a50429a );
 a50431a <=( a50430a  and  a50425a );
 a50435a <=( (not A269)  and  (not A267) );
 a50436a <=( (not A266)  and  a50435a );
 a50439a <=( A299  and  A298 );
 a50442a <=( (not A302)  and  A301 );
 a50443a <=( a50442a  and  a50439a );
 a50444a <=( a50443a  and  a50436a );
 a50448a <=( (not A199)  and  (not A166) );
 a50449a <=( A167  and  a50448a );
 a50453a <=( A265  and  A203 );
 a50454a <=( (not A200)  and  a50453a );
 a50455a <=( a50454a  and  a50449a );
 a50459a <=( (not A269)  and  (not A267) );
 a50460a <=( (not A266)  and  a50459a );
 a50463a <=( (not A299)  and  A298 );
 a50466a <=( A302  and  (not A301) );
 a50467a <=( a50466a  and  a50463a );
 a50468a <=( a50467a  and  a50460a );
 a50472a <=( (not A199)  and  (not A166) );
 a50473a <=( A167  and  a50472a );
 a50477a <=( A265  and  A203 );
 a50478a <=( (not A200)  and  a50477a );
 a50479a <=( a50478a  and  a50473a );
 a50483a <=( (not A269)  and  (not A267) );
 a50484a <=( (not A266)  and  a50483a );
 a50487a <=( A299  and  (not A298) );
 a50490a <=( A302  and  (not A301) );
 a50491a <=( a50490a  and  a50487a );
 a50492a <=( a50491a  and  a50484a );
 a50496a <=( (not A199)  and  (not A166) );
 a50497a <=( A167  and  a50496a );
 a50501a <=( A265  and  A203 );
 a50502a <=( (not A200)  and  a50501a );
 a50503a <=( a50502a  and  a50497a );
 a50507a <=( (not A269)  and  (not A267) );
 a50508a <=( (not A266)  and  a50507a );
 a50511a <=( (not A299)  and  (not A298) );
 a50514a <=( (not A302)  and  A301 );
 a50515a <=( a50514a  and  a50511a );
 a50516a <=( a50515a  and  a50508a );
 a50520a <=( (not A199)  and  (not A166) );
 a50521a <=( A167  and  a50520a );
 a50525a <=( (not A203)  and  A202 );
 a50526a <=( (not A200)  and  a50525a );
 a50527a <=( a50526a  and  a50521a );
 a50531a <=( A268  and  A266 );
 a50532a <=( A265  and  a50531a );
 a50535a <=( (not A298)  and  (not A269) );
 a50538a <=( (not A301)  and  (not A299) );
 a50539a <=( a50538a  and  a50535a );
 a50540a <=( a50539a  and  a50532a );
 a50544a <=( (not A199)  and  (not A166) );
 a50545a <=( A167  and  a50544a );
 a50549a <=( (not A203)  and  A202 );
 a50550a <=( (not A200)  and  a50549a );
 a50551a <=( a50550a  and  a50545a );
 a50555a <=( A268  and  A266 );
 a50556a <=( A265  and  a50555a );
 a50559a <=( (not A298)  and  (not A269) );
 a50562a <=( A302  and  (not A299) );
 a50563a <=( a50562a  and  a50559a );
 a50564a <=( a50563a  and  a50556a );
 a50568a <=( (not A199)  and  (not A166) );
 a50569a <=( A167  and  a50568a );
 a50573a <=( (not A203)  and  A202 );
 a50574a <=( (not A200)  and  a50573a );
 a50575a <=( a50574a  and  a50569a );
 a50579a <=( (not A268)  and  A266 );
 a50580a <=( (not A265)  and  a50579a );
 a50583a <=( (not A298)  and  A269 );
 a50586a <=( (not A301)  and  (not A299) );
 a50587a <=( a50586a  and  a50583a );
 a50588a <=( a50587a  and  a50580a );
 a50592a <=( (not A199)  and  (not A166) );
 a50593a <=( A167  and  a50592a );
 a50597a <=( (not A203)  and  A202 );
 a50598a <=( (not A200)  and  a50597a );
 a50599a <=( a50598a  and  a50593a );
 a50603a <=( (not A268)  and  A266 );
 a50604a <=( (not A265)  and  a50603a );
 a50607a <=( (not A298)  and  A269 );
 a50610a <=( A302  and  (not A299) );
 a50611a <=( a50610a  and  a50607a );
 a50612a <=( a50611a  and  a50604a );
 a50616a <=( (not A199)  and  (not A166) );
 a50617a <=( A167  and  a50616a );
 a50621a <=( (not A203)  and  A202 );
 a50622a <=( (not A200)  and  a50621a );
 a50623a <=( a50622a  and  a50617a );
 a50627a <=( (not A268)  and  (not A266) );
 a50628a <=( A265  and  a50627a );
 a50631a <=( (not A298)  and  A269 );
 a50634a <=( (not A301)  and  (not A299) );
 a50635a <=( a50634a  and  a50631a );
 a50636a <=( a50635a  and  a50628a );
 a50640a <=( (not A199)  and  (not A166) );
 a50641a <=( A167  and  a50640a );
 a50645a <=( (not A203)  and  A202 );
 a50646a <=( (not A200)  and  a50645a );
 a50647a <=( a50646a  and  a50641a );
 a50651a <=( (not A268)  and  (not A266) );
 a50652a <=( A265  and  a50651a );
 a50655a <=( (not A298)  and  A269 );
 a50658a <=( A302  and  (not A299) );
 a50659a <=( a50658a  and  a50655a );
 a50660a <=( a50659a  and  a50652a );
 a50664a <=( (not A199)  and  (not A166) );
 a50665a <=( A167  and  a50664a );
 a50669a <=( (not A203)  and  A202 );
 a50670a <=( (not A200)  and  a50669a );
 a50671a <=( a50670a  and  a50665a );
 a50675a <=( A268  and  (not A266) );
 a50676a <=( (not A265)  and  a50675a );
 a50679a <=( (not A298)  and  (not A269) );
 a50682a <=( (not A301)  and  (not A299) );
 a50683a <=( a50682a  and  a50679a );
 a50684a <=( a50683a  and  a50676a );
 a50688a <=( (not A199)  and  (not A166) );
 a50689a <=( A167  and  a50688a );
 a50693a <=( (not A203)  and  A202 );
 a50694a <=( (not A200)  and  a50693a );
 a50695a <=( a50694a  and  a50689a );
 a50699a <=( A268  and  (not A266) );
 a50700a <=( (not A265)  and  a50699a );
 a50703a <=( (not A298)  and  (not A269) );
 a50706a <=( A302  and  (not A299) );
 a50707a <=( a50706a  and  a50703a );
 a50708a <=( a50707a  and  a50700a );
 a50712a <=( A199  and  (not A166) );
 a50713a <=( (not A167)  and  a50712a );
 a50717a <=( (not A203)  and  A202 );
 a50718a <=( A200  and  a50717a );
 a50719a <=( a50718a  and  a50713a );
 a50723a <=( (not A268)  and  (not A266) );
 a50724a <=( (not A265)  and  a50723a );
 a50727a <=( A299  and  A298 );
 a50730a <=( (not A302)  and  A301 );
 a50731a <=( a50730a  and  a50727a );
 a50732a <=( a50731a  and  a50724a );
 a50736a <=( A199  and  (not A166) );
 a50737a <=( (not A167)  and  a50736a );
 a50741a <=( (not A203)  and  A202 );
 a50742a <=( A200  and  a50741a );
 a50743a <=( a50742a  and  a50737a );
 a50747a <=( (not A268)  and  (not A266) );
 a50748a <=( (not A265)  and  a50747a );
 a50751a <=( (not A299)  and  A298 );
 a50754a <=( A302  and  (not A301) );
 a50755a <=( a50754a  and  a50751a );
 a50756a <=( a50755a  and  a50748a );
 a50760a <=( A199  and  (not A166) );
 a50761a <=( (not A167)  and  a50760a );
 a50765a <=( (not A203)  and  A202 );
 a50766a <=( A200  and  a50765a );
 a50767a <=( a50766a  and  a50761a );
 a50771a <=( (not A268)  and  (not A266) );
 a50772a <=( (not A265)  and  a50771a );
 a50775a <=( A299  and  (not A298) );
 a50778a <=( A302  and  (not A301) );
 a50779a <=( a50778a  and  a50775a );
 a50780a <=( a50779a  and  a50772a );
 a50784a <=( A199  and  (not A166) );
 a50785a <=( (not A167)  and  a50784a );
 a50789a <=( (not A203)  and  A202 );
 a50790a <=( A200  and  a50789a );
 a50791a <=( a50790a  and  a50785a );
 a50795a <=( (not A268)  and  (not A266) );
 a50796a <=( (not A265)  and  a50795a );
 a50799a <=( (not A299)  and  (not A298) );
 a50802a <=( (not A302)  and  A301 );
 a50803a <=( a50802a  and  a50799a );
 a50804a <=( a50803a  and  a50796a );
 a50808a <=( A199  and  (not A166) );
 a50809a <=( (not A167)  and  a50808a );
 a50813a <=( (not A203)  and  A202 );
 a50814a <=( A200  and  a50813a );
 a50815a <=( a50814a  and  a50809a );
 a50819a <=( A269  and  (not A266) );
 a50820a <=( (not A265)  and  a50819a );
 a50823a <=( A299  and  A298 );
 a50826a <=( (not A302)  and  A301 );
 a50827a <=( a50826a  and  a50823a );
 a50828a <=( a50827a  and  a50820a );
 a50832a <=( A199  and  (not A166) );
 a50833a <=( (not A167)  and  a50832a );
 a50837a <=( (not A203)  and  A202 );
 a50838a <=( A200  and  a50837a );
 a50839a <=( a50838a  and  a50833a );
 a50843a <=( A269  and  (not A266) );
 a50844a <=( (not A265)  and  a50843a );
 a50847a <=( (not A299)  and  A298 );
 a50850a <=( A302  and  (not A301) );
 a50851a <=( a50850a  and  a50847a );
 a50852a <=( a50851a  and  a50844a );
 a50856a <=( A199  and  (not A166) );
 a50857a <=( (not A167)  and  a50856a );
 a50861a <=( (not A203)  and  A202 );
 a50862a <=( A200  and  a50861a );
 a50863a <=( a50862a  and  a50857a );
 a50867a <=( A269  and  (not A266) );
 a50868a <=( (not A265)  and  a50867a );
 a50871a <=( A299  and  (not A298) );
 a50874a <=( A302  and  (not A301) );
 a50875a <=( a50874a  and  a50871a );
 a50876a <=( a50875a  and  a50868a );
 a50880a <=( A199  and  (not A166) );
 a50881a <=( (not A167)  and  a50880a );
 a50885a <=( (not A203)  and  A202 );
 a50886a <=( A200  and  a50885a );
 a50887a <=( a50886a  and  a50881a );
 a50891a <=( A269  and  (not A266) );
 a50892a <=( (not A265)  and  a50891a );
 a50895a <=( (not A299)  and  (not A298) );
 a50898a <=( (not A302)  and  A301 );
 a50899a <=( a50898a  and  a50895a );
 a50900a <=( a50899a  and  a50892a );
 a50904a <=( A199  and  (not A166) );
 a50905a <=( (not A167)  and  a50904a );
 a50909a <=( (not A202)  and  (not A201) );
 a50910a <=( A200  and  a50909a );
 a50911a <=( a50910a  and  a50905a );
 a50915a <=( A268  and  A266 );
 a50916a <=( A265  and  a50915a );
 a50919a <=( (not A298)  and  (not A269) );
 a50922a <=( (not A301)  and  (not A299) );
 a50923a <=( a50922a  and  a50919a );
 a50924a <=( a50923a  and  a50916a );
 a50928a <=( A199  and  (not A166) );
 a50929a <=( (not A167)  and  a50928a );
 a50933a <=( (not A202)  and  (not A201) );
 a50934a <=( A200  and  a50933a );
 a50935a <=( a50934a  and  a50929a );
 a50939a <=( A268  and  A266 );
 a50940a <=( A265  and  a50939a );
 a50943a <=( (not A298)  and  (not A269) );
 a50946a <=( A302  and  (not A299) );
 a50947a <=( a50946a  and  a50943a );
 a50948a <=( a50947a  and  a50940a );
 a50952a <=( A199  and  (not A166) );
 a50953a <=( (not A167)  and  a50952a );
 a50957a <=( (not A202)  and  (not A201) );
 a50958a <=( A200  and  a50957a );
 a50959a <=( a50958a  and  a50953a );
 a50963a <=( (not A268)  and  A266 );
 a50964a <=( (not A265)  and  a50963a );
 a50967a <=( (not A298)  and  A269 );
 a50970a <=( (not A301)  and  (not A299) );
 a50971a <=( a50970a  and  a50967a );
 a50972a <=( a50971a  and  a50964a );
 a50976a <=( A199  and  (not A166) );
 a50977a <=( (not A167)  and  a50976a );
 a50981a <=( (not A202)  and  (not A201) );
 a50982a <=( A200  and  a50981a );
 a50983a <=( a50982a  and  a50977a );
 a50987a <=( (not A268)  and  A266 );
 a50988a <=( (not A265)  and  a50987a );
 a50991a <=( (not A298)  and  A269 );
 a50994a <=( A302  and  (not A299) );
 a50995a <=( a50994a  and  a50991a );
 a50996a <=( a50995a  and  a50988a );
 a51000a <=( A199  and  (not A166) );
 a51001a <=( (not A167)  and  a51000a );
 a51005a <=( (not A202)  and  (not A201) );
 a51006a <=( A200  and  a51005a );
 a51007a <=( a51006a  and  a51001a );
 a51011a <=( (not A268)  and  (not A266) );
 a51012a <=( A265  and  a51011a );
 a51015a <=( (not A298)  and  A269 );
 a51018a <=( (not A301)  and  (not A299) );
 a51019a <=( a51018a  and  a51015a );
 a51020a <=( a51019a  and  a51012a );
 a51024a <=( A199  and  (not A166) );
 a51025a <=( (not A167)  and  a51024a );
 a51029a <=( (not A202)  and  (not A201) );
 a51030a <=( A200  and  a51029a );
 a51031a <=( a51030a  and  a51025a );
 a51035a <=( (not A268)  and  (not A266) );
 a51036a <=( A265  and  a51035a );
 a51039a <=( (not A298)  and  A269 );
 a51042a <=( A302  and  (not A299) );
 a51043a <=( a51042a  and  a51039a );
 a51044a <=( a51043a  and  a51036a );
 a51048a <=( A199  and  (not A166) );
 a51049a <=( (not A167)  and  a51048a );
 a51053a <=( (not A202)  and  (not A201) );
 a51054a <=( A200  and  a51053a );
 a51055a <=( a51054a  and  a51049a );
 a51059a <=( A268  and  (not A266) );
 a51060a <=( (not A265)  and  a51059a );
 a51063a <=( (not A298)  and  (not A269) );
 a51066a <=( (not A301)  and  (not A299) );
 a51067a <=( a51066a  and  a51063a );
 a51068a <=( a51067a  and  a51060a );
 a51072a <=( A199  and  (not A166) );
 a51073a <=( (not A167)  and  a51072a );
 a51077a <=( (not A202)  and  (not A201) );
 a51078a <=( A200  and  a51077a );
 a51079a <=( a51078a  and  a51073a );
 a51083a <=( A268  and  (not A266) );
 a51084a <=( (not A265)  and  a51083a );
 a51087a <=( (not A298)  and  (not A269) );
 a51090a <=( A302  and  (not A299) );
 a51091a <=( a51090a  and  a51087a );
 a51092a <=( a51091a  and  a51084a );
 a51096a <=( A199  and  (not A166) );
 a51097a <=( (not A167)  and  a51096a );
 a51101a <=( A203  and  (not A201) );
 a51102a <=( A200  and  a51101a );
 a51103a <=( a51102a  and  a51097a );
 a51107a <=( A268  and  A266 );
 a51108a <=( A265  and  a51107a );
 a51111a <=( (not A298)  and  (not A269) );
 a51114a <=( (not A301)  and  (not A299) );
 a51115a <=( a51114a  and  a51111a );
 a51116a <=( a51115a  and  a51108a );
 a51120a <=( A199  and  (not A166) );
 a51121a <=( (not A167)  and  a51120a );
 a51125a <=( A203  and  (not A201) );
 a51126a <=( A200  and  a51125a );
 a51127a <=( a51126a  and  a51121a );
 a51131a <=( A268  and  A266 );
 a51132a <=( A265  and  a51131a );
 a51135a <=( (not A298)  and  (not A269) );
 a51138a <=( A302  and  (not A299) );
 a51139a <=( a51138a  and  a51135a );
 a51140a <=( a51139a  and  a51132a );
 a51144a <=( A199  and  (not A166) );
 a51145a <=( (not A167)  and  a51144a );
 a51149a <=( A203  and  (not A201) );
 a51150a <=( A200  and  a51149a );
 a51151a <=( a51150a  and  a51145a );
 a51155a <=( (not A268)  and  A266 );
 a51156a <=( (not A265)  and  a51155a );
 a51159a <=( (not A298)  and  A269 );
 a51162a <=( (not A301)  and  (not A299) );
 a51163a <=( a51162a  and  a51159a );
 a51164a <=( a51163a  and  a51156a );
 a51168a <=( A199  and  (not A166) );
 a51169a <=( (not A167)  and  a51168a );
 a51173a <=( A203  and  (not A201) );
 a51174a <=( A200  and  a51173a );
 a51175a <=( a51174a  and  a51169a );
 a51179a <=( (not A268)  and  A266 );
 a51180a <=( (not A265)  and  a51179a );
 a51183a <=( (not A298)  and  A269 );
 a51186a <=( A302  and  (not A299) );
 a51187a <=( a51186a  and  a51183a );
 a51188a <=( a51187a  and  a51180a );
 a51192a <=( A199  and  (not A166) );
 a51193a <=( (not A167)  and  a51192a );
 a51197a <=( A203  and  (not A201) );
 a51198a <=( A200  and  a51197a );
 a51199a <=( a51198a  and  a51193a );
 a51203a <=( (not A268)  and  (not A266) );
 a51204a <=( A265  and  a51203a );
 a51207a <=( (not A298)  and  A269 );
 a51210a <=( (not A301)  and  (not A299) );
 a51211a <=( a51210a  and  a51207a );
 a51212a <=( a51211a  and  a51204a );
 a51216a <=( A199  and  (not A166) );
 a51217a <=( (not A167)  and  a51216a );
 a51221a <=( A203  and  (not A201) );
 a51222a <=( A200  and  a51221a );
 a51223a <=( a51222a  and  a51217a );
 a51227a <=( (not A268)  and  (not A266) );
 a51228a <=( A265  and  a51227a );
 a51231a <=( (not A298)  and  A269 );
 a51234a <=( A302  and  (not A299) );
 a51235a <=( a51234a  and  a51231a );
 a51236a <=( a51235a  and  a51228a );
 a51240a <=( A199  and  (not A166) );
 a51241a <=( (not A167)  and  a51240a );
 a51245a <=( A203  and  (not A201) );
 a51246a <=( A200  and  a51245a );
 a51247a <=( a51246a  and  a51241a );
 a51251a <=( A268  and  (not A266) );
 a51252a <=( (not A265)  and  a51251a );
 a51255a <=( (not A298)  and  (not A269) );
 a51258a <=( (not A301)  and  (not A299) );
 a51259a <=( a51258a  and  a51255a );
 a51260a <=( a51259a  and  a51252a );
 a51264a <=( A199  and  (not A166) );
 a51265a <=( (not A167)  and  a51264a );
 a51269a <=( A203  and  (not A201) );
 a51270a <=( A200  and  a51269a );
 a51271a <=( a51270a  and  a51265a );
 a51275a <=( A268  and  (not A266) );
 a51276a <=( (not A265)  and  a51275a );
 a51279a <=( (not A298)  and  (not A269) );
 a51282a <=( A302  and  (not A299) );
 a51283a <=( a51282a  and  a51279a );
 a51284a <=( a51283a  and  a51276a );
 a51288a <=( (not A199)  and  (not A166) );
 a51289a <=( (not A167)  and  a51288a );
 a51293a <=( A203  and  (not A202) );
 a51294a <=( A200  and  a51293a );
 a51295a <=( a51294a  and  a51289a );
 a51299a <=( (not A268)  and  (not A266) );
 a51300a <=( (not A265)  and  a51299a );
 a51303a <=( A299  and  A298 );
 a51306a <=( (not A302)  and  A301 );
 a51307a <=( a51306a  and  a51303a );
 a51308a <=( a51307a  and  a51300a );
 a51312a <=( (not A199)  and  (not A166) );
 a51313a <=( (not A167)  and  a51312a );
 a51317a <=( A203  and  (not A202) );
 a51318a <=( A200  and  a51317a );
 a51319a <=( a51318a  and  a51313a );
 a51323a <=( (not A268)  and  (not A266) );
 a51324a <=( (not A265)  and  a51323a );
 a51327a <=( (not A299)  and  A298 );
 a51330a <=( A302  and  (not A301) );
 a51331a <=( a51330a  and  a51327a );
 a51332a <=( a51331a  and  a51324a );
 a51336a <=( (not A199)  and  (not A166) );
 a51337a <=( (not A167)  and  a51336a );
 a51341a <=( A203  and  (not A202) );
 a51342a <=( A200  and  a51341a );
 a51343a <=( a51342a  and  a51337a );
 a51347a <=( (not A268)  and  (not A266) );
 a51348a <=( (not A265)  and  a51347a );
 a51351a <=( A299  and  (not A298) );
 a51354a <=( A302  and  (not A301) );
 a51355a <=( a51354a  and  a51351a );
 a51356a <=( a51355a  and  a51348a );
 a51360a <=( (not A199)  and  (not A166) );
 a51361a <=( (not A167)  and  a51360a );
 a51365a <=( A203  and  (not A202) );
 a51366a <=( A200  and  a51365a );
 a51367a <=( a51366a  and  a51361a );
 a51371a <=( (not A268)  and  (not A266) );
 a51372a <=( (not A265)  and  a51371a );
 a51375a <=( (not A299)  and  (not A298) );
 a51378a <=( (not A302)  and  A301 );
 a51379a <=( a51378a  and  a51375a );
 a51380a <=( a51379a  and  a51372a );
 a51384a <=( (not A199)  and  (not A166) );
 a51385a <=( (not A167)  and  a51384a );
 a51389a <=( A203  and  (not A202) );
 a51390a <=( A200  and  a51389a );
 a51391a <=( a51390a  and  a51385a );
 a51395a <=( A269  and  (not A266) );
 a51396a <=( (not A265)  and  a51395a );
 a51399a <=( A299  and  A298 );
 a51402a <=( (not A302)  and  A301 );
 a51403a <=( a51402a  and  a51399a );
 a51404a <=( a51403a  and  a51396a );
 a51408a <=( (not A199)  and  (not A166) );
 a51409a <=( (not A167)  and  a51408a );
 a51413a <=( A203  and  (not A202) );
 a51414a <=( A200  and  a51413a );
 a51415a <=( a51414a  and  a51409a );
 a51419a <=( A269  and  (not A266) );
 a51420a <=( (not A265)  and  a51419a );
 a51423a <=( (not A299)  and  A298 );
 a51426a <=( A302  and  (not A301) );
 a51427a <=( a51426a  and  a51423a );
 a51428a <=( a51427a  and  a51420a );
 a51432a <=( (not A199)  and  (not A166) );
 a51433a <=( (not A167)  and  a51432a );
 a51437a <=( A203  and  (not A202) );
 a51438a <=( A200  and  a51437a );
 a51439a <=( a51438a  and  a51433a );
 a51443a <=( A269  and  (not A266) );
 a51444a <=( (not A265)  and  a51443a );
 a51447a <=( A299  and  (not A298) );
 a51450a <=( A302  and  (not A301) );
 a51451a <=( a51450a  and  a51447a );
 a51452a <=( a51451a  and  a51444a );
 a51456a <=( (not A199)  and  (not A166) );
 a51457a <=( (not A167)  and  a51456a );
 a51461a <=( A203  and  (not A202) );
 a51462a <=( A200  and  a51461a );
 a51463a <=( a51462a  and  a51457a );
 a51467a <=( A269  and  (not A266) );
 a51468a <=( (not A265)  and  a51467a );
 a51471a <=( (not A299)  and  (not A298) );
 a51474a <=( (not A302)  and  A301 );
 a51475a <=( a51474a  and  a51471a );
 a51476a <=( a51475a  and  a51468a );
 a51480a <=( (not A199)  and  (not A166) );
 a51481a <=( (not A167)  and  a51480a );
 a51485a <=( A202  and  (not A201) );
 a51486a <=( A200  and  a51485a );
 a51487a <=( a51486a  and  a51481a );
 a51491a <=( A268  and  A266 );
 a51492a <=( A265  and  a51491a );
 a51495a <=( (not A298)  and  (not A269) );
 a51498a <=( (not A301)  and  (not A299) );
 a51499a <=( a51498a  and  a51495a );
 a51500a <=( a51499a  and  a51492a );
 a51504a <=( (not A199)  and  (not A166) );
 a51505a <=( (not A167)  and  a51504a );
 a51509a <=( A202  and  (not A201) );
 a51510a <=( A200  and  a51509a );
 a51511a <=( a51510a  and  a51505a );
 a51515a <=( A268  and  A266 );
 a51516a <=( A265  and  a51515a );
 a51519a <=( (not A298)  and  (not A269) );
 a51522a <=( A302  and  (not A299) );
 a51523a <=( a51522a  and  a51519a );
 a51524a <=( a51523a  and  a51516a );
 a51528a <=( (not A199)  and  (not A166) );
 a51529a <=( (not A167)  and  a51528a );
 a51533a <=( A202  and  (not A201) );
 a51534a <=( A200  and  a51533a );
 a51535a <=( a51534a  and  a51529a );
 a51539a <=( (not A268)  and  A266 );
 a51540a <=( (not A265)  and  a51539a );
 a51543a <=( (not A298)  and  A269 );
 a51546a <=( (not A301)  and  (not A299) );
 a51547a <=( a51546a  and  a51543a );
 a51548a <=( a51547a  and  a51540a );
 a51552a <=( (not A199)  and  (not A166) );
 a51553a <=( (not A167)  and  a51552a );
 a51557a <=( A202  and  (not A201) );
 a51558a <=( A200  and  a51557a );
 a51559a <=( a51558a  and  a51553a );
 a51563a <=( (not A268)  and  A266 );
 a51564a <=( (not A265)  and  a51563a );
 a51567a <=( (not A298)  and  A269 );
 a51570a <=( A302  and  (not A299) );
 a51571a <=( a51570a  and  a51567a );
 a51572a <=( a51571a  and  a51564a );
 a51576a <=( (not A199)  and  (not A166) );
 a51577a <=( (not A167)  and  a51576a );
 a51581a <=( A202  and  (not A201) );
 a51582a <=( A200  and  a51581a );
 a51583a <=( a51582a  and  a51577a );
 a51587a <=( (not A268)  and  (not A266) );
 a51588a <=( A265  and  a51587a );
 a51591a <=( (not A298)  and  A269 );
 a51594a <=( (not A301)  and  (not A299) );
 a51595a <=( a51594a  and  a51591a );
 a51596a <=( a51595a  and  a51588a );
 a51600a <=( (not A199)  and  (not A166) );
 a51601a <=( (not A167)  and  a51600a );
 a51605a <=( A202  and  (not A201) );
 a51606a <=( A200  and  a51605a );
 a51607a <=( a51606a  and  a51601a );
 a51611a <=( (not A268)  and  (not A266) );
 a51612a <=( A265  and  a51611a );
 a51615a <=( (not A298)  and  A269 );
 a51618a <=( A302  and  (not A299) );
 a51619a <=( a51618a  and  a51615a );
 a51620a <=( a51619a  and  a51612a );
 a51624a <=( (not A199)  and  (not A166) );
 a51625a <=( (not A167)  and  a51624a );
 a51629a <=( A202  and  (not A201) );
 a51630a <=( A200  and  a51629a );
 a51631a <=( a51630a  and  a51625a );
 a51635a <=( A268  and  (not A266) );
 a51636a <=( (not A265)  and  a51635a );
 a51639a <=( (not A298)  and  (not A269) );
 a51642a <=( (not A301)  and  (not A299) );
 a51643a <=( a51642a  and  a51639a );
 a51644a <=( a51643a  and  a51636a );
 a51648a <=( (not A199)  and  (not A166) );
 a51649a <=( (not A167)  and  a51648a );
 a51653a <=( A202  and  (not A201) );
 a51654a <=( A200  and  a51653a );
 a51655a <=( a51654a  and  a51649a );
 a51659a <=( A268  and  (not A266) );
 a51660a <=( (not A265)  and  a51659a );
 a51663a <=( (not A298)  and  (not A269) );
 a51666a <=( A302  and  (not A299) );
 a51667a <=( a51666a  and  a51663a );
 a51668a <=( a51667a  and  a51660a );
 a51672a <=( (not A199)  and  (not A166) );
 a51673a <=( (not A167)  and  a51672a );
 a51677a <=( (not A203)  and  (not A201) );
 a51678a <=( A200  and  a51677a );
 a51679a <=( a51678a  and  a51673a );
 a51683a <=( A268  and  A266 );
 a51684a <=( A265  and  a51683a );
 a51687a <=( (not A298)  and  (not A269) );
 a51690a <=( (not A301)  and  (not A299) );
 a51691a <=( a51690a  and  a51687a );
 a51692a <=( a51691a  and  a51684a );
 a51696a <=( (not A199)  and  (not A166) );
 a51697a <=( (not A167)  and  a51696a );
 a51701a <=( (not A203)  and  (not A201) );
 a51702a <=( A200  and  a51701a );
 a51703a <=( a51702a  and  a51697a );
 a51707a <=( A268  and  A266 );
 a51708a <=( A265  and  a51707a );
 a51711a <=( (not A298)  and  (not A269) );
 a51714a <=( A302  and  (not A299) );
 a51715a <=( a51714a  and  a51711a );
 a51716a <=( a51715a  and  a51708a );
 a51720a <=( (not A199)  and  (not A166) );
 a51721a <=( (not A167)  and  a51720a );
 a51725a <=( (not A203)  and  (not A201) );
 a51726a <=( A200  and  a51725a );
 a51727a <=( a51726a  and  a51721a );
 a51731a <=( (not A268)  and  A266 );
 a51732a <=( (not A265)  and  a51731a );
 a51735a <=( (not A298)  and  A269 );
 a51738a <=( (not A301)  and  (not A299) );
 a51739a <=( a51738a  and  a51735a );
 a51740a <=( a51739a  and  a51732a );
 a51744a <=( (not A199)  and  (not A166) );
 a51745a <=( (not A167)  and  a51744a );
 a51749a <=( (not A203)  and  (not A201) );
 a51750a <=( A200  and  a51749a );
 a51751a <=( a51750a  and  a51745a );
 a51755a <=( (not A268)  and  A266 );
 a51756a <=( (not A265)  and  a51755a );
 a51759a <=( (not A298)  and  A269 );
 a51762a <=( A302  and  (not A299) );
 a51763a <=( a51762a  and  a51759a );
 a51764a <=( a51763a  and  a51756a );
 a51768a <=( (not A199)  and  (not A166) );
 a51769a <=( (not A167)  and  a51768a );
 a51773a <=( (not A203)  and  (not A201) );
 a51774a <=( A200  and  a51773a );
 a51775a <=( a51774a  and  a51769a );
 a51779a <=( (not A268)  and  (not A266) );
 a51780a <=( A265  and  a51779a );
 a51783a <=( (not A298)  and  A269 );
 a51786a <=( (not A301)  and  (not A299) );
 a51787a <=( a51786a  and  a51783a );
 a51788a <=( a51787a  and  a51780a );
 a51792a <=( (not A199)  and  (not A166) );
 a51793a <=( (not A167)  and  a51792a );
 a51797a <=( (not A203)  and  (not A201) );
 a51798a <=( A200  and  a51797a );
 a51799a <=( a51798a  and  a51793a );
 a51803a <=( (not A268)  and  (not A266) );
 a51804a <=( A265  and  a51803a );
 a51807a <=( (not A298)  and  A269 );
 a51810a <=( A302  and  (not A299) );
 a51811a <=( a51810a  and  a51807a );
 a51812a <=( a51811a  and  a51804a );
 a51816a <=( (not A199)  and  (not A166) );
 a51817a <=( (not A167)  and  a51816a );
 a51821a <=( (not A203)  and  (not A201) );
 a51822a <=( A200  and  a51821a );
 a51823a <=( a51822a  and  a51817a );
 a51827a <=( A268  and  (not A266) );
 a51828a <=( (not A265)  and  a51827a );
 a51831a <=( (not A298)  and  (not A269) );
 a51834a <=( (not A301)  and  (not A299) );
 a51835a <=( a51834a  and  a51831a );
 a51836a <=( a51835a  and  a51828a );
 a51840a <=( (not A199)  and  (not A166) );
 a51841a <=( (not A167)  and  a51840a );
 a51845a <=( (not A203)  and  (not A201) );
 a51846a <=( A200  and  a51845a );
 a51847a <=( a51846a  and  a51841a );
 a51851a <=( A268  and  (not A266) );
 a51852a <=( (not A265)  and  a51851a );
 a51855a <=( (not A298)  and  (not A269) );
 a51858a <=( A302  and  (not A299) );
 a51859a <=( a51858a  and  a51855a );
 a51860a <=( a51859a  and  a51852a );
 a51864a <=( A199  and  (not A166) );
 a51865a <=( (not A167)  and  a51864a );
 a51869a <=( A203  and  (not A202) );
 a51870a <=( (not A200)  and  a51869a );
 a51871a <=( a51870a  and  a51865a );
 a51875a <=( (not A268)  and  (not A266) );
 a51876a <=( (not A265)  and  a51875a );
 a51879a <=( A299  and  A298 );
 a51882a <=( (not A302)  and  A301 );
 a51883a <=( a51882a  and  a51879a );
 a51884a <=( a51883a  and  a51876a );
 a51888a <=( A199  and  (not A166) );
 a51889a <=( (not A167)  and  a51888a );
 a51893a <=( A203  and  (not A202) );
 a51894a <=( (not A200)  and  a51893a );
 a51895a <=( a51894a  and  a51889a );
 a51899a <=( (not A268)  and  (not A266) );
 a51900a <=( (not A265)  and  a51899a );
 a51903a <=( (not A299)  and  A298 );
 a51906a <=( A302  and  (not A301) );
 a51907a <=( a51906a  and  a51903a );
 a51908a <=( a51907a  and  a51900a );
 a51912a <=( A199  and  (not A166) );
 a51913a <=( (not A167)  and  a51912a );
 a51917a <=( A203  and  (not A202) );
 a51918a <=( (not A200)  and  a51917a );
 a51919a <=( a51918a  and  a51913a );
 a51923a <=( (not A268)  and  (not A266) );
 a51924a <=( (not A265)  and  a51923a );
 a51927a <=( A299  and  (not A298) );
 a51930a <=( A302  and  (not A301) );
 a51931a <=( a51930a  and  a51927a );
 a51932a <=( a51931a  and  a51924a );
 a51936a <=( A199  and  (not A166) );
 a51937a <=( (not A167)  and  a51936a );
 a51941a <=( A203  and  (not A202) );
 a51942a <=( (not A200)  and  a51941a );
 a51943a <=( a51942a  and  a51937a );
 a51947a <=( (not A268)  and  (not A266) );
 a51948a <=( (not A265)  and  a51947a );
 a51951a <=( (not A299)  and  (not A298) );
 a51954a <=( (not A302)  and  A301 );
 a51955a <=( a51954a  and  a51951a );
 a51956a <=( a51955a  and  a51948a );
 a51960a <=( A199  and  (not A166) );
 a51961a <=( (not A167)  and  a51960a );
 a51965a <=( A203  and  (not A202) );
 a51966a <=( (not A200)  and  a51965a );
 a51967a <=( a51966a  and  a51961a );
 a51971a <=( A269  and  (not A266) );
 a51972a <=( (not A265)  and  a51971a );
 a51975a <=( A299  and  A298 );
 a51978a <=( (not A302)  and  A301 );
 a51979a <=( a51978a  and  a51975a );
 a51980a <=( a51979a  and  a51972a );
 a51984a <=( A199  and  (not A166) );
 a51985a <=( (not A167)  and  a51984a );
 a51989a <=( A203  and  (not A202) );
 a51990a <=( (not A200)  and  a51989a );
 a51991a <=( a51990a  and  a51985a );
 a51995a <=( A269  and  (not A266) );
 a51996a <=( (not A265)  and  a51995a );
 a51999a <=( (not A299)  and  A298 );
 a52002a <=( A302  and  (not A301) );
 a52003a <=( a52002a  and  a51999a );
 a52004a <=( a52003a  and  a51996a );
 a52008a <=( A199  and  (not A166) );
 a52009a <=( (not A167)  and  a52008a );
 a52013a <=( A203  and  (not A202) );
 a52014a <=( (not A200)  and  a52013a );
 a52015a <=( a52014a  and  a52009a );
 a52019a <=( A269  and  (not A266) );
 a52020a <=( (not A265)  and  a52019a );
 a52023a <=( A299  and  (not A298) );
 a52026a <=( A302  and  (not A301) );
 a52027a <=( a52026a  and  a52023a );
 a52028a <=( a52027a  and  a52020a );
 a52032a <=( A199  and  (not A166) );
 a52033a <=( (not A167)  and  a52032a );
 a52037a <=( A203  and  (not A202) );
 a52038a <=( (not A200)  and  a52037a );
 a52039a <=( a52038a  and  a52033a );
 a52043a <=( A269  and  (not A266) );
 a52044a <=( (not A265)  and  a52043a );
 a52047a <=( (not A299)  and  (not A298) );
 a52050a <=( (not A302)  and  A301 );
 a52051a <=( a52050a  and  a52047a );
 a52052a <=( a52051a  and  a52044a );
 a52056a <=( A199  and  (not A166) );
 a52057a <=( (not A167)  and  a52056a );
 a52061a <=( A202  and  (not A201) );
 a52062a <=( (not A200)  and  a52061a );
 a52063a <=( a52062a  and  a52057a );
 a52067a <=( A268  and  A266 );
 a52068a <=( A265  and  a52067a );
 a52071a <=( (not A298)  and  (not A269) );
 a52074a <=( (not A301)  and  (not A299) );
 a52075a <=( a52074a  and  a52071a );
 a52076a <=( a52075a  and  a52068a );
 a52080a <=( A199  and  (not A166) );
 a52081a <=( (not A167)  and  a52080a );
 a52085a <=( A202  and  (not A201) );
 a52086a <=( (not A200)  and  a52085a );
 a52087a <=( a52086a  and  a52081a );
 a52091a <=( A268  and  A266 );
 a52092a <=( A265  and  a52091a );
 a52095a <=( (not A298)  and  (not A269) );
 a52098a <=( A302  and  (not A299) );
 a52099a <=( a52098a  and  a52095a );
 a52100a <=( a52099a  and  a52092a );
 a52104a <=( A199  and  (not A166) );
 a52105a <=( (not A167)  and  a52104a );
 a52109a <=( A202  and  (not A201) );
 a52110a <=( (not A200)  and  a52109a );
 a52111a <=( a52110a  and  a52105a );
 a52115a <=( (not A268)  and  A266 );
 a52116a <=( (not A265)  and  a52115a );
 a52119a <=( (not A298)  and  A269 );
 a52122a <=( (not A301)  and  (not A299) );
 a52123a <=( a52122a  and  a52119a );
 a52124a <=( a52123a  and  a52116a );
 a52128a <=( A199  and  (not A166) );
 a52129a <=( (not A167)  and  a52128a );
 a52133a <=( A202  and  (not A201) );
 a52134a <=( (not A200)  and  a52133a );
 a52135a <=( a52134a  and  a52129a );
 a52139a <=( (not A268)  and  A266 );
 a52140a <=( (not A265)  and  a52139a );
 a52143a <=( (not A298)  and  A269 );
 a52146a <=( A302  and  (not A299) );
 a52147a <=( a52146a  and  a52143a );
 a52148a <=( a52147a  and  a52140a );
 a52152a <=( A199  and  (not A166) );
 a52153a <=( (not A167)  and  a52152a );
 a52157a <=( A202  and  (not A201) );
 a52158a <=( (not A200)  and  a52157a );
 a52159a <=( a52158a  and  a52153a );
 a52163a <=( (not A268)  and  (not A266) );
 a52164a <=( A265  and  a52163a );
 a52167a <=( (not A298)  and  A269 );
 a52170a <=( (not A301)  and  (not A299) );
 a52171a <=( a52170a  and  a52167a );
 a52172a <=( a52171a  and  a52164a );
 a52176a <=( A199  and  (not A166) );
 a52177a <=( (not A167)  and  a52176a );
 a52181a <=( A202  and  (not A201) );
 a52182a <=( (not A200)  and  a52181a );
 a52183a <=( a52182a  and  a52177a );
 a52187a <=( (not A268)  and  (not A266) );
 a52188a <=( A265  and  a52187a );
 a52191a <=( (not A298)  and  A269 );
 a52194a <=( A302  and  (not A299) );
 a52195a <=( a52194a  and  a52191a );
 a52196a <=( a52195a  and  a52188a );
 a52200a <=( A199  and  (not A166) );
 a52201a <=( (not A167)  and  a52200a );
 a52205a <=( A202  and  (not A201) );
 a52206a <=( (not A200)  and  a52205a );
 a52207a <=( a52206a  and  a52201a );
 a52211a <=( A268  and  (not A266) );
 a52212a <=( (not A265)  and  a52211a );
 a52215a <=( (not A298)  and  (not A269) );
 a52218a <=( (not A301)  and  (not A299) );
 a52219a <=( a52218a  and  a52215a );
 a52220a <=( a52219a  and  a52212a );
 a52224a <=( A199  and  (not A166) );
 a52225a <=( (not A167)  and  a52224a );
 a52229a <=( A202  and  (not A201) );
 a52230a <=( (not A200)  and  a52229a );
 a52231a <=( a52230a  and  a52225a );
 a52235a <=( A268  and  (not A266) );
 a52236a <=( (not A265)  and  a52235a );
 a52239a <=( (not A298)  and  (not A269) );
 a52242a <=( A302  and  (not A299) );
 a52243a <=( a52242a  and  a52239a );
 a52244a <=( a52243a  and  a52236a );
 a52248a <=( A199  and  (not A166) );
 a52249a <=( (not A167)  and  a52248a );
 a52253a <=( (not A203)  and  (not A201) );
 a52254a <=( (not A200)  and  a52253a );
 a52255a <=( a52254a  and  a52249a );
 a52259a <=( A268  and  A266 );
 a52260a <=( A265  and  a52259a );
 a52263a <=( (not A298)  and  (not A269) );
 a52266a <=( (not A301)  and  (not A299) );
 a52267a <=( a52266a  and  a52263a );
 a52268a <=( a52267a  and  a52260a );
 a52272a <=( A199  and  (not A166) );
 a52273a <=( (not A167)  and  a52272a );
 a52277a <=( (not A203)  and  (not A201) );
 a52278a <=( (not A200)  and  a52277a );
 a52279a <=( a52278a  and  a52273a );
 a52283a <=( A268  and  A266 );
 a52284a <=( A265  and  a52283a );
 a52287a <=( (not A298)  and  (not A269) );
 a52290a <=( A302  and  (not A299) );
 a52291a <=( a52290a  and  a52287a );
 a52292a <=( a52291a  and  a52284a );
 a52296a <=( A199  and  (not A166) );
 a52297a <=( (not A167)  and  a52296a );
 a52301a <=( (not A203)  and  (not A201) );
 a52302a <=( (not A200)  and  a52301a );
 a52303a <=( a52302a  and  a52297a );
 a52307a <=( (not A268)  and  A266 );
 a52308a <=( (not A265)  and  a52307a );
 a52311a <=( (not A298)  and  A269 );
 a52314a <=( (not A301)  and  (not A299) );
 a52315a <=( a52314a  and  a52311a );
 a52316a <=( a52315a  and  a52308a );
 a52320a <=( A199  and  (not A166) );
 a52321a <=( (not A167)  and  a52320a );
 a52325a <=( (not A203)  and  (not A201) );
 a52326a <=( (not A200)  and  a52325a );
 a52327a <=( a52326a  and  a52321a );
 a52331a <=( (not A268)  and  A266 );
 a52332a <=( (not A265)  and  a52331a );
 a52335a <=( (not A298)  and  A269 );
 a52338a <=( A302  and  (not A299) );
 a52339a <=( a52338a  and  a52335a );
 a52340a <=( a52339a  and  a52332a );
 a52344a <=( A199  and  (not A166) );
 a52345a <=( (not A167)  and  a52344a );
 a52349a <=( (not A203)  and  (not A201) );
 a52350a <=( (not A200)  and  a52349a );
 a52351a <=( a52350a  and  a52345a );
 a52355a <=( (not A268)  and  (not A266) );
 a52356a <=( A265  and  a52355a );
 a52359a <=( (not A298)  and  A269 );
 a52362a <=( (not A301)  and  (not A299) );
 a52363a <=( a52362a  and  a52359a );
 a52364a <=( a52363a  and  a52356a );
 a52368a <=( A199  and  (not A166) );
 a52369a <=( (not A167)  and  a52368a );
 a52373a <=( (not A203)  and  (not A201) );
 a52374a <=( (not A200)  and  a52373a );
 a52375a <=( a52374a  and  a52369a );
 a52379a <=( (not A268)  and  (not A266) );
 a52380a <=( A265  and  a52379a );
 a52383a <=( (not A298)  and  A269 );
 a52386a <=( A302  and  (not A299) );
 a52387a <=( a52386a  and  a52383a );
 a52388a <=( a52387a  and  a52380a );
 a52392a <=( A199  and  (not A166) );
 a52393a <=( (not A167)  and  a52392a );
 a52397a <=( (not A203)  and  (not A201) );
 a52398a <=( (not A200)  and  a52397a );
 a52399a <=( a52398a  and  a52393a );
 a52403a <=( A268  and  (not A266) );
 a52404a <=( (not A265)  and  a52403a );
 a52407a <=( (not A298)  and  (not A269) );
 a52410a <=( (not A301)  and  (not A299) );
 a52411a <=( a52410a  and  a52407a );
 a52412a <=( a52411a  and  a52404a );
 a52416a <=( A199  and  (not A166) );
 a52417a <=( (not A167)  and  a52416a );
 a52421a <=( (not A203)  and  (not A201) );
 a52422a <=( (not A200)  and  a52421a );
 a52423a <=( a52422a  and  a52417a );
 a52427a <=( A268  and  (not A266) );
 a52428a <=( (not A265)  and  a52427a );
 a52431a <=( (not A298)  and  (not A269) );
 a52434a <=( A302  and  (not A299) );
 a52435a <=( a52434a  and  a52431a );
 a52436a <=( a52435a  and  a52428a );
 a52440a <=( (not A199)  and  (not A166) );
 a52441a <=( (not A167)  and  a52440a );
 a52445a <=( A265  and  (not A202) );
 a52446a <=( (not A200)  and  a52445a );
 a52447a <=( a52446a  and  a52441a );
 a52451a <=( (not A269)  and  A268 );
 a52452a <=( A266  and  a52451a );
 a52455a <=( A299  and  A298 );
 a52458a <=( (not A301)  and  (not A300) );
 a52459a <=( a52458a  and  a52455a );
 a52460a <=( a52459a  and  a52452a );
 a52464a <=( (not A199)  and  (not A166) );
 a52465a <=( (not A167)  and  a52464a );
 a52469a <=( A265  and  (not A202) );
 a52470a <=( (not A200)  and  a52469a );
 a52471a <=( a52470a  and  a52465a );
 a52475a <=( (not A269)  and  A268 );
 a52476a <=( A266  and  a52475a );
 a52479a <=( A299  and  A298 );
 a52482a <=( A302  and  (not A300) );
 a52483a <=( a52482a  and  a52479a );
 a52484a <=( a52483a  and  a52476a );
 a52488a <=( (not A199)  and  (not A166) );
 a52489a <=( (not A167)  and  a52488a );
 a52493a <=( A265  and  (not A202) );
 a52494a <=( (not A200)  and  a52493a );
 a52495a <=( a52494a  and  a52489a );
 a52499a <=( (not A269)  and  A268 );
 a52500a <=( A266  and  a52499a );
 a52503a <=( (not A299)  and  A298 );
 a52506a <=( A301  and  (not A300) );
 a52507a <=( a52506a  and  a52503a );
 a52508a <=( a52507a  and  a52500a );
 a52512a <=( (not A199)  and  (not A166) );
 a52513a <=( (not A167)  and  a52512a );
 a52517a <=( A265  and  (not A202) );
 a52518a <=( (not A200)  and  a52517a );
 a52519a <=( a52518a  and  a52513a );
 a52523a <=( (not A269)  and  A268 );
 a52524a <=( A266  and  a52523a );
 a52527a <=( (not A299)  and  A298 );
 a52530a <=( (not A302)  and  (not A300) );
 a52531a <=( a52530a  and  a52527a );
 a52532a <=( a52531a  and  a52524a );
 a52536a <=( (not A199)  and  (not A166) );
 a52537a <=( (not A167)  and  a52536a );
 a52541a <=( A265  and  (not A202) );
 a52542a <=( (not A200)  and  a52541a );
 a52543a <=( a52542a  and  a52537a );
 a52547a <=( (not A269)  and  A268 );
 a52548a <=( A266  and  a52547a );
 a52551a <=( A299  and  (not A298) );
 a52554a <=( A301  and  (not A300) );
 a52555a <=( a52554a  and  a52551a );
 a52556a <=( a52555a  and  a52548a );
 a52560a <=( (not A199)  and  (not A166) );
 a52561a <=( (not A167)  and  a52560a );
 a52565a <=( A265  and  (not A202) );
 a52566a <=( (not A200)  and  a52565a );
 a52567a <=( a52566a  and  a52561a );
 a52571a <=( (not A269)  and  A268 );
 a52572a <=( A266  and  a52571a );
 a52575a <=( A299  and  (not A298) );
 a52578a <=( (not A302)  and  (not A300) );
 a52579a <=( a52578a  and  a52575a );
 a52580a <=( a52579a  and  a52572a );
 a52584a <=( (not A199)  and  (not A166) );
 a52585a <=( (not A167)  and  a52584a );
 a52589a <=( (not A265)  and  (not A202) );
 a52590a <=( (not A200)  and  a52589a );
 a52591a <=( a52590a  and  a52585a );
 a52595a <=( A269  and  (not A268) );
 a52596a <=( A266  and  a52595a );
 a52599a <=( A299  and  A298 );
 a52602a <=( (not A301)  and  (not A300) );
 a52603a <=( a52602a  and  a52599a );
 a52604a <=( a52603a  and  a52596a );
 a52608a <=( (not A199)  and  (not A166) );
 a52609a <=( (not A167)  and  a52608a );
 a52613a <=( (not A265)  and  (not A202) );
 a52614a <=( (not A200)  and  a52613a );
 a52615a <=( a52614a  and  a52609a );
 a52619a <=( A269  and  (not A268) );
 a52620a <=( A266  and  a52619a );
 a52623a <=( A299  and  A298 );
 a52626a <=( A302  and  (not A300) );
 a52627a <=( a52626a  and  a52623a );
 a52628a <=( a52627a  and  a52620a );
 a52632a <=( (not A199)  and  (not A166) );
 a52633a <=( (not A167)  and  a52632a );
 a52637a <=( (not A265)  and  (not A202) );
 a52638a <=( (not A200)  and  a52637a );
 a52639a <=( a52638a  and  a52633a );
 a52643a <=( A269  and  (not A268) );
 a52644a <=( A266  and  a52643a );
 a52647a <=( (not A299)  and  A298 );
 a52650a <=( A301  and  (not A300) );
 a52651a <=( a52650a  and  a52647a );
 a52652a <=( a52651a  and  a52644a );
 a52656a <=( (not A199)  and  (not A166) );
 a52657a <=( (not A167)  and  a52656a );
 a52661a <=( (not A265)  and  (not A202) );
 a52662a <=( (not A200)  and  a52661a );
 a52663a <=( a52662a  and  a52657a );
 a52667a <=( A269  and  (not A268) );
 a52668a <=( A266  and  a52667a );
 a52671a <=( (not A299)  and  A298 );
 a52674a <=( (not A302)  and  (not A300) );
 a52675a <=( a52674a  and  a52671a );
 a52676a <=( a52675a  and  a52668a );
 a52680a <=( (not A199)  and  (not A166) );
 a52681a <=( (not A167)  and  a52680a );
 a52685a <=( (not A265)  and  (not A202) );
 a52686a <=( (not A200)  and  a52685a );
 a52687a <=( a52686a  and  a52681a );
 a52691a <=( A269  and  (not A268) );
 a52692a <=( A266  and  a52691a );
 a52695a <=( A299  and  (not A298) );
 a52698a <=( A301  and  (not A300) );
 a52699a <=( a52698a  and  a52695a );
 a52700a <=( a52699a  and  a52692a );
 a52704a <=( (not A199)  and  (not A166) );
 a52705a <=( (not A167)  and  a52704a );
 a52709a <=( (not A265)  and  (not A202) );
 a52710a <=( (not A200)  and  a52709a );
 a52711a <=( a52710a  and  a52705a );
 a52715a <=( A269  and  (not A268) );
 a52716a <=( A266  and  a52715a );
 a52719a <=( A299  and  (not A298) );
 a52722a <=( (not A302)  and  (not A300) );
 a52723a <=( a52722a  and  a52719a );
 a52724a <=( a52723a  and  a52716a );
 a52728a <=( (not A199)  and  (not A166) );
 a52729a <=( (not A167)  and  a52728a );
 a52733a <=( A265  and  (not A202) );
 a52734a <=( (not A200)  and  a52733a );
 a52735a <=( a52734a  and  a52729a );
 a52739a <=( A269  and  (not A268) );
 a52740a <=( (not A266)  and  a52739a );
 a52743a <=( A299  and  A298 );
 a52746a <=( (not A301)  and  (not A300) );
 a52747a <=( a52746a  and  a52743a );
 a52748a <=( a52747a  and  a52740a );
 a52752a <=( (not A199)  and  (not A166) );
 a52753a <=( (not A167)  and  a52752a );
 a52757a <=( A265  and  (not A202) );
 a52758a <=( (not A200)  and  a52757a );
 a52759a <=( a52758a  and  a52753a );
 a52763a <=( A269  and  (not A268) );
 a52764a <=( (not A266)  and  a52763a );
 a52767a <=( A299  and  A298 );
 a52770a <=( A302  and  (not A300) );
 a52771a <=( a52770a  and  a52767a );
 a52772a <=( a52771a  and  a52764a );
 a52776a <=( (not A199)  and  (not A166) );
 a52777a <=( (not A167)  and  a52776a );
 a52781a <=( A265  and  (not A202) );
 a52782a <=( (not A200)  and  a52781a );
 a52783a <=( a52782a  and  a52777a );
 a52787a <=( A269  and  (not A268) );
 a52788a <=( (not A266)  and  a52787a );
 a52791a <=( (not A299)  and  A298 );
 a52794a <=( A301  and  (not A300) );
 a52795a <=( a52794a  and  a52791a );
 a52796a <=( a52795a  and  a52788a );
 a52800a <=( (not A199)  and  (not A166) );
 a52801a <=( (not A167)  and  a52800a );
 a52805a <=( A265  and  (not A202) );
 a52806a <=( (not A200)  and  a52805a );
 a52807a <=( a52806a  and  a52801a );
 a52811a <=( A269  and  (not A268) );
 a52812a <=( (not A266)  and  a52811a );
 a52815a <=( (not A299)  and  A298 );
 a52818a <=( (not A302)  and  (not A300) );
 a52819a <=( a52818a  and  a52815a );
 a52820a <=( a52819a  and  a52812a );
 a52824a <=( (not A199)  and  (not A166) );
 a52825a <=( (not A167)  and  a52824a );
 a52829a <=( A265  and  (not A202) );
 a52830a <=( (not A200)  and  a52829a );
 a52831a <=( a52830a  and  a52825a );
 a52835a <=( A269  and  (not A268) );
 a52836a <=( (not A266)  and  a52835a );
 a52839a <=( A299  and  (not A298) );
 a52842a <=( A301  and  (not A300) );
 a52843a <=( a52842a  and  a52839a );
 a52844a <=( a52843a  and  a52836a );
 a52848a <=( (not A199)  and  (not A166) );
 a52849a <=( (not A167)  and  a52848a );
 a52853a <=( A265  and  (not A202) );
 a52854a <=( (not A200)  and  a52853a );
 a52855a <=( a52854a  and  a52849a );
 a52859a <=( A269  and  (not A268) );
 a52860a <=( (not A266)  and  a52859a );
 a52863a <=( A299  and  (not A298) );
 a52866a <=( (not A302)  and  (not A300) );
 a52867a <=( a52866a  and  a52863a );
 a52868a <=( a52867a  and  a52860a );
 a52872a <=( (not A199)  and  (not A166) );
 a52873a <=( (not A167)  and  a52872a );
 a52877a <=( (not A265)  and  (not A202) );
 a52878a <=( (not A200)  and  a52877a );
 a52879a <=( a52878a  and  a52873a );
 a52883a <=( (not A269)  and  A268 );
 a52884a <=( (not A266)  and  a52883a );
 a52887a <=( A299  and  A298 );
 a52890a <=( (not A301)  and  (not A300) );
 a52891a <=( a52890a  and  a52887a );
 a52892a <=( a52891a  and  a52884a );
 a52896a <=( (not A199)  and  (not A166) );
 a52897a <=( (not A167)  and  a52896a );
 a52901a <=( (not A265)  and  (not A202) );
 a52902a <=( (not A200)  and  a52901a );
 a52903a <=( a52902a  and  a52897a );
 a52907a <=( (not A269)  and  A268 );
 a52908a <=( (not A266)  and  a52907a );
 a52911a <=( A299  and  A298 );
 a52914a <=( A302  and  (not A300) );
 a52915a <=( a52914a  and  a52911a );
 a52916a <=( a52915a  and  a52908a );
 a52920a <=( (not A199)  and  (not A166) );
 a52921a <=( (not A167)  and  a52920a );
 a52925a <=( (not A265)  and  (not A202) );
 a52926a <=( (not A200)  and  a52925a );
 a52927a <=( a52926a  and  a52921a );
 a52931a <=( (not A269)  and  A268 );
 a52932a <=( (not A266)  and  a52931a );
 a52935a <=( (not A299)  and  A298 );
 a52938a <=( A301  and  (not A300) );
 a52939a <=( a52938a  and  a52935a );
 a52940a <=( a52939a  and  a52932a );
 a52944a <=( (not A199)  and  (not A166) );
 a52945a <=( (not A167)  and  a52944a );
 a52949a <=( (not A265)  and  (not A202) );
 a52950a <=( (not A200)  and  a52949a );
 a52951a <=( a52950a  and  a52945a );
 a52955a <=( (not A269)  and  A268 );
 a52956a <=( (not A266)  and  a52955a );
 a52959a <=( (not A299)  and  A298 );
 a52962a <=( (not A302)  and  (not A300) );
 a52963a <=( a52962a  and  a52959a );
 a52964a <=( a52963a  and  a52956a );
 a52968a <=( (not A199)  and  (not A166) );
 a52969a <=( (not A167)  and  a52968a );
 a52973a <=( (not A265)  and  (not A202) );
 a52974a <=( (not A200)  and  a52973a );
 a52975a <=( a52974a  and  a52969a );
 a52979a <=( (not A269)  and  A268 );
 a52980a <=( (not A266)  and  a52979a );
 a52983a <=( A299  and  (not A298) );
 a52986a <=( A301  and  (not A300) );
 a52987a <=( a52986a  and  a52983a );
 a52988a <=( a52987a  and  a52980a );
 a52992a <=( (not A199)  and  (not A166) );
 a52993a <=( (not A167)  and  a52992a );
 a52997a <=( (not A265)  and  (not A202) );
 a52998a <=( (not A200)  and  a52997a );
 a52999a <=( a52998a  and  a52993a );
 a53003a <=( (not A269)  and  A268 );
 a53004a <=( (not A266)  and  a53003a );
 a53007a <=( A299  and  (not A298) );
 a53010a <=( (not A302)  and  (not A300) );
 a53011a <=( a53010a  and  a53007a );
 a53012a <=( a53011a  and  a53004a );
 a53016a <=( (not A199)  and  (not A166) );
 a53017a <=( (not A167)  and  a53016a );
 a53021a <=( A265  and  A203 );
 a53022a <=( (not A200)  and  a53021a );
 a53023a <=( a53022a  and  a53017a );
 a53027a <=( (not A269)  and  A268 );
 a53028a <=( A266  and  a53027a );
 a53031a <=( A299  and  A298 );
 a53034a <=( (not A301)  and  (not A300) );
 a53035a <=( a53034a  and  a53031a );
 a53036a <=( a53035a  and  a53028a );
 a53040a <=( (not A199)  and  (not A166) );
 a53041a <=( (not A167)  and  a53040a );
 a53045a <=( A265  and  A203 );
 a53046a <=( (not A200)  and  a53045a );
 a53047a <=( a53046a  and  a53041a );
 a53051a <=( (not A269)  and  A268 );
 a53052a <=( A266  and  a53051a );
 a53055a <=( A299  and  A298 );
 a53058a <=( A302  and  (not A300) );
 a53059a <=( a53058a  and  a53055a );
 a53060a <=( a53059a  and  a53052a );
 a53064a <=( (not A199)  and  (not A166) );
 a53065a <=( (not A167)  and  a53064a );
 a53069a <=( A265  and  A203 );
 a53070a <=( (not A200)  and  a53069a );
 a53071a <=( a53070a  and  a53065a );
 a53075a <=( (not A269)  and  A268 );
 a53076a <=( A266  and  a53075a );
 a53079a <=( (not A299)  and  A298 );
 a53082a <=( A301  and  (not A300) );
 a53083a <=( a53082a  and  a53079a );
 a53084a <=( a53083a  and  a53076a );
 a53088a <=( (not A199)  and  (not A166) );
 a53089a <=( (not A167)  and  a53088a );
 a53093a <=( A265  and  A203 );
 a53094a <=( (not A200)  and  a53093a );
 a53095a <=( a53094a  and  a53089a );
 a53099a <=( (not A269)  and  A268 );
 a53100a <=( A266  and  a53099a );
 a53103a <=( (not A299)  and  A298 );
 a53106a <=( (not A302)  and  (not A300) );
 a53107a <=( a53106a  and  a53103a );
 a53108a <=( a53107a  and  a53100a );
 a53112a <=( (not A199)  and  (not A166) );
 a53113a <=( (not A167)  and  a53112a );
 a53117a <=( A265  and  A203 );
 a53118a <=( (not A200)  and  a53117a );
 a53119a <=( a53118a  and  a53113a );
 a53123a <=( (not A269)  and  A268 );
 a53124a <=( A266  and  a53123a );
 a53127a <=( A299  and  (not A298) );
 a53130a <=( A301  and  (not A300) );
 a53131a <=( a53130a  and  a53127a );
 a53132a <=( a53131a  and  a53124a );
 a53136a <=( (not A199)  and  (not A166) );
 a53137a <=( (not A167)  and  a53136a );
 a53141a <=( A265  and  A203 );
 a53142a <=( (not A200)  and  a53141a );
 a53143a <=( a53142a  and  a53137a );
 a53147a <=( (not A269)  and  A268 );
 a53148a <=( A266  and  a53147a );
 a53151a <=( A299  and  (not A298) );
 a53154a <=( (not A302)  and  (not A300) );
 a53155a <=( a53154a  and  a53151a );
 a53156a <=( a53155a  and  a53148a );
 a53160a <=( (not A199)  and  (not A166) );
 a53161a <=( (not A167)  and  a53160a );
 a53165a <=( (not A265)  and  A203 );
 a53166a <=( (not A200)  and  a53165a );
 a53167a <=( a53166a  and  a53161a );
 a53171a <=( A269  and  (not A268) );
 a53172a <=( A266  and  a53171a );
 a53175a <=( A299  and  A298 );
 a53178a <=( (not A301)  and  (not A300) );
 a53179a <=( a53178a  and  a53175a );
 a53180a <=( a53179a  and  a53172a );
 a53184a <=( (not A199)  and  (not A166) );
 a53185a <=( (not A167)  and  a53184a );
 a53189a <=( (not A265)  and  A203 );
 a53190a <=( (not A200)  and  a53189a );
 a53191a <=( a53190a  and  a53185a );
 a53195a <=( A269  and  (not A268) );
 a53196a <=( A266  and  a53195a );
 a53199a <=( A299  and  A298 );
 a53202a <=( A302  and  (not A300) );
 a53203a <=( a53202a  and  a53199a );
 a53204a <=( a53203a  and  a53196a );
 a53208a <=( (not A199)  and  (not A166) );
 a53209a <=( (not A167)  and  a53208a );
 a53213a <=( (not A265)  and  A203 );
 a53214a <=( (not A200)  and  a53213a );
 a53215a <=( a53214a  and  a53209a );
 a53219a <=( A269  and  (not A268) );
 a53220a <=( A266  and  a53219a );
 a53223a <=( (not A299)  and  A298 );
 a53226a <=( A301  and  (not A300) );
 a53227a <=( a53226a  and  a53223a );
 a53228a <=( a53227a  and  a53220a );
 a53232a <=( (not A199)  and  (not A166) );
 a53233a <=( (not A167)  and  a53232a );
 a53237a <=( (not A265)  and  A203 );
 a53238a <=( (not A200)  and  a53237a );
 a53239a <=( a53238a  and  a53233a );
 a53243a <=( A269  and  (not A268) );
 a53244a <=( A266  and  a53243a );
 a53247a <=( (not A299)  and  A298 );
 a53250a <=( (not A302)  and  (not A300) );
 a53251a <=( a53250a  and  a53247a );
 a53252a <=( a53251a  and  a53244a );
 a53256a <=( (not A199)  and  (not A166) );
 a53257a <=( (not A167)  and  a53256a );
 a53261a <=( (not A265)  and  A203 );
 a53262a <=( (not A200)  and  a53261a );
 a53263a <=( a53262a  and  a53257a );
 a53267a <=( A269  and  (not A268) );
 a53268a <=( A266  and  a53267a );
 a53271a <=( A299  and  (not A298) );
 a53274a <=( A301  and  (not A300) );
 a53275a <=( a53274a  and  a53271a );
 a53276a <=( a53275a  and  a53268a );
 a53280a <=( (not A199)  and  (not A166) );
 a53281a <=( (not A167)  and  a53280a );
 a53285a <=( (not A265)  and  A203 );
 a53286a <=( (not A200)  and  a53285a );
 a53287a <=( a53286a  and  a53281a );
 a53291a <=( A269  and  (not A268) );
 a53292a <=( A266  and  a53291a );
 a53295a <=( A299  and  (not A298) );
 a53298a <=( (not A302)  and  (not A300) );
 a53299a <=( a53298a  and  a53295a );
 a53300a <=( a53299a  and  a53292a );
 a53304a <=( (not A199)  and  (not A166) );
 a53305a <=( (not A167)  and  a53304a );
 a53309a <=( A265  and  A203 );
 a53310a <=( (not A200)  and  a53309a );
 a53311a <=( a53310a  and  a53305a );
 a53315a <=( A269  and  (not A268) );
 a53316a <=( (not A266)  and  a53315a );
 a53319a <=( A299  and  A298 );
 a53322a <=( (not A301)  and  (not A300) );
 a53323a <=( a53322a  and  a53319a );
 a53324a <=( a53323a  and  a53316a );
 a53328a <=( (not A199)  and  (not A166) );
 a53329a <=( (not A167)  and  a53328a );
 a53333a <=( A265  and  A203 );
 a53334a <=( (not A200)  and  a53333a );
 a53335a <=( a53334a  and  a53329a );
 a53339a <=( A269  and  (not A268) );
 a53340a <=( (not A266)  and  a53339a );
 a53343a <=( A299  and  A298 );
 a53346a <=( A302  and  (not A300) );
 a53347a <=( a53346a  and  a53343a );
 a53348a <=( a53347a  and  a53340a );
 a53352a <=( (not A199)  and  (not A166) );
 a53353a <=( (not A167)  and  a53352a );
 a53357a <=( A265  and  A203 );
 a53358a <=( (not A200)  and  a53357a );
 a53359a <=( a53358a  and  a53353a );
 a53363a <=( A269  and  (not A268) );
 a53364a <=( (not A266)  and  a53363a );
 a53367a <=( (not A299)  and  A298 );
 a53370a <=( A301  and  (not A300) );
 a53371a <=( a53370a  and  a53367a );
 a53372a <=( a53371a  and  a53364a );
 a53376a <=( (not A199)  and  (not A166) );
 a53377a <=( (not A167)  and  a53376a );
 a53381a <=( A265  and  A203 );
 a53382a <=( (not A200)  and  a53381a );
 a53383a <=( a53382a  and  a53377a );
 a53387a <=( A269  and  (not A268) );
 a53388a <=( (not A266)  and  a53387a );
 a53391a <=( (not A299)  and  A298 );
 a53394a <=( (not A302)  and  (not A300) );
 a53395a <=( a53394a  and  a53391a );
 a53396a <=( a53395a  and  a53388a );
 a53400a <=( (not A199)  and  (not A166) );
 a53401a <=( (not A167)  and  a53400a );
 a53405a <=( A265  and  A203 );
 a53406a <=( (not A200)  and  a53405a );
 a53407a <=( a53406a  and  a53401a );
 a53411a <=( A269  and  (not A268) );
 a53412a <=( (not A266)  and  a53411a );
 a53415a <=( A299  and  (not A298) );
 a53418a <=( A301  and  (not A300) );
 a53419a <=( a53418a  and  a53415a );
 a53420a <=( a53419a  and  a53412a );
 a53424a <=( (not A199)  and  (not A166) );
 a53425a <=( (not A167)  and  a53424a );
 a53429a <=( A265  and  A203 );
 a53430a <=( (not A200)  and  a53429a );
 a53431a <=( a53430a  and  a53425a );
 a53435a <=( A269  and  (not A268) );
 a53436a <=( (not A266)  and  a53435a );
 a53439a <=( A299  and  (not A298) );
 a53442a <=( (not A302)  and  (not A300) );
 a53443a <=( a53442a  and  a53439a );
 a53444a <=( a53443a  and  a53436a );
 a53448a <=( (not A199)  and  (not A166) );
 a53449a <=( (not A167)  and  a53448a );
 a53453a <=( (not A265)  and  A203 );
 a53454a <=( (not A200)  and  a53453a );
 a53455a <=( a53454a  and  a53449a );
 a53459a <=( (not A269)  and  A268 );
 a53460a <=( (not A266)  and  a53459a );
 a53463a <=( A299  and  A298 );
 a53466a <=( (not A301)  and  (not A300) );
 a53467a <=( a53466a  and  a53463a );
 a53468a <=( a53467a  and  a53460a );
 a53472a <=( (not A199)  and  (not A166) );
 a53473a <=( (not A167)  and  a53472a );
 a53477a <=( (not A265)  and  A203 );
 a53478a <=( (not A200)  and  a53477a );
 a53479a <=( a53478a  and  a53473a );
 a53483a <=( (not A269)  and  A268 );
 a53484a <=( (not A266)  and  a53483a );
 a53487a <=( A299  and  A298 );
 a53490a <=( A302  and  (not A300) );
 a53491a <=( a53490a  and  a53487a );
 a53492a <=( a53491a  and  a53484a );
 a53496a <=( (not A199)  and  (not A166) );
 a53497a <=( (not A167)  and  a53496a );
 a53501a <=( (not A265)  and  A203 );
 a53502a <=( (not A200)  and  a53501a );
 a53503a <=( a53502a  and  a53497a );
 a53507a <=( (not A269)  and  A268 );
 a53508a <=( (not A266)  and  a53507a );
 a53511a <=( (not A299)  and  A298 );
 a53514a <=( A301  and  (not A300) );
 a53515a <=( a53514a  and  a53511a );
 a53516a <=( a53515a  and  a53508a );
 a53520a <=( (not A199)  and  (not A166) );
 a53521a <=( (not A167)  and  a53520a );
 a53525a <=( (not A265)  and  A203 );
 a53526a <=( (not A200)  and  a53525a );
 a53527a <=( a53526a  and  a53521a );
 a53531a <=( (not A269)  and  A268 );
 a53532a <=( (not A266)  and  a53531a );
 a53535a <=( (not A299)  and  A298 );
 a53538a <=( (not A302)  and  (not A300) );
 a53539a <=( a53538a  and  a53535a );
 a53540a <=( a53539a  and  a53532a );
 a53544a <=( (not A199)  and  (not A166) );
 a53545a <=( (not A167)  and  a53544a );
 a53549a <=( (not A265)  and  A203 );
 a53550a <=( (not A200)  and  a53549a );
 a53551a <=( a53550a  and  a53545a );
 a53555a <=( (not A269)  and  A268 );
 a53556a <=( (not A266)  and  a53555a );
 a53559a <=( A299  and  (not A298) );
 a53562a <=( A301  and  (not A300) );
 a53563a <=( a53562a  and  a53559a );
 a53564a <=( a53563a  and  a53556a );
 a53568a <=( (not A199)  and  (not A166) );
 a53569a <=( (not A167)  and  a53568a );
 a53573a <=( (not A265)  and  A203 );
 a53574a <=( (not A200)  and  a53573a );
 a53575a <=( a53574a  and  a53569a );
 a53579a <=( (not A269)  and  A268 );
 a53580a <=( (not A266)  and  a53579a );
 a53583a <=( A299  and  (not A298) );
 a53586a <=( (not A302)  and  (not A300) );
 a53587a <=( a53586a  and  a53583a );
 a53588a <=( a53587a  and  a53580a );
 a53592a <=( (not A199)  and  (not A166) );
 a53593a <=( (not A167)  and  a53592a );
 a53597a <=( (not A203)  and  A202 );
 a53598a <=( (not A200)  and  a53597a );
 a53599a <=( a53598a  and  a53593a );
 a53603a <=( (not A268)  and  (not A266) );
 a53604a <=( (not A265)  and  a53603a );
 a53607a <=( A299  and  A298 );
 a53610a <=( (not A302)  and  A301 );
 a53611a <=( a53610a  and  a53607a );
 a53612a <=( a53611a  and  a53604a );
 a53616a <=( (not A199)  and  (not A166) );
 a53617a <=( (not A167)  and  a53616a );
 a53621a <=( (not A203)  and  A202 );
 a53622a <=( (not A200)  and  a53621a );
 a53623a <=( a53622a  and  a53617a );
 a53627a <=( (not A268)  and  (not A266) );
 a53628a <=( (not A265)  and  a53627a );
 a53631a <=( (not A299)  and  A298 );
 a53634a <=( A302  and  (not A301) );
 a53635a <=( a53634a  and  a53631a );
 a53636a <=( a53635a  and  a53628a );
 a53640a <=( (not A199)  and  (not A166) );
 a53641a <=( (not A167)  and  a53640a );
 a53645a <=( (not A203)  and  A202 );
 a53646a <=( (not A200)  and  a53645a );
 a53647a <=( a53646a  and  a53641a );
 a53651a <=( (not A268)  and  (not A266) );
 a53652a <=( (not A265)  and  a53651a );
 a53655a <=( A299  and  (not A298) );
 a53658a <=( A302  and  (not A301) );
 a53659a <=( a53658a  and  a53655a );
 a53660a <=( a53659a  and  a53652a );
 a53664a <=( (not A199)  and  (not A166) );
 a53665a <=( (not A167)  and  a53664a );
 a53669a <=( (not A203)  and  A202 );
 a53670a <=( (not A200)  and  a53669a );
 a53671a <=( a53670a  and  a53665a );
 a53675a <=( (not A268)  and  (not A266) );
 a53676a <=( (not A265)  and  a53675a );
 a53679a <=( (not A299)  and  (not A298) );
 a53682a <=( (not A302)  and  A301 );
 a53683a <=( a53682a  and  a53679a );
 a53684a <=( a53683a  and  a53676a );
 a53688a <=( (not A199)  and  (not A166) );
 a53689a <=( (not A167)  and  a53688a );
 a53693a <=( (not A203)  and  A202 );
 a53694a <=( (not A200)  and  a53693a );
 a53695a <=( a53694a  and  a53689a );
 a53699a <=( A269  and  (not A266) );
 a53700a <=( (not A265)  and  a53699a );
 a53703a <=( A299  and  A298 );
 a53706a <=( (not A302)  and  A301 );
 a53707a <=( a53706a  and  a53703a );
 a53708a <=( a53707a  and  a53700a );
 a53712a <=( (not A199)  and  (not A166) );
 a53713a <=( (not A167)  and  a53712a );
 a53717a <=( (not A203)  and  A202 );
 a53718a <=( (not A200)  and  a53717a );
 a53719a <=( a53718a  and  a53713a );
 a53723a <=( A269  and  (not A266) );
 a53724a <=( (not A265)  and  a53723a );
 a53727a <=( (not A299)  and  A298 );
 a53730a <=( A302  and  (not A301) );
 a53731a <=( a53730a  and  a53727a );
 a53732a <=( a53731a  and  a53724a );
 a53736a <=( (not A199)  and  (not A166) );
 a53737a <=( (not A167)  and  a53736a );
 a53741a <=( (not A203)  and  A202 );
 a53742a <=( (not A200)  and  a53741a );
 a53743a <=( a53742a  and  a53737a );
 a53747a <=( A269  and  (not A266) );
 a53748a <=( (not A265)  and  a53747a );
 a53751a <=( A299  and  (not A298) );
 a53754a <=( A302  and  (not A301) );
 a53755a <=( a53754a  and  a53751a );
 a53756a <=( a53755a  and  a53748a );
 a53760a <=( (not A199)  and  (not A166) );
 a53761a <=( (not A167)  and  a53760a );
 a53765a <=( (not A203)  and  A202 );
 a53766a <=( (not A200)  and  a53765a );
 a53767a <=( a53766a  and  a53761a );
 a53771a <=( A269  and  (not A266) );
 a53772a <=( (not A265)  and  a53771a );
 a53775a <=( (not A299)  and  (not A298) );
 a53778a <=( (not A302)  and  A301 );
 a53779a <=( a53778a  and  a53775a );
 a53780a <=( a53779a  and  a53772a );
 a53784a <=( A199  and  (not A167) );
 a53785a <=( (not A168)  and  a53784a );
 a53789a <=( (not A203)  and  A202 );
 a53790a <=( A200  and  a53789a );
 a53791a <=( a53790a  and  a53785a );
 a53795a <=( (not A268)  and  (not A266) );
 a53796a <=( (not A265)  and  a53795a );
 a53799a <=( A299  and  A298 );
 a53802a <=( (not A302)  and  A301 );
 a53803a <=( a53802a  and  a53799a );
 a53804a <=( a53803a  and  a53796a );
 a53808a <=( A199  and  (not A167) );
 a53809a <=( (not A168)  and  a53808a );
 a53813a <=( (not A203)  and  A202 );
 a53814a <=( A200  and  a53813a );
 a53815a <=( a53814a  and  a53809a );
 a53819a <=( (not A268)  and  (not A266) );
 a53820a <=( (not A265)  and  a53819a );
 a53823a <=( (not A299)  and  A298 );
 a53826a <=( A302  and  (not A301) );
 a53827a <=( a53826a  and  a53823a );
 a53828a <=( a53827a  and  a53820a );
 a53832a <=( A199  and  (not A167) );
 a53833a <=( (not A168)  and  a53832a );
 a53837a <=( (not A203)  and  A202 );
 a53838a <=( A200  and  a53837a );
 a53839a <=( a53838a  and  a53833a );
 a53843a <=( (not A268)  and  (not A266) );
 a53844a <=( (not A265)  and  a53843a );
 a53847a <=( A299  and  (not A298) );
 a53850a <=( A302  and  (not A301) );
 a53851a <=( a53850a  and  a53847a );
 a53852a <=( a53851a  and  a53844a );
 a53856a <=( A199  and  (not A167) );
 a53857a <=( (not A168)  and  a53856a );
 a53861a <=( (not A203)  and  A202 );
 a53862a <=( A200  and  a53861a );
 a53863a <=( a53862a  and  a53857a );
 a53867a <=( (not A268)  and  (not A266) );
 a53868a <=( (not A265)  and  a53867a );
 a53871a <=( (not A299)  and  (not A298) );
 a53874a <=( (not A302)  and  A301 );
 a53875a <=( a53874a  and  a53871a );
 a53876a <=( a53875a  and  a53868a );
 a53880a <=( A199  and  (not A167) );
 a53881a <=( (not A168)  and  a53880a );
 a53885a <=( (not A203)  and  A202 );
 a53886a <=( A200  and  a53885a );
 a53887a <=( a53886a  and  a53881a );
 a53891a <=( A269  and  (not A266) );
 a53892a <=( (not A265)  and  a53891a );
 a53895a <=( A299  and  A298 );
 a53898a <=( (not A302)  and  A301 );
 a53899a <=( a53898a  and  a53895a );
 a53900a <=( a53899a  and  a53892a );
 a53904a <=( A199  and  (not A167) );
 a53905a <=( (not A168)  and  a53904a );
 a53909a <=( (not A203)  and  A202 );
 a53910a <=( A200  and  a53909a );
 a53911a <=( a53910a  and  a53905a );
 a53915a <=( A269  and  (not A266) );
 a53916a <=( (not A265)  and  a53915a );
 a53919a <=( (not A299)  and  A298 );
 a53922a <=( A302  and  (not A301) );
 a53923a <=( a53922a  and  a53919a );
 a53924a <=( a53923a  and  a53916a );
 a53928a <=( A199  and  (not A167) );
 a53929a <=( (not A168)  and  a53928a );
 a53933a <=( (not A203)  and  A202 );
 a53934a <=( A200  and  a53933a );
 a53935a <=( a53934a  and  a53929a );
 a53939a <=( A269  and  (not A266) );
 a53940a <=( (not A265)  and  a53939a );
 a53943a <=( A299  and  (not A298) );
 a53946a <=( A302  and  (not A301) );
 a53947a <=( a53946a  and  a53943a );
 a53948a <=( a53947a  and  a53940a );
 a53952a <=( A199  and  (not A167) );
 a53953a <=( (not A168)  and  a53952a );
 a53957a <=( (not A203)  and  A202 );
 a53958a <=( A200  and  a53957a );
 a53959a <=( a53958a  and  a53953a );
 a53963a <=( A269  and  (not A266) );
 a53964a <=( (not A265)  and  a53963a );
 a53967a <=( (not A299)  and  (not A298) );
 a53970a <=( (not A302)  and  A301 );
 a53971a <=( a53970a  and  a53967a );
 a53972a <=( a53971a  and  a53964a );
 a53976a <=( A199  and  (not A167) );
 a53977a <=( (not A168)  and  a53976a );
 a53981a <=( (not A202)  and  (not A201) );
 a53982a <=( A200  and  a53981a );
 a53983a <=( a53982a  and  a53977a );
 a53987a <=( A268  and  A266 );
 a53988a <=( A265  and  a53987a );
 a53991a <=( (not A298)  and  (not A269) );
 a53994a <=( (not A301)  and  (not A299) );
 a53995a <=( a53994a  and  a53991a );
 a53996a <=( a53995a  and  a53988a );
 a54000a <=( A199  and  (not A167) );
 a54001a <=( (not A168)  and  a54000a );
 a54005a <=( (not A202)  and  (not A201) );
 a54006a <=( A200  and  a54005a );
 a54007a <=( a54006a  and  a54001a );
 a54011a <=( A268  and  A266 );
 a54012a <=( A265  and  a54011a );
 a54015a <=( (not A298)  and  (not A269) );
 a54018a <=( A302  and  (not A299) );
 a54019a <=( a54018a  and  a54015a );
 a54020a <=( a54019a  and  a54012a );
 a54024a <=( A199  and  (not A167) );
 a54025a <=( (not A168)  and  a54024a );
 a54029a <=( (not A202)  and  (not A201) );
 a54030a <=( A200  and  a54029a );
 a54031a <=( a54030a  and  a54025a );
 a54035a <=( (not A268)  and  A266 );
 a54036a <=( (not A265)  and  a54035a );
 a54039a <=( (not A298)  and  A269 );
 a54042a <=( (not A301)  and  (not A299) );
 a54043a <=( a54042a  and  a54039a );
 a54044a <=( a54043a  and  a54036a );
 a54048a <=( A199  and  (not A167) );
 a54049a <=( (not A168)  and  a54048a );
 a54053a <=( (not A202)  and  (not A201) );
 a54054a <=( A200  and  a54053a );
 a54055a <=( a54054a  and  a54049a );
 a54059a <=( (not A268)  and  A266 );
 a54060a <=( (not A265)  and  a54059a );
 a54063a <=( (not A298)  and  A269 );
 a54066a <=( A302  and  (not A299) );
 a54067a <=( a54066a  and  a54063a );
 a54068a <=( a54067a  and  a54060a );
 a54072a <=( A199  and  (not A167) );
 a54073a <=( (not A168)  and  a54072a );
 a54077a <=( (not A202)  and  (not A201) );
 a54078a <=( A200  and  a54077a );
 a54079a <=( a54078a  and  a54073a );
 a54083a <=( (not A268)  and  (not A266) );
 a54084a <=( A265  and  a54083a );
 a54087a <=( (not A298)  and  A269 );
 a54090a <=( (not A301)  and  (not A299) );
 a54091a <=( a54090a  and  a54087a );
 a54092a <=( a54091a  and  a54084a );
 a54096a <=( A199  and  (not A167) );
 a54097a <=( (not A168)  and  a54096a );
 a54101a <=( (not A202)  and  (not A201) );
 a54102a <=( A200  and  a54101a );
 a54103a <=( a54102a  and  a54097a );
 a54107a <=( (not A268)  and  (not A266) );
 a54108a <=( A265  and  a54107a );
 a54111a <=( (not A298)  and  A269 );
 a54114a <=( A302  and  (not A299) );
 a54115a <=( a54114a  and  a54111a );
 a54116a <=( a54115a  and  a54108a );
 a54120a <=( A199  and  (not A167) );
 a54121a <=( (not A168)  and  a54120a );
 a54125a <=( (not A202)  and  (not A201) );
 a54126a <=( A200  and  a54125a );
 a54127a <=( a54126a  and  a54121a );
 a54131a <=( A268  and  (not A266) );
 a54132a <=( (not A265)  and  a54131a );
 a54135a <=( (not A298)  and  (not A269) );
 a54138a <=( (not A301)  and  (not A299) );
 a54139a <=( a54138a  and  a54135a );
 a54140a <=( a54139a  and  a54132a );
 a54144a <=( A199  and  (not A167) );
 a54145a <=( (not A168)  and  a54144a );
 a54149a <=( (not A202)  and  (not A201) );
 a54150a <=( A200  and  a54149a );
 a54151a <=( a54150a  and  a54145a );
 a54155a <=( A268  and  (not A266) );
 a54156a <=( (not A265)  and  a54155a );
 a54159a <=( (not A298)  and  (not A269) );
 a54162a <=( A302  and  (not A299) );
 a54163a <=( a54162a  and  a54159a );
 a54164a <=( a54163a  and  a54156a );
 a54168a <=( A199  and  (not A167) );
 a54169a <=( (not A168)  and  a54168a );
 a54173a <=( A203  and  (not A201) );
 a54174a <=( A200  and  a54173a );
 a54175a <=( a54174a  and  a54169a );
 a54179a <=( A268  and  A266 );
 a54180a <=( A265  and  a54179a );
 a54183a <=( (not A298)  and  (not A269) );
 a54186a <=( (not A301)  and  (not A299) );
 a54187a <=( a54186a  and  a54183a );
 a54188a <=( a54187a  and  a54180a );
 a54192a <=( A199  and  (not A167) );
 a54193a <=( (not A168)  and  a54192a );
 a54197a <=( A203  and  (not A201) );
 a54198a <=( A200  and  a54197a );
 a54199a <=( a54198a  and  a54193a );
 a54203a <=( A268  and  A266 );
 a54204a <=( A265  and  a54203a );
 a54207a <=( (not A298)  and  (not A269) );
 a54210a <=( A302  and  (not A299) );
 a54211a <=( a54210a  and  a54207a );
 a54212a <=( a54211a  and  a54204a );
 a54216a <=( A199  and  (not A167) );
 a54217a <=( (not A168)  and  a54216a );
 a54221a <=( A203  and  (not A201) );
 a54222a <=( A200  and  a54221a );
 a54223a <=( a54222a  and  a54217a );
 a54227a <=( (not A268)  and  A266 );
 a54228a <=( (not A265)  and  a54227a );
 a54231a <=( (not A298)  and  A269 );
 a54234a <=( (not A301)  and  (not A299) );
 a54235a <=( a54234a  and  a54231a );
 a54236a <=( a54235a  and  a54228a );
 a54240a <=( A199  and  (not A167) );
 a54241a <=( (not A168)  and  a54240a );
 a54245a <=( A203  and  (not A201) );
 a54246a <=( A200  and  a54245a );
 a54247a <=( a54246a  and  a54241a );
 a54251a <=( (not A268)  and  A266 );
 a54252a <=( (not A265)  and  a54251a );
 a54255a <=( (not A298)  and  A269 );
 a54258a <=( A302  and  (not A299) );
 a54259a <=( a54258a  and  a54255a );
 a54260a <=( a54259a  and  a54252a );
 a54264a <=( A199  and  (not A167) );
 a54265a <=( (not A168)  and  a54264a );
 a54269a <=( A203  and  (not A201) );
 a54270a <=( A200  and  a54269a );
 a54271a <=( a54270a  and  a54265a );
 a54275a <=( (not A268)  and  (not A266) );
 a54276a <=( A265  and  a54275a );
 a54279a <=( (not A298)  and  A269 );
 a54282a <=( (not A301)  and  (not A299) );
 a54283a <=( a54282a  and  a54279a );
 a54284a <=( a54283a  and  a54276a );
 a54288a <=( A199  and  (not A167) );
 a54289a <=( (not A168)  and  a54288a );
 a54293a <=( A203  and  (not A201) );
 a54294a <=( A200  and  a54293a );
 a54295a <=( a54294a  and  a54289a );
 a54299a <=( (not A268)  and  (not A266) );
 a54300a <=( A265  and  a54299a );
 a54303a <=( (not A298)  and  A269 );
 a54306a <=( A302  and  (not A299) );
 a54307a <=( a54306a  and  a54303a );
 a54308a <=( a54307a  and  a54300a );
 a54312a <=( A199  and  (not A167) );
 a54313a <=( (not A168)  and  a54312a );
 a54317a <=( A203  and  (not A201) );
 a54318a <=( A200  and  a54317a );
 a54319a <=( a54318a  and  a54313a );
 a54323a <=( A268  and  (not A266) );
 a54324a <=( (not A265)  and  a54323a );
 a54327a <=( (not A298)  and  (not A269) );
 a54330a <=( (not A301)  and  (not A299) );
 a54331a <=( a54330a  and  a54327a );
 a54332a <=( a54331a  and  a54324a );
 a54336a <=( A199  and  (not A167) );
 a54337a <=( (not A168)  and  a54336a );
 a54341a <=( A203  and  (not A201) );
 a54342a <=( A200  and  a54341a );
 a54343a <=( a54342a  and  a54337a );
 a54347a <=( A268  and  (not A266) );
 a54348a <=( (not A265)  and  a54347a );
 a54351a <=( (not A298)  and  (not A269) );
 a54354a <=( A302  and  (not A299) );
 a54355a <=( a54354a  and  a54351a );
 a54356a <=( a54355a  and  a54348a );
 a54360a <=( (not A199)  and  (not A167) );
 a54361a <=( (not A168)  and  a54360a );
 a54365a <=( A203  and  (not A202) );
 a54366a <=( A200  and  a54365a );
 a54367a <=( a54366a  and  a54361a );
 a54371a <=( (not A268)  and  (not A266) );
 a54372a <=( (not A265)  and  a54371a );
 a54375a <=( A299  and  A298 );
 a54378a <=( (not A302)  and  A301 );
 a54379a <=( a54378a  and  a54375a );
 a54380a <=( a54379a  and  a54372a );
 a54384a <=( (not A199)  and  (not A167) );
 a54385a <=( (not A168)  and  a54384a );
 a54389a <=( A203  and  (not A202) );
 a54390a <=( A200  and  a54389a );
 a54391a <=( a54390a  and  a54385a );
 a54395a <=( (not A268)  and  (not A266) );
 a54396a <=( (not A265)  and  a54395a );
 a54399a <=( (not A299)  and  A298 );
 a54402a <=( A302  and  (not A301) );
 a54403a <=( a54402a  and  a54399a );
 a54404a <=( a54403a  and  a54396a );
 a54408a <=( (not A199)  and  (not A167) );
 a54409a <=( (not A168)  and  a54408a );
 a54413a <=( A203  and  (not A202) );
 a54414a <=( A200  and  a54413a );
 a54415a <=( a54414a  and  a54409a );
 a54419a <=( (not A268)  and  (not A266) );
 a54420a <=( (not A265)  and  a54419a );
 a54423a <=( A299  and  (not A298) );
 a54426a <=( A302  and  (not A301) );
 a54427a <=( a54426a  and  a54423a );
 a54428a <=( a54427a  and  a54420a );
 a54432a <=( (not A199)  and  (not A167) );
 a54433a <=( (not A168)  and  a54432a );
 a54437a <=( A203  and  (not A202) );
 a54438a <=( A200  and  a54437a );
 a54439a <=( a54438a  and  a54433a );
 a54443a <=( (not A268)  and  (not A266) );
 a54444a <=( (not A265)  and  a54443a );
 a54447a <=( (not A299)  and  (not A298) );
 a54450a <=( (not A302)  and  A301 );
 a54451a <=( a54450a  and  a54447a );
 a54452a <=( a54451a  and  a54444a );
 a54456a <=( (not A199)  and  (not A167) );
 a54457a <=( (not A168)  and  a54456a );
 a54461a <=( A203  and  (not A202) );
 a54462a <=( A200  and  a54461a );
 a54463a <=( a54462a  and  a54457a );
 a54467a <=( A269  and  (not A266) );
 a54468a <=( (not A265)  and  a54467a );
 a54471a <=( A299  and  A298 );
 a54474a <=( (not A302)  and  A301 );
 a54475a <=( a54474a  and  a54471a );
 a54476a <=( a54475a  and  a54468a );
 a54480a <=( (not A199)  and  (not A167) );
 a54481a <=( (not A168)  and  a54480a );
 a54485a <=( A203  and  (not A202) );
 a54486a <=( A200  and  a54485a );
 a54487a <=( a54486a  and  a54481a );
 a54491a <=( A269  and  (not A266) );
 a54492a <=( (not A265)  and  a54491a );
 a54495a <=( (not A299)  and  A298 );
 a54498a <=( A302  and  (not A301) );
 a54499a <=( a54498a  and  a54495a );
 a54500a <=( a54499a  and  a54492a );
 a54504a <=( (not A199)  and  (not A167) );
 a54505a <=( (not A168)  and  a54504a );
 a54509a <=( A203  and  (not A202) );
 a54510a <=( A200  and  a54509a );
 a54511a <=( a54510a  and  a54505a );
 a54515a <=( A269  and  (not A266) );
 a54516a <=( (not A265)  and  a54515a );
 a54519a <=( A299  and  (not A298) );
 a54522a <=( A302  and  (not A301) );
 a54523a <=( a54522a  and  a54519a );
 a54524a <=( a54523a  and  a54516a );
 a54528a <=( (not A199)  and  (not A167) );
 a54529a <=( (not A168)  and  a54528a );
 a54533a <=( A203  and  (not A202) );
 a54534a <=( A200  and  a54533a );
 a54535a <=( a54534a  and  a54529a );
 a54539a <=( A269  and  (not A266) );
 a54540a <=( (not A265)  and  a54539a );
 a54543a <=( (not A299)  and  (not A298) );
 a54546a <=( (not A302)  and  A301 );
 a54547a <=( a54546a  and  a54543a );
 a54548a <=( a54547a  and  a54540a );
 a54552a <=( (not A199)  and  (not A167) );
 a54553a <=( (not A168)  and  a54552a );
 a54557a <=( A202  and  (not A201) );
 a54558a <=( A200  and  a54557a );
 a54559a <=( a54558a  and  a54553a );
 a54563a <=( A268  and  A266 );
 a54564a <=( A265  and  a54563a );
 a54567a <=( (not A298)  and  (not A269) );
 a54570a <=( (not A301)  and  (not A299) );
 a54571a <=( a54570a  and  a54567a );
 a54572a <=( a54571a  and  a54564a );
 a54576a <=( (not A199)  and  (not A167) );
 a54577a <=( (not A168)  and  a54576a );
 a54581a <=( A202  and  (not A201) );
 a54582a <=( A200  and  a54581a );
 a54583a <=( a54582a  and  a54577a );
 a54587a <=( A268  and  A266 );
 a54588a <=( A265  and  a54587a );
 a54591a <=( (not A298)  and  (not A269) );
 a54594a <=( A302  and  (not A299) );
 a54595a <=( a54594a  and  a54591a );
 a54596a <=( a54595a  and  a54588a );
 a54600a <=( (not A199)  and  (not A167) );
 a54601a <=( (not A168)  and  a54600a );
 a54605a <=( A202  and  (not A201) );
 a54606a <=( A200  and  a54605a );
 a54607a <=( a54606a  and  a54601a );
 a54611a <=( (not A268)  and  A266 );
 a54612a <=( (not A265)  and  a54611a );
 a54615a <=( (not A298)  and  A269 );
 a54618a <=( (not A301)  and  (not A299) );
 a54619a <=( a54618a  and  a54615a );
 a54620a <=( a54619a  and  a54612a );
 a54624a <=( (not A199)  and  (not A167) );
 a54625a <=( (not A168)  and  a54624a );
 a54629a <=( A202  and  (not A201) );
 a54630a <=( A200  and  a54629a );
 a54631a <=( a54630a  and  a54625a );
 a54635a <=( (not A268)  and  A266 );
 a54636a <=( (not A265)  and  a54635a );
 a54639a <=( (not A298)  and  A269 );
 a54642a <=( A302  and  (not A299) );
 a54643a <=( a54642a  and  a54639a );
 a54644a <=( a54643a  and  a54636a );
 a54648a <=( (not A199)  and  (not A167) );
 a54649a <=( (not A168)  and  a54648a );
 a54653a <=( A202  and  (not A201) );
 a54654a <=( A200  and  a54653a );
 a54655a <=( a54654a  and  a54649a );
 a54659a <=( (not A268)  and  (not A266) );
 a54660a <=( A265  and  a54659a );
 a54663a <=( (not A298)  and  A269 );
 a54666a <=( (not A301)  and  (not A299) );
 a54667a <=( a54666a  and  a54663a );
 a54668a <=( a54667a  and  a54660a );
 a54672a <=( (not A199)  and  (not A167) );
 a54673a <=( (not A168)  and  a54672a );
 a54677a <=( A202  and  (not A201) );
 a54678a <=( A200  and  a54677a );
 a54679a <=( a54678a  and  a54673a );
 a54683a <=( (not A268)  and  (not A266) );
 a54684a <=( A265  and  a54683a );
 a54687a <=( (not A298)  and  A269 );
 a54690a <=( A302  and  (not A299) );
 a54691a <=( a54690a  and  a54687a );
 a54692a <=( a54691a  and  a54684a );
 a54696a <=( (not A199)  and  (not A167) );
 a54697a <=( (not A168)  and  a54696a );
 a54701a <=( A202  and  (not A201) );
 a54702a <=( A200  and  a54701a );
 a54703a <=( a54702a  and  a54697a );
 a54707a <=( A268  and  (not A266) );
 a54708a <=( (not A265)  and  a54707a );
 a54711a <=( (not A298)  and  (not A269) );
 a54714a <=( (not A301)  and  (not A299) );
 a54715a <=( a54714a  and  a54711a );
 a54716a <=( a54715a  and  a54708a );
 a54720a <=( (not A199)  and  (not A167) );
 a54721a <=( (not A168)  and  a54720a );
 a54725a <=( A202  and  (not A201) );
 a54726a <=( A200  and  a54725a );
 a54727a <=( a54726a  and  a54721a );
 a54731a <=( A268  and  (not A266) );
 a54732a <=( (not A265)  and  a54731a );
 a54735a <=( (not A298)  and  (not A269) );
 a54738a <=( A302  and  (not A299) );
 a54739a <=( a54738a  and  a54735a );
 a54740a <=( a54739a  and  a54732a );
 a54744a <=( (not A199)  and  (not A167) );
 a54745a <=( (not A168)  and  a54744a );
 a54749a <=( (not A203)  and  (not A201) );
 a54750a <=( A200  and  a54749a );
 a54751a <=( a54750a  and  a54745a );
 a54755a <=( A268  and  A266 );
 a54756a <=( A265  and  a54755a );
 a54759a <=( (not A298)  and  (not A269) );
 a54762a <=( (not A301)  and  (not A299) );
 a54763a <=( a54762a  and  a54759a );
 a54764a <=( a54763a  and  a54756a );
 a54768a <=( (not A199)  and  (not A167) );
 a54769a <=( (not A168)  and  a54768a );
 a54773a <=( (not A203)  and  (not A201) );
 a54774a <=( A200  and  a54773a );
 a54775a <=( a54774a  and  a54769a );
 a54779a <=( A268  and  A266 );
 a54780a <=( A265  and  a54779a );
 a54783a <=( (not A298)  and  (not A269) );
 a54786a <=( A302  and  (not A299) );
 a54787a <=( a54786a  and  a54783a );
 a54788a <=( a54787a  and  a54780a );
 a54792a <=( (not A199)  and  (not A167) );
 a54793a <=( (not A168)  and  a54792a );
 a54797a <=( (not A203)  and  (not A201) );
 a54798a <=( A200  and  a54797a );
 a54799a <=( a54798a  and  a54793a );
 a54803a <=( (not A268)  and  A266 );
 a54804a <=( (not A265)  and  a54803a );
 a54807a <=( (not A298)  and  A269 );
 a54810a <=( (not A301)  and  (not A299) );
 a54811a <=( a54810a  and  a54807a );
 a54812a <=( a54811a  and  a54804a );
 a54816a <=( (not A199)  and  (not A167) );
 a54817a <=( (not A168)  and  a54816a );
 a54821a <=( (not A203)  and  (not A201) );
 a54822a <=( A200  and  a54821a );
 a54823a <=( a54822a  and  a54817a );
 a54827a <=( (not A268)  and  A266 );
 a54828a <=( (not A265)  and  a54827a );
 a54831a <=( (not A298)  and  A269 );
 a54834a <=( A302  and  (not A299) );
 a54835a <=( a54834a  and  a54831a );
 a54836a <=( a54835a  and  a54828a );
 a54840a <=( (not A199)  and  (not A167) );
 a54841a <=( (not A168)  and  a54840a );
 a54845a <=( (not A203)  and  (not A201) );
 a54846a <=( A200  and  a54845a );
 a54847a <=( a54846a  and  a54841a );
 a54851a <=( (not A268)  and  (not A266) );
 a54852a <=( A265  and  a54851a );
 a54855a <=( (not A298)  and  A269 );
 a54858a <=( (not A301)  and  (not A299) );
 a54859a <=( a54858a  and  a54855a );
 a54860a <=( a54859a  and  a54852a );
 a54864a <=( (not A199)  and  (not A167) );
 a54865a <=( (not A168)  and  a54864a );
 a54869a <=( (not A203)  and  (not A201) );
 a54870a <=( A200  and  a54869a );
 a54871a <=( a54870a  and  a54865a );
 a54875a <=( (not A268)  and  (not A266) );
 a54876a <=( A265  and  a54875a );
 a54879a <=( (not A298)  and  A269 );
 a54882a <=( A302  and  (not A299) );
 a54883a <=( a54882a  and  a54879a );
 a54884a <=( a54883a  and  a54876a );
 a54888a <=( (not A199)  and  (not A167) );
 a54889a <=( (not A168)  and  a54888a );
 a54893a <=( (not A203)  and  (not A201) );
 a54894a <=( A200  and  a54893a );
 a54895a <=( a54894a  and  a54889a );
 a54899a <=( A268  and  (not A266) );
 a54900a <=( (not A265)  and  a54899a );
 a54903a <=( (not A298)  and  (not A269) );
 a54906a <=( (not A301)  and  (not A299) );
 a54907a <=( a54906a  and  a54903a );
 a54908a <=( a54907a  and  a54900a );
 a54912a <=( (not A199)  and  (not A167) );
 a54913a <=( (not A168)  and  a54912a );
 a54917a <=( (not A203)  and  (not A201) );
 a54918a <=( A200  and  a54917a );
 a54919a <=( a54918a  and  a54913a );
 a54923a <=( A268  and  (not A266) );
 a54924a <=( (not A265)  and  a54923a );
 a54927a <=( (not A298)  and  (not A269) );
 a54930a <=( A302  and  (not A299) );
 a54931a <=( a54930a  and  a54927a );
 a54932a <=( a54931a  and  a54924a );
 a54936a <=( A199  and  (not A167) );
 a54937a <=( (not A168)  and  a54936a );
 a54941a <=( A203  and  (not A202) );
 a54942a <=( (not A200)  and  a54941a );
 a54943a <=( a54942a  and  a54937a );
 a54947a <=( (not A268)  and  (not A266) );
 a54948a <=( (not A265)  and  a54947a );
 a54951a <=( A299  and  A298 );
 a54954a <=( (not A302)  and  A301 );
 a54955a <=( a54954a  and  a54951a );
 a54956a <=( a54955a  and  a54948a );
 a54960a <=( A199  and  (not A167) );
 a54961a <=( (not A168)  and  a54960a );
 a54965a <=( A203  and  (not A202) );
 a54966a <=( (not A200)  and  a54965a );
 a54967a <=( a54966a  and  a54961a );
 a54971a <=( (not A268)  and  (not A266) );
 a54972a <=( (not A265)  and  a54971a );
 a54975a <=( (not A299)  and  A298 );
 a54978a <=( A302  and  (not A301) );
 a54979a <=( a54978a  and  a54975a );
 a54980a <=( a54979a  and  a54972a );
 a54984a <=( A199  and  (not A167) );
 a54985a <=( (not A168)  and  a54984a );
 a54989a <=( A203  and  (not A202) );
 a54990a <=( (not A200)  and  a54989a );
 a54991a <=( a54990a  and  a54985a );
 a54995a <=( (not A268)  and  (not A266) );
 a54996a <=( (not A265)  and  a54995a );
 a54999a <=( A299  and  (not A298) );
 a55002a <=( A302  and  (not A301) );
 a55003a <=( a55002a  and  a54999a );
 a55004a <=( a55003a  and  a54996a );
 a55008a <=( A199  and  (not A167) );
 a55009a <=( (not A168)  and  a55008a );
 a55013a <=( A203  and  (not A202) );
 a55014a <=( (not A200)  and  a55013a );
 a55015a <=( a55014a  and  a55009a );
 a55019a <=( (not A268)  and  (not A266) );
 a55020a <=( (not A265)  and  a55019a );
 a55023a <=( (not A299)  and  (not A298) );
 a55026a <=( (not A302)  and  A301 );
 a55027a <=( a55026a  and  a55023a );
 a55028a <=( a55027a  and  a55020a );
 a55032a <=( A199  and  (not A167) );
 a55033a <=( (not A168)  and  a55032a );
 a55037a <=( A203  and  (not A202) );
 a55038a <=( (not A200)  and  a55037a );
 a55039a <=( a55038a  and  a55033a );
 a55043a <=( A269  and  (not A266) );
 a55044a <=( (not A265)  and  a55043a );
 a55047a <=( A299  and  A298 );
 a55050a <=( (not A302)  and  A301 );
 a55051a <=( a55050a  and  a55047a );
 a55052a <=( a55051a  and  a55044a );
 a55056a <=( A199  and  (not A167) );
 a55057a <=( (not A168)  and  a55056a );
 a55061a <=( A203  and  (not A202) );
 a55062a <=( (not A200)  and  a55061a );
 a55063a <=( a55062a  and  a55057a );
 a55067a <=( A269  and  (not A266) );
 a55068a <=( (not A265)  and  a55067a );
 a55071a <=( (not A299)  and  A298 );
 a55074a <=( A302  and  (not A301) );
 a55075a <=( a55074a  and  a55071a );
 a55076a <=( a55075a  and  a55068a );
 a55080a <=( A199  and  (not A167) );
 a55081a <=( (not A168)  and  a55080a );
 a55085a <=( A203  and  (not A202) );
 a55086a <=( (not A200)  and  a55085a );
 a55087a <=( a55086a  and  a55081a );
 a55091a <=( A269  and  (not A266) );
 a55092a <=( (not A265)  and  a55091a );
 a55095a <=( A299  and  (not A298) );
 a55098a <=( A302  and  (not A301) );
 a55099a <=( a55098a  and  a55095a );
 a55100a <=( a55099a  and  a55092a );
 a55104a <=( A199  and  (not A167) );
 a55105a <=( (not A168)  and  a55104a );
 a55109a <=( A203  and  (not A202) );
 a55110a <=( (not A200)  and  a55109a );
 a55111a <=( a55110a  and  a55105a );
 a55115a <=( A269  and  (not A266) );
 a55116a <=( (not A265)  and  a55115a );
 a55119a <=( (not A299)  and  (not A298) );
 a55122a <=( (not A302)  and  A301 );
 a55123a <=( a55122a  and  a55119a );
 a55124a <=( a55123a  and  a55116a );
 a55128a <=( A199  and  (not A167) );
 a55129a <=( (not A168)  and  a55128a );
 a55133a <=( A202  and  (not A201) );
 a55134a <=( (not A200)  and  a55133a );
 a55135a <=( a55134a  and  a55129a );
 a55139a <=( A268  and  A266 );
 a55140a <=( A265  and  a55139a );
 a55143a <=( (not A298)  and  (not A269) );
 a55146a <=( (not A301)  and  (not A299) );
 a55147a <=( a55146a  and  a55143a );
 a55148a <=( a55147a  and  a55140a );
 a55152a <=( A199  and  (not A167) );
 a55153a <=( (not A168)  and  a55152a );
 a55157a <=( A202  and  (not A201) );
 a55158a <=( (not A200)  and  a55157a );
 a55159a <=( a55158a  and  a55153a );
 a55163a <=( A268  and  A266 );
 a55164a <=( A265  and  a55163a );
 a55167a <=( (not A298)  and  (not A269) );
 a55170a <=( A302  and  (not A299) );
 a55171a <=( a55170a  and  a55167a );
 a55172a <=( a55171a  and  a55164a );
 a55176a <=( A199  and  (not A167) );
 a55177a <=( (not A168)  and  a55176a );
 a55181a <=( A202  and  (not A201) );
 a55182a <=( (not A200)  and  a55181a );
 a55183a <=( a55182a  and  a55177a );
 a55187a <=( (not A268)  and  A266 );
 a55188a <=( (not A265)  and  a55187a );
 a55191a <=( (not A298)  and  A269 );
 a55194a <=( (not A301)  and  (not A299) );
 a55195a <=( a55194a  and  a55191a );
 a55196a <=( a55195a  and  a55188a );
 a55200a <=( A199  and  (not A167) );
 a55201a <=( (not A168)  and  a55200a );
 a55205a <=( A202  and  (not A201) );
 a55206a <=( (not A200)  and  a55205a );
 a55207a <=( a55206a  and  a55201a );
 a55211a <=( (not A268)  and  A266 );
 a55212a <=( (not A265)  and  a55211a );
 a55215a <=( (not A298)  and  A269 );
 a55218a <=( A302  and  (not A299) );
 a55219a <=( a55218a  and  a55215a );
 a55220a <=( a55219a  and  a55212a );
 a55224a <=( A199  and  (not A167) );
 a55225a <=( (not A168)  and  a55224a );
 a55229a <=( A202  and  (not A201) );
 a55230a <=( (not A200)  and  a55229a );
 a55231a <=( a55230a  and  a55225a );
 a55235a <=( (not A268)  and  (not A266) );
 a55236a <=( A265  and  a55235a );
 a55239a <=( (not A298)  and  A269 );
 a55242a <=( (not A301)  and  (not A299) );
 a55243a <=( a55242a  and  a55239a );
 a55244a <=( a55243a  and  a55236a );
 a55248a <=( A199  and  (not A167) );
 a55249a <=( (not A168)  and  a55248a );
 a55253a <=( A202  and  (not A201) );
 a55254a <=( (not A200)  and  a55253a );
 a55255a <=( a55254a  and  a55249a );
 a55259a <=( (not A268)  and  (not A266) );
 a55260a <=( A265  and  a55259a );
 a55263a <=( (not A298)  and  A269 );
 a55266a <=( A302  and  (not A299) );
 a55267a <=( a55266a  and  a55263a );
 a55268a <=( a55267a  and  a55260a );
 a55272a <=( A199  and  (not A167) );
 a55273a <=( (not A168)  and  a55272a );
 a55277a <=( A202  and  (not A201) );
 a55278a <=( (not A200)  and  a55277a );
 a55279a <=( a55278a  and  a55273a );
 a55283a <=( A268  and  (not A266) );
 a55284a <=( (not A265)  and  a55283a );
 a55287a <=( (not A298)  and  (not A269) );
 a55290a <=( (not A301)  and  (not A299) );
 a55291a <=( a55290a  and  a55287a );
 a55292a <=( a55291a  and  a55284a );
 a55296a <=( A199  and  (not A167) );
 a55297a <=( (not A168)  and  a55296a );
 a55301a <=( A202  and  (not A201) );
 a55302a <=( (not A200)  and  a55301a );
 a55303a <=( a55302a  and  a55297a );
 a55307a <=( A268  and  (not A266) );
 a55308a <=( (not A265)  and  a55307a );
 a55311a <=( (not A298)  and  (not A269) );
 a55314a <=( A302  and  (not A299) );
 a55315a <=( a55314a  and  a55311a );
 a55316a <=( a55315a  and  a55308a );
 a55320a <=( A199  and  (not A167) );
 a55321a <=( (not A168)  and  a55320a );
 a55325a <=( (not A203)  and  (not A201) );
 a55326a <=( (not A200)  and  a55325a );
 a55327a <=( a55326a  and  a55321a );
 a55331a <=( A268  and  A266 );
 a55332a <=( A265  and  a55331a );
 a55335a <=( (not A298)  and  (not A269) );
 a55338a <=( (not A301)  and  (not A299) );
 a55339a <=( a55338a  and  a55335a );
 a55340a <=( a55339a  and  a55332a );
 a55344a <=( A199  and  (not A167) );
 a55345a <=( (not A168)  and  a55344a );
 a55349a <=( (not A203)  and  (not A201) );
 a55350a <=( (not A200)  and  a55349a );
 a55351a <=( a55350a  and  a55345a );
 a55355a <=( A268  and  A266 );
 a55356a <=( A265  and  a55355a );
 a55359a <=( (not A298)  and  (not A269) );
 a55362a <=( A302  and  (not A299) );
 a55363a <=( a55362a  and  a55359a );
 a55364a <=( a55363a  and  a55356a );
 a55368a <=( A199  and  (not A167) );
 a55369a <=( (not A168)  and  a55368a );
 a55373a <=( (not A203)  and  (not A201) );
 a55374a <=( (not A200)  and  a55373a );
 a55375a <=( a55374a  and  a55369a );
 a55379a <=( (not A268)  and  A266 );
 a55380a <=( (not A265)  and  a55379a );
 a55383a <=( (not A298)  and  A269 );
 a55386a <=( (not A301)  and  (not A299) );
 a55387a <=( a55386a  and  a55383a );
 a55388a <=( a55387a  and  a55380a );
 a55392a <=( A199  and  (not A167) );
 a55393a <=( (not A168)  and  a55392a );
 a55397a <=( (not A203)  and  (not A201) );
 a55398a <=( (not A200)  and  a55397a );
 a55399a <=( a55398a  and  a55393a );
 a55403a <=( (not A268)  and  A266 );
 a55404a <=( (not A265)  and  a55403a );
 a55407a <=( (not A298)  and  A269 );
 a55410a <=( A302  and  (not A299) );
 a55411a <=( a55410a  and  a55407a );
 a55412a <=( a55411a  and  a55404a );
 a55416a <=( A199  and  (not A167) );
 a55417a <=( (not A168)  and  a55416a );
 a55421a <=( (not A203)  and  (not A201) );
 a55422a <=( (not A200)  and  a55421a );
 a55423a <=( a55422a  and  a55417a );
 a55427a <=( (not A268)  and  (not A266) );
 a55428a <=( A265  and  a55427a );
 a55431a <=( (not A298)  and  A269 );
 a55434a <=( (not A301)  and  (not A299) );
 a55435a <=( a55434a  and  a55431a );
 a55436a <=( a55435a  and  a55428a );
 a55440a <=( A199  and  (not A167) );
 a55441a <=( (not A168)  and  a55440a );
 a55445a <=( (not A203)  and  (not A201) );
 a55446a <=( (not A200)  and  a55445a );
 a55447a <=( a55446a  and  a55441a );
 a55451a <=( (not A268)  and  (not A266) );
 a55452a <=( A265  and  a55451a );
 a55455a <=( (not A298)  and  A269 );
 a55458a <=( A302  and  (not A299) );
 a55459a <=( a55458a  and  a55455a );
 a55460a <=( a55459a  and  a55452a );
 a55464a <=( A199  and  (not A167) );
 a55465a <=( (not A168)  and  a55464a );
 a55469a <=( (not A203)  and  (not A201) );
 a55470a <=( (not A200)  and  a55469a );
 a55471a <=( a55470a  and  a55465a );
 a55475a <=( A268  and  (not A266) );
 a55476a <=( (not A265)  and  a55475a );
 a55479a <=( (not A298)  and  (not A269) );
 a55482a <=( (not A301)  and  (not A299) );
 a55483a <=( a55482a  and  a55479a );
 a55484a <=( a55483a  and  a55476a );
 a55488a <=( A199  and  (not A167) );
 a55489a <=( (not A168)  and  a55488a );
 a55493a <=( (not A203)  and  (not A201) );
 a55494a <=( (not A200)  and  a55493a );
 a55495a <=( a55494a  and  a55489a );
 a55499a <=( A268  and  (not A266) );
 a55500a <=( (not A265)  and  a55499a );
 a55503a <=( (not A298)  and  (not A269) );
 a55506a <=( A302  and  (not A299) );
 a55507a <=( a55506a  and  a55503a );
 a55508a <=( a55507a  and  a55500a );
 a55512a <=( (not A199)  and  (not A167) );
 a55513a <=( (not A168)  and  a55512a );
 a55517a <=( A265  and  (not A202) );
 a55518a <=( (not A200)  and  a55517a );
 a55519a <=( a55518a  and  a55513a );
 a55523a <=( (not A269)  and  A268 );
 a55524a <=( A266  and  a55523a );
 a55527a <=( A299  and  A298 );
 a55530a <=( (not A301)  and  (not A300) );
 a55531a <=( a55530a  and  a55527a );
 a55532a <=( a55531a  and  a55524a );
 a55536a <=( (not A199)  and  (not A167) );
 a55537a <=( (not A168)  and  a55536a );
 a55541a <=( A265  and  (not A202) );
 a55542a <=( (not A200)  and  a55541a );
 a55543a <=( a55542a  and  a55537a );
 a55547a <=( (not A269)  and  A268 );
 a55548a <=( A266  and  a55547a );
 a55551a <=( A299  and  A298 );
 a55554a <=( A302  and  (not A300) );
 a55555a <=( a55554a  and  a55551a );
 a55556a <=( a55555a  and  a55548a );
 a55560a <=( (not A199)  and  (not A167) );
 a55561a <=( (not A168)  and  a55560a );
 a55565a <=( A265  and  (not A202) );
 a55566a <=( (not A200)  and  a55565a );
 a55567a <=( a55566a  and  a55561a );
 a55571a <=( (not A269)  and  A268 );
 a55572a <=( A266  and  a55571a );
 a55575a <=( (not A299)  and  A298 );
 a55578a <=( A301  and  (not A300) );
 a55579a <=( a55578a  and  a55575a );
 a55580a <=( a55579a  and  a55572a );
 a55584a <=( (not A199)  and  (not A167) );
 a55585a <=( (not A168)  and  a55584a );
 a55589a <=( A265  and  (not A202) );
 a55590a <=( (not A200)  and  a55589a );
 a55591a <=( a55590a  and  a55585a );
 a55595a <=( (not A269)  and  A268 );
 a55596a <=( A266  and  a55595a );
 a55599a <=( (not A299)  and  A298 );
 a55602a <=( (not A302)  and  (not A300) );
 a55603a <=( a55602a  and  a55599a );
 a55604a <=( a55603a  and  a55596a );
 a55608a <=( (not A199)  and  (not A167) );
 a55609a <=( (not A168)  and  a55608a );
 a55613a <=( A265  and  (not A202) );
 a55614a <=( (not A200)  and  a55613a );
 a55615a <=( a55614a  and  a55609a );
 a55619a <=( (not A269)  and  A268 );
 a55620a <=( A266  and  a55619a );
 a55623a <=( A299  and  (not A298) );
 a55626a <=( A301  and  (not A300) );
 a55627a <=( a55626a  and  a55623a );
 a55628a <=( a55627a  and  a55620a );
 a55632a <=( (not A199)  and  (not A167) );
 a55633a <=( (not A168)  and  a55632a );
 a55637a <=( A265  and  (not A202) );
 a55638a <=( (not A200)  and  a55637a );
 a55639a <=( a55638a  and  a55633a );
 a55643a <=( (not A269)  and  A268 );
 a55644a <=( A266  and  a55643a );
 a55647a <=( A299  and  (not A298) );
 a55650a <=( (not A302)  and  (not A300) );
 a55651a <=( a55650a  and  a55647a );
 a55652a <=( a55651a  and  a55644a );
 a55656a <=( (not A199)  and  (not A167) );
 a55657a <=( (not A168)  and  a55656a );
 a55661a <=( (not A265)  and  (not A202) );
 a55662a <=( (not A200)  and  a55661a );
 a55663a <=( a55662a  and  a55657a );
 a55667a <=( A269  and  (not A268) );
 a55668a <=( A266  and  a55667a );
 a55671a <=( A299  and  A298 );
 a55674a <=( (not A301)  and  (not A300) );
 a55675a <=( a55674a  and  a55671a );
 a55676a <=( a55675a  and  a55668a );
 a55680a <=( (not A199)  and  (not A167) );
 a55681a <=( (not A168)  and  a55680a );
 a55685a <=( (not A265)  and  (not A202) );
 a55686a <=( (not A200)  and  a55685a );
 a55687a <=( a55686a  and  a55681a );
 a55691a <=( A269  and  (not A268) );
 a55692a <=( A266  and  a55691a );
 a55695a <=( A299  and  A298 );
 a55698a <=( A302  and  (not A300) );
 a55699a <=( a55698a  and  a55695a );
 a55700a <=( a55699a  and  a55692a );
 a55704a <=( (not A199)  and  (not A167) );
 a55705a <=( (not A168)  and  a55704a );
 a55709a <=( (not A265)  and  (not A202) );
 a55710a <=( (not A200)  and  a55709a );
 a55711a <=( a55710a  and  a55705a );
 a55715a <=( A269  and  (not A268) );
 a55716a <=( A266  and  a55715a );
 a55719a <=( (not A299)  and  A298 );
 a55722a <=( A301  and  (not A300) );
 a55723a <=( a55722a  and  a55719a );
 a55724a <=( a55723a  and  a55716a );
 a55728a <=( (not A199)  and  (not A167) );
 a55729a <=( (not A168)  and  a55728a );
 a55733a <=( (not A265)  and  (not A202) );
 a55734a <=( (not A200)  and  a55733a );
 a55735a <=( a55734a  and  a55729a );
 a55739a <=( A269  and  (not A268) );
 a55740a <=( A266  and  a55739a );
 a55743a <=( (not A299)  and  A298 );
 a55746a <=( (not A302)  and  (not A300) );
 a55747a <=( a55746a  and  a55743a );
 a55748a <=( a55747a  and  a55740a );
 a55752a <=( (not A199)  and  (not A167) );
 a55753a <=( (not A168)  and  a55752a );
 a55757a <=( (not A265)  and  (not A202) );
 a55758a <=( (not A200)  and  a55757a );
 a55759a <=( a55758a  and  a55753a );
 a55763a <=( A269  and  (not A268) );
 a55764a <=( A266  and  a55763a );
 a55767a <=( A299  and  (not A298) );
 a55770a <=( A301  and  (not A300) );
 a55771a <=( a55770a  and  a55767a );
 a55772a <=( a55771a  and  a55764a );
 a55776a <=( (not A199)  and  (not A167) );
 a55777a <=( (not A168)  and  a55776a );
 a55781a <=( (not A265)  and  (not A202) );
 a55782a <=( (not A200)  and  a55781a );
 a55783a <=( a55782a  and  a55777a );
 a55787a <=( A269  and  (not A268) );
 a55788a <=( A266  and  a55787a );
 a55791a <=( A299  and  (not A298) );
 a55794a <=( (not A302)  and  (not A300) );
 a55795a <=( a55794a  and  a55791a );
 a55796a <=( a55795a  and  a55788a );
 a55800a <=( (not A199)  and  (not A167) );
 a55801a <=( (not A168)  and  a55800a );
 a55805a <=( A265  and  (not A202) );
 a55806a <=( (not A200)  and  a55805a );
 a55807a <=( a55806a  and  a55801a );
 a55811a <=( A269  and  (not A268) );
 a55812a <=( (not A266)  and  a55811a );
 a55815a <=( A299  and  A298 );
 a55818a <=( (not A301)  and  (not A300) );
 a55819a <=( a55818a  and  a55815a );
 a55820a <=( a55819a  and  a55812a );
 a55824a <=( (not A199)  and  (not A167) );
 a55825a <=( (not A168)  and  a55824a );
 a55829a <=( A265  and  (not A202) );
 a55830a <=( (not A200)  and  a55829a );
 a55831a <=( a55830a  and  a55825a );
 a55835a <=( A269  and  (not A268) );
 a55836a <=( (not A266)  and  a55835a );
 a55839a <=( A299  and  A298 );
 a55842a <=( A302  and  (not A300) );
 a55843a <=( a55842a  and  a55839a );
 a55844a <=( a55843a  and  a55836a );
 a55848a <=( (not A199)  and  (not A167) );
 a55849a <=( (not A168)  and  a55848a );
 a55853a <=( A265  and  (not A202) );
 a55854a <=( (not A200)  and  a55853a );
 a55855a <=( a55854a  and  a55849a );
 a55859a <=( A269  and  (not A268) );
 a55860a <=( (not A266)  and  a55859a );
 a55863a <=( (not A299)  and  A298 );
 a55866a <=( A301  and  (not A300) );
 a55867a <=( a55866a  and  a55863a );
 a55868a <=( a55867a  and  a55860a );
 a55872a <=( (not A199)  and  (not A167) );
 a55873a <=( (not A168)  and  a55872a );
 a55877a <=( A265  and  (not A202) );
 a55878a <=( (not A200)  and  a55877a );
 a55879a <=( a55878a  and  a55873a );
 a55883a <=( A269  and  (not A268) );
 a55884a <=( (not A266)  and  a55883a );
 a55887a <=( (not A299)  and  A298 );
 a55890a <=( (not A302)  and  (not A300) );
 a55891a <=( a55890a  and  a55887a );
 a55892a <=( a55891a  and  a55884a );
 a55896a <=( (not A199)  and  (not A167) );
 a55897a <=( (not A168)  and  a55896a );
 a55901a <=( A265  and  (not A202) );
 a55902a <=( (not A200)  and  a55901a );
 a55903a <=( a55902a  and  a55897a );
 a55907a <=( A269  and  (not A268) );
 a55908a <=( (not A266)  and  a55907a );
 a55911a <=( A299  and  (not A298) );
 a55914a <=( A301  and  (not A300) );
 a55915a <=( a55914a  and  a55911a );
 a55916a <=( a55915a  and  a55908a );
 a55920a <=( (not A199)  and  (not A167) );
 a55921a <=( (not A168)  and  a55920a );
 a55925a <=( A265  and  (not A202) );
 a55926a <=( (not A200)  and  a55925a );
 a55927a <=( a55926a  and  a55921a );
 a55931a <=( A269  and  (not A268) );
 a55932a <=( (not A266)  and  a55931a );
 a55935a <=( A299  and  (not A298) );
 a55938a <=( (not A302)  and  (not A300) );
 a55939a <=( a55938a  and  a55935a );
 a55940a <=( a55939a  and  a55932a );
 a55944a <=( (not A199)  and  (not A167) );
 a55945a <=( (not A168)  and  a55944a );
 a55949a <=( (not A265)  and  (not A202) );
 a55950a <=( (not A200)  and  a55949a );
 a55951a <=( a55950a  and  a55945a );
 a55955a <=( (not A269)  and  A268 );
 a55956a <=( (not A266)  and  a55955a );
 a55959a <=( A299  and  A298 );
 a55962a <=( (not A301)  and  (not A300) );
 a55963a <=( a55962a  and  a55959a );
 a55964a <=( a55963a  and  a55956a );
 a55968a <=( (not A199)  and  (not A167) );
 a55969a <=( (not A168)  and  a55968a );
 a55973a <=( (not A265)  and  (not A202) );
 a55974a <=( (not A200)  and  a55973a );
 a55975a <=( a55974a  and  a55969a );
 a55979a <=( (not A269)  and  A268 );
 a55980a <=( (not A266)  and  a55979a );
 a55983a <=( A299  and  A298 );
 a55986a <=( A302  and  (not A300) );
 a55987a <=( a55986a  and  a55983a );
 a55988a <=( a55987a  and  a55980a );
 a55992a <=( (not A199)  and  (not A167) );
 a55993a <=( (not A168)  and  a55992a );
 a55997a <=( (not A265)  and  (not A202) );
 a55998a <=( (not A200)  and  a55997a );
 a55999a <=( a55998a  and  a55993a );
 a56003a <=( (not A269)  and  A268 );
 a56004a <=( (not A266)  and  a56003a );
 a56007a <=( (not A299)  and  A298 );
 a56010a <=( A301  and  (not A300) );
 a56011a <=( a56010a  and  a56007a );
 a56012a <=( a56011a  and  a56004a );
 a56016a <=( (not A199)  and  (not A167) );
 a56017a <=( (not A168)  and  a56016a );
 a56021a <=( (not A265)  and  (not A202) );
 a56022a <=( (not A200)  and  a56021a );
 a56023a <=( a56022a  and  a56017a );
 a56027a <=( (not A269)  and  A268 );
 a56028a <=( (not A266)  and  a56027a );
 a56031a <=( (not A299)  and  A298 );
 a56034a <=( (not A302)  and  (not A300) );
 a56035a <=( a56034a  and  a56031a );
 a56036a <=( a56035a  and  a56028a );
 a56040a <=( (not A199)  and  (not A167) );
 a56041a <=( (not A168)  and  a56040a );
 a56045a <=( (not A265)  and  (not A202) );
 a56046a <=( (not A200)  and  a56045a );
 a56047a <=( a56046a  and  a56041a );
 a56051a <=( (not A269)  and  A268 );
 a56052a <=( (not A266)  and  a56051a );
 a56055a <=( A299  and  (not A298) );
 a56058a <=( A301  and  (not A300) );
 a56059a <=( a56058a  and  a56055a );
 a56060a <=( a56059a  and  a56052a );
 a56064a <=( (not A199)  and  (not A167) );
 a56065a <=( (not A168)  and  a56064a );
 a56069a <=( (not A265)  and  (not A202) );
 a56070a <=( (not A200)  and  a56069a );
 a56071a <=( a56070a  and  a56065a );
 a56075a <=( (not A269)  and  A268 );
 a56076a <=( (not A266)  and  a56075a );
 a56079a <=( A299  and  (not A298) );
 a56082a <=( (not A302)  and  (not A300) );
 a56083a <=( a56082a  and  a56079a );
 a56084a <=( a56083a  and  a56076a );
 a56088a <=( (not A199)  and  (not A167) );
 a56089a <=( (not A168)  and  a56088a );
 a56093a <=( A265  and  A203 );
 a56094a <=( (not A200)  and  a56093a );
 a56095a <=( a56094a  and  a56089a );
 a56099a <=( (not A269)  and  A268 );
 a56100a <=( A266  and  a56099a );
 a56103a <=( A299  and  A298 );
 a56106a <=( (not A301)  and  (not A300) );
 a56107a <=( a56106a  and  a56103a );
 a56108a <=( a56107a  and  a56100a );
 a56112a <=( (not A199)  and  (not A167) );
 a56113a <=( (not A168)  and  a56112a );
 a56117a <=( A265  and  A203 );
 a56118a <=( (not A200)  and  a56117a );
 a56119a <=( a56118a  and  a56113a );
 a56123a <=( (not A269)  and  A268 );
 a56124a <=( A266  and  a56123a );
 a56127a <=( A299  and  A298 );
 a56130a <=( A302  and  (not A300) );
 a56131a <=( a56130a  and  a56127a );
 a56132a <=( a56131a  and  a56124a );
 a56136a <=( (not A199)  and  (not A167) );
 a56137a <=( (not A168)  and  a56136a );
 a56141a <=( A265  and  A203 );
 a56142a <=( (not A200)  and  a56141a );
 a56143a <=( a56142a  and  a56137a );
 a56147a <=( (not A269)  and  A268 );
 a56148a <=( A266  and  a56147a );
 a56151a <=( (not A299)  and  A298 );
 a56154a <=( A301  and  (not A300) );
 a56155a <=( a56154a  and  a56151a );
 a56156a <=( a56155a  and  a56148a );
 a56160a <=( (not A199)  and  (not A167) );
 a56161a <=( (not A168)  and  a56160a );
 a56165a <=( A265  and  A203 );
 a56166a <=( (not A200)  and  a56165a );
 a56167a <=( a56166a  and  a56161a );
 a56171a <=( (not A269)  and  A268 );
 a56172a <=( A266  and  a56171a );
 a56175a <=( (not A299)  and  A298 );
 a56178a <=( (not A302)  and  (not A300) );
 a56179a <=( a56178a  and  a56175a );
 a56180a <=( a56179a  and  a56172a );
 a56184a <=( (not A199)  and  (not A167) );
 a56185a <=( (not A168)  and  a56184a );
 a56189a <=( A265  and  A203 );
 a56190a <=( (not A200)  and  a56189a );
 a56191a <=( a56190a  and  a56185a );
 a56195a <=( (not A269)  and  A268 );
 a56196a <=( A266  and  a56195a );
 a56199a <=( A299  and  (not A298) );
 a56202a <=( A301  and  (not A300) );
 a56203a <=( a56202a  and  a56199a );
 a56204a <=( a56203a  and  a56196a );
 a56208a <=( (not A199)  and  (not A167) );
 a56209a <=( (not A168)  and  a56208a );
 a56213a <=( A265  and  A203 );
 a56214a <=( (not A200)  and  a56213a );
 a56215a <=( a56214a  and  a56209a );
 a56219a <=( (not A269)  and  A268 );
 a56220a <=( A266  and  a56219a );
 a56223a <=( A299  and  (not A298) );
 a56226a <=( (not A302)  and  (not A300) );
 a56227a <=( a56226a  and  a56223a );
 a56228a <=( a56227a  and  a56220a );
 a56232a <=( (not A199)  and  (not A167) );
 a56233a <=( (not A168)  and  a56232a );
 a56237a <=( (not A265)  and  A203 );
 a56238a <=( (not A200)  and  a56237a );
 a56239a <=( a56238a  and  a56233a );
 a56243a <=( A269  and  (not A268) );
 a56244a <=( A266  and  a56243a );
 a56247a <=( A299  and  A298 );
 a56250a <=( (not A301)  and  (not A300) );
 a56251a <=( a56250a  and  a56247a );
 a56252a <=( a56251a  and  a56244a );
 a56256a <=( (not A199)  and  (not A167) );
 a56257a <=( (not A168)  and  a56256a );
 a56261a <=( (not A265)  and  A203 );
 a56262a <=( (not A200)  and  a56261a );
 a56263a <=( a56262a  and  a56257a );
 a56267a <=( A269  and  (not A268) );
 a56268a <=( A266  and  a56267a );
 a56271a <=( A299  and  A298 );
 a56274a <=( A302  and  (not A300) );
 a56275a <=( a56274a  and  a56271a );
 a56276a <=( a56275a  and  a56268a );
 a56280a <=( (not A199)  and  (not A167) );
 a56281a <=( (not A168)  and  a56280a );
 a56285a <=( (not A265)  and  A203 );
 a56286a <=( (not A200)  and  a56285a );
 a56287a <=( a56286a  and  a56281a );
 a56291a <=( A269  and  (not A268) );
 a56292a <=( A266  and  a56291a );
 a56295a <=( (not A299)  and  A298 );
 a56298a <=( A301  and  (not A300) );
 a56299a <=( a56298a  and  a56295a );
 a56300a <=( a56299a  and  a56292a );
 a56304a <=( (not A199)  and  (not A167) );
 a56305a <=( (not A168)  and  a56304a );
 a56309a <=( (not A265)  and  A203 );
 a56310a <=( (not A200)  and  a56309a );
 a56311a <=( a56310a  and  a56305a );
 a56315a <=( A269  and  (not A268) );
 a56316a <=( A266  and  a56315a );
 a56319a <=( (not A299)  and  A298 );
 a56322a <=( (not A302)  and  (not A300) );
 a56323a <=( a56322a  and  a56319a );
 a56324a <=( a56323a  and  a56316a );
 a56328a <=( (not A199)  and  (not A167) );
 a56329a <=( (not A168)  and  a56328a );
 a56333a <=( (not A265)  and  A203 );
 a56334a <=( (not A200)  and  a56333a );
 a56335a <=( a56334a  and  a56329a );
 a56339a <=( A269  and  (not A268) );
 a56340a <=( A266  and  a56339a );
 a56343a <=( A299  and  (not A298) );
 a56346a <=( A301  and  (not A300) );
 a56347a <=( a56346a  and  a56343a );
 a56348a <=( a56347a  and  a56340a );
 a56352a <=( (not A199)  and  (not A167) );
 a56353a <=( (not A168)  and  a56352a );
 a56357a <=( (not A265)  and  A203 );
 a56358a <=( (not A200)  and  a56357a );
 a56359a <=( a56358a  and  a56353a );
 a56363a <=( A269  and  (not A268) );
 a56364a <=( A266  and  a56363a );
 a56367a <=( A299  and  (not A298) );
 a56370a <=( (not A302)  and  (not A300) );
 a56371a <=( a56370a  and  a56367a );
 a56372a <=( a56371a  and  a56364a );
 a56376a <=( (not A199)  and  (not A167) );
 a56377a <=( (not A168)  and  a56376a );
 a56381a <=( A265  and  A203 );
 a56382a <=( (not A200)  and  a56381a );
 a56383a <=( a56382a  and  a56377a );
 a56387a <=( A269  and  (not A268) );
 a56388a <=( (not A266)  and  a56387a );
 a56391a <=( A299  and  A298 );
 a56394a <=( (not A301)  and  (not A300) );
 a56395a <=( a56394a  and  a56391a );
 a56396a <=( a56395a  and  a56388a );
 a56400a <=( (not A199)  and  (not A167) );
 a56401a <=( (not A168)  and  a56400a );
 a56405a <=( A265  and  A203 );
 a56406a <=( (not A200)  and  a56405a );
 a56407a <=( a56406a  and  a56401a );
 a56411a <=( A269  and  (not A268) );
 a56412a <=( (not A266)  and  a56411a );
 a56415a <=( A299  and  A298 );
 a56418a <=( A302  and  (not A300) );
 a56419a <=( a56418a  and  a56415a );
 a56420a <=( a56419a  and  a56412a );
 a56424a <=( (not A199)  and  (not A167) );
 a56425a <=( (not A168)  and  a56424a );
 a56429a <=( A265  and  A203 );
 a56430a <=( (not A200)  and  a56429a );
 a56431a <=( a56430a  and  a56425a );
 a56435a <=( A269  and  (not A268) );
 a56436a <=( (not A266)  and  a56435a );
 a56439a <=( (not A299)  and  A298 );
 a56442a <=( A301  and  (not A300) );
 a56443a <=( a56442a  and  a56439a );
 a56444a <=( a56443a  and  a56436a );
 a56448a <=( (not A199)  and  (not A167) );
 a56449a <=( (not A168)  and  a56448a );
 a56453a <=( A265  and  A203 );
 a56454a <=( (not A200)  and  a56453a );
 a56455a <=( a56454a  and  a56449a );
 a56459a <=( A269  and  (not A268) );
 a56460a <=( (not A266)  and  a56459a );
 a56463a <=( (not A299)  and  A298 );
 a56466a <=( (not A302)  and  (not A300) );
 a56467a <=( a56466a  and  a56463a );
 a56468a <=( a56467a  and  a56460a );
 a56472a <=( (not A199)  and  (not A167) );
 a56473a <=( (not A168)  and  a56472a );
 a56477a <=( A265  and  A203 );
 a56478a <=( (not A200)  and  a56477a );
 a56479a <=( a56478a  and  a56473a );
 a56483a <=( A269  and  (not A268) );
 a56484a <=( (not A266)  and  a56483a );
 a56487a <=( A299  and  (not A298) );
 a56490a <=( A301  and  (not A300) );
 a56491a <=( a56490a  and  a56487a );
 a56492a <=( a56491a  and  a56484a );
 a56496a <=( (not A199)  and  (not A167) );
 a56497a <=( (not A168)  and  a56496a );
 a56501a <=( A265  and  A203 );
 a56502a <=( (not A200)  and  a56501a );
 a56503a <=( a56502a  and  a56497a );
 a56507a <=( A269  and  (not A268) );
 a56508a <=( (not A266)  and  a56507a );
 a56511a <=( A299  and  (not A298) );
 a56514a <=( (not A302)  and  (not A300) );
 a56515a <=( a56514a  and  a56511a );
 a56516a <=( a56515a  and  a56508a );
 a56520a <=( (not A199)  and  (not A167) );
 a56521a <=( (not A168)  and  a56520a );
 a56525a <=( (not A265)  and  A203 );
 a56526a <=( (not A200)  and  a56525a );
 a56527a <=( a56526a  and  a56521a );
 a56531a <=( (not A269)  and  A268 );
 a56532a <=( (not A266)  and  a56531a );
 a56535a <=( A299  and  A298 );
 a56538a <=( (not A301)  and  (not A300) );
 a56539a <=( a56538a  and  a56535a );
 a56540a <=( a56539a  and  a56532a );
 a56544a <=( (not A199)  and  (not A167) );
 a56545a <=( (not A168)  and  a56544a );
 a56549a <=( (not A265)  and  A203 );
 a56550a <=( (not A200)  and  a56549a );
 a56551a <=( a56550a  and  a56545a );
 a56555a <=( (not A269)  and  A268 );
 a56556a <=( (not A266)  and  a56555a );
 a56559a <=( A299  and  A298 );
 a56562a <=( A302  and  (not A300) );
 a56563a <=( a56562a  and  a56559a );
 a56564a <=( a56563a  and  a56556a );
 a56568a <=( (not A199)  and  (not A167) );
 a56569a <=( (not A168)  and  a56568a );
 a56573a <=( (not A265)  and  A203 );
 a56574a <=( (not A200)  and  a56573a );
 a56575a <=( a56574a  and  a56569a );
 a56579a <=( (not A269)  and  A268 );
 a56580a <=( (not A266)  and  a56579a );
 a56583a <=( (not A299)  and  A298 );
 a56586a <=( A301  and  (not A300) );
 a56587a <=( a56586a  and  a56583a );
 a56588a <=( a56587a  and  a56580a );
 a56592a <=( (not A199)  and  (not A167) );
 a56593a <=( (not A168)  and  a56592a );
 a56597a <=( (not A265)  and  A203 );
 a56598a <=( (not A200)  and  a56597a );
 a56599a <=( a56598a  and  a56593a );
 a56603a <=( (not A269)  and  A268 );
 a56604a <=( (not A266)  and  a56603a );
 a56607a <=( (not A299)  and  A298 );
 a56610a <=( (not A302)  and  (not A300) );
 a56611a <=( a56610a  and  a56607a );
 a56612a <=( a56611a  and  a56604a );
 a56616a <=( (not A199)  and  (not A167) );
 a56617a <=( (not A168)  and  a56616a );
 a56621a <=( (not A265)  and  A203 );
 a56622a <=( (not A200)  and  a56621a );
 a56623a <=( a56622a  and  a56617a );
 a56627a <=( (not A269)  and  A268 );
 a56628a <=( (not A266)  and  a56627a );
 a56631a <=( A299  and  (not A298) );
 a56634a <=( A301  and  (not A300) );
 a56635a <=( a56634a  and  a56631a );
 a56636a <=( a56635a  and  a56628a );
 a56640a <=( (not A199)  and  (not A167) );
 a56641a <=( (not A168)  and  a56640a );
 a56645a <=( (not A265)  and  A203 );
 a56646a <=( (not A200)  and  a56645a );
 a56647a <=( a56646a  and  a56641a );
 a56651a <=( (not A269)  and  A268 );
 a56652a <=( (not A266)  and  a56651a );
 a56655a <=( A299  and  (not A298) );
 a56658a <=( (not A302)  and  (not A300) );
 a56659a <=( a56658a  and  a56655a );
 a56660a <=( a56659a  and  a56652a );
 a56664a <=( (not A199)  and  (not A167) );
 a56665a <=( (not A168)  and  a56664a );
 a56669a <=( (not A203)  and  A202 );
 a56670a <=( (not A200)  and  a56669a );
 a56671a <=( a56670a  and  a56665a );
 a56675a <=( (not A268)  and  (not A266) );
 a56676a <=( (not A265)  and  a56675a );
 a56679a <=( A299  and  A298 );
 a56682a <=( (not A302)  and  A301 );
 a56683a <=( a56682a  and  a56679a );
 a56684a <=( a56683a  and  a56676a );
 a56688a <=( (not A199)  and  (not A167) );
 a56689a <=( (not A168)  and  a56688a );
 a56693a <=( (not A203)  and  A202 );
 a56694a <=( (not A200)  and  a56693a );
 a56695a <=( a56694a  and  a56689a );
 a56699a <=( (not A268)  and  (not A266) );
 a56700a <=( (not A265)  and  a56699a );
 a56703a <=( (not A299)  and  A298 );
 a56706a <=( A302  and  (not A301) );
 a56707a <=( a56706a  and  a56703a );
 a56708a <=( a56707a  and  a56700a );
 a56712a <=( (not A199)  and  (not A167) );
 a56713a <=( (not A168)  and  a56712a );
 a56717a <=( (not A203)  and  A202 );
 a56718a <=( (not A200)  and  a56717a );
 a56719a <=( a56718a  and  a56713a );
 a56723a <=( (not A268)  and  (not A266) );
 a56724a <=( (not A265)  and  a56723a );
 a56727a <=( A299  and  (not A298) );
 a56730a <=( A302  and  (not A301) );
 a56731a <=( a56730a  and  a56727a );
 a56732a <=( a56731a  and  a56724a );
 a56736a <=( (not A199)  and  (not A167) );
 a56737a <=( (not A168)  and  a56736a );
 a56741a <=( (not A203)  and  A202 );
 a56742a <=( (not A200)  and  a56741a );
 a56743a <=( a56742a  and  a56737a );
 a56747a <=( (not A268)  and  (not A266) );
 a56748a <=( (not A265)  and  a56747a );
 a56751a <=( (not A299)  and  (not A298) );
 a56754a <=( (not A302)  and  A301 );
 a56755a <=( a56754a  and  a56751a );
 a56756a <=( a56755a  and  a56748a );
 a56760a <=( (not A199)  and  (not A167) );
 a56761a <=( (not A168)  and  a56760a );
 a56765a <=( (not A203)  and  A202 );
 a56766a <=( (not A200)  and  a56765a );
 a56767a <=( a56766a  and  a56761a );
 a56771a <=( A269  and  (not A266) );
 a56772a <=( (not A265)  and  a56771a );
 a56775a <=( A299  and  A298 );
 a56778a <=( (not A302)  and  A301 );
 a56779a <=( a56778a  and  a56775a );
 a56780a <=( a56779a  and  a56772a );
 a56784a <=( (not A199)  and  (not A167) );
 a56785a <=( (not A168)  and  a56784a );
 a56789a <=( (not A203)  and  A202 );
 a56790a <=( (not A200)  and  a56789a );
 a56791a <=( a56790a  and  a56785a );
 a56795a <=( A269  and  (not A266) );
 a56796a <=( (not A265)  and  a56795a );
 a56799a <=( (not A299)  and  A298 );
 a56802a <=( A302  and  (not A301) );
 a56803a <=( a56802a  and  a56799a );
 a56804a <=( a56803a  and  a56796a );
 a56808a <=( (not A199)  and  (not A167) );
 a56809a <=( (not A168)  and  a56808a );
 a56813a <=( (not A203)  and  A202 );
 a56814a <=( (not A200)  and  a56813a );
 a56815a <=( a56814a  and  a56809a );
 a56819a <=( A269  and  (not A266) );
 a56820a <=( (not A265)  and  a56819a );
 a56823a <=( A299  and  (not A298) );
 a56826a <=( A302  and  (not A301) );
 a56827a <=( a56826a  and  a56823a );
 a56828a <=( a56827a  and  a56820a );
 a56832a <=( (not A199)  and  (not A167) );
 a56833a <=( (not A168)  and  a56832a );
 a56837a <=( (not A203)  and  A202 );
 a56838a <=( (not A200)  and  a56837a );
 a56839a <=( a56838a  and  a56833a );
 a56843a <=( A269  and  (not A266) );
 a56844a <=( (not A265)  and  a56843a );
 a56847a <=( (not A299)  and  (not A298) );
 a56850a <=( (not A302)  and  A301 );
 a56851a <=( a56850a  and  a56847a );
 a56852a <=( a56851a  and  a56844a );
 a56856a <=( (not A167)  and  A168 );
 a56857a <=( A170  and  a56856a );
 a56861a <=( A201  and  A199 );
 a56862a <=( A166  and  a56861a );
 a56863a <=( a56862a  and  a56857a );
 a56867a <=( A268  and  A266 );
 a56868a <=( A265  and  a56867a );
 a56871a <=( (not A298)  and  (not A269) );
 a56874a <=( (not A301)  and  (not A299) );
 a56875a <=( a56874a  and  a56871a );
 a56876a <=( a56875a  and  a56868a );
 a56880a <=( (not A167)  and  A168 );
 a56881a <=( A170  and  a56880a );
 a56885a <=( A201  and  A199 );
 a56886a <=( A166  and  a56885a );
 a56887a <=( a56886a  and  a56881a );
 a56891a <=( A268  and  A266 );
 a56892a <=( A265  and  a56891a );
 a56895a <=( (not A298)  and  (not A269) );
 a56898a <=( A302  and  (not A299) );
 a56899a <=( a56898a  and  a56895a );
 a56900a <=( a56899a  and  a56892a );
 a56904a <=( (not A167)  and  A168 );
 a56905a <=( A170  and  a56904a );
 a56909a <=( A201  and  A199 );
 a56910a <=( A166  and  a56909a );
 a56911a <=( a56910a  and  a56905a );
 a56915a <=( (not A268)  and  A266 );
 a56916a <=( (not A265)  and  a56915a );
 a56919a <=( (not A298)  and  A269 );
 a56922a <=( (not A301)  and  (not A299) );
 a56923a <=( a56922a  and  a56919a );
 a56924a <=( a56923a  and  a56916a );
 a56928a <=( (not A167)  and  A168 );
 a56929a <=( A170  and  a56928a );
 a56933a <=( A201  and  A199 );
 a56934a <=( A166  and  a56933a );
 a56935a <=( a56934a  and  a56929a );
 a56939a <=( (not A268)  and  A266 );
 a56940a <=( (not A265)  and  a56939a );
 a56943a <=( (not A298)  and  A269 );
 a56946a <=( A302  and  (not A299) );
 a56947a <=( a56946a  and  a56943a );
 a56948a <=( a56947a  and  a56940a );
 a56952a <=( (not A167)  and  A168 );
 a56953a <=( A170  and  a56952a );
 a56957a <=( A201  and  A199 );
 a56958a <=( A166  and  a56957a );
 a56959a <=( a56958a  and  a56953a );
 a56963a <=( (not A268)  and  (not A266) );
 a56964a <=( A265  and  a56963a );
 a56967a <=( (not A298)  and  A269 );
 a56970a <=( (not A301)  and  (not A299) );
 a56971a <=( a56970a  and  a56967a );
 a56972a <=( a56971a  and  a56964a );
 a56976a <=( (not A167)  and  A168 );
 a56977a <=( A170  and  a56976a );
 a56981a <=( A201  and  A199 );
 a56982a <=( A166  and  a56981a );
 a56983a <=( a56982a  and  a56977a );
 a56987a <=( (not A268)  and  (not A266) );
 a56988a <=( A265  and  a56987a );
 a56991a <=( (not A298)  and  A269 );
 a56994a <=( A302  and  (not A299) );
 a56995a <=( a56994a  and  a56991a );
 a56996a <=( a56995a  and  a56988a );
 a57000a <=( (not A167)  and  A168 );
 a57001a <=( A170  and  a57000a );
 a57005a <=( A201  and  A199 );
 a57006a <=( A166  and  a57005a );
 a57007a <=( a57006a  and  a57001a );
 a57011a <=( A268  and  (not A266) );
 a57012a <=( (not A265)  and  a57011a );
 a57015a <=( (not A298)  and  (not A269) );
 a57018a <=( (not A301)  and  (not A299) );
 a57019a <=( a57018a  and  a57015a );
 a57020a <=( a57019a  and  a57012a );
 a57024a <=( (not A167)  and  A168 );
 a57025a <=( A170  and  a57024a );
 a57029a <=( A201  and  A199 );
 a57030a <=( A166  and  a57029a );
 a57031a <=( a57030a  and  a57025a );
 a57035a <=( A268  and  (not A266) );
 a57036a <=( (not A265)  and  a57035a );
 a57039a <=( (not A298)  and  (not A269) );
 a57042a <=( A302  and  (not A299) );
 a57043a <=( a57042a  and  a57039a );
 a57044a <=( a57043a  and  a57036a );
 a57048a <=( (not A167)  and  A168 );
 a57049a <=( A170  and  a57048a );
 a57053a <=( A201  and  A200 );
 a57054a <=( A166  and  a57053a );
 a57055a <=( a57054a  and  a57049a );
 a57059a <=( A268  and  A266 );
 a57060a <=( A265  and  a57059a );
 a57063a <=( (not A298)  and  (not A269) );
 a57066a <=( (not A301)  and  (not A299) );
 a57067a <=( a57066a  and  a57063a );
 a57068a <=( a57067a  and  a57060a );
 a57072a <=( (not A167)  and  A168 );
 a57073a <=( A170  and  a57072a );
 a57077a <=( A201  and  A200 );
 a57078a <=( A166  and  a57077a );
 a57079a <=( a57078a  and  a57073a );
 a57083a <=( A268  and  A266 );
 a57084a <=( A265  and  a57083a );
 a57087a <=( (not A298)  and  (not A269) );
 a57090a <=( A302  and  (not A299) );
 a57091a <=( a57090a  and  a57087a );
 a57092a <=( a57091a  and  a57084a );
 a57096a <=( (not A167)  and  A168 );
 a57097a <=( A170  and  a57096a );
 a57101a <=( A201  and  A200 );
 a57102a <=( A166  and  a57101a );
 a57103a <=( a57102a  and  a57097a );
 a57107a <=( (not A268)  and  A266 );
 a57108a <=( (not A265)  and  a57107a );
 a57111a <=( (not A298)  and  A269 );
 a57114a <=( (not A301)  and  (not A299) );
 a57115a <=( a57114a  and  a57111a );
 a57116a <=( a57115a  and  a57108a );
 a57120a <=( (not A167)  and  A168 );
 a57121a <=( A170  and  a57120a );
 a57125a <=( A201  and  A200 );
 a57126a <=( A166  and  a57125a );
 a57127a <=( a57126a  and  a57121a );
 a57131a <=( (not A268)  and  A266 );
 a57132a <=( (not A265)  and  a57131a );
 a57135a <=( (not A298)  and  A269 );
 a57138a <=( A302  and  (not A299) );
 a57139a <=( a57138a  and  a57135a );
 a57140a <=( a57139a  and  a57132a );
 a57144a <=( (not A167)  and  A168 );
 a57145a <=( A170  and  a57144a );
 a57149a <=( A201  and  A200 );
 a57150a <=( A166  and  a57149a );
 a57151a <=( a57150a  and  a57145a );
 a57155a <=( (not A268)  and  (not A266) );
 a57156a <=( A265  and  a57155a );
 a57159a <=( (not A298)  and  A269 );
 a57162a <=( (not A301)  and  (not A299) );
 a57163a <=( a57162a  and  a57159a );
 a57164a <=( a57163a  and  a57156a );
 a57168a <=( (not A167)  and  A168 );
 a57169a <=( A170  and  a57168a );
 a57173a <=( A201  and  A200 );
 a57174a <=( A166  and  a57173a );
 a57175a <=( a57174a  and  a57169a );
 a57179a <=( (not A268)  and  (not A266) );
 a57180a <=( A265  and  a57179a );
 a57183a <=( (not A298)  and  A269 );
 a57186a <=( A302  and  (not A299) );
 a57187a <=( a57186a  and  a57183a );
 a57188a <=( a57187a  and  a57180a );
 a57192a <=( (not A167)  and  A168 );
 a57193a <=( A170  and  a57192a );
 a57197a <=( A201  and  A200 );
 a57198a <=( A166  and  a57197a );
 a57199a <=( a57198a  and  a57193a );
 a57203a <=( A268  and  (not A266) );
 a57204a <=( (not A265)  and  a57203a );
 a57207a <=( (not A298)  and  (not A269) );
 a57210a <=( (not A301)  and  (not A299) );
 a57211a <=( a57210a  and  a57207a );
 a57212a <=( a57211a  and  a57204a );
 a57216a <=( (not A167)  and  A168 );
 a57217a <=( A170  and  a57216a );
 a57221a <=( A201  and  A200 );
 a57222a <=( A166  and  a57221a );
 a57223a <=( a57222a  and  a57217a );
 a57227a <=( A268  and  (not A266) );
 a57228a <=( (not A265)  and  a57227a );
 a57231a <=( (not A298)  and  (not A269) );
 a57234a <=( A302  and  (not A299) );
 a57235a <=( a57234a  and  a57231a );
 a57236a <=( a57235a  and  a57228a );
 a57240a <=( (not A167)  and  A168 );
 a57241a <=( A170  and  a57240a );
 a57245a <=( A200  and  A199 );
 a57246a <=( A166  and  a57245a );
 a57247a <=( a57246a  and  a57241a );
 a57251a <=( A265  and  (not A203) );
 a57252a <=( A202  and  a57251a );
 a57255a <=( (not A298)  and  A267 );
 a57258a <=( (not A301)  and  (not A299) );
 a57259a <=( a57258a  and  a57255a );
 a57260a <=( a57259a  and  a57252a );
 a57264a <=( (not A167)  and  A168 );
 a57265a <=( A170  and  a57264a );
 a57269a <=( A200  and  A199 );
 a57270a <=( A166  and  a57269a );
 a57271a <=( a57270a  and  a57265a );
 a57275a <=( A265  and  (not A203) );
 a57276a <=( A202  and  a57275a );
 a57279a <=( (not A298)  and  A267 );
 a57282a <=( A302  and  (not A299) );
 a57283a <=( a57282a  and  a57279a );
 a57284a <=( a57283a  and  a57276a );
 a57288a <=( (not A167)  and  A168 );
 a57289a <=( A170  and  a57288a );
 a57293a <=( A200  and  A199 );
 a57294a <=( A166  and  a57293a );
 a57295a <=( a57294a  and  a57289a );
 a57299a <=( A266  and  (not A203) );
 a57300a <=( A202  and  a57299a );
 a57303a <=( (not A298)  and  A267 );
 a57306a <=( (not A301)  and  (not A299) );
 a57307a <=( a57306a  and  a57303a );
 a57308a <=( a57307a  and  a57300a );
 a57312a <=( (not A167)  and  A168 );
 a57313a <=( A170  and  a57312a );
 a57317a <=( A200  and  A199 );
 a57318a <=( A166  and  a57317a );
 a57319a <=( a57318a  and  a57313a );
 a57323a <=( A266  and  (not A203) );
 a57324a <=( A202  and  a57323a );
 a57327a <=( (not A298)  and  A267 );
 a57330a <=( A302  and  (not A299) );
 a57331a <=( a57330a  and  a57327a );
 a57332a <=( a57331a  and  a57324a );
 a57336a <=( (not A167)  and  A168 );
 a57337a <=( A170  and  a57336a );
 a57341a <=( A200  and  A199 );
 a57342a <=( A166  and  a57341a );
 a57343a <=( a57342a  and  a57337a );
 a57347a <=( (not A265)  and  (not A202) );
 a57348a <=( (not A201)  and  a57347a );
 a57351a <=( (not A268)  and  (not A266) );
 a57354a <=( A300  and  A299 );
 a57355a <=( a57354a  and  a57351a );
 a57356a <=( a57355a  and  a57348a );
 a57360a <=( (not A167)  and  A168 );
 a57361a <=( A170  and  a57360a );
 a57365a <=( A200  and  A199 );
 a57366a <=( A166  and  a57365a );
 a57367a <=( a57366a  and  a57361a );
 a57371a <=( (not A265)  and  (not A202) );
 a57372a <=( (not A201)  and  a57371a );
 a57375a <=( (not A268)  and  (not A266) );
 a57378a <=( A300  and  A298 );
 a57379a <=( a57378a  and  a57375a );
 a57380a <=( a57379a  and  a57372a );
 a57384a <=( (not A167)  and  A168 );
 a57385a <=( A170  and  a57384a );
 a57389a <=( A200  and  A199 );
 a57390a <=( A166  and  a57389a );
 a57391a <=( a57390a  and  a57385a );
 a57395a <=( (not A265)  and  (not A202) );
 a57396a <=( (not A201)  and  a57395a );
 a57399a <=( A269  and  (not A266) );
 a57402a <=( A300  and  A299 );
 a57403a <=( a57402a  and  a57399a );
 a57404a <=( a57403a  and  a57396a );
 a57408a <=( (not A167)  and  A168 );
 a57409a <=( A170  and  a57408a );
 a57413a <=( A200  and  A199 );
 a57414a <=( A166  and  a57413a );
 a57415a <=( a57414a  and  a57409a );
 a57419a <=( (not A265)  and  (not A202) );
 a57420a <=( (not A201)  and  a57419a );
 a57423a <=( A269  and  (not A266) );
 a57426a <=( A300  and  A298 );
 a57427a <=( a57426a  and  a57423a );
 a57428a <=( a57427a  and  a57420a );
 a57432a <=( (not A167)  and  A168 );
 a57433a <=( A170  and  a57432a );
 a57437a <=( A200  and  A199 );
 a57438a <=( A166  and  a57437a );
 a57439a <=( a57438a  and  a57433a );
 a57443a <=( (not A265)  and  A203 );
 a57444a <=( (not A201)  and  a57443a );
 a57447a <=( (not A268)  and  (not A266) );
 a57450a <=( A300  and  A299 );
 a57451a <=( a57450a  and  a57447a );
 a57452a <=( a57451a  and  a57444a );
 a57456a <=( (not A167)  and  A168 );
 a57457a <=( A170  and  a57456a );
 a57461a <=( A200  and  A199 );
 a57462a <=( A166  and  a57461a );
 a57463a <=( a57462a  and  a57457a );
 a57467a <=( (not A265)  and  A203 );
 a57468a <=( (not A201)  and  a57467a );
 a57471a <=( (not A268)  and  (not A266) );
 a57474a <=( A300  and  A298 );
 a57475a <=( a57474a  and  a57471a );
 a57476a <=( a57475a  and  a57468a );
 a57480a <=( (not A167)  and  A168 );
 a57481a <=( A170  and  a57480a );
 a57485a <=( A200  and  A199 );
 a57486a <=( A166  and  a57485a );
 a57487a <=( a57486a  and  a57481a );
 a57491a <=( (not A265)  and  A203 );
 a57492a <=( (not A201)  and  a57491a );
 a57495a <=( A269  and  (not A266) );
 a57498a <=( A300  and  A299 );
 a57499a <=( a57498a  and  a57495a );
 a57500a <=( a57499a  and  a57492a );
 a57504a <=( (not A167)  and  A168 );
 a57505a <=( A170  and  a57504a );
 a57509a <=( A200  and  A199 );
 a57510a <=( A166  and  a57509a );
 a57511a <=( a57510a  and  a57505a );
 a57515a <=( (not A265)  and  A203 );
 a57516a <=( (not A201)  and  a57515a );
 a57519a <=( A269  and  (not A266) );
 a57522a <=( A300  and  A298 );
 a57523a <=( a57522a  and  a57519a );
 a57524a <=( a57523a  and  a57516a );
 a57528a <=( (not A167)  and  A168 );
 a57529a <=( A170  and  a57528a );
 a57533a <=( A200  and  (not A199) );
 a57534a <=( A166  and  a57533a );
 a57535a <=( a57534a  and  a57529a );
 a57539a <=( A265  and  A203 );
 a57540a <=( (not A202)  and  a57539a );
 a57543a <=( (not A298)  and  A267 );
 a57546a <=( (not A301)  and  (not A299) );
 a57547a <=( a57546a  and  a57543a );
 a57548a <=( a57547a  and  a57540a );
 a57552a <=( (not A167)  and  A168 );
 a57553a <=( A170  and  a57552a );
 a57557a <=( A200  and  (not A199) );
 a57558a <=( A166  and  a57557a );
 a57559a <=( a57558a  and  a57553a );
 a57563a <=( A265  and  A203 );
 a57564a <=( (not A202)  and  a57563a );
 a57567a <=( (not A298)  and  A267 );
 a57570a <=( A302  and  (not A299) );
 a57571a <=( a57570a  and  a57567a );
 a57572a <=( a57571a  and  a57564a );
 a57576a <=( (not A167)  and  A168 );
 a57577a <=( A170  and  a57576a );
 a57581a <=( A200  and  (not A199) );
 a57582a <=( A166  and  a57581a );
 a57583a <=( a57582a  and  a57577a );
 a57587a <=( A266  and  A203 );
 a57588a <=( (not A202)  and  a57587a );
 a57591a <=( (not A298)  and  A267 );
 a57594a <=( (not A301)  and  (not A299) );
 a57595a <=( a57594a  and  a57591a );
 a57596a <=( a57595a  and  a57588a );
 a57600a <=( (not A167)  and  A168 );
 a57601a <=( A170  and  a57600a );
 a57605a <=( A200  and  (not A199) );
 a57606a <=( A166  and  a57605a );
 a57607a <=( a57606a  and  a57601a );
 a57611a <=( A266  and  A203 );
 a57612a <=( (not A202)  and  a57611a );
 a57615a <=( (not A298)  and  A267 );
 a57618a <=( A302  and  (not A299) );
 a57619a <=( a57618a  and  a57615a );
 a57620a <=( a57619a  and  a57612a );
 a57624a <=( (not A167)  and  A168 );
 a57625a <=( A170  and  a57624a );
 a57629a <=( A200  and  (not A199) );
 a57630a <=( A166  and  a57629a );
 a57631a <=( a57630a  and  a57625a );
 a57635a <=( (not A265)  and  A202 );
 a57636a <=( (not A201)  and  a57635a );
 a57639a <=( (not A268)  and  (not A266) );
 a57642a <=( A300  and  A299 );
 a57643a <=( a57642a  and  a57639a );
 a57644a <=( a57643a  and  a57636a );
 a57648a <=( (not A167)  and  A168 );
 a57649a <=( A170  and  a57648a );
 a57653a <=( A200  and  (not A199) );
 a57654a <=( A166  and  a57653a );
 a57655a <=( a57654a  and  a57649a );
 a57659a <=( (not A265)  and  A202 );
 a57660a <=( (not A201)  and  a57659a );
 a57663a <=( (not A268)  and  (not A266) );
 a57666a <=( A300  and  A298 );
 a57667a <=( a57666a  and  a57663a );
 a57668a <=( a57667a  and  a57660a );
 a57672a <=( (not A167)  and  A168 );
 a57673a <=( A170  and  a57672a );
 a57677a <=( A200  and  (not A199) );
 a57678a <=( A166  and  a57677a );
 a57679a <=( a57678a  and  a57673a );
 a57683a <=( (not A265)  and  A202 );
 a57684a <=( (not A201)  and  a57683a );
 a57687a <=( A269  and  (not A266) );
 a57690a <=( A300  and  A299 );
 a57691a <=( a57690a  and  a57687a );
 a57692a <=( a57691a  and  a57684a );
 a57696a <=( (not A167)  and  A168 );
 a57697a <=( A170  and  a57696a );
 a57701a <=( A200  and  (not A199) );
 a57702a <=( A166  and  a57701a );
 a57703a <=( a57702a  and  a57697a );
 a57707a <=( (not A265)  and  A202 );
 a57708a <=( (not A201)  and  a57707a );
 a57711a <=( A269  and  (not A266) );
 a57714a <=( A300  and  A298 );
 a57715a <=( a57714a  and  a57711a );
 a57716a <=( a57715a  and  a57708a );
 a57720a <=( (not A167)  and  A168 );
 a57721a <=( A170  and  a57720a );
 a57725a <=( A200  and  (not A199) );
 a57726a <=( A166  and  a57725a );
 a57727a <=( a57726a  and  a57721a );
 a57731a <=( (not A265)  and  (not A203) );
 a57732a <=( (not A201)  and  a57731a );
 a57735a <=( (not A268)  and  (not A266) );
 a57738a <=( A300  and  A299 );
 a57739a <=( a57738a  and  a57735a );
 a57740a <=( a57739a  and  a57732a );
 a57744a <=( (not A167)  and  A168 );
 a57745a <=( A170  and  a57744a );
 a57749a <=( A200  and  (not A199) );
 a57750a <=( A166  and  a57749a );
 a57751a <=( a57750a  and  a57745a );
 a57755a <=( (not A265)  and  (not A203) );
 a57756a <=( (not A201)  and  a57755a );
 a57759a <=( (not A268)  and  (not A266) );
 a57762a <=( A300  and  A298 );
 a57763a <=( a57762a  and  a57759a );
 a57764a <=( a57763a  and  a57756a );
 a57768a <=( (not A167)  and  A168 );
 a57769a <=( A170  and  a57768a );
 a57773a <=( A200  and  (not A199) );
 a57774a <=( A166  and  a57773a );
 a57775a <=( a57774a  and  a57769a );
 a57779a <=( (not A265)  and  (not A203) );
 a57780a <=( (not A201)  and  a57779a );
 a57783a <=( A269  and  (not A266) );
 a57786a <=( A300  and  A299 );
 a57787a <=( a57786a  and  a57783a );
 a57788a <=( a57787a  and  a57780a );
 a57792a <=( (not A167)  and  A168 );
 a57793a <=( A170  and  a57792a );
 a57797a <=( A200  and  (not A199) );
 a57798a <=( A166  and  a57797a );
 a57799a <=( a57798a  and  a57793a );
 a57803a <=( (not A265)  and  (not A203) );
 a57804a <=( (not A201)  and  a57803a );
 a57807a <=( A269  and  (not A266) );
 a57810a <=( A300  and  A298 );
 a57811a <=( a57810a  and  a57807a );
 a57812a <=( a57811a  and  a57804a );
 a57816a <=( (not A167)  and  A168 );
 a57817a <=( A170  and  a57816a );
 a57821a <=( (not A200)  and  A199 );
 a57822a <=( A166  and  a57821a );
 a57823a <=( a57822a  and  a57817a );
 a57827a <=( A265  and  A203 );
 a57828a <=( (not A202)  and  a57827a );
 a57831a <=( (not A298)  and  A267 );
 a57834a <=( (not A301)  and  (not A299) );
 a57835a <=( a57834a  and  a57831a );
 a57836a <=( a57835a  and  a57828a );
 a57840a <=( (not A167)  and  A168 );
 a57841a <=( A170  and  a57840a );
 a57845a <=( (not A200)  and  A199 );
 a57846a <=( A166  and  a57845a );
 a57847a <=( a57846a  and  a57841a );
 a57851a <=( A265  and  A203 );
 a57852a <=( (not A202)  and  a57851a );
 a57855a <=( (not A298)  and  A267 );
 a57858a <=( A302  and  (not A299) );
 a57859a <=( a57858a  and  a57855a );
 a57860a <=( a57859a  and  a57852a );
 a57864a <=( (not A167)  and  A168 );
 a57865a <=( A170  and  a57864a );
 a57869a <=( (not A200)  and  A199 );
 a57870a <=( A166  and  a57869a );
 a57871a <=( a57870a  and  a57865a );
 a57875a <=( A266  and  A203 );
 a57876a <=( (not A202)  and  a57875a );
 a57879a <=( (not A298)  and  A267 );
 a57882a <=( (not A301)  and  (not A299) );
 a57883a <=( a57882a  and  a57879a );
 a57884a <=( a57883a  and  a57876a );
 a57888a <=( (not A167)  and  A168 );
 a57889a <=( A170  and  a57888a );
 a57893a <=( (not A200)  and  A199 );
 a57894a <=( A166  and  a57893a );
 a57895a <=( a57894a  and  a57889a );
 a57899a <=( A266  and  A203 );
 a57900a <=( (not A202)  and  a57899a );
 a57903a <=( (not A298)  and  A267 );
 a57906a <=( A302  and  (not A299) );
 a57907a <=( a57906a  and  a57903a );
 a57908a <=( a57907a  and  a57900a );
 a57912a <=( (not A167)  and  A168 );
 a57913a <=( A170  and  a57912a );
 a57917a <=( (not A200)  and  A199 );
 a57918a <=( A166  and  a57917a );
 a57919a <=( a57918a  and  a57913a );
 a57923a <=( (not A265)  and  A202 );
 a57924a <=( (not A201)  and  a57923a );
 a57927a <=( (not A268)  and  (not A266) );
 a57930a <=( A300  and  A299 );
 a57931a <=( a57930a  and  a57927a );
 a57932a <=( a57931a  and  a57924a );
 a57936a <=( (not A167)  and  A168 );
 a57937a <=( A170  and  a57936a );
 a57941a <=( (not A200)  and  A199 );
 a57942a <=( A166  and  a57941a );
 a57943a <=( a57942a  and  a57937a );
 a57947a <=( (not A265)  and  A202 );
 a57948a <=( (not A201)  and  a57947a );
 a57951a <=( (not A268)  and  (not A266) );
 a57954a <=( A300  and  A298 );
 a57955a <=( a57954a  and  a57951a );
 a57956a <=( a57955a  and  a57948a );
 a57960a <=( (not A167)  and  A168 );
 a57961a <=( A170  and  a57960a );
 a57965a <=( (not A200)  and  A199 );
 a57966a <=( A166  and  a57965a );
 a57967a <=( a57966a  and  a57961a );
 a57971a <=( (not A265)  and  A202 );
 a57972a <=( (not A201)  and  a57971a );
 a57975a <=( A269  and  (not A266) );
 a57978a <=( A300  and  A299 );
 a57979a <=( a57978a  and  a57975a );
 a57980a <=( a57979a  and  a57972a );
 a57984a <=( (not A167)  and  A168 );
 a57985a <=( A170  and  a57984a );
 a57989a <=( (not A200)  and  A199 );
 a57990a <=( A166  and  a57989a );
 a57991a <=( a57990a  and  a57985a );
 a57995a <=( (not A265)  and  A202 );
 a57996a <=( (not A201)  and  a57995a );
 a57999a <=( A269  and  (not A266) );
 a58002a <=( A300  and  A298 );
 a58003a <=( a58002a  and  a57999a );
 a58004a <=( a58003a  and  a57996a );
 a58008a <=( (not A167)  and  A168 );
 a58009a <=( A170  and  a58008a );
 a58013a <=( (not A200)  and  A199 );
 a58014a <=( A166  and  a58013a );
 a58015a <=( a58014a  and  a58009a );
 a58019a <=( (not A265)  and  (not A203) );
 a58020a <=( (not A201)  and  a58019a );
 a58023a <=( (not A268)  and  (not A266) );
 a58026a <=( A300  and  A299 );
 a58027a <=( a58026a  and  a58023a );
 a58028a <=( a58027a  and  a58020a );
 a58032a <=( (not A167)  and  A168 );
 a58033a <=( A170  and  a58032a );
 a58037a <=( (not A200)  and  A199 );
 a58038a <=( A166  and  a58037a );
 a58039a <=( a58038a  and  a58033a );
 a58043a <=( (not A265)  and  (not A203) );
 a58044a <=( (not A201)  and  a58043a );
 a58047a <=( (not A268)  and  (not A266) );
 a58050a <=( A300  and  A298 );
 a58051a <=( a58050a  and  a58047a );
 a58052a <=( a58051a  and  a58044a );
 a58056a <=( (not A167)  and  A168 );
 a58057a <=( A170  and  a58056a );
 a58061a <=( (not A200)  and  A199 );
 a58062a <=( A166  and  a58061a );
 a58063a <=( a58062a  and  a58057a );
 a58067a <=( (not A265)  and  (not A203) );
 a58068a <=( (not A201)  and  a58067a );
 a58071a <=( A269  and  (not A266) );
 a58074a <=( A300  and  A299 );
 a58075a <=( a58074a  and  a58071a );
 a58076a <=( a58075a  and  a58068a );
 a58080a <=( (not A167)  and  A168 );
 a58081a <=( A170  and  a58080a );
 a58085a <=( (not A200)  and  A199 );
 a58086a <=( A166  and  a58085a );
 a58087a <=( a58086a  and  a58081a );
 a58091a <=( (not A265)  and  (not A203) );
 a58092a <=( (not A201)  and  a58091a );
 a58095a <=( A269  and  (not A266) );
 a58098a <=( A300  and  A298 );
 a58099a <=( a58098a  and  a58095a );
 a58100a <=( a58099a  and  a58092a );
 a58104a <=( (not A167)  and  A168 );
 a58105a <=( A170  and  a58104a );
 a58109a <=( (not A200)  and  (not A199) );
 a58110a <=( A166  and  a58109a );
 a58111a <=( a58110a  and  a58105a );
 a58115a <=( A266  and  A265 );
 a58116a <=( (not A202)  and  a58115a );
 a58119a <=( (not A268)  and  (not A267) );
 a58122a <=( A300  and  A299 );
 a58123a <=( a58122a  and  a58119a );
 a58124a <=( a58123a  and  a58116a );
 a58128a <=( (not A167)  and  A168 );
 a58129a <=( A170  and  a58128a );
 a58133a <=( (not A200)  and  (not A199) );
 a58134a <=( A166  and  a58133a );
 a58135a <=( a58134a  and  a58129a );
 a58139a <=( A266  and  A265 );
 a58140a <=( (not A202)  and  a58139a );
 a58143a <=( (not A268)  and  (not A267) );
 a58146a <=( A300  and  A298 );
 a58147a <=( a58146a  and  a58143a );
 a58148a <=( a58147a  and  a58140a );
 a58152a <=( (not A167)  and  A168 );
 a58153a <=( A170  and  a58152a );
 a58157a <=( (not A200)  and  (not A199) );
 a58158a <=( A166  and  a58157a );
 a58159a <=( a58158a  and  a58153a );
 a58163a <=( A266  and  A265 );
 a58164a <=( (not A202)  and  a58163a );
 a58167a <=( A269  and  (not A267) );
 a58170a <=( A300  and  A299 );
 a58171a <=( a58170a  and  a58167a );
 a58172a <=( a58171a  and  a58164a );
 a58176a <=( (not A167)  and  A168 );
 a58177a <=( A170  and  a58176a );
 a58181a <=( (not A200)  and  (not A199) );
 a58182a <=( A166  and  a58181a );
 a58183a <=( a58182a  and  a58177a );
 a58187a <=( A266  and  A265 );
 a58188a <=( (not A202)  and  a58187a );
 a58191a <=( A269  and  (not A267) );
 a58194a <=( A300  and  A298 );
 a58195a <=( a58194a  and  a58191a );
 a58196a <=( a58195a  and  a58188a );
 a58200a <=( (not A167)  and  A168 );
 a58201a <=( A170  and  a58200a );
 a58205a <=( (not A200)  and  (not A199) );
 a58206a <=( A166  and  a58205a );
 a58207a <=( a58206a  and  a58201a );
 a58211a <=( A266  and  (not A265) );
 a58212a <=( (not A202)  and  a58211a );
 a58215a <=( A268  and  (not A267) );
 a58218a <=( A300  and  A299 );
 a58219a <=( a58218a  and  a58215a );
 a58220a <=( a58219a  and  a58212a );
 a58224a <=( (not A167)  and  A168 );
 a58225a <=( A170  and  a58224a );
 a58229a <=( (not A200)  and  (not A199) );
 a58230a <=( A166  and  a58229a );
 a58231a <=( a58230a  and  a58225a );
 a58235a <=( A266  and  (not A265) );
 a58236a <=( (not A202)  and  a58235a );
 a58239a <=( A268  and  (not A267) );
 a58242a <=( A300  and  A298 );
 a58243a <=( a58242a  and  a58239a );
 a58244a <=( a58243a  and  a58236a );
 a58248a <=( (not A167)  and  A168 );
 a58249a <=( A170  and  a58248a );
 a58253a <=( (not A200)  and  (not A199) );
 a58254a <=( A166  and  a58253a );
 a58255a <=( a58254a  and  a58249a );
 a58259a <=( A266  and  (not A265) );
 a58260a <=( (not A202)  and  a58259a );
 a58263a <=( (not A269)  and  (not A267) );
 a58266a <=( A300  and  A299 );
 a58267a <=( a58266a  and  a58263a );
 a58268a <=( a58267a  and  a58260a );
 a58272a <=( (not A167)  and  A168 );
 a58273a <=( A170  and  a58272a );
 a58277a <=( (not A200)  and  (not A199) );
 a58278a <=( A166  and  a58277a );
 a58279a <=( a58278a  and  a58273a );
 a58283a <=( A266  and  (not A265) );
 a58284a <=( (not A202)  and  a58283a );
 a58287a <=( (not A269)  and  (not A267) );
 a58290a <=( A300  and  A298 );
 a58291a <=( a58290a  and  a58287a );
 a58292a <=( a58291a  and  a58284a );
 a58296a <=( (not A167)  and  A168 );
 a58297a <=( A170  and  a58296a );
 a58301a <=( (not A200)  and  (not A199) );
 a58302a <=( A166  and  a58301a );
 a58303a <=( a58302a  and  a58297a );
 a58307a <=( (not A266)  and  A265 );
 a58308a <=( (not A202)  and  a58307a );
 a58311a <=( A268  and  (not A267) );
 a58314a <=( A300  and  A299 );
 a58315a <=( a58314a  and  a58311a );
 a58316a <=( a58315a  and  a58308a );
 a58320a <=( (not A167)  and  A168 );
 a58321a <=( A170  and  a58320a );
 a58325a <=( (not A200)  and  (not A199) );
 a58326a <=( A166  and  a58325a );
 a58327a <=( a58326a  and  a58321a );
 a58331a <=( (not A266)  and  A265 );
 a58332a <=( (not A202)  and  a58331a );
 a58335a <=( A268  and  (not A267) );
 a58338a <=( A300  and  A298 );
 a58339a <=( a58338a  and  a58335a );
 a58340a <=( a58339a  and  a58332a );
 a58344a <=( (not A167)  and  A168 );
 a58345a <=( A170  and  a58344a );
 a58349a <=( (not A200)  and  (not A199) );
 a58350a <=( A166  and  a58349a );
 a58351a <=( a58350a  and  a58345a );
 a58355a <=( (not A266)  and  A265 );
 a58356a <=( (not A202)  and  a58355a );
 a58359a <=( (not A269)  and  (not A267) );
 a58362a <=( A300  and  A299 );
 a58363a <=( a58362a  and  a58359a );
 a58364a <=( a58363a  and  a58356a );
 a58368a <=( (not A167)  and  A168 );
 a58369a <=( A170  and  a58368a );
 a58373a <=( (not A200)  and  (not A199) );
 a58374a <=( A166  and  a58373a );
 a58375a <=( a58374a  and  a58369a );
 a58379a <=( (not A266)  and  A265 );
 a58380a <=( (not A202)  and  a58379a );
 a58383a <=( (not A269)  and  (not A267) );
 a58386a <=( A300  and  A298 );
 a58387a <=( a58386a  and  a58383a );
 a58388a <=( a58387a  and  a58380a );
 a58392a <=( (not A167)  and  A168 );
 a58393a <=( A170  and  a58392a );
 a58397a <=( (not A200)  and  (not A199) );
 a58398a <=( A166  and  a58397a );
 a58399a <=( a58398a  and  a58393a );
 a58403a <=( A266  and  A265 );
 a58404a <=( A203  and  a58403a );
 a58407a <=( (not A268)  and  (not A267) );
 a58410a <=( A300  and  A299 );
 a58411a <=( a58410a  and  a58407a );
 a58412a <=( a58411a  and  a58404a );
 a58416a <=( (not A167)  and  A168 );
 a58417a <=( A170  and  a58416a );
 a58421a <=( (not A200)  and  (not A199) );
 a58422a <=( A166  and  a58421a );
 a58423a <=( a58422a  and  a58417a );
 a58427a <=( A266  and  A265 );
 a58428a <=( A203  and  a58427a );
 a58431a <=( (not A268)  and  (not A267) );
 a58434a <=( A300  and  A298 );
 a58435a <=( a58434a  and  a58431a );
 a58436a <=( a58435a  and  a58428a );
 a58440a <=( (not A167)  and  A168 );
 a58441a <=( A170  and  a58440a );
 a58445a <=( (not A200)  and  (not A199) );
 a58446a <=( A166  and  a58445a );
 a58447a <=( a58446a  and  a58441a );
 a58451a <=( A266  and  A265 );
 a58452a <=( A203  and  a58451a );
 a58455a <=( A269  and  (not A267) );
 a58458a <=( A300  and  A299 );
 a58459a <=( a58458a  and  a58455a );
 a58460a <=( a58459a  and  a58452a );
 a58464a <=( (not A167)  and  A168 );
 a58465a <=( A170  and  a58464a );
 a58469a <=( (not A200)  and  (not A199) );
 a58470a <=( A166  and  a58469a );
 a58471a <=( a58470a  and  a58465a );
 a58475a <=( A266  and  A265 );
 a58476a <=( A203  and  a58475a );
 a58479a <=( A269  and  (not A267) );
 a58482a <=( A300  and  A298 );
 a58483a <=( a58482a  and  a58479a );
 a58484a <=( a58483a  and  a58476a );
 a58488a <=( (not A167)  and  A168 );
 a58489a <=( A170  and  a58488a );
 a58493a <=( (not A200)  and  (not A199) );
 a58494a <=( A166  and  a58493a );
 a58495a <=( a58494a  and  a58489a );
 a58499a <=( A266  and  (not A265) );
 a58500a <=( A203  and  a58499a );
 a58503a <=( A268  and  (not A267) );
 a58506a <=( A300  and  A299 );
 a58507a <=( a58506a  and  a58503a );
 a58508a <=( a58507a  and  a58500a );
 a58512a <=( (not A167)  and  A168 );
 a58513a <=( A170  and  a58512a );
 a58517a <=( (not A200)  and  (not A199) );
 a58518a <=( A166  and  a58517a );
 a58519a <=( a58518a  and  a58513a );
 a58523a <=( A266  and  (not A265) );
 a58524a <=( A203  and  a58523a );
 a58527a <=( A268  and  (not A267) );
 a58530a <=( A300  and  A298 );
 a58531a <=( a58530a  and  a58527a );
 a58532a <=( a58531a  and  a58524a );
 a58536a <=( (not A167)  and  A168 );
 a58537a <=( A170  and  a58536a );
 a58541a <=( (not A200)  and  (not A199) );
 a58542a <=( A166  and  a58541a );
 a58543a <=( a58542a  and  a58537a );
 a58547a <=( A266  and  (not A265) );
 a58548a <=( A203  and  a58547a );
 a58551a <=( (not A269)  and  (not A267) );
 a58554a <=( A300  and  A299 );
 a58555a <=( a58554a  and  a58551a );
 a58556a <=( a58555a  and  a58548a );
 a58560a <=( (not A167)  and  A168 );
 a58561a <=( A170  and  a58560a );
 a58565a <=( (not A200)  and  (not A199) );
 a58566a <=( A166  and  a58565a );
 a58567a <=( a58566a  and  a58561a );
 a58571a <=( A266  and  (not A265) );
 a58572a <=( A203  and  a58571a );
 a58575a <=( (not A269)  and  (not A267) );
 a58578a <=( A300  and  A298 );
 a58579a <=( a58578a  and  a58575a );
 a58580a <=( a58579a  and  a58572a );
 a58584a <=( (not A167)  and  A168 );
 a58585a <=( A170  and  a58584a );
 a58589a <=( (not A200)  and  (not A199) );
 a58590a <=( A166  and  a58589a );
 a58591a <=( a58590a  and  a58585a );
 a58595a <=( (not A266)  and  A265 );
 a58596a <=( A203  and  a58595a );
 a58599a <=( A268  and  (not A267) );
 a58602a <=( A300  and  A299 );
 a58603a <=( a58602a  and  a58599a );
 a58604a <=( a58603a  and  a58596a );
 a58608a <=( (not A167)  and  A168 );
 a58609a <=( A170  and  a58608a );
 a58613a <=( (not A200)  and  (not A199) );
 a58614a <=( A166  and  a58613a );
 a58615a <=( a58614a  and  a58609a );
 a58619a <=( (not A266)  and  A265 );
 a58620a <=( A203  and  a58619a );
 a58623a <=( A268  and  (not A267) );
 a58626a <=( A300  and  A298 );
 a58627a <=( a58626a  and  a58623a );
 a58628a <=( a58627a  and  a58620a );
 a58632a <=( (not A167)  and  A168 );
 a58633a <=( A170  and  a58632a );
 a58637a <=( (not A200)  and  (not A199) );
 a58638a <=( A166  and  a58637a );
 a58639a <=( a58638a  and  a58633a );
 a58643a <=( (not A266)  and  A265 );
 a58644a <=( A203  and  a58643a );
 a58647a <=( (not A269)  and  (not A267) );
 a58650a <=( A300  and  A299 );
 a58651a <=( a58650a  and  a58647a );
 a58652a <=( a58651a  and  a58644a );
 a58656a <=( (not A167)  and  A168 );
 a58657a <=( A170  and  a58656a );
 a58661a <=( (not A200)  and  (not A199) );
 a58662a <=( A166  and  a58661a );
 a58663a <=( a58662a  and  a58657a );
 a58667a <=( (not A266)  and  A265 );
 a58668a <=( A203  and  a58667a );
 a58671a <=( (not A269)  and  (not A267) );
 a58674a <=( A300  and  A298 );
 a58675a <=( a58674a  and  a58671a );
 a58676a <=( a58675a  and  a58668a );
 a58680a <=( (not A167)  and  A168 );
 a58681a <=( A170  and  a58680a );
 a58685a <=( (not A200)  and  (not A199) );
 a58686a <=( A166  and  a58685a );
 a58687a <=( a58686a  and  a58681a );
 a58691a <=( A265  and  (not A203) );
 a58692a <=( A202  and  a58691a );
 a58695a <=( (not A298)  and  A267 );
 a58698a <=( (not A301)  and  (not A299) );
 a58699a <=( a58698a  and  a58695a );
 a58700a <=( a58699a  and  a58692a );
 a58704a <=( (not A167)  and  A168 );
 a58705a <=( A170  and  a58704a );
 a58709a <=( (not A200)  and  (not A199) );
 a58710a <=( A166  and  a58709a );
 a58711a <=( a58710a  and  a58705a );
 a58715a <=( A265  and  (not A203) );
 a58716a <=( A202  and  a58715a );
 a58719a <=( (not A298)  and  A267 );
 a58722a <=( A302  and  (not A299) );
 a58723a <=( a58722a  and  a58719a );
 a58724a <=( a58723a  and  a58716a );
 a58728a <=( (not A167)  and  A168 );
 a58729a <=( A170  and  a58728a );
 a58733a <=( (not A200)  and  (not A199) );
 a58734a <=( A166  and  a58733a );
 a58735a <=( a58734a  and  a58729a );
 a58739a <=( A266  and  (not A203) );
 a58740a <=( A202  and  a58739a );
 a58743a <=( (not A298)  and  A267 );
 a58746a <=( (not A301)  and  (not A299) );
 a58747a <=( a58746a  and  a58743a );
 a58748a <=( a58747a  and  a58740a );
 a58752a <=( (not A167)  and  A168 );
 a58753a <=( A170  and  a58752a );
 a58757a <=( (not A200)  and  (not A199) );
 a58758a <=( A166  and  a58757a );
 a58759a <=( a58758a  and  a58753a );
 a58763a <=( A266  and  (not A203) );
 a58764a <=( A202  and  a58763a );
 a58767a <=( (not A298)  and  A267 );
 a58770a <=( A302  and  (not A299) );
 a58771a <=( a58770a  and  a58767a );
 a58772a <=( a58771a  and  a58764a );
 a58776a <=( (not A167)  and  A168 );
 a58777a <=( A169  and  a58776a );
 a58781a <=( A201  and  A199 );
 a58782a <=( A166  and  a58781a );
 a58783a <=( a58782a  and  a58777a );
 a58787a <=( A268  and  A266 );
 a58788a <=( A265  and  a58787a );
 a58791a <=( (not A298)  and  (not A269) );
 a58794a <=( (not A301)  and  (not A299) );
 a58795a <=( a58794a  and  a58791a );
 a58796a <=( a58795a  and  a58788a );
 a58800a <=( (not A167)  and  A168 );
 a58801a <=( A169  and  a58800a );
 a58805a <=( A201  and  A199 );
 a58806a <=( A166  and  a58805a );
 a58807a <=( a58806a  and  a58801a );
 a58811a <=( A268  and  A266 );
 a58812a <=( A265  and  a58811a );
 a58815a <=( (not A298)  and  (not A269) );
 a58818a <=( A302  and  (not A299) );
 a58819a <=( a58818a  and  a58815a );
 a58820a <=( a58819a  and  a58812a );
 a58824a <=( (not A167)  and  A168 );
 a58825a <=( A169  and  a58824a );
 a58829a <=( A201  and  A199 );
 a58830a <=( A166  and  a58829a );
 a58831a <=( a58830a  and  a58825a );
 a58835a <=( (not A268)  and  A266 );
 a58836a <=( (not A265)  and  a58835a );
 a58839a <=( (not A298)  and  A269 );
 a58842a <=( (not A301)  and  (not A299) );
 a58843a <=( a58842a  and  a58839a );
 a58844a <=( a58843a  and  a58836a );
 a58848a <=( (not A167)  and  A168 );
 a58849a <=( A169  and  a58848a );
 a58853a <=( A201  and  A199 );
 a58854a <=( A166  and  a58853a );
 a58855a <=( a58854a  and  a58849a );
 a58859a <=( (not A268)  and  A266 );
 a58860a <=( (not A265)  and  a58859a );
 a58863a <=( (not A298)  and  A269 );
 a58866a <=( A302  and  (not A299) );
 a58867a <=( a58866a  and  a58863a );
 a58868a <=( a58867a  and  a58860a );
 a58872a <=( (not A167)  and  A168 );
 a58873a <=( A169  and  a58872a );
 a58877a <=( A201  and  A199 );
 a58878a <=( A166  and  a58877a );
 a58879a <=( a58878a  and  a58873a );
 a58883a <=( (not A268)  and  (not A266) );
 a58884a <=( A265  and  a58883a );
 a58887a <=( (not A298)  and  A269 );
 a58890a <=( (not A301)  and  (not A299) );
 a58891a <=( a58890a  and  a58887a );
 a58892a <=( a58891a  and  a58884a );
 a58896a <=( (not A167)  and  A168 );
 a58897a <=( A169  and  a58896a );
 a58901a <=( A201  and  A199 );
 a58902a <=( A166  and  a58901a );
 a58903a <=( a58902a  and  a58897a );
 a58907a <=( (not A268)  and  (not A266) );
 a58908a <=( A265  and  a58907a );
 a58911a <=( (not A298)  and  A269 );
 a58914a <=( A302  and  (not A299) );
 a58915a <=( a58914a  and  a58911a );
 a58916a <=( a58915a  and  a58908a );
 a58920a <=( (not A167)  and  A168 );
 a58921a <=( A169  and  a58920a );
 a58925a <=( A201  and  A199 );
 a58926a <=( A166  and  a58925a );
 a58927a <=( a58926a  and  a58921a );
 a58931a <=( A268  and  (not A266) );
 a58932a <=( (not A265)  and  a58931a );
 a58935a <=( (not A298)  and  (not A269) );
 a58938a <=( (not A301)  and  (not A299) );
 a58939a <=( a58938a  and  a58935a );
 a58940a <=( a58939a  and  a58932a );
 a58944a <=( (not A167)  and  A168 );
 a58945a <=( A169  and  a58944a );
 a58949a <=( A201  and  A199 );
 a58950a <=( A166  and  a58949a );
 a58951a <=( a58950a  and  a58945a );
 a58955a <=( A268  and  (not A266) );
 a58956a <=( (not A265)  and  a58955a );
 a58959a <=( (not A298)  and  (not A269) );
 a58962a <=( A302  and  (not A299) );
 a58963a <=( a58962a  and  a58959a );
 a58964a <=( a58963a  and  a58956a );
 a58968a <=( (not A167)  and  A168 );
 a58969a <=( A169  and  a58968a );
 a58973a <=( A201  and  A200 );
 a58974a <=( A166  and  a58973a );
 a58975a <=( a58974a  and  a58969a );
 a58979a <=( A268  and  A266 );
 a58980a <=( A265  and  a58979a );
 a58983a <=( (not A298)  and  (not A269) );
 a58986a <=( (not A301)  and  (not A299) );
 a58987a <=( a58986a  and  a58983a );
 a58988a <=( a58987a  and  a58980a );
 a58992a <=( (not A167)  and  A168 );
 a58993a <=( A169  and  a58992a );
 a58997a <=( A201  and  A200 );
 a58998a <=( A166  and  a58997a );
 a58999a <=( a58998a  and  a58993a );
 a59003a <=( A268  and  A266 );
 a59004a <=( A265  and  a59003a );
 a59007a <=( (not A298)  and  (not A269) );
 a59010a <=( A302  and  (not A299) );
 a59011a <=( a59010a  and  a59007a );
 a59012a <=( a59011a  and  a59004a );
 a59016a <=( (not A167)  and  A168 );
 a59017a <=( A169  and  a59016a );
 a59021a <=( A201  and  A200 );
 a59022a <=( A166  and  a59021a );
 a59023a <=( a59022a  and  a59017a );
 a59027a <=( (not A268)  and  A266 );
 a59028a <=( (not A265)  and  a59027a );
 a59031a <=( (not A298)  and  A269 );
 a59034a <=( (not A301)  and  (not A299) );
 a59035a <=( a59034a  and  a59031a );
 a59036a <=( a59035a  and  a59028a );
 a59040a <=( (not A167)  and  A168 );
 a59041a <=( A169  and  a59040a );
 a59045a <=( A201  and  A200 );
 a59046a <=( A166  and  a59045a );
 a59047a <=( a59046a  and  a59041a );
 a59051a <=( (not A268)  and  A266 );
 a59052a <=( (not A265)  and  a59051a );
 a59055a <=( (not A298)  and  A269 );
 a59058a <=( A302  and  (not A299) );
 a59059a <=( a59058a  and  a59055a );
 a59060a <=( a59059a  and  a59052a );
 a59064a <=( (not A167)  and  A168 );
 a59065a <=( A169  and  a59064a );
 a59069a <=( A201  and  A200 );
 a59070a <=( A166  and  a59069a );
 a59071a <=( a59070a  and  a59065a );
 a59075a <=( (not A268)  and  (not A266) );
 a59076a <=( A265  and  a59075a );
 a59079a <=( (not A298)  and  A269 );
 a59082a <=( (not A301)  and  (not A299) );
 a59083a <=( a59082a  and  a59079a );
 a59084a <=( a59083a  and  a59076a );
 a59088a <=( (not A167)  and  A168 );
 a59089a <=( A169  and  a59088a );
 a59093a <=( A201  and  A200 );
 a59094a <=( A166  and  a59093a );
 a59095a <=( a59094a  and  a59089a );
 a59099a <=( (not A268)  and  (not A266) );
 a59100a <=( A265  and  a59099a );
 a59103a <=( (not A298)  and  A269 );
 a59106a <=( A302  and  (not A299) );
 a59107a <=( a59106a  and  a59103a );
 a59108a <=( a59107a  and  a59100a );
 a59112a <=( (not A167)  and  A168 );
 a59113a <=( A169  and  a59112a );
 a59117a <=( A201  and  A200 );
 a59118a <=( A166  and  a59117a );
 a59119a <=( a59118a  and  a59113a );
 a59123a <=( A268  and  (not A266) );
 a59124a <=( (not A265)  and  a59123a );
 a59127a <=( (not A298)  and  (not A269) );
 a59130a <=( (not A301)  and  (not A299) );
 a59131a <=( a59130a  and  a59127a );
 a59132a <=( a59131a  and  a59124a );
 a59136a <=( (not A167)  and  A168 );
 a59137a <=( A169  and  a59136a );
 a59141a <=( A201  and  A200 );
 a59142a <=( A166  and  a59141a );
 a59143a <=( a59142a  and  a59137a );
 a59147a <=( A268  and  (not A266) );
 a59148a <=( (not A265)  and  a59147a );
 a59151a <=( (not A298)  and  (not A269) );
 a59154a <=( A302  and  (not A299) );
 a59155a <=( a59154a  and  a59151a );
 a59156a <=( a59155a  and  a59148a );
 a59160a <=( (not A167)  and  A168 );
 a59161a <=( A169  and  a59160a );
 a59165a <=( A200  and  A199 );
 a59166a <=( A166  and  a59165a );
 a59167a <=( a59166a  and  a59161a );
 a59171a <=( A265  and  (not A203) );
 a59172a <=( A202  and  a59171a );
 a59175a <=( (not A298)  and  A267 );
 a59178a <=( (not A301)  and  (not A299) );
 a59179a <=( a59178a  and  a59175a );
 a59180a <=( a59179a  and  a59172a );
 a59184a <=( (not A167)  and  A168 );
 a59185a <=( A169  and  a59184a );
 a59189a <=( A200  and  A199 );
 a59190a <=( A166  and  a59189a );
 a59191a <=( a59190a  and  a59185a );
 a59195a <=( A265  and  (not A203) );
 a59196a <=( A202  and  a59195a );
 a59199a <=( (not A298)  and  A267 );
 a59202a <=( A302  and  (not A299) );
 a59203a <=( a59202a  and  a59199a );
 a59204a <=( a59203a  and  a59196a );
 a59208a <=( (not A167)  and  A168 );
 a59209a <=( A169  and  a59208a );
 a59213a <=( A200  and  A199 );
 a59214a <=( A166  and  a59213a );
 a59215a <=( a59214a  and  a59209a );
 a59219a <=( A266  and  (not A203) );
 a59220a <=( A202  and  a59219a );
 a59223a <=( (not A298)  and  A267 );
 a59226a <=( (not A301)  and  (not A299) );
 a59227a <=( a59226a  and  a59223a );
 a59228a <=( a59227a  and  a59220a );
 a59232a <=( (not A167)  and  A168 );
 a59233a <=( A169  and  a59232a );
 a59237a <=( A200  and  A199 );
 a59238a <=( A166  and  a59237a );
 a59239a <=( a59238a  and  a59233a );
 a59243a <=( A266  and  (not A203) );
 a59244a <=( A202  and  a59243a );
 a59247a <=( (not A298)  and  A267 );
 a59250a <=( A302  and  (not A299) );
 a59251a <=( a59250a  and  a59247a );
 a59252a <=( a59251a  and  a59244a );
 a59256a <=( (not A167)  and  A168 );
 a59257a <=( A169  and  a59256a );
 a59261a <=( A200  and  A199 );
 a59262a <=( A166  and  a59261a );
 a59263a <=( a59262a  and  a59257a );
 a59267a <=( (not A265)  and  (not A202) );
 a59268a <=( (not A201)  and  a59267a );
 a59271a <=( (not A268)  and  (not A266) );
 a59274a <=( A300  and  A299 );
 a59275a <=( a59274a  and  a59271a );
 a59276a <=( a59275a  and  a59268a );
 a59280a <=( (not A167)  and  A168 );
 a59281a <=( A169  and  a59280a );
 a59285a <=( A200  and  A199 );
 a59286a <=( A166  and  a59285a );
 a59287a <=( a59286a  and  a59281a );
 a59291a <=( (not A265)  and  (not A202) );
 a59292a <=( (not A201)  and  a59291a );
 a59295a <=( (not A268)  and  (not A266) );
 a59298a <=( A300  and  A298 );
 a59299a <=( a59298a  and  a59295a );
 a59300a <=( a59299a  and  a59292a );
 a59304a <=( (not A167)  and  A168 );
 a59305a <=( A169  and  a59304a );
 a59309a <=( A200  and  A199 );
 a59310a <=( A166  and  a59309a );
 a59311a <=( a59310a  and  a59305a );
 a59315a <=( (not A265)  and  (not A202) );
 a59316a <=( (not A201)  and  a59315a );
 a59319a <=( A269  and  (not A266) );
 a59322a <=( A300  and  A299 );
 a59323a <=( a59322a  and  a59319a );
 a59324a <=( a59323a  and  a59316a );
 a59328a <=( (not A167)  and  A168 );
 a59329a <=( A169  and  a59328a );
 a59333a <=( A200  and  A199 );
 a59334a <=( A166  and  a59333a );
 a59335a <=( a59334a  and  a59329a );
 a59339a <=( (not A265)  and  (not A202) );
 a59340a <=( (not A201)  and  a59339a );
 a59343a <=( A269  and  (not A266) );
 a59346a <=( A300  and  A298 );
 a59347a <=( a59346a  and  a59343a );
 a59348a <=( a59347a  and  a59340a );
 a59352a <=( (not A167)  and  A168 );
 a59353a <=( A169  and  a59352a );
 a59357a <=( A200  and  A199 );
 a59358a <=( A166  and  a59357a );
 a59359a <=( a59358a  and  a59353a );
 a59363a <=( (not A265)  and  A203 );
 a59364a <=( (not A201)  and  a59363a );
 a59367a <=( (not A268)  and  (not A266) );
 a59370a <=( A300  and  A299 );
 a59371a <=( a59370a  and  a59367a );
 a59372a <=( a59371a  and  a59364a );
 a59376a <=( (not A167)  and  A168 );
 a59377a <=( A169  and  a59376a );
 a59381a <=( A200  and  A199 );
 a59382a <=( A166  and  a59381a );
 a59383a <=( a59382a  and  a59377a );
 a59387a <=( (not A265)  and  A203 );
 a59388a <=( (not A201)  and  a59387a );
 a59391a <=( (not A268)  and  (not A266) );
 a59394a <=( A300  and  A298 );
 a59395a <=( a59394a  and  a59391a );
 a59396a <=( a59395a  and  a59388a );
 a59400a <=( (not A167)  and  A168 );
 a59401a <=( A169  and  a59400a );
 a59405a <=( A200  and  A199 );
 a59406a <=( A166  and  a59405a );
 a59407a <=( a59406a  and  a59401a );
 a59411a <=( (not A265)  and  A203 );
 a59412a <=( (not A201)  and  a59411a );
 a59415a <=( A269  and  (not A266) );
 a59418a <=( A300  and  A299 );
 a59419a <=( a59418a  and  a59415a );
 a59420a <=( a59419a  and  a59412a );
 a59424a <=( (not A167)  and  A168 );
 a59425a <=( A169  and  a59424a );
 a59429a <=( A200  and  A199 );
 a59430a <=( A166  and  a59429a );
 a59431a <=( a59430a  and  a59425a );
 a59435a <=( (not A265)  and  A203 );
 a59436a <=( (not A201)  and  a59435a );
 a59439a <=( A269  and  (not A266) );
 a59442a <=( A300  and  A298 );
 a59443a <=( a59442a  and  a59439a );
 a59444a <=( a59443a  and  a59436a );
 a59448a <=( (not A167)  and  A168 );
 a59449a <=( A169  and  a59448a );
 a59453a <=( A200  and  (not A199) );
 a59454a <=( A166  and  a59453a );
 a59455a <=( a59454a  and  a59449a );
 a59459a <=( A265  and  A203 );
 a59460a <=( (not A202)  and  a59459a );
 a59463a <=( (not A298)  and  A267 );
 a59466a <=( (not A301)  and  (not A299) );
 a59467a <=( a59466a  and  a59463a );
 a59468a <=( a59467a  and  a59460a );
 a59472a <=( (not A167)  and  A168 );
 a59473a <=( A169  and  a59472a );
 a59477a <=( A200  and  (not A199) );
 a59478a <=( A166  and  a59477a );
 a59479a <=( a59478a  and  a59473a );
 a59483a <=( A265  and  A203 );
 a59484a <=( (not A202)  and  a59483a );
 a59487a <=( (not A298)  and  A267 );
 a59490a <=( A302  and  (not A299) );
 a59491a <=( a59490a  and  a59487a );
 a59492a <=( a59491a  and  a59484a );
 a59496a <=( (not A167)  and  A168 );
 a59497a <=( A169  and  a59496a );
 a59501a <=( A200  and  (not A199) );
 a59502a <=( A166  and  a59501a );
 a59503a <=( a59502a  and  a59497a );
 a59507a <=( A266  and  A203 );
 a59508a <=( (not A202)  and  a59507a );
 a59511a <=( (not A298)  and  A267 );
 a59514a <=( (not A301)  and  (not A299) );
 a59515a <=( a59514a  and  a59511a );
 a59516a <=( a59515a  and  a59508a );
 a59520a <=( (not A167)  and  A168 );
 a59521a <=( A169  and  a59520a );
 a59525a <=( A200  and  (not A199) );
 a59526a <=( A166  and  a59525a );
 a59527a <=( a59526a  and  a59521a );
 a59531a <=( A266  and  A203 );
 a59532a <=( (not A202)  and  a59531a );
 a59535a <=( (not A298)  and  A267 );
 a59538a <=( A302  and  (not A299) );
 a59539a <=( a59538a  and  a59535a );
 a59540a <=( a59539a  and  a59532a );
 a59544a <=( (not A167)  and  A168 );
 a59545a <=( A169  and  a59544a );
 a59549a <=( A200  and  (not A199) );
 a59550a <=( A166  and  a59549a );
 a59551a <=( a59550a  and  a59545a );
 a59555a <=( (not A265)  and  A202 );
 a59556a <=( (not A201)  and  a59555a );
 a59559a <=( (not A268)  and  (not A266) );
 a59562a <=( A300  and  A299 );
 a59563a <=( a59562a  and  a59559a );
 a59564a <=( a59563a  and  a59556a );
 a59568a <=( (not A167)  and  A168 );
 a59569a <=( A169  and  a59568a );
 a59573a <=( A200  and  (not A199) );
 a59574a <=( A166  and  a59573a );
 a59575a <=( a59574a  and  a59569a );
 a59579a <=( (not A265)  and  A202 );
 a59580a <=( (not A201)  and  a59579a );
 a59583a <=( (not A268)  and  (not A266) );
 a59586a <=( A300  and  A298 );
 a59587a <=( a59586a  and  a59583a );
 a59588a <=( a59587a  and  a59580a );
 a59592a <=( (not A167)  and  A168 );
 a59593a <=( A169  and  a59592a );
 a59597a <=( A200  and  (not A199) );
 a59598a <=( A166  and  a59597a );
 a59599a <=( a59598a  and  a59593a );
 a59603a <=( (not A265)  and  A202 );
 a59604a <=( (not A201)  and  a59603a );
 a59607a <=( A269  and  (not A266) );
 a59610a <=( A300  and  A299 );
 a59611a <=( a59610a  and  a59607a );
 a59612a <=( a59611a  and  a59604a );
 a59616a <=( (not A167)  and  A168 );
 a59617a <=( A169  and  a59616a );
 a59621a <=( A200  and  (not A199) );
 a59622a <=( A166  and  a59621a );
 a59623a <=( a59622a  and  a59617a );
 a59627a <=( (not A265)  and  A202 );
 a59628a <=( (not A201)  and  a59627a );
 a59631a <=( A269  and  (not A266) );
 a59634a <=( A300  and  A298 );
 a59635a <=( a59634a  and  a59631a );
 a59636a <=( a59635a  and  a59628a );
 a59640a <=( (not A167)  and  A168 );
 a59641a <=( A169  and  a59640a );
 a59645a <=( A200  and  (not A199) );
 a59646a <=( A166  and  a59645a );
 a59647a <=( a59646a  and  a59641a );
 a59651a <=( (not A265)  and  (not A203) );
 a59652a <=( (not A201)  and  a59651a );
 a59655a <=( (not A268)  and  (not A266) );
 a59658a <=( A300  and  A299 );
 a59659a <=( a59658a  and  a59655a );
 a59660a <=( a59659a  and  a59652a );
 a59664a <=( (not A167)  and  A168 );
 a59665a <=( A169  and  a59664a );
 a59669a <=( A200  and  (not A199) );
 a59670a <=( A166  and  a59669a );
 a59671a <=( a59670a  and  a59665a );
 a59675a <=( (not A265)  and  (not A203) );
 a59676a <=( (not A201)  and  a59675a );
 a59679a <=( (not A268)  and  (not A266) );
 a59682a <=( A300  and  A298 );
 a59683a <=( a59682a  and  a59679a );
 a59684a <=( a59683a  and  a59676a );
 a59688a <=( (not A167)  and  A168 );
 a59689a <=( A169  and  a59688a );
 a59693a <=( A200  and  (not A199) );
 a59694a <=( A166  and  a59693a );
 a59695a <=( a59694a  and  a59689a );
 a59699a <=( (not A265)  and  (not A203) );
 a59700a <=( (not A201)  and  a59699a );
 a59703a <=( A269  and  (not A266) );
 a59706a <=( A300  and  A299 );
 a59707a <=( a59706a  and  a59703a );
 a59708a <=( a59707a  and  a59700a );
 a59712a <=( (not A167)  and  A168 );
 a59713a <=( A169  and  a59712a );
 a59717a <=( A200  and  (not A199) );
 a59718a <=( A166  and  a59717a );
 a59719a <=( a59718a  and  a59713a );
 a59723a <=( (not A265)  and  (not A203) );
 a59724a <=( (not A201)  and  a59723a );
 a59727a <=( A269  and  (not A266) );
 a59730a <=( A300  and  A298 );
 a59731a <=( a59730a  and  a59727a );
 a59732a <=( a59731a  and  a59724a );
 a59736a <=( (not A167)  and  A168 );
 a59737a <=( A169  and  a59736a );
 a59741a <=( (not A200)  and  A199 );
 a59742a <=( A166  and  a59741a );
 a59743a <=( a59742a  and  a59737a );
 a59747a <=( A265  and  A203 );
 a59748a <=( (not A202)  and  a59747a );
 a59751a <=( (not A298)  and  A267 );
 a59754a <=( (not A301)  and  (not A299) );
 a59755a <=( a59754a  and  a59751a );
 a59756a <=( a59755a  and  a59748a );
 a59760a <=( (not A167)  and  A168 );
 a59761a <=( A169  and  a59760a );
 a59765a <=( (not A200)  and  A199 );
 a59766a <=( A166  and  a59765a );
 a59767a <=( a59766a  and  a59761a );
 a59771a <=( A265  and  A203 );
 a59772a <=( (not A202)  and  a59771a );
 a59775a <=( (not A298)  and  A267 );
 a59778a <=( A302  and  (not A299) );
 a59779a <=( a59778a  and  a59775a );
 a59780a <=( a59779a  and  a59772a );
 a59784a <=( (not A167)  and  A168 );
 a59785a <=( A169  and  a59784a );
 a59789a <=( (not A200)  and  A199 );
 a59790a <=( A166  and  a59789a );
 a59791a <=( a59790a  and  a59785a );
 a59795a <=( A266  and  A203 );
 a59796a <=( (not A202)  and  a59795a );
 a59799a <=( (not A298)  and  A267 );
 a59802a <=( (not A301)  and  (not A299) );
 a59803a <=( a59802a  and  a59799a );
 a59804a <=( a59803a  and  a59796a );
 a59808a <=( (not A167)  and  A168 );
 a59809a <=( A169  and  a59808a );
 a59813a <=( (not A200)  and  A199 );
 a59814a <=( A166  and  a59813a );
 a59815a <=( a59814a  and  a59809a );
 a59819a <=( A266  and  A203 );
 a59820a <=( (not A202)  and  a59819a );
 a59823a <=( (not A298)  and  A267 );
 a59826a <=( A302  and  (not A299) );
 a59827a <=( a59826a  and  a59823a );
 a59828a <=( a59827a  and  a59820a );
 a59832a <=( (not A167)  and  A168 );
 a59833a <=( A169  and  a59832a );
 a59837a <=( (not A200)  and  A199 );
 a59838a <=( A166  and  a59837a );
 a59839a <=( a59838a  and  a59833a );
 a59843a <=( (not A265)  and  A202 );
 a59844a <=( (not A201)  and  a59843a );
 a59847a <=( (not A268)  and  (not A266) );
 a59850a <=( A300  and  A299 );
 a59851a <=( a59850a  and  a59847a );
 a59852a <=( a59851a  and  a59844a );
 a59856a <=( (not A167)  and  A168 );
 a59857a <=( A169  and  a59856a );
 a59861a <=( (not A200)  and  A199 );
 a59862a <=( A166  and  a59861a );
 a59863a <=( a59862a  and  a59857a );
 a59867a <=( (not A265)  and  A202 );
 a59868a <=( (not A201)  and  a59867a );
 a59871a <=( (not A268)  and  (not A266) );
 a59874a <=( A300  and  A298 );
 a59875a <=( a59874a  and  a59871a );
 a59876a <=( a59875a  and  a59868a );
 a59880a <=( (not A167)  and  A168 );
 a59881a <=( A169  and  a59880a );
 a59885a <=( (not A200)  and  A199 );
 a59886a <=( A166  and  a59885a );
 a59887a <=( a59886a  and  a59881a );
 a59891a <=( (not A265)  and  A202 );
 a59892a <=( (not A201)  and  a59891a );
 a59895a <=( A269  and  (not A266) );
 a59898a <=( A300  and  A299 );
 a59899a <=( a59898a  and  a59895a );
 a59900a <=( a59899a  and  a59892a );
 a59904a <=( (not A167)  and  A168 );
 a59905a <=( A169  and  a59904a );
 a59909a <=( (not A200)  and  A199 );
 a59910a <=( A166  and  a59909a );
 a59911a <=( a59910a  and  a59905a );
 a59915a <=( (not A265)  and  A202 );
 a59916a <=( (not A201)  and  a59915a );
 a59919a <=( A269  and  (not A266) );
 a59922a <=( A300  and  A298 );
 a59923a <=( a59922a  and  a59919a );
 a59924a <=( a59923a  and  a59916a );
 a59928a <=( (not A167)  and  A168 );
 a59929a <=( A169  and  a59928a );
 a59933a <=( (not A200)  and  A199 );
 a59934a <=( A166  and  a59933a );
 a59935a <=( a59934a  and  a59929a );
 a59939a <=( (not A265)  and  (not A203) );
 a59940a <=( (not A201)  and  a59939a );
 a59943a <=( (not A268)  and  (not A266) );
 a59946a <=( A300  and  A299 );
 a59947a <=( a59946a  and  a59943a );
 a59948a <=( a59947a  and  a59940a );
 a59952a <=( (not A167)  and  A168 );
 a59953a <=( A169  and  a59952a );
 a59957a <=( (not A200)  and  A199 );
 a59958a <=( A166  and  a59957a );
 a59959a <=( a59958a  and  a59953a );
 a59963a <=( (not A265)  and  (not A203) );
 a59964a <=( (not A201)  and  a59963a );
 a59967a <=( (not A268)  and  (not A266) );
 a59970a <=( A300  and  A298 );
 a59971a <=( a59970a  and  a59967a );
 a59972a <=( a59971a  and  a59964a );
 a59976a <=( (not A167)  and  A168 );
 a59977a <=( A169  and  a59976a );
 a59981a <=( (not A200)  and  A199 );
 a59982a <=( A166  and  a59981a );
 a59983a <=( a59982a  and  a59977a );
 a59987a <=( (not A265)  and  (not A203) );
 a59988a <=( (not A201)  and  a59987a );
 a59991a <=( A269  and  (not A266) );
 a59994a <=( A300  and  A299 );
 a59995a <=( a59994a  and  a59991a );
 a59996a <=( a59995a  and  a59988a );
 a60000a <=( (not A167)  and  A168 );
 a60001a <=( A169  and  a60000a );
 a60005a <=( (not A200)  and  A199 );
 a60006a <=( A166  and  a60005a );
 a60007a <=( a60006a  and  a60001a );
 a60011a <=( (not A265)  and  (not A203) );
 a60012a <=( (not A201)  and  a60011a );
 a60015a <=( A269  and  (not A266) );
 a60018a <=( A300  and  A298 );
 a60019a <=( a60018a  and  a60015a );
 a60020a <=( a60019a  and  a60012a );
 a60024a <=( (not A167)  and  A168 );
 a60025a <=( A169  and  a60024a );
 a60029a <=( (not A200)  and  (not A199) );
 a60030a <=( A166  and  a60029a );
 a60031a <=( a60030a  and  a60025a );
 a60035a <=( A266  and  A265 );
 a60036a <=( (not A202)  and  a60035a );
 a60039a <=( (not A268)  and  (not A267) );
 a60042a <=( A300  and  A299 );
 a60043a <=( a60042a  and  a60039a );
 a60044a <=( a60043a  and  a60036a );
 a60048a <=( (not A167)  and  A168 );
 a60049a <=( A169  and  a60048a );
 a60053a <=( (not A200)  and  (not A199) );
 a60054a <=( A166  and  a60053a );
 a60055a <=( a60054a  and  a60049a );
 a60059a <=( A266  and  A265 );
 a60060a <=( (not A202)  and  a60059a );
 a60063a <=( (not A268)  and  (not A267) );
 a60066a <=( A300  and  A298 );
 a60067a <=( a60066a  and  a60063a );
 a60068a <=( a60067a  and  a60060a );
 a60072a <=( (not A167)  and  A168 );
 a60073a <=( A169  and  a60072a );
 a60077a <=( (not A200)  and  (not A199) );
 a60078a <=( A166  and  a60077a );
 a60079a <=( a60078a  and  a60073a );
 a60083a <=( A266  and  A265 );
 a60084a <=( (not A202)  and  a60083a );
 a60087a <=( A269  and  (not A267) );
 a60090a <=( A300  and  A299 );
 a60091a <=( a60090a  and  a60087a );
 a60092a <=( a60091a  and  a60084a );
 a60096a <=( (not A167)  and  A168 );
 a60097a <=( A169  and  a60096a );
 a60101a <=( (not A200)  and  (not A199) );
 a60102a <=( A166  and  a60101a );
 a60103a <=( a60102a  and  a60097a );
 a60107a <=( A266  and  A265 );
 a60108a <=( (not A202)  and  a60107a );
 a60111a <=( A269  and  (not A267) );
 a60114a <=( A300  and  A298 );
 a60115a <=( a60114a  and  a60111a );
 a60116a <=( a60115a  and  a60108a );
 a60120a <=( (not A167)  and  A168 );
 a60121a <=( A169  and  a60120a );
 a60125a <=( (not A200)  and  (not A199) );
 a60126a <=( A166  and  a60125a );
 a60127a <=( a60126a  and  a60121a );
 a60131a <=( A266  and  (not A265) );
 a60132a <=( (not A202)  and  a60131a );
 a60135a <=( A268  and  (not A267) );
 a60138a <=( A300  and  A299 );
 a60139a <=( a60138a  and  a60135a );
 a60140a <=( a60139a  and  a60132a );
 a60144a <=( (not A167)  and  A168 );
 a60145a <=( A169  and  a60144a );
 a60149a <=( (not A200)  and  (not A199) );
 a60150a <=( A166  and  a60149a );
 a60151a <=( a60150a  and  a60145a );
 a60155a <=( A266  and  (not A265) );
 a60156a <=( (not A202)  and  a60155a );
 a60159a <=( A268  and  (not A267) );
 a60162a <=( A300  and  A298 );
 a60163a <=( a60162a  and  a60159a );
 a60164a <=( a60163a  and  a60156a );
 a60168a <=( (not A167)  and  A168 );
 a60169a <=( A169  and  a60168a );
 a60173a <=( (not A200)  and  (not A199) );
 a60174a <=( A166  and  a60173a );
 a60175a <=( a60174a  and  a60169a );
 a60179a <=( A266  and  (not A265) );
 a60180a <=( (not A202)  and  a60179a );
 a60183a <=( (not A269)  and  (not A267) );
 a60186a <=( A300  and  A299 );
 a60187a <=( a60186a  and  a60183a );
 a60188a <=( a60187a  and  a60180a );
 a60192a <=( (not A167)  and  A168 );
 a60193a <=( A169  and  a60192a );
 a60197a <=( (not A200)  and  (not A199) );
 a60198a <=( A166  and  a60197a );
 a60199a <=( a60198a  and  a60193a );
 a60203a <=( A266  and  (not A265) );
 a60204a <=( (not A202)  and  a60203a );
 a60207a <=( (not A269)  and  (not A267) );
 a60210a <=( A300  and  A298 );
 a60211a <=( a60210a  and  a60207a );
 a60212a <=( a60211a  and  a60204a );
 a60216a <=( (not A167)  and  A168 );
 a60217a <=( A169  and  a60216a );
 a60221a <=( (not A200)  and  (not A199) );
 a60222a <=( A166  and  a60221a );
 a60223a <=( a60222a  and  a60217a );
 a60227a <=( (not A266)  and  A265 );
 a60228a <=( (not A202)  and  a60227a );
 a60231a <=( A268  and  (not A267) );
 a60234a <=( A300  and  A299 );
 a60235a <=( a60234a  and  a60231a );
 a60236a <=( a60235a  and  a60228a );
 a60240a <=( (not A167)  and  A168 );
 a60241a <=( A169  and  a60240a );
 a60245a <=( (not A200)  and  (not A199) );
 a60246a <=( A166  and  a60245a );
 a60247a <=( a60246a  and  a60241a );
 a60251a <=( (not A266)  and  A265 );
 a60252a <=( (not A202)  and  a60251a );
 a60255a <=( A268  and  (not A267) );
 a60258a <=( A300  and  A298 );
 a60259a <=( a60258a  and  a60255a );
 a60260a <=( a60259a  and  a60252a );
 a60264a <=( (not A167)  and  A168 );
 a60265a <=( A169  and  a60264a );
 a60269a <=( (not A200)  and  (not A199) );
 a60270a <=( A166  and  a60269a );
 a60271a <=( a60270a  and  a60265a );
 a60275a <=( (not A266)  and  A265 );
 a60276a <=( (not A202)  and  a60275a );
 a60279a <=( (not A269)  and  (not A267) );
 a60282a <=( A300  and  A299 );
 a60283a <=( a60282a  and  a60279a );
 a60284a <=( a60283a  and  a60276a );
 a60288a <=( (not A167)  and  A168 );
 a60289a <=( A169  and  a60288a );
 a60293a <=( (not A200)  and  (not A199) );
 a60294a <=( A166  and  a60293a );
 a60295a <=( a60294a  and  a60289a );
 a60299a <=( (not A266)  and  A265 );
 a60300a <=( (not A202)  and  a60299a );
 a60303a <=( (not A269)  and  (not A267) );
 a60306a <=( A300  and  A298 );
 a60307a <=( a60306a  and  a60303a );
 a60308a <=( a60307a  and  a60300a );
 a60312a <=( (not A167)  and  A168 );
 a60313a <=( A169  and  a60312a );
 a60317a <=( (not A200)  and  (not A199) );
 a60318a <=( A166  and  a60317a );
 a60319a <=( a60318a  and  a60313a );
 a60323a <=( A266  and  A265 );
 a60324a <=( A203  and  a60323a );
 a60327a <=( (not A268)  and  (not A267) );
 a60330a <=( A300  and  A299 );
 a60331a <=( a60330a  and  a60327a );
 a60332a <=( a60331a  and  a60324a );
 a60336a <=( (not A167)  and  A168 );
 a60337a <=( A169  and  a60336a );
 a60341a <=( (not A200)  and  (not A199) );
 a60342a <=( A166  and  a60341a );
 a60343a <=( a60342a  and  a60337a );
 a60347a <=( A266  and  A265 );
 a60348a <=( A203  and  a60347a );
 a60351a <=( (not A268)  and  (not A267) );
 a60354a <=( A300  and  A298 );
 a60355a <=( a60354a  and  a60351a );
 a60356a <=( a60355a  and  a60348a );
 a60360a <=( (not A167)  and  A168 );
 a60361a <=( A169  and  a60360a );
 a60365a <=( (not A200)  and  (not A199) );
 a60366a <=( A166  and  a60365a );
 a60367a <=( a60366a  and  a60361a );
 a60371a <=( A266  and  A265 );
 a60372a <=( A203  and  a60371a );
 a60375a <=( A269  and  (not A267) );
 a60378a <=( A300  and  A299 );
 a60379a <=( a60378a  and  a60375a );
 a60380a <=( a60379a  and  a60372a );
 a60384a <=( (not A167)  and  A168 );
 a60385a <=( A169  and  a60384a );
 a60389a <=( (not A200)  and  (not A199) );
 a60390a <=( A166  and  a60389a );
 a60391a <=( a60390a  and  a60385a );
 a60395a <=( A266  and  A265 );
 a60396a <=( A203  and  a60395a );
 a60399a <=( A269  and  (not A267) );
 a60402a <=( A300  and  A298 );
 a60403a <=( a60402a  and  a60399a );
 a60404a <=( a60403a  and  a60396a );
 a60408a <=( (not A167)  and  A168 );
 a60409a <=( A169  and  a60408a );
 a60413a <=( (not A200)  and  (not A199) );
 a60414a <=( A166  and  a60413a );
 a60415a <=( a60414a  and  a60409a );
 a60419a <=( A266  and  (not A265) );
 a60420a <=( A203  and  a60419a );
 a60423a <=( A268  and  (not A267) );
 a60426a <=( A300  and  A299 );
 a60427a <=( a60426a  and  a60423a );
 a60428a <=( a60427a  and  a60420a );
 a60432a <=( (not A167)  and  A168 );
 a60433a <=( A169  and  a60432a );
 a60437a <=( (not A200)  and  (not A199) );
 a60438a <=( A166  and  a60437a );
 a60439a <=( a60438a  and  a60433a );
 a60443a <=( A266  and  (not A265) );
 a60444a <=( A203  and  a60443a );
 a60447a <=( A268  and  (not A267) );
 a60450a <=( A300  and  A298 );
 a60451a <=( a60450a  and  a60447a );
 a60452a <=( a60451a  and  a60444a );
 a60456a <=( (not A167)  and  A168 );
 a60457a <=( A169  and  a60456a );
 a60461a <=( (not A200)  and  (not A199) );
 a60462a <=( A166  and  a60461a );
 a60463a <=( a60462a  and  a60457a );
 a60467a <=( A266  and  (not A265) );
 a60468a <=( A203  and  a60467a );
 a60471a <=( (not A269)  and  (not A267) );
 a60474a <=( A300  and  A299 );
 a60475a <=( a60474a  and  a60471a );
 a60476a <=( a60475a  and  a60468a );
 a60480a <=( (not A167)  and  A168 );
 a60481a <=( A169  and  a60480a );
 a60485a <=( (not A200)  and  (not A199) );
 a60486a <=( A166  and  a60485a );
 a60487a <=( a60486a  and  a60481a );
 a60491a <=( A266  and  (not A265) );
 a60492a <=( A203  and  a60491a );
 a60495a <=( (not A269)  and  (not A267) );
 a60498a <=( A300  and  A298 );
 a60499a <=( a60498a  and  a60495a );
 a60500a <=( a60499a  and  a60492a );
 a60504a <=( (not A167)  and  A168 );
 a60505a <=( A169  and  a60504a );
 a60509a <=( (not A200)  and  (not A199) );
 a60510a <=( A166  and  a60509a );
 a60511a <=( a60510a  and  a60505a );
 a60515a <=( (not A266)  and  A265 );
 a60516a <=( A203  and  a60515a );
 a60519a <=( A268  and  (not A267) );
 a60522a <=( A300  and  A299 );
 a60523a <=( a60522a  and  a60519a );
 a60524a <=( a60523a  and  a60516a );
 a60528a <=( (not A167)  and  A168 );
 a60529a <=( A169  and  a60528a );
 a60533a <=( (not A200)  and  (not A199) );
 a60534a <=( A166  and  a60533a );
 a60535a <=( a60534a  and  a60529a );
 a60539a <=( (not A266)  and  A265 );
 a60540a <=( A203  and  a60539a );
 a60543a <=( A268  and  (not A267) );
 a60546a <=( A300  and  A298 );
 a60547a <=( a60546a  and  a60543a );
 a60548a <=( a60547a  and  a60540a );
 a60552a <=( (not A167)  and  A168 );
 a60553a <=( A169  and  a60552a );
 a60557a <=( (not A200)  and  (not A199) );
 a60558a <=( A166  and  a60557a );
 a60559a <=( a60558a  and  a60553a );
 a60563a <=( (not A266)  and  A265 );
 a60564a <=( A203  and  a60563a );
 a60567a <=( (not A269)  and  (not A267) );
 a60570a <=( A300  and  A299 );
 a60571a <=( a60570a  and  a60567a );
 a60572a <=( a60571a  and  a60564a );
 a60576a <=( (not A167)  and  A168 );
 a60577a <=( A169  and  a60576a );
 a60581a <=( (not A200)  and  (not A199) );
 a60582a <=( A166  and  a60581a );
 a60583a <=( a60582a  and  a60577a );
 a60587a <=( (not A266)  and  A265 );
 a60588a <=( A203  and  a60587a );
 a60591a <=( (not A269)  and  (not A267) );
 a60594a <=( A300  and  A298 );
 a60595a <=( a60594a  and  a60591a );
 a60596a <=( a60595a  and  a60588a );
 a60600a <=( (not A167)  and  A168 );
 a60601a <=( A169  and  a60600a );
 a60605a <=( (not A200)  and  (not A199) );
 a60606a <=( A166  and  a60605a );
 a60607a <=( a60606a  and  a60601a );
 a60611a <=( A265  and  (not A203) );
 a60612a <=( A202  and  a60611a );
 a60615a <=( (not A298)  and  A267 );
 a60618a <=( (not A301)  and  (not A299) );
 a60619a <=( a60618a  and  a60615a );
 a60620a <=( a60619a  and  a60612a );
 a60624a <=( (not A167)  and  A168 );
 a60625a <=( A169  and  a60624a );
 a60629a <=( (not A200)  and  (not A199) );
 a60630a <=( A166  and  a60629a );
 a60631a <=( a60630a  and  a60625a );
 a60635a <=( A265  and  (not A203) );
 a60636a <=( A202  and  a60635a );
 a60639a <=( (not A298)  and  A267 );
 a60642a <=( A302  and  (not A299) );
 a60643a <=( a60642a  and  a60639a );
 a60644a <=( a60643a  and  a60636a );
 a60648a <=( (not A167)  and  A168 );
 a60649a <=( A169  and  a60648a );
 a60653a <=( (not A200)  and  (not A199) );
 a60654a <=( A166  and  a60653a );
 a60655a <=( a60654a  and  a60649a );
 a60659a <=( A266  and  (not A203) );
 a60660a <=( A202  and  a60659a );
 a60663a <=( (not A298)  and  A267 );
 a60666a <=( (not A301)  and  (not A299) );
 a60667a <=( a60666a  and  a60663a );
 a60668a <=( a60667a  and  a60660a );
 a60672a <=( (not A167)  and  A168 );
 a60673a <=( A169  and  a60672a );
 a60677a <=( (not A200)  and  (not A199) );
 a60678a <=( A166  and  a60677a );
 a60679a <=( a60678a  and  a60673a );
 a60683a <=( A266  and  (not A203) );
 a60684a <=( A202  and  a60683a );
 a60687a <=( (not A298)  and  A267 );
 a60690a <=( A302  and  (not A299) );
 a60691a <=( a60690a  and  a60687a );
 a60692a <=( a60691a  and  a60684a );
 a60696a <=( (not A167)  and  (not A169) );
 a60697a <=( (not A170)  and  a60696a );
 a60701a <=( A265  and  A201 );
 a60702a <=( A199  and  a60701a );
 a60703a <=( a60702a  and  a60697a );
 a60707a <=( (not A268)  and  (not A267) );
 a60708a <=( A266  and  a60707a );
 a60711a <=( A299  and  A298 );
 a60714a <=( (not A302)  and  A301 );
 a60715a <=( a60714a  and  a60711a );
 a60716a <=( a60715a  and  a60708a );
 a60720a <=( (not A167)  and  (not A169) );
 a60721a <=( (not A170)  and  a60720a );
 a60725a <=( A265  and  A201 );
 a60726a <=( A199  and  a60725a );
 a60727a <=( a60726a  and  a60721a );
 a60731a <=( (not A268)  and  (not A267) );
 a60732a <=( A266  and  a60731a );
 a60735a <=( (not A299)  and  A298 );
 a60738a <=( A302  and  (not A301) );
 a60739a <=( a60738a  and  a60735a );
 a60740a <=( a60739a  and  a60732a );
 a60744a <=( (not A167)  and  (not A169) );
 a60745a <=( (not A170)  and  a60744a );
 a60749a <=( A265  and  A201 );
 a60750a <=( A199  and  a60749a );
 a60751a <=( a60750a  and  a60745a );
 a60755a <=( (not A268)  and  (not A267) );
 a60756a <=( A266  and  a60755a );
 a60759a <=( A299  and  (not A298) );
 a60762a <=( A302  and  (not A301) );
 a60763a <=( a60762a  and  a60759a );
 a60764a <=( a60763a  and  a60756a );
 a60768a <=( (not A167)  and  (not A169) );
 a60769a <=( (not A170)  and  a60768a );
 a60773a <=( A265  and  A201 );
 a60774a <=( A199  and  a60773a );
 a60775a <=( a60774a  and  a60769a );
 a60779a <=( (not A268)  and  (not A267) );
 a60780a <=( A266  and  a60779a );
 a60783a <=( (not A299)  and  (not A298) );
 a60786a <=( (not A302)  and  A301 );
 a60787a <=( a60786a  and  a60783a );
 a60788a <=( a60787a  and  a60780a );
 a60792a <=( (not A167)  and  (not A169) );
 a60793a <=( (not A170)  and  a60792a );
 a60797a <=( A265  and  A201 );
 a60798a <=( A199  and  a60797a );
 a60799a <=( a60798a  and  a60793a );
 a60803a <=( A269  and  (not A267) );
 a60804a <=( A266  and  a60803a );
 a60807a <=( A299  and  A298 );
 a60810a <=( (not A302)  and  A301 );
 a60811a <=( a60810a  and  a60807a );
 a60812a <=( a60811a  and  a60804a );
 a60816a <=( (not A167)  and  (not A169) );
 a60817a <=( (not A170)  and  a60816a );
 a60821a <=( A265  and  A201 );
 a60822a <=( A199  and  a60821a );
 a60823a <=( a60822a  and  a60817a );
 a60827a <=( A269  and  (not A267) );
 a60828a <=( A266  and  a60827a );
 a60831a <=( (not A299)  and  A298 );
 a60834a <=( A302  and  (not A301) );
 a60835a <=( a60834a  and  a60831a );
 a60836a <=( a60835a  and  a60828a );
 a60840a <=( (not A167)  and  (not A169) );
 a60841a <=( (not A170)  and  a60840a );
 a60845a <=( A265  and  A201 );
 a60846a <=( A199  and  a60845a );
 a60847a <=( a60846a  and  a60841a );
 a60851a <=( A269  and  (not A267) );
 a60852a <=( A266  and  a60851a );
 a60855a <=( A299  and  (not A298) );
 a60858a <=( A302  and  (not A301) );
 a60859a <=( a60858a  and  a60855a );
 a60860a <=( a60859a  and  a60852a );
 a60864a <=( (not A167)  and  (not A169) );
 a60865a <=( (not A170)  and  a60864a );
 a60869a <=( A265  and  A201 );
 a60870a <=( A199  and  a60869a );
 a60871a <=( a60870a  and  a60865a );
 a60875a <=( A269  and  (not A267) );
 a60876a <=( A266  and  a60875a );
 a60879a <=( (not A299)  and  (not A298) );
 a60882a <=( (not A302)  and  A301 );
 a60883a <=( a60882a  and  a60879a );
 a60884a <=( a60883a  and  a60876a );
 a60888a <=( (not A167)  and  (not A169) );
 a60889a <=( (not A170)  and  a60888a );
 a60893a <=( (not A265)  and  A201 );
 a60894a <=( A199  and  a60893a );
 a60895a <=( a60894a  and  a60889a );
 a60899a <=( A268  and  (not A267) );
 a60900a <=( A266  and  a60899a );
 a60903a <=( A299  and  A298 );
 a60906a <=( (not A302)  and  A301 );
 a60907a <=( a60906a  and  a60903a );
 a60908a <=( a60907a  and  a60900a );
 a60912a <=( (not A167)  and  (not A169) );
 a60913a <=( (not A170)  and  a60912a );
 a60917a <=( (not A265)  and  A201 );
 a60918a <=( A199  and  a60917a );
 a60919a <=( a60918a  and  a60913a );
 a60923a <=( A268  and  (not A267) );
 a60924a <=( A266  and  a60923a );
 a60927a <=( (not A299)  and  A298 );
 a60930a <=( A302  and  (not A301) );
 a60931a <=( a60930a  and  a60927a );
 a60932a <=( a60931a  and  a60924a );
 a60936a <=( (not A167)  and  (not A169) );
 a60937a <=( (not A170)  and  a60936a );
 a60941a <=( (not A265)  and  A201 );
 a60942a <=( A199  and  a60941a );
 a60943a <=( a60942a  and  a60937a );
 a60947a <=( A268  and  (not A267) );
 a60948a <=( A266  and  a60947a );
 a60951a <=( A299  and  (not A298) );
 a60954a <=( A302  and  (not A301) );
 a60955a <=( a60954a  and  a60951a );
 a60956a <=( a60955a  and  a60948a );
 a60960a <=( (not A167)  and  (not A169) );
 a60961a <=( (not A170)  and  a60960a );
 a60965a <=( (not A265)  and  A201 );
 a60966a <=( A199  and  a60965a );
 a60967a <=( a60966a  and  a60961a );
 a60971a <=( A268  and  (not A267) );
 a60972a <=( A266  and  a60971a );
 a60975a <=( (not A299)  and  (not A298) );
 a60978a <=( (not A302)  and  A301 );
 a60979a <=( a60978a  and  a60975a );
 a60980a <=( a60979a  and  a60972a );
 a60984a <=( (not A167)  and  (not A169) );
 a60985a <=( (not A170)  and  a60984a );
 a60989a <=( (not A265)  and  A201 );
 a60990a <=( A199  and  a60989a );
 a60991a <=( a60990a  and  a60985a );
 a60995a <=( (not A269)  and  (not A267) );
 a60996a <=( A266  and  a60995a );
 a60999a <=( A299  and  A298 );
 a61002a <=( (not A302)  and  A301 );
 a61003a <=( a61002a  and  a60999a );
 a61004a <=( a61003a  and  a60996a );
 a61008a <=( (not A167)  and  (not A169) );
 a61009a <=( (not A170)  and  a61008a );
 a61013a <=( (not A265)  and  A201 );
 a61014a <=( A199  and  a61013a );
 a61015a <=( a61014a  and  a61009a );
 a61019a <=( (not A269)  and  (not A267) );
 a61020a <=( A266  and  a61019a );
 a61023a <=( (not A299)  and  A298 );
 a61026a <=( A302  and  (not A301) );
 a61027a <=( a61026a  and  a61023a );
 a61028a <=( a61027a  and  a61020a );
 a61032a <=( (not A167)  and  (not A169) );
 a61033a <=( (not A170)  and  a61032a );
 a61037a <=( (not A265)  and  A201 );
 a61038a <=( A199  and  a61037a );
 a61039a <=( a61038a  and  a61033a );
 a61043a <=( (not A269)  and  (not A267) );
 a61044a <=( A266  and  a61043a );
 a61047a <=( A299  and  (not A298) );
 a61050a <=( A302  and  (not A301) );
 a61051a <=( a61050a  and  a61047a );
 a61052a <=( a61051a  and  a61044a );
 a61056a <=( (not A167)  and  (not A169) );
 a61057a <=( (not A170)  and  a61056a );
 a61061a <=( (not A265)  and  A201 );
 a61062a <=( A199  and  a61061a );
 a61063a <=( a61062a  and  a61057a );
 a61067a <=( (not A269)  and  (not A267) );
 a61068a <=( A266  and  a61067a );
 a61071a <=( (not A299)  and  (not A298) );
 a61074a <=( (not A302)  and  A301 );
 a61075a <=( a61074a  and  a61071a );
 a61076a <=( a61075a  and  a61068a );
 a61080a <=( (not A167)  and  (not A169) );
 a61081a <=( (not A170)  and  a61080a );
 a61085a <=( A265  and  A201 );
 a61086a <=( A199  and  a61085a );
 a61087a <=( a61086a  and  a61081a );
 a61091a <=( A268  and  (not A267) );
 a61092a <=( (not A266)  and  a61091a );
 a61095a <=( A299  and  A298 );
 a61098a <=( (not A302)  and  A301 );
 a61099a <=( a61098a  and  a61095a );
 a61100a <=( a61099a  and  a61092a );
 a61104a <=( (not A167)  and  (not A169) );
 a61105a <=( (not A170)  and  a61104a );
 a61109a <=( A265  and  A201 );
 a61110a <=( A199  and  a61109a );
 a61111a <=( a61110a  and  a61105a );
 a61115a <=( A268  and  (not A267) );
 a61116a <=( (not A266)  and  a61115a );
 a61119a <=( (not A299)  and  A298 );
 a61122a <=( A302  and  (not A301) );
 a61123a <=( a61122a  and  a61119a );
 a61124a <=( a61123a  and  a61116a );
 a61128a <=( (not A167)  and  (not A169) );
 a61129a <=( (not A170)  and  a61128a );
 a61133a <=( A265  and  A201 );
 a61134a <=( A199  and  a61133a );
 a61135a <=( a61134a  and  a61129a );
 a61139a <=( A268  and  (not A267) );
 a61140a <=( (not A266)  and  a61139a );
 a61143a <=( A299  and  (not A298) );
 a61146a <=( A302  and  (not A301) );
 a61147a <=( a61146a  and  a61143a );
 a61148a <=( a61147a  and  a61140a );
 a61152a <=( (not A167)  and  (not A169) );
 a61153a <=( (not A170)  and  a61152a );
 a61157a <=( A265  and  A201 );
 a61158a <=( A199  and  a61157a );
 a61159a <=( a61158a  and  a61153a );
 a61163a <=( A268  and  (not A267) );
 a61164a <=( (not A266)  and  a61163a );
 a61167a <=( (not A299)  and  (not A298) );
 a61170a <=( (not A302)  and  A301 );
 a61171a <=( a61170a  and  a61167a );
 a61172a <=( a61171a  and  a61164a );
 a61176a <=( (not A167)  and  (not A169) );
 a61177a <=( (not A170)  and  a61176a );
 a61181a <=( A265  and  A201 );
 a61182a <=( A199  and  a61181a );
 a61183a <=( a61182a  and  a61177a );
 a61187a <=( (not A269)  and  (not A267) );
 a61188a <=( (not A266)  and  a61187a );
 a61191a <=( A299  and  A298 );
 a61194a <=( (not A302)  and  A301 );
 a61195a <=( a61194a  and  a61191a );
 a61196a <=( a61195a  and  a61188a );
 a61200a <=( (not A167)  and  (not A169) );
 a61201a <=( (not A170)  and  a61200a );
 a61205a <=( A265  and  A201 );
 a61206a <=( A199  and  a61205a );
 a61207a <=( a61206a  and  a61201a );
 a61211a <=( (not A269)  and  (not A267) );
 a61212a <=( (not A266)  and  a61211a );
 a61215a <=( (not A299)  and  A298 );
 a61218a <=( A302  and  (not A301) );
 a61219a <=( a61218a  and  a61215a );
 a61220a <=( a61219a  and  a61212a );
 a61224a <=( (not A167)  and  (not A169) );
 a61225a <=( (not A170)  and  a61224a );
 a61229a <=( A265  and  A201 );
 a61230a <=( A199  and  a61229a );
 a61231a <=( a61230a  and  a61225a );
 a61235a <=( (not A269)  and  (not A267) );
 a61236a <=( (not A266)  and  a61235a );
 a61239a <=( A299  and  (not A298) );
 a61242a <=( A302  and  (not A301) );
 a61243a <=( a61242a  and  a61239a );
 a61244a <=( a61243a  and  a61236a );
 a61248a <=( (not A167)  and  (not A169) );
 a61249a <=( (not A170)  and  a61248a );
 a61253a <=( A265  and  A201 );
 a61254a <=( A199  and  a61253a );
 a61255a <=( a61254a  and  a61249a );
 a61259a <=( (not A269)  and  (not A267) );
 a61260a <=( (not A266)  and  a61259a );
 a61263a <=( (not A299)  and  (not A298) );
 a61266a <=( (not A302)  and  A301 );
 a61267a <=( a61266a  and  a61263a );
 a61268a <=( a61267a  and  a61260a );
 a61272a <=( (not A167)  and  (not A169) );
 a61273a <=( (not A170)  and  a61272a );
 a61277a <=( A265  and  A201 );
 a61278a <=( A200  and  a61277a );
 a61279a <=( a61278a  and  a61273a );
 a61283a <=( (not A268)  and  (not A267) );
 a61284a <=( A266  and  a61283a );
 a61287a <=( A299  and  A298 );
 a61290a <=( (not A302)  and  A301 );
 a61291a <=( a61290a  and  a61287a );
 a61292a <=( a61291a  and  a61284a );
 a61296a <=( (not A167)  and  (not A169) );
 a61297a <=( (not A170)  and  a61296a );
 a61301a <=( A265  and  A201 );
 a61302a <=( A200  and  a61301a );
 a61303a <=( a61302a  and  a61297a );
 a61307a <=( (not A268)  and  (not A267) );
 a61308a <=( A266  and  a61307a );
 a61311a <=( (not A299)  and  A298 );
 a61314a <=( A302  and  (not A301) );
 a61315a <=( a61314a  and  a61311a );
 a61316a <=( a61315a  and  a61308a );
 a61320a <=( (not A167)  and  (not A169) );
 a61321a <=( (not A170)  and  a61320a );
 a61325a <=( A265  and  A201 );
 a61326a <=( A200  and  a61325a );
 a61327a <=( a61326a  and  a61321a );
 a61331a <=( (not A268)  and  (not A267) );
 a61332a <=( A266  and  a61331a );
 a61335a <=( A299  and  (not A298) );
 a61338a <=( A302  and  (not A301) );
 a61339a <=( a61338a  and  a61335a );
 a61340a <=( a61339a  and  a61332a );
 a61344a <=( (not A167)  and  (not A169) );
 a61345a <=( (not A170)  and  a61344a );
 a61349a <=( A265  and  A201 );
 a61350a <=( A200  and  a61349a );
 a61351a <=( a61350a  and  a61345a );
 a61355a <=( (not A268)  and  (not A267) );
 a61356a <=( A266  and  a61355a );
 a61359a <=( (not A299)  and  (not A298) );
 a61362a <=( (not A302)  and  A301 );
 a61363a <=( a61362a  and  a61359a );
 a61364a <=( a61363a  and  a61356a );
 a61368a <=( (not A167)  and  (not A169) );
 a61369a <=( (not A170)  and  a61368a );
 a61373a <=( A265  and  A201 );
 a61374a <=( A200  and  a61373a );
 a61375a <=( a61374a  and  a61369a );
 a61379a <=( A269  and  (not A267) );
 a61380a <=( A266  and  a61379a );
 a61383a <=( A299  and  A298 );
 a61386a <=( (not A302)  and  A301 );
 a61387a <=( a61386a  and  a61383a );
 a61388a <=( a61387a  and  a61380a );
 a61392a <=( (not A167)  and  (not A169) );
 a61393a <=( (not A170)  and  a61392a );
 a61397a <=( A265  and  A201 );
 a61398a <=( A200  and  a61397a );
 a61399a <=( a61398a  and  a61393a );
 a61403a <=( A269  and  (not A267) );
 a61404a <=( A266  and  a61403a );
 a61407a <=( (not A299)  and  A298 );
 a61410a <=( A302  and  (not A301) );
 a61411a <=( a61410a  and  a61407a );
 a61412a <=( a61411a  and  a61404a );
 a61416a <=( (not A167)  and  (not A169) );
 a61417a <=( (not A170)  and  a61416a );
 a61421a <=( A265  and  A201 );
 a61422a <=( A200  and  a61421a );
 a61423a <=( a61422a  and  a61417a );
 a61427a <=( A269  and  (not A267) );
 a61428a <=( A266  and  a61427a );
 a61431a <=( A299  and  (not A298) );
 a61434a <=( A302  and  (not A301) );
 a61435a <=( a61434a  and  a61431a );
 a61436a <=( a61435a  and  a61428a );
 a61440a <=( (not A167)  and  (not A169) );
 a61441a <=( (not A170)  and  a61440a );
 a61445a <=( A265  and  A201 );
 a61446a <=( A200  and  a61445a );
 a61447a <=( a61446a  and  a61441a );
 a61451a <=( A269  and  (not A267) );
 a61452a <=( A266  and  a61451a );
 a61455a <=( (not A299)  and  (not A298) );
 a61458a <=( (not A302)  and  A301 );
 a61459a <=( a61458a  and  a61455a );
 a61460a <=( a61459a  and  a61452a );
 a61464a <=( (not A167)  and  (not A169) );
 a61465a <=( (not A170)  and  a61464a );
 a61469a <=( (not A265)  and  A201 );
 a61470a <=( A200  and  a61469a );
 a61471a <=( a61470a  and  a61465a );
 a61475a <=( A268  and  (not A267) );
 a61476a <=( A266  and  a61475a );
 a61479a <=( A299  and  A298 );
 a61482a <=( (not A302)  and  A301 );
 a61483a <=( a61482a  and  a61479a );
 a61484a <=( a61483a  and  a61476a );
 a61488a <=( (not A167)  and  (not A169) );
 a61489a <=( (not A170)  and  a61488a );
 a61493a <=( (not A265)  and  A201 );
 a61494a <=( A200  and  a61493a );
 a61495a <=( a61494a  and  a61489a );
 a61499a <=( A268  and  (not A267) );
 a61500a <=( A266  and  a61499a );
 a61503a <=( (not A299)  and  A298 );
 a61506a <=( A302  and  (not A301) );
 a61507a <=( a61506a  and  a61503a );
 a61508a <=( a61507a  and  a61500a );
 a61512a <=( (not A167)  and  (not A169) );
 a61513a <=( (not A170)  and  a61512a );
 a61517a <=( (not A265)  and  A201 );
 a61518a <=( A200  and  a61517a );
 a61519a <=( a61518a  and  a61513a );
 a61523a <=( A268  and  (not A267) );
 a61524a <=( A266  and  a61523a );
 a61527a <=( A299  and  (not A298) );
 a61530a <=( A302  and  (not A301) );
 a61531a <=( a61530a  and  a61527a );
 a61532a <=( a61531a  and  a61524a );
 a61536a <=( (not A167)  and  (not A169) );
 a61537a <=( (not A170)  and  a61536a );
 a61541a <=( (not A265)  and  A201 );
 a61542a <=( A200  and  a61541a );
 a61543a <=( a61542a  and  a61537a );
 a61547a <=( A268  and  (not A267) );
 a61548a <=( A266  and  a61547a );
 a61551a <=( (not A299)  and  (not A298) );
 a61554a <=( (not A302)  and  A301 );
 a61555a <=( a61554a  and  a61551a );
 a61556a <=( a61555a  and  a61548a );
 a61560a <=( (not A167)  and  (not A169) );
 a61561a <=( (not A170)  and  a61560a );
 a61565a <=( (not A265)  and  A201 );
 a61566a <=( A200  and  a61565a );
 a61567a <=( a61566a  and  a61561a );
 a61571a <=( (not A269)  and  (not A267) );
 a61572a <=( A266  and  a61571a );
 a61575a <=( A299  and  A298 );
 a61578a <=( (not A302)  and  A301 );
 a61579a <=( a61578a  and  a61575a );
 a61580a <=( a61579a  and  a61572a );
 a61584a <=( (not A167)  and  (not A169) );
 a61585a <=( (not A170)  and  a61584a );
 a61589a <=( (not A265)  and  A201 );
 a61590a <=( A200  and  a61589a );
 a61591a <=( a61590a  and  a61585a );
 a61595a <=( (not A269)  and  (not A267) );
 a61596a <=( A266  and  a61595a );
 a61599a <=( (not A299)  and  A298 );
 a61602a <=( A302  and  (not A301) );
 a61603a <=( a61602a  and  a61599a );
 a61604a <=( a61603a  and  a61596a );
 a61608a <=( (not A167)  and  (not A169) );
 a61609a <=( (not A170)  and  a61608a );
 a61613a <=( (not A265)  and  A201 );
 a61614a <=( A200  and  a61613a );
 a61615a <=( a61614a  and  a61609a );
 a61619a <=( (not A269)  and  (not A267) );
 a61620a <=( A266  and  a61619a );
 a61623a <=( A299  and  (not A298) );
 a61626a <=( A302  and  (not A301) );
 a61627a <=( a61626a  and  a61623a );
 a61628a <=( a61627a  and  a61620a );
 a61632a <=( (not A167)  and  (not A169) );
 a61633a <=( (not A170)  and  a61632a );
 a61637a <=( (not A265)  and  A201 );
 a61638a <=( A200  and  a61637a );
 a61639a <=( a61638a  and  a61633a );
 a61643a <=( (not A269)  and  (not A267) );
 a61644a <=( A266  and  a61643a );
 a61647a <=( (not A299)  and  (not A298) );
 a61650a <=( (not A302)  and  A301 );
 a61651a <=( a61650a  and  a61647a );
 a61652a <=( a61651a  and  a61644a );
 a61656a <=( (not A167)  and  (not A169) );
 a61657a <=( (not A170)  and  a61656a );
 a61661a <=( A265  and  A201 );
 a61662a <=( A200  and  a61661a );
 a61663a <=( a61662a  and  a61657a );
 a61667a <=( A268  and  (not A267) );
 a61668a <=( (not A266)  and  a61667a );
 a61671a <=( A299  and  A298 );
 a61674a <=( (not A302)  and  A301 );
 a61675a <=( a61674a  and  a61671a );
 a61676a <=( a61675a  and  a61668a );
 a61680a <=( (not A167)  and  (not A169) );
 a61681a <=( (not A170)  and  a61680a );
 a61685a <=( A265  and  A201 );
 a61686a <=( A200  and  a61685a );
 a61687a <=( a61686a  and  a61681a );
 a61691a <=( A268  and  (not A267) );
 a61692a <=( (not A266)  and  a61691a );
 a61695a <=( (not A299)  and  A298 );
 a61698a <=( A302  and  (not A301) );
 a61699a <=( a61698a  and  a61695a );
 a61700a <=( a61699a  and  a61692a );
 a61704a <=( (not A167)  and  (not A169) );
 a61705a <=( (not A170)  and  a61704a );
 a61709a <=( A265  and  A201 );
 a61710a <=( A200  and  a61709a );
 a61711a <=( a61710a  and  a61705a );
 a61715a <=( A268  and  (not A267) );
 a61716a <=( (not A266)  and  a61715a );
 a61719a <=( A299  and  (not A298) );
 a61722a <=( A302  and  (not A301) );
 a61723a <=( a61722a  and  a61719a );
 a61724a <=( a61723a  and  a61716a );
 a61728a <=( (not A167)  and  (not A169) );
 a61729a <=( (not A170)  and  a61728a );
 a61733a <=( A265  and  A201 );
 a61734a <=( A200  and  a61733a );
 a61735a <=( a61734a  and  a61729a );
 a61739a <=( A268  and  (not A267) );
 a61740a <=( (not A266)  and  a61739a );
 a61743a <=( (not A299)  and  (not A298) );
 a61746a <=( (not A302)  and  A301 );
 a61747a <=( a61746a  and  a61743a );
 a61748a <=( a61747a  and  a61740a );
 a61752a <=( (not A167)  and  (not A169) );
 a61753a <=( (not A170)  and  a61752a );
 a61757a <=( A265  and  A201 );
 a61758a <=( A200  and  a61757a );
 a61759a <=( a61758a  and  a61753a );
 a61763a <=( (not A269)  and  (not A267) );
 a61764a <=( (not A266)  and  a61763a );
 a61767a <=( A299  and  A298 );
 a61770a <=( (not A302)  and  A301 );
 a61771a <=( a61770a  and  a61767a );
 a61772a <=( a61771a  and  a61764a );
 a61776a <=( (not A167)  and  (not A169) );
 a61777a <=( (not A170)  and  a61776a );
 a61781a <=( A265  and  A201 );
 a61782a <=( A200  and  a61781a );
 a61783a <=( a61782a  and  a61777a );
 a61787a <=( (not A269)  and  (not A267) );
 a61788a <=( (not A266)  and  a61787a );
 a61791a <=( (not A299)  and  A298 );
 a61794a <=( A302  and  (not A301) );
 a61795a <=( a61794a  and  a61791a );
 a61796a <=( a61795a  and  a61788a );
 a61800a <=( (not A167)  and  (not A169) );
 a61801a <=( (not A170)  and  a61800a );
 a61805a <=( A265  and  A201 );
 a61806a <=( A200  and  a61805a );
 a61807a <=( a61806a  and  a61801a );
 a61811a <=( (not A269)  and  (not A267) );
 a61812a <=( (not A266)  and  a61811a );
 a61815a <=( A299  and  (not A298) );
 a61818a <=( A302  and  (not A301) );
 a61819a <=( a61818a  and  a61815a );
 a61820a <=( a61819a  and  a61812a );
 a61824a <=( (not A167)  and  (not A169) );
 a61825a <=( (not A170)  and  a61824a );
 a61829a <=( A265  and  A201 );
 a61830a <=( A200  and  a61829a );
 a61831a <=( a61830a  and  a61825a );
 a61835a <=( (not A269)  and  (not A267) );
 a61836a <=( (not A266)  and  a61835a );
 a61839a <=( (not A299)  and  (not A298) );
 a61842a <=( (not A302)  and  A301 );
 a61843a <=( a61842a  and  a61839a );
 a61844a <=( a61843a  and  a61836a );
 a61848a <=( (not A167)  and  (not A169) );
 a61849a <=( (not A170)  and  a61848a );
 a61853a <=( A202  and  A200 );
 a61854a <=( A199  and  a61853a );
 a61855a <=( a61854a  and  a61849a );
 a61859a <=( A266  and  A265 );
 a61860a <=( (not A203)  and  a61859a );
 a61863a <=( (not A268)  and  (not A267) );
 a61866a <=( A300  and  A299 );
 a61867a <=( a61866a  and  a61863a );
 a61868a <=( a61867a  and  a61860a );
 a61872a <=( (not A167)  and  (not A169) );
 a61873a <=( (not A170)  and  a61872a );
 a61877a <=( A202  and  A200 );
 a61878a <=( A199  and  a61877a );
 a61879a <=( a61878a  and  a61873a );
 a61883a <=( A266  and  A265 );
 a61884a <=( (not A203)  and  a61883a );
 a61887a <=( (not A268)  and  (not A267) );
 a61890a <=( A300  and  A298 );
 a61891a <=( a61890a  and  a61887a );
 a61892a <=( a61891a  and  a61884a );
 a61896a <=( (not A167)  and  (not A169) );
 a61897a <=( (not A170)  and  a61896a );
 a61901a <=( A202  and  A200 );
 a61902a <=( A199  and  a61901a );
 a61903a <=( a61902a  and  a61897a );
 a61907a <=( A266  and  A265 );
 a61908a <=( (not A203)  and  a61907a );
 a61911a <=( A269  and  (not A267) );
 a61914a <=( A300  and  A299 );
 a61915a <=( a61914a  and  a61911a );
 a61916a <=( a61915a  and  a61908a );
 a61920a <=( (not A167)  and  (not A169) );
 a61921a <=( (not A170)  and  a61920a );
 a61925a <=( A202  and  A200 );
 a61926a <=( A199  and  a61925a );
 a61927a <=( a61926a  and  a61921a );
 a61931a <=( A266  and  A265 );
 a61932a <=( (not A203)  and  a61931a );
 a61935a <=( A269  and  (not A267) );
 a61938a <=( A300  and  A298 );
 a61939a <=( a61938a  and  a61935a );
 a61940a <=( a61939a  and  a61932a );
 a61944a <=( (not A167)  and  (not A169) );
 a61945a <=( (not A170)  and  a61944a );
 a61949a <=( A202  and  A200 );
 a61950a <=( A199  and  a61949a );
 a61951a <=( a61950a  and  a61945a );
 a61955a <=( A266  and  (not A265) );
 a61956a <=( (not A203)  and  a61955a );
 a61959a <=( A268  and  (not A267) );
 a61962a <=( A300  and  A299 );
 a61963a <=( a61962a  and  a61959a );
 a61964a <=( a61963a  and  a61956a );
 a61968a <=( (not A167)  and  (not A169) );
 a61969a <=( (not A170)  and  a61968a );
 a61973a <=( A202  and  A200 );
 a61974a <=( A199  and  a61973a );
 a61975a <=( a61974a  and  a61969a );
 a61979a <=( A266  and  (not A265) );
 a61980a <=( (not A203)  and  a61979a );
 a61983a <=( A268  and  (not A267) );
 a61986a <=( A300  and  A298 );
 a61987a <=( a61986a  and  a61983a );
 a61988a <=( a61987a  and  a61980a );
 a61992a <=( (not A167)  and  (not A169) );
 a61993a <=( (not A170)  and  a61992a );
 a61997a <=( A202  and  A200 );
 a61998a <=( A199  and  a61997a );
 a61999a <=( a61998a  and  a61993a );
 a62003a <=( A266  and  (not A265) );
 a62004a <=( (not A203)  and  a62003a );
 a62007a <=( (not A269)  and  (not A267) );
 a62010a <=( A300  and  A299 );
 a62011a <=( a62010a  and  a62007a );
 a62012a <=( a62011a  and  a62004a );
 a62016a <=( (not A167)  and  (not A169) );
 a62017a <=( (not A170)  and  a62016a );
 a62021a <=( A202  and  A200 );
 a62022a <=( A199  and  a62021a );
 a62023a <=( a62022a  and  a62017a );
 a62027a <=( A266  and  (not A265) );
 a62028a <=( (not A203)  and  a62027a );
 a62031a <=( (not A269)  and  (not A267) );
 a62034a <=( A300  and  A298 );
 a62035a <=( a62034a  and  a62031a );
 a62036a <=( a62035a  and  a62028a );
 a62040a <=( (not A167)  and  (not A169) );
 a62041a <=( (not A170)  and  a62040a );
 a62045a <=( A202  and  A200 );
 a62046a <=( A199  and  a62045a );
 a62047a <=( a62046a  and  a62041a );
 a62051a <=( (not A266)  and  A265 );
 a62052a <=( (not A203)  and  a62051a );
 a62055a <=( A268  and  (not A267) );
 a62058a <=( A300  and  A299 );
 a62059a <=( a62058a  and  a62055a );
 a62060a <=( a62059a  and  a62052a );
 a62064a <=( (not A167)  and  (not A169) );
 a62065a <=( (not A170)  and  a62064a );
 a62069a <=( A202  and  A200 );
 a62070a <=( A199  and  a62069a );
 a62071a <=( a62070a  and  a62065a );
 a62075a <=( (not A266)  and  A265 );
 a62076a <=( (not A203)  and  a62075a );
 a62079a <=( A268  and  (not A267) );
 a62082a <=( A300  and  A298 );
 a62083a <=( a62082a  and  a62079a );
 a62084a <=( a62083a  and  a62076a );
 a62088a <=( (not A167)  and  (not A169) );
 a62089a <=( (not A170)  and  a62088a );
 a62093a <=( A202  and  A200 );
 a62094a <=( A199  and  a62093a );
 a62095a <=( a62094a  and  a62089a );
 a62099a <=( (not A266)  and  A265 );
 a62100a <=( (not A203)  and  a62099a );
 a62103a <=( (not A269)  and  (not A267) );
 a62106a <=( A300  and  A299 );
 a62107a <=( a62106a  and  a62103a );
 a62108a <=( a62107a  and  a62100a );
 a62112a <=( (not A167)  and  (not A169) );
 a62113a <=( (not A170)  and  a62112a );
 a62117a <=( A202  and  A200 );
 a62118a <=( A199  and  a62117a );
 a62119a <=( a62118a  and  a62113a );
 a62123a <=( (not A266)  and  A265 );
 a62124a <=( (not A203)  and  a62123a );
 a62127a <=( (not A269)  and  (not A267) );
 a62130a <=( A300  and  A298 );
 a62131a <=( a62130a  and  a62127a );
 a62132a <=( a62131a  and  a62124a );
 a62136a <=( (not A167)  and  (not A169) );
 a62137a <=( (not A170)  and  a62136a );
 a62141a <=( (not A201)  and  A200 );
 a62142a <=( A199  and  a62141a );
 a62143a <=( a62142a  and  a62137a );
 a62147a <=( A267  and  A265 );
 a62148a <=( (not A202)  and  a62147a );
 a62151a <=( A299  and  A298 );
 a62154a <=( (not A301)  and  (not A300) );
 a62155a <=( a62154a  and  a62151a );
 a62156a <=( a62155a  and  a62148a );
 a62160a <=( (not A167)  and  (not A169) );
 a62161a <=( (not A170)  and  a62160a );
 a62165a <=( (not A201)  and  A200 );
 a62166a <=( A199  and  a62165a );
 a62167a <=( a62166a  and  a62161a );
 a62171a <=( A267  and  A265 );
 a62172a <=( (not A202)  and  a62171a );
 a62175a <=( A299  and  A298 );
 a62178a <=( A302  and  (not A300) );
 a62179a <=( a62178a  and  a62175a );
 a62180a <=( a62179a  and  a62172a );
 a62184a <=( (not A167)  and  (not A169) );
 a62185a <=( (not A170)  and  a62184a );
 a62189a <=( (not A201)  and  A200 );
 a62190a <=( A199  and  a62189a );
 a62191a <=( a62190a  and  a62185a );
 a62195a <=( A267  and  A265 );
 a62196a <=( (not A202)  and  a62195a );
 a62199a <=( (not A299)  and  A298 );
 a62202a <=( A301  and  (not A300) );
 a62203a <=( a62202a  and  a62199a );
 a62204a <=( a62203a  and  a62196a );
 a62208a <=( (not A167)  and  (not A169) );
 a62209a <=( (not A170)  and  a62208a );
 a62213a <=( (not A201)  and  A200 );
 a62214a <=( A199  and  a62213a );
 a62215a <=( a62214a  and  a62209a );
 a62219a <=( A267  and  A265 );
 a62220a <=( (not A202)  and  a62219a );
 a62223a <=( (not A299)  and  A298 );
 a62226a <=( (not A302)  and  (not A300) );
 a62227a <=( a62226a  and  a62223a );
 a62228a <=( a62227a  and  a62220a );
 a62232a <=( (not A167)  and  (not A169) );
 a62233a <=( (not A170)  and  a62232a );
 a62237a <=( (not A201)  and  A200 );
 a62238a <=( A199  and  a62237a );
 a62239a <=( a62238a  and  a62233a );
 a62243a <=( A267  and  A265 );
 a62244a <=( (not A202)  and  a62243a );
 a62247a <=( A299  and  (not A298) );
 a62250a <=( A301  and  (not A300) );
 a62251a <=( a62250a  and  a62247a );
 a62252a <=( a62251a  and  a62244a );
 a62256a <=( (not A167)  and  (not A169) );
 a62257a <=( (not A170)  and  a62256a );
 a62261a <=( (not A201)  and  A200 );
 a62262a <=( A199  and  a62261a );
 a62263a <=( a62262a  and  a62257a );
 a62267a <=( A267  and  A265 );
 a62268a <=( (not A202)  and  a62267a );
 a62271a <=( A299  and  (not A298) );
 a62274a <=( (not A302)  and  (not A300) );
 a62275a <=( a62274a  and  a62271a );
 a62276a <=( a62275a  and  a62268a );
 a62280a <=( (not A167)  and  (not A169) );
 a62281a <=( (not A170)  and  a62280a );
 a62285a <=( (not A201)  and  A200 );
 a62286a <=( A199  and  a62285a );
 a62287a <=( a62286a  and  a62281a );
 a62291a <=( A267  and  A266 );
 a62292a <=( (not A202)  and  a62291a );
 a62295a <=( A299  and  A298 );
 a62298a <=( (not A301)  and  (not A300) );
 a62299a <=( a62298a  and  a62295a );
 a62300a <=( a62299a  and  a62292a );
 a62304a <=( (not A167)  and  (not A169) );
 a62305a <=( (not A170)  and  a62304a );
 a62309a <=( (not A201)  and  A200 );
 a62310a <=( A199  and  a62309a );
 a62311a <=( a62310a  and  a62305a );
 a62315a <=( A267  and  A266 );
 a62316a <=( (not A202)  and  a62315a );
 a62319a <=( A299  and  A298 );
 a62322a <=( A302  and  (not A300) );
 a62323a <=( a62322a  and  a62319a );
 a62324a <=( a62323a  and  a62316a );
 a62328a <=( (not A167)  and  (not A169) );
 a62329a <=( (not A170)  and  a62328a );
 a62333a <=( (not A201)  and  A200 );
 a62334a <=( A199  and  a62333a );
 a62335a <=( a62334a  and  a62329a );
 a62339a <=( A267  and  A266 );
 a62340a <=( (not A202)  and  a62339a );
 a62343a <=( (not A299)  and  A298 );
 a62346a <=( A301  and  (not A300) );
 a62347a <=( a62346a  and  a62343a );
 a62348a <=( a62347a  and  a62340a );
 a62352a <=( (not A167)  and  (not A169) );
 a62353a <=( (not A170)  and  a62352a );
 a62357a <=( (not A201)  and  A200 );
 a62358a <=( A199  and  a62357a );
 a62359a <=( a62358a  and  a62353a );
 a62363a <=( A267  and  A266 );
 a62364a <=( (not A202)  and  a62363a );
 a62367a <=( (not A299)  and  A298 );
 a62370a <=( (not A302)  and  (not A300) );
 a62371a <=( a62370a  and  a62367a );
 a62372a <=( a62371a  and  a62364a );
 a62376a <=( (not A167)  and  (not A169) );
 a62377a <=( (not A170)  and  a62376a );
 a62381a <=( (not A201)  and  A200 );
 a62382a <=( A199  and  a62381a );
 a62383a <=( a62382a  and  a62377a );
 a62387a <=( A267  and  A266 );
 a62388a <=( (not A202)  and  a62387a );
 a62391a <=( A299  and  (not A298) );
 a62394a <=( A301  and  (not A300) );
 a62395a <=( a62394a  and  a62391a );
 a62396a <=( a62395a  and  a62388a );
 a62400a <=( (not A167)  and  (not A169) );
 a62401a <=( (not A170)  and  a62400a );
 a62405a <=( (not A201)  and  A200 );
 a62406a <=( A199  and  a62405a );
 a62407a <=( a62406a  and  a62401a );
 a62411a <=( A267  and  A266 );
 a62412a <=( (not A202)  and  a62411a );
 a62415a <=( A299  and  (not A298) );
 a62418a <=( (not A302)  and  (not A300) );
 a62419a <=( a62418a  and  a62415a );
 a62420a <=( a62419a  and  a62412a );
 a62424a <=( (not A167)  and  (not A169) );
 a62425a <=( (not A170)  and  a62424a );
 a62429a <=( (not A201)  and  A200 );
 a62430a <=( A199  and  a62429a );
 a62431a <=( a62430a  and  a62425a );
 a62435a <=( A267  and  A265 );
 a62436a <=( A203  and  a62435a );
 a62439a <=( A299  and  A298 );
 a62442a <=( (not A301)  and  (not A300) );
 a62443a <=( a62442a  and  a62439a );
 a62444a <=( a62443a  and  a62436a );
 a62448a <=( (not A167)  and  (not A169) );
 a62449a <=( (not A170)  and  a62448a );
 a62453a <=( (not A201)  and  A200 );
 a62454a <=( A199  and  a62453a );
 a62455a <=( a62454a  and  a62449a );
 a62459a <=( A267  and  A265 );
 a62460a <=( A203  and  a62459a );
 a62463a <=( A299  and  A298 );
 a62466a <=( A302  and  (not A300) );
 a62467a <=( a62466a  and  a62463a );
 a62468a <=( a62467a  and  a62460a );
 a62472a <=( (not A167)  and  (not A169) );
 a62473a <=( (not A170)  and  a62472a );
 a62477a <=( (not A201)  and  A200 );
 a62478a <=( A199  and  a62477a );
 a62479a <=( a62478a  and  a62473a );
 a62483a <=( A267  and  A265 );
 a62484a <=( A203  and  a62483a );
 a62487a <=( (not A299)  and  A298 );
 a62490a <=( A301  and  (not A300) );
 a62491a <=( a62490a  and  a62487a );
 a62492a <=( a62491a  and  a62484a );
 a62496a <=( (not A167)  and  (not A169) );
 a62497a <=( (not A170)  and  a62496a );
 a62501a <=( (not A201)  and  A200 );
 a62502a <=( A199  and  a62501a );
 a62503a <=( a62502a  and  a62497a );
 a62507a <=( A267  and  A265 );
 a62508a <=( A203  and  a62507a );
 a62511a <=( (not A299)  and  A298 );
 a62514a <=( (not A302)  and  (not A300) );
 a62515a <=( a62514a  and  a62511a );
 a62516a <=( a62515a  and  a62508a );
 a62520a <=( (not A167)  and  (not A169) );
 a62521a <=( (not A170)  and  a62520a );
 a62525a <=( (not A201)  and  A200 );
 a62526a <=( A199  and  a62525a );
 a62527a <=( a62526a  and  a62521a );
 a62531a <=( A267  and  A265 );
 a62532a <=( A203  and  a62531a );
 a62535a <=( A299  and  (not A298) );
 a62538a <=( A301  and  (not A300) );
 a62539a <=( a62538a  and  a62535a );
 a62540a <=( a62539a  and  a62532a );
 a62544a <=( (not A167)  and  (not A169) );
 a62545a <=( (not A170)  and  a62544a );
 a62549a <=( (not A201)  and  A200 );
 a62550a <=( A199  and  a62549a );
 a62551a <=( a62550a  and  a62545a );
 a62555a <=( A267  and  A265 );
 a62556a <=( A203  and  a62555a );
 a62559a <=( A299  and  (not A298) );
 a62562a <=( (not A302)  and  (not A300) );
 a62563a <=( a62562a  and  a62559a );
 a62564a <=( a62563a  and  a62556a );
 a62568a <=( (not A167)  and  (not A169) );
 a62569a <=( (not A170)  and  a62568a );
 a62573a <=( (not A201)  and  A200 );
 a62574a <=( A199  and  a62573a );
 a62575a <=( a62574a  and  a62569a );
 a62579a <=( A267  and  A266 );
 a62580a <=( A203  and  a62579a );
 a62583a <=( A299  and  A298 );
 a62586a <=( (not A301)  and  (not A300) );
 a62587a <=( a62586a  and  a62583a );
 a62588a <=( a62587a  and  a62580a );
 a62592a <=( (not A167)  and  (not A169) );
 a62593a <=( (not A170)  and  a62592a );
 a62597a <=( (not A201)  and  A200 );
 a62598a <=( A199  and  a62597a );
 a62599a <=( a62598a  and  a62593a );
 a62603a <=( A267  and  A266 );
 a62604a <=( A203  and  a62603a );
 a62607a <=( A299  and  A298 );
 a62610a <=( A302  and  (not A300) );
 a62611a <=( a62610a  and  a62607a );
 a62612a <=( a62611a  and  a62604a );
 a62616a <=( (not A167)  and  (not A169) );
 a62617a <=( (not A170)  and  a62616a );
 a62621a <=( (not A201)  and  A200 );
 a62622a <=( A199  and  a62621a );
 a62623a <=( a62622a  and  a62617a );
 a62627a <=( A267  and  A266 );
 a62628a <=( A203  and  a62627a );
 a62631a <=( (not A299)  and  A298 );
 a62634a <=( A301  and  (not A300) );
 a62635a <=( a62634a  and  a62631a );
 a62636a <=( a62635a  and  a62628a );
 a62640a <=( (not A167)  and  (not A169) );
 a62641a <=( (not A170)  and  a62640a );
 a62645a <=( (not A201)  and  A200 );
 a62646a <=( A199  and  a62645a );
 a62647a <=( a62646a  and  a62641a );
 a62651a <=( A267  and  A266 );
 a62652a <=( A203  and  a62651a );
 a62655a <=( (not A299)  and  A298 );
 a62658a <=( (not A302)  and  (not A300) );
 a62659a <=( a62658a  and  a62655a );
 a62660a <=( a62659a  and  a62652a );
 a62664a <=( (not A167)  and  (not A169) );
 a62665a <=( (not A170)  and  a62664a );
 a62669a <=( (not A201)  and  A200 );
 a62670a <=( A199  and  a62669a );
 a62671a <=( a62670a  and  a62665a );
 a62675a <=( A267  and  A266 );
 a62676a <=( A203  and  a62675a );
 a62679a <=( A299  and  (not A298) );
 a62682a <=( A301  and  (not A300) );
 a62683a <=( a62682a  and  a62679a );
 a62684a <=( a62683a  and  a62676a );
 a62688a <=( (not A167)  and  (not A169) );
 a62689a <=( (not A170)  and  a62688a );
 a62693a <=( (not A201)  and  A200 );
 a62694a <=( A199  and  a62693a );
 a62695a <=( a62694a  and  a62689a );
 a62699a <=( A267  and  A266 );
 a62700a <=( A203  and  a62699a );
 a62703a <=( A299  and  (not A298) );
 a62706a <=( (not A302)  and  (not A300) );
 a62707a <=( a62706a  and  a62703a );
 a62708a <=( a62707a  and  a62700a );
 a62712a <=( (not A167)  and  (not A169) );
 a62713a <=( (not A170)  and  a62712a );
 a62717a <=( (not A202)  and  A200 );
 a62718a <=( (not A199)  and  a62717a );
 a62719a <=( a62718a  and  a62713a );
 a62723a <=( A266  and  A265 );
 a62724a <=( A203  and  a62723a );
 a62727a <=( (not A268)  and  (not A267) );
 a62730a <=( A300  and  A299 );
 a62731a <=( a62730a  and  a62727a );
 a62732a <=( a62731a  and  a62724a );
 a62736a <=( (not A167)  and  (not A169) );
 a62737a <=( (not A170)  and  a62736a );
 a62741a <=( (not A202)  and  A200 );
 a62742a <=( (not A199)  and  a62741a );
 a62743a <=( a62742a  and  a62737a );
 a62747a <=( A266  and  A265 );
 a62748a <=( A203  and  a62747a );
 a62751a <=( (not A268)  and  (not A267) );
 a62754a <=( A300  and  A298 );
 a62755a <=( a62754a  and  a62751a );
 a62756a <=( a62755a  and  a62748a );
 a62760a <=( (not A167)  and  (not A169) );
 a62761a <=( (not A170)  and  a62760a );
 a62765a <=( (not A202)  and  A200 );
 a62766a <=( (not A199)  and  a62765a );
 a62767a <=( a62766a  and  a62761a );
 a62771a <=( A266  and  A265 );
 a62772a <=( A203  and  a62771a );
 a62775a <=( A269  and  (not A267) );
 a62778a <=( A300  and  A299 );
 a62779a <=( a62778a  and  a62775a );
 a62780a <=( a62779a  and  a62772a );
 a62784a <=( (not A167)  and  (not A169) );
 a62785a <=( (not A170)  and  a62784a );
 a62789a <=( (not A202)  and  A200 );
 a62790a <=( (not A199)  and  a62789a );
 a62791a <=( a62790a  and  a62785a );
 a62795a <=( A266  and  A265 );
 a62796a <=( A203  and  a62795a );
 a62799a <=( A269  and  (not A267) );
 a62802a <=( A300  and  A298 );
 a62803a <=( a62802a  and  a62799a );
 a62804a <=( a62803a  and  a62796a );
 a62808a <=( (not A167)  and  (not A169) );
 a62809a <=( (not A170)  and  a62808a );
 a62813a <=( (not A202)  and  A200 );
 a62814a <=( (not A199)  and  a62813a );
 a62815a <=( a62814a  and  a62809a );
 a62819a <=( A266  and  (not A265) );
 a62820a <=( A203  and  a62819a );
 a62823a <=( A268  and  (not A267) );
 a62826a <=( A300  and  A299 );
 a62827a <=( a62826a  and  a62823a );
 a62828a <=( a62827a  and  a62820a );
 a62832a <=( (not A167)  and  (not A169) );
 a62833a <=( (not A170)  and  a62832a );
 a62837a <=( (not A202)  and  A200 );
 a62838a <=( (not A199)  and  a62837a );
 a62839a <=( a62838a  and  a62833a );
 a62843a <=( A266  and  (not A265) );
 a62844a <=( A203  and  a62843a );
 a62847a <=( A268  and  (not A267) );
 a62850a <=( A300  and  A298 );
 a62851a <=( a62850a  and  a62847a );
 a62852a <=( a62851a  and  a62844a );
 a62856a <=( (not A167)  and  (not A169) );
 a62857a <=( (not A170)  and  a62856a );
 a62861a <=( (not A202)  and  A200 );
 a62862a <=( (not A199)  and  a62861a );
 a62863a <=( a62862a  and  a62857a );
 a62867a <=( A266  and  (not A265) );
 a62868a <=( A203  and  a62867a );
 a62871a <=( (not A269)  and  (not A267) );
 a62874a <=( A300  and  A299 );
 a62875a <=( a62874a  and  a62871a );
 a62876a <=( a62875a  and  a62868a );
 a62880a <=( (not A167)  and  (not A169) );
 a62881a <=( (not A170)  and  a62880a );
 a62885a <=( (not A202)  and  A200 );
 a62886a <=( (not A199)  and  a62885a );
 a62887a <=( a62886a  and  a62881a );
 a62891a <=( A266  and  (not A265) );
 a62892a <=( A203  and  a62891a );
 a62895a <=( (not A269)  and  (not A267) );
 a62898a <=( A300  and  A298 );
 a62899a <=( a62898a  and  a62895a );
 a62900a <=( a62899a  and  a62892a );
 a62904a <=( (not A167)  and  (not A169) );
 a62905a <=( (not A170)  and  a62904a );
 a62909a <=( (not A202)  and  A200 );
 a62910a <=( (not A199)  and  a62909a );
 a62911a <=( a62910a  and  a62905a );
 a62915a <=( (not A266)  and  A265 );
 a62916a <=( A203  and  a62915a );
 a62919a <=( A268  and  (not A267) );
 a62922a <=( A300  and  A299 );
 a62923a <=( a62922a  and  a62919a );
 a62924a <=( a62923a  and  a62916a );
 a62928a <=( (not A167)  and  (not A169) );
 a62929a <=( (not A170)  and  a62928a );
 a62933a <=( (not A202)  and  A200 );
 a62934a <=( (not A199)  and  a62933a );
 a62935a <=( a62934a  and  a62929a );
 a62939a <=( (not A266)  and  A265 );
 a62940a <=( A203  and  a62939a );
 a62943a <=( A268  and  (not A267) );
 a62946a <=( A300  and  A298 );
 a62947a <=( a62946a  and  a62943a );
 a62948a <=( a62947a  and  a62940a );
 a62952a <=( (not A167)  and  (not A169) );
 a62953a <=( (not A170)  and  a62952a );
 a62957a <=( (not A202)  and  A200 );
 a62958a <=( (not A199)  and  a62957a );
 a62959a <=( a62958a  and  a62953a );
 a62963a <=( (not A266)  and  A265 );
 a62964a <=( A203  and  a62963a );
 a62967a <=( (not A269)  and  (not A267) );
 a62970a <=( A300  and  A299 );
 a62971a <=( a62970a  and  a62967a );
 a62972a <=( a62971a  and  a62964a );
 a62976a <=( (not A167)  and  (not A169) );
 a62977a <=( (not A170)  and  a62976a );
 a62981a <=( (not A202)  and  A200 );
 a62982a <=( (not A199)  and  a62981a );
 a62983a <=( a62982a  and  a62977a );
 a62987a <=( (not A266)  and  A265 );
 a62988a <=( A203  and  a62987a );
 a62991a <=( (not A269)  and  (not A267) );
 a62994a <=( A300  and  A298 );
 a62995a <=( a62994a  and  a62991a );
 a62996a <=( a62995a  and  a62988a );
 a63000a <=( (not A167)  and  (not A169) );
 a63001a <=( (not A170)  and  a63000a );
 a63005a <=( (not A201)  and  A200 );
 a63006a <=( (not A199)  and  a63005a );
 a63007a <=( a63006a  and  a63001a );
 a63011a <=( A267  and  A265 );
 a63012a <=( A202  and  a63011a );
 a63015a <=( A299  and  A298 );
 a63018a <=( (not A301)  and  (not A300) );
 a63019a <=( a63018a  and  a63015a );
 a63020a <=( a63019a  and  a63012a );
 a63024a <=( (not A167)  and  (not A169) );
 a63025a <=( (not A170)  and  a63024a );
 a63029a <=( (not A201)  and  A200 );
 a63030a <=( (not A199)  and  a63029a );
 a63031a <=( a63030a  and  a63025a );
 a63035a <=( A267  and  A265 );
 a63036a <=( A202  and  a63035a );
 a63039a <=( A299  and  A298 );
 a63042a <=( A302  and  (not A300) );
 a63043a <=( a63042a  and  a63039a );
 a63044a <=( a63043a  and  a63036a );
 a63048a <=( (not A167)  and  (not A169) );
 a63049a <=( (not A170)  and  a63048a );
 a63053a <=( (not A201)  and  A200 );
 a63054a <=( (not A199)  and  a63053a );
 a63055a <=( a63054a  and  a63049a );
 a63059a <=( A267  and  A265 );
 a63060a <=( A202  and  a63059a );
 a63063a <=( (not A299)  and  A298 );
 a63066a <=( A301  and  (not A300) );
 a63067a <=( a63066a  and  a63063a );
 a63068a <=( a63067a  and  a63060a );
 a63072a <=( (not A167)  and  (not A169) );
 a63073a <=( (not A170)  and  a63072a );
 a63077a <=( (not A201)  and  A200 );
 a63078a <=( (not A199)  and  a63077a );
 a63079a <=( a63078a  and  a63073a );
 a63083a <=( A267  and  A265 );
 a63084a <=( A202  and  a63083a );
 a63087a <=( (not A299)  and  A298 );
 a63090a <=( (not A302)  and  (not A300) );
 a63091a <=( a63090a  and  a63087a );
 a63092a <=( a63091a  and  a63084a );
 a63096a <=( (not A167)  and  (not A169) );
 a63097a <=( (not A170)  and  a63096a );
 a63101a <=( (not A201)  and  A200 );
 a63102a <=( (not A199)  and  a63101a );
 a63103a <=( a63102a  and  a63097a );
 a63107a <=( A267  and  A265 );
 a63108a <=( A202  and  a63107a );
 a63111a <=( A299  and  (not A298) );
 a63114a <=( A301  and  (not A300) );
 a63115a <=( a63114a  and  a63111a );
 a63116a <=( a63115a  and  a63108a );
 a63120a <=( (not A167)  and  (not A169) );
 a63121a <=( (not A170)  and  a63120a );
 a63125a <=( (not A201)  and  A200 );
 a63126a <=( (not A199)  and  a63125a );
 a63127a <=( a63126a  and  a63121a );
 a63131a <=( A267  and  A265 );
 a63132a <=( A202  and  a63131a );
 a63135a <=( A299  and  (not A298) );
 a63138a <=( (not A302)  and  (not A300) );
 a63139a <=( a63138a  and  a63135a );
 a63140a <=( a63139a  and  a63132a );
 a63144a <=( (not A167)  and  (not A169) );
 a63145a <=( (not A170)  and  a63144a );
 a63149a <=( (not A201)  and  A200 );
 a63150a <=( (not A199)  and  a63149a );
 a63151a <=( a63150a  and  a63145a );
 a63155a <=( A267  and  A266 );
 a63156a <=( A202  and  a63155a );
 a63159a <=( A299  and  A298 );
 a63162a <=( (not A301)  and  (not A300) );
 a63163a <=( a63162a  and  a63159a );
 a63164a <=( a63163a  and  a63156a );
 a63168a <=( (not A167)  and  (not A169) );
 a63169a <=( (not A170)  and  a63168a );
 a63173a <=( (not A201)  and  A200 );
 a63174a <=( (not A199)  and  a63173a );
 a63175a <=( a63174a  and  a63169a );
 a63179a <=( A267  and  A266 );
 a63180a <=( A202  and  a63179a );
 a63183a <=( A299  and  A298 );
 a63186a <=( A302  and  (not A300) );
 a63187a <=( a63186a  and  a63183a );
 a63188a <=( a63187a  and  a63180a );
 a63192a <=( (not A167)  and  (not A169) );
 a63193a <=( (not A170)  and  a63192a );
 a63197a <=( (not A201)  and  A200 );
 a63198a <=( (not A199)  and  a63197a );
 a63199a <=( a63198a  and  a63193a );
 a63203a <=( A267  and  A266 );
 a63204a <=( A202  and  a63203a );
 a63207a <=( (not A299)  and  A298 );
 a63210a <=( A301  and  (not A300) );
 a63211a <=( a63210a  and  a63207a );
 a63212a <=( a63211a  and  a63204a );
 a63216a <=( (not A167)  and  (not A169) );
 a63217a <=( (not A170)  and  a63216a );
 a63221a <=( (not A201)  and  A200 );
 a63222a <=( (not A199)  and  a63221a );
 a63223a <=( a63222a  and  a63217a );
 a63227a <=( A267  and  A266 );
 a63228a <=( A202  and  a63227a );
 a63231a <=( (not A299)  and  A298 );
 a63234a <=( (not A302)  and  (not A300) );
 a63235a <=( a63234a  and  a63231a );
 a63236a <=( a63235a  and  a63228a );
 a63240a <=( (not A167)  and  (not A169) );
 a63241a <=( (not A170)  and  a63240a );
 a63245a <=( (not A201)  and  A200 );
 a63246a <=( (not A199)  and  a63245a );
 a63247a <=( a63246a  and  a63241a );
 a63251a <=( A267  and  A266 );
 a63252a <=( A202  and  a63251a );
 a63255a <=( A299  and  (not A298) );
 a63258a <=( A301  and  (not A300) );
 a63259a <=( a63258a  and  a63255a );
 a63260a <=( a63259a  and  a63252a );
 a63264a <=( (not A167)  and  (not A169) );
 a63265a <=( (not A170)  and  a63264a );
 a63269a <=( (not A201)  and  A200 );
 a63270a <=( (not A199)  and  a63269a );
 a63271a <=( a63270a  and  a63265a );
 a63275a <=( A267  and  A266 );
 a63276a <=( A202  and  a63275a );
 a63279a <=( A299  and  (not A298) );
 a63282a <=( (not A302)  and  (not A300) );
 a63283a <=( a63282a  and  a63279a );
 a63284a <=( a63283a  and  a63276a );
 a63288a <=( (not A167)  and  (not A169) );
 a63289a <=( (not A170)  and  a63288a );
 a63293a <=( (not A201)  and  A200 );
 a63294a <=( (not A199)  and  a63293a );
 a63295a <=( a63294a  and  a63289a );
 a63299a <=( A267  and  A265 );
 a63300a <=( (not A203)  and  a63299a );
 a63303a <=( A299  and  A298 );
 a63306a <=( (not A301)  and  (not A300) );
 a63307a <=( a63306a  and  a63303a );
 a63308a <=( a63307a  and  a63300a );
 a63312a <=( (not A167)  and  (not A169) );
 a63313a <=( (not A170)  and  a63312a );
 a63317a <=( (not A201)  and  A200 );
 a63318a <=( (not A199)  and  a63317a );
 a63319a <=( a63318a  and  a63313a );
 a63323a <=( A267  and  A265 );
 a63324a <=( (not A203)  and  a63323a );
 a63327a <=( A299  and  A298 );
 a63330a <=( A302  and  (not A300) );
 a63331a <=( a63330a  and  a63327a );
 a63332a <=( a63331a  and  a63324a );
 a63336a <=( (not A167)  and  (not A169) );
 a63337a <=( (not A170)  and  a63336a );
 a63341a <=( (not A201)  and  A200 );
 a63342a <=( (not A199)  and  a63341a );
 a63343a <=( a63342a  and  a63337a );
 a63347a <=( A267  and  A265 );
 a63348a <=( (not A203)  and  a63347a );
 a63351a <=( (not A299)  and  A298 );
 a63354a <=( A301  and  (not A300) );
 a63355a <=( a63354a  and  a63351a );
 a63356a <=( a63355a  and  a63348a );
 a63360a <=( (not A167)  and  (not A169) );
 a63361a <=( (not A170)  and  a63360a );
 a63365a <=( (not A201)  and  A200 );
 a63366a <=( (not A199)  and  a63365a );
 a63367a <=( a63366a  and  a63361a );
 a63371a <=( A267  and  A265 );
 a63372a <=( (not A203)  and  a63371a );
 a63375a <=( (not A299)  and  A298 );
 a63378a <=( (not A302)  and  (not A300) );
 a63379a <=( a63378a  and  a63375a );
 a63380a <=( a63379a  and  a63372a );
 a63384a <=( (not A167)  and  (not A169) );
 a63385a <=( (not A170)  and  a63384a );
 a63389a <=( (not A201)  and  A200 );
 a63390a <=( (not A199)  and  a63389a );
 a63391a <=( a63390a  and  a63385a );
 a63395a <=( A267  and  A265 );
 a63396a <=( (not A203)  and  a63395a );
 a63399a <=( A299  and  (not A298) );
 a63402a <=( A301  and  (not A300) );
 a63403a <=( a63402a  and  a63399a );
 a63404a <=( a63403a  and  a63396a );
 a63408a <=( (not A167)  and  (not A169) );
 a63409a <=( (not A170)  and  a63408a );
 a63413a <=( (not A201)  and  A200 );
 a63414a <=( (not A199)  and  a63413a );
 a63415a <=( a63414a  and  a63409a );
 a63419a <=( A267  and  A265 );
 a63420a <=( (not A203)  and  a63419a );
 a63423a <=( A299  and  (not A298) );
 a63426a <=( (not A302)  and  (not A300) );
 a63427a <=( a63426a  and  a63423a );
 a63428a <=( a63427a  and  a63420a );
 a63432a <=( (not A167)  and  (not A169) );
 a63433a <=( (not A170)  and  a63432a );
 a63437a <=( (not A201)  and  A200 );
 a63438a <=( (not A199)  and  a63437a );
 a63439a <=( a63438a  and  a63433a );
 a63443a <=( A267  and  A266 );
 a63444a <=( (not A203)  and  a63443a );
 a63447a <=( A299  and  A298 );
 a63450a <=( (not A301)  and  (not A300) );
 a63451a <=( a63450a  and  a63447a );
 a63452a <=( a63451a  and  a63444a );
 a63456a <=( (not A167)  and  (not A169) );
 a63457a <=( (not A170)  and  a63456a );
 a63461a <=( (not A201)  and  A200 );
 a63462a <=( (not A199)  and  a63461a );
 a63463a <=( a63462a  and  a63457a );
 a63467a <=( A267  and  A266 );
 a63468a <=( (not A203)  and  a63467a );
 a63471a <=( A299  and  A298 );
 a63474a <=( A302  and  (not A300) );
 a63475a <=( a63474a  and  a63471a );
 a63476a <=( a63475a  and  a63468a );
 a63480a <=( (not A167)  and  (not A169) );
 a63481a <=( (not A170)  and  a63480a );
 a63485a <=( (not A201)  and  A200 );
 a63486a <=( (not A199)  and  a63485a );
 a63487a <=( a63486a  and  a63481a );
 a63491a <=( A267  and  A266 );
 a63492a <=( (not A203)  and  a63491a );
 a63495a <=( (not A299)  and  A298 );
 a63498a <=( A301  and  (not A300) );
 a63499a <=( a63498a  and  a63495a );
 a63500a <=( a63499a  and  a63492a );
 a63504a <=( (not A167)  and  (not A169) );
 a63505a <=( (not A170)  and  a63504a );
 a63509a <=( (not A201)  and  A200 );
 a63510a <=( (not A199)  and  a63509a );
 a63511a <=( a63510a  and  a63505a );
 a63515a <=( A267  and  A266 );
 a63516a <=( (not A203)  and  a63515a );
 a63519a <=( (not A299)  and  A298 );
 a63522a <=( (not A302)  and  (not A300) );
 a63523a <=( a63522a  and  a63519a );
 a63524a <=( a63523a  and  a63516a );
 a63528a <=( (not A167)  and  (not A169) );
 a63529a <=( (not A170)  and  a63528a );
 a63533a <=( (not A201)  and  A200 );
 a63534a <=( (not A199)  and  a63533a );
 a63535a <=( a63534a  and  a63529a );
 a63539a <=( A267  and  A266 );
 a63540a <=( (not A203)  and  a63539a );
 a63543a <=( A299  and  (not A298) );
 a63546a <=( A301  and  (not A300) );
 a63547a <=( a63546a  and  a63543a );
 a63548a <=( a63547a  and  a63540a );
 a63552a <=( (not A167)  and  (not A169) );
 a63553a <=( (not A170)  and  a63552a );
 a63557a <=( (not A201)  and  A200 );
 a63558a <=( (not A199)  and  a63557a );
 a63559a <=( a63558a  and  a63553a );
 a63563a <=( A267  and  A266 );
 a63564a <=( (not A203)  and  a63563a );
 a63567a <=( A299  and  (not A298) );
 a63570a <=( (not A302)  and  (not A300) );
 a63571a <=( a63570a  and  a63567a );
 a63572a <=( a63571a  and  a63564a );
 a63576a <=( (not A167)  and  (not A169) );
 a63577a <=( (not A170)  and  a63576a );
 a63581a <=( (not A202)  and  (not A200) );
 a63582a <=( A199  and  a63581a );
 a63583a <=( a63582a  and  a63577a );
 a63587a <=( A266  and  A265 );
 a63588a <=( A203  and  a63587a );
 a63591a <=( (not A268)  and  (not A267) );
 a63594a <=( A300  and  A299 );
 a63595a <=( a63594a  and  a63591a );
 a63596a <=( a63595a  and  a63588a );
 a63600a <=( (not A167)  and  (not A169) );
 a63601a <=( (not A170)  and  a63600a );
 a63605a <=( (not A202)  and  (not A200) );
 a63606a <=( A199  and  a63605a );
 a63607a <=( a63606a  and  a63601a );
 a63611a <=( A266  and  A265 );
 a63612a <=( A203  and  a63611a );
 a63615a <=( (not A268)  and  (not A267) );
 a63618a <=( A300  and  A298 );
 a63619a <=( a63618a  and  a63615a );
 a63620a <=( a63619a  and  a63612a );
 a63624a <=( (not A167)  and  (not A169) );
 a63625a <=( (not A170)  and  a63624a );
 a63629a <=( (not A202)  and  (not A200) );
 a63630a <=( A199  and  a63629a );
 a63631a <=( a63630a  and  a63625a );
 a63635a <=( A266  and  A265 );
 a63636a <=( A203  and  a63635a );
 a63639a <=( A269  and  (not A267) );
 a63642a <=( A300  and  A299 );
 a63643a <=( a63642a  and  a63639a );
 a63644a <=( a63643a  and  a63636a );
 a63648a <=( (not A167)  and  (not A169) );
 a63649a <=( (not A170)  and  a63648a );
 a63653a <=( (not A202)  and  (not A200) );
 a63654a <=( A199  and  a63653a );
 a63655a <=( a63654a  and  a63649a );
 a63659a <=( A266  and  A265 );
 a63660a <=( A203  and  a63659a );
 a63663a <=( A269  and  (not A267) );
 a63666a <=( A300  and  A298 );
 a63667a <=( a63666a  and  a63663a );
 a63668a <=( a63667a  and  a63660a );
 a63672a <=( (not A167)  and  (not A169) );
 a63673a <=( (not A170)  and  a63672a );
 a63677a <=( (not A202)  and  (not A200) );
 a63678a <=( A199  and  a63677a );
 a63679a <=( a63678a  and  a63673a );
 a63683a <=( A266  and  (not A265) );
 a63684a <=( A203  and  a63683a );
 a63687a <=( A268  and  (not A267) );
 a63690a <=( A300  and  A299 );
 a63691a <=( a63690a  and  a63687a );
 a63692a <=( a63691a  and  a63684a );
 a63696a <=( (not A167)  and  (not A169) );
 a63697a <=( (not A170)  and  a63696a );
 a63701a <=( (not A202)  and  (not A200) );
 a63702a <=( A199  and  a63701a );
 a63703a <=( a63702a  and  a63697a );
 a63707a <=( A266  and  (not A265) );
 a63708a <=( A203  and  a63707a );
 a63711a <=( A268  and  (not A267) );
 a63714a <=( A300  and  A298 );
 a63715a <=( a63714a  and  a63711a );
 a63716a <=( a63715a  and  a63708a );
 a63720a <=( (not A167)  and  (not A169) );
 a63721a <=( (not A170)  and  a63720a );
 a63725a <=( (not A202)  and  (not A200) );
 a63726a <=( A199  and  a63725a );
 a63727a <=( a63726a  and  a63721a );
 a63731a <=( A266  and  (not A265) );
 a63732a <=( A203  and  a63731a );
 a63735a <=( (not A269)  and  (not A267) );
 a63738a <=( A300  and  A299 );
 a63739a <=( a63738a  and  a63735a );
 a63740a <=( a63739a  and  a63732a );
 a63744a <=( (not A167)  and  (not A169) );
 a63745a <=( (not A170)  and  a63744a );
 a63749a <=( (not A202)  and  (not A200) );
 a63750a <=( A199  and  a63749a );
 a63751a <=( a63750a  and  a63745a );
 a63755a <=( A266  and  (not A265) );
 a63756a <=( A203  and  a63755a );
 a63759a <=( (not A269)  and  (not A267) );
 a63762a <=( A300  and  A298 );
 a63763a <=( a63762a  and  a63759a );
 a63764a <=( a63763a  and  a63756a );
 a63768a <=( (not A167)  and  (not A169) );
 a63769a <=( (not A170)  and  a63768a );
 a63773a <=( (not A202)  and  (not A200) );
 a63774a <=( A199  and  a63773a );
 a63775a <=( a63774a  and  a63769a );
 a63779a <=( (not A266)  and  A265 );
 a63780a <=( A203  and  a63779a );
 a63783a <=( A268  and  (not A267) );
 a63786a <=( A300  and  A299 );
 a63787a <=( a63786a  and  a63783a );
 a63788a <=( a63787a  and  a63780a );
 a63792a <=( (not A167)  and  (not A169) );
 a63793a <=( (not A170)  and  a63792a );
 a63797a <=( (not A202)  and  (not A200) );
 a63798a <=( A199  and  a63797a );
 a63799a <=( a63798a  and  a63793a );
 a63803a <=( (not A266)  and  A265 );
 a63804a <=( A203  and  a63803a );
 a63807a <=( A268  and  (not A267) );
 a63810a <=( A300  and  A298 );
 a63811a <=( a63810a  and  a63807a );
 a63812a <=( a63811a  and  a63804a );
 a63816a <=( (not A167)  and  (not A169) );
 a63817a <=( (not A170)  and  a63816a );
 a63821a <=( (not A202)  and  (not A200) );
 a63822a <=( A199  and  a63821a );
 a63823a <=( a63822a  and  a63817a );
 a63827a <=( (not A266)  and  A265 );
 a63828a <=( A203  and  a63827a );
 a63831a <=( (not A269)  and  (not A267) );
 a63834a <=( A300  and  A299 );
 a63835a <=( a63834a  and  a63831a );
 a63836a <=( a63835a  and  a63828a );
 a63840a <=( (not A167)  and  (not A169) );
 a63841a <=( (not A170)  and  a63840a );
 a63845a <=( (not A202)  and  (not A200) );
 a63846a <=( A199  and  a63845a );
 a63847a <=( a63846a  and  a63841a );
 a63851a <=( (not A266)  and  A265 );
 a63852a <=( A203  and  a63851a );
 a63855a <=( (not A269)  and  (not A267) );
 a63858a <=( A300  and  A298 );
 a63859a <=( a63858a  and  a63855a );
 a63860a <=( a63859a  and  a63852a );
 a63864a <=( (not A167)  and  (not A169) );
 a63865a <=( (not A170)  and  a63864a );
 a63869a <=( (not A201)  and  (not A200) );
 a63870a <=( A199  and  a63869a );
 a63871a <=( a63870a  and  a63865a );
 a63875a <=( A267  and  A265 );
 a63876a <=( A202  and  a63875a );
 a63879a <=( A299  and  A298 );
 a63882a <=( (not A301)  and  (not A300) );
 a63883a <=( a63882a  and  a63879a );
 a63884a <=( a63883a  and  a63876a );
 a63888a <=( (not A167)  and  (not A169) );
 a63889a <=( (not A170)  and  a63888a );
 a63893a <=( (not A201)  and  (not A200) );
 a63894a <=( A199  and  a63893a );
 a63895a <=( a63894a  and  a63889a );
 a63899a <=( A267  and  A265 );
 a63900a <=( A202  and  a63899a );
 a63903a <=( A299  and  A298 );
 a63906a <=( A302  and  (not A300) );
 a63907a <=( a63906a  and  a63903a );
 a63908a <=( a63907a  and  a63900a );
 a63912a <=( (not A167)  and  (not A169) );
 a63913a <=( (not A170)  and  a63912a );
 a63917a <=( (not A201)  and  (not A200) );
 a63918a <=( A199  and  a63917a );
 a63919a <=( a63918a  and  a63913a );
 a63923a <=( A267  and  A265 );
 a63924a <=( A202  and  a63923a );
 a63927a <=( (not A299)  and  A298 );
 a63930a <=( A301  and  (not A300) );
 a63931a <=( a63930a  and  a63927a );
 a63932a <=( a63931a  and  a63924a );
 a63936a <=( (not A167)  and  (not A169) );
 a63937a <=( (not A170)  and  a63936a );
 a63941a <=( (not A201)  and  (not A200) );
 a63942a <=( A199  and  a63941a );
 a63943a <=( a63942a  and  a63937a );
 a63947a <=( A267  and  A265 );
 a63948a <=( A202  and  a63947a );
 a63951a <=( (not A299)  and  A298 );
 a63954a <=( (not A302)  and  (not A300) );
 a63955a <=( a63954a  and  a63951a );
 a63956a <=( a63955a  and  a63948a );
 a63960a <=( (not A167)  and  (not A169) );
 a63961a <=( (not A170)  and  a63960a );
 a63965a <=( (not A201)  and  (not A200) );
 a63966a <=( A199  and  a63965a );
 a63967a <=( a63966a  and  a63961a );
 a63971a <=( A267  and  A265 );
 a63972a <=( A202  and  a63971a );
 a63975a <=( A299  and  (not A298) );
 a63978a <=( A301  and  (not A300) );
 a63979a <=( a63978a  and  a63975a );
 a63980a <=( a63979a  and  a63972a );
 a63984a <=( (not A167)  and  (not A169) );
 a63985a <=( (not A170)  and  a63984a );
 a63989a <=( (not A201)  and  (not A200) );
 a63990a <=( A199  and  a63989a );
 a63991a <=( a63990a  and  a63985a );
 a63995a <=( A267  and  A265 );
 a63996a <=( A202  and  a63995a );
 a63999a <=( A299  and  (not A298) );
 a64002a <=( (not A302)  and  (not A300) );
 a64003a <=( a64002a  and  a63999a );
 a64004a <=( a64003a  and  a63996a );
 a64008a <=( (not A167)  and  (not A169) );
 a64009a <=( (not A170)  and  a64008a );
 a64013a <=( (not A201)  and  (not A200) );
 a64014a <=( A199  and  a64013a );
 a64015a <=( a64014a  and  a64009a );
 a64019a <=( A267  and  A266 );
 a64020a <=( A202  and  a64019a );
 a64023a <=( A299  and  A298 );
 a64026a <=( (not A301)  and  (not A300) );
 a64027a <=( a64026a  and  a64023a );
 a64028a <=( a64027a  and  a64020a );
 a64032a <=( (not A167)  and  (not A169) );
 a64033a <=( (not A170)  and  a64032a );
 a64037a <=( (not A201)  and  (not A200) );
 a64038a <=( A199  and  a64037a );
 a64039a <=( a64038a  and  a64033a );
 a64043a <=( A267  and  A266 );
 a64044a <=( A202  and  a64043a );
 a64047a <=( A299  and  A298 );
 a64050a <=( A302  and  (not A300) );
 a64051a <=( a64050a  and  a64047a );
 a64052a <=( a64051a  and  a64044a );
 a64056a <=( (not A167)  and  (not A169) );
 a64057a <=( (not A170)  and  a64056a );
 a64061a <=( (not A201)  and  (not A200) );
 a64062a <=( A199  and  a64061a );
 a64063a <=( a64062a  and  a64057a );
 a64067a <=( A267  and  A266 );
 a64068a <=( A202  and  a64067a );
 a64071a <=( (not A299)  and  A298 );
 a64074a <=( A301  and  (not A300) );
 a64075a <=( a64074a  and  a64071a );
 a64076a <=( a64075a  and  a64068a );
 a64080a <=( (not A167)  and  (not A169) );
 a64081a <=( (not A170)  and  a64080a );
 a64085a <=( (not A201)  and  (not A200) );
 a64086a <=( A199  and  a64085a );
 a64087a <=( a64086a  and  a64081a );
 a64091a <=( A267  and  A266 );
 a64092a <=( A202  and  a64091a );
 a64095a <=( (not A299)  and  A298 );
 a64098a <=( (not A302)  and  (not A300) );
 a64099a <=( a64098a  and  a64095a );
 a64100a <=( a64099a  and  a64092a );
 a64104a <=( (not A167)  and  (not A169) );
 a64105a <=( (not A170)  and  a64104a );
 a64109a <=( (not A201)  and  (not A200) );
 a64110a <=( A199  and  a64109a );
 a64111a <=( a64110a  and  a64105a );
 a64115a <=( A267  and  A266 );
 a64116a <=( A202  and  a64115a );
 a64119a <=( A299  and  (not A298) );
 a64122a <=( A301  and  (not A300) );
 a64123a <=( a64122a  and  a64119a );
 a64124a <=( a64123a  and  a64116a );
 a64128a <=( (not A167)  and  (not A169) );
 a64129a <=( (not A170)  and  a64128a );
 a64133a <=( (not A201)  and  (not A200) );
 a64134a <=( A199  and  a64133a );
 a64135a <=( a64134a  and  a64129a );
 a64139a <=( A267  and  A266 );
 a64140a <=( A202  and  a64139a );
 a64143a <=( A299  and  (not A298) );
 a64146a <=( (not A302)  and  (not A300) );
 a64147a <=( a64146a  and  a64143a );
 a64148a <=( a64147a  and  a64140a );
 a64152a <=( (not A167)  and  (not A169) );
 a64153a <=( (not A170)  and  a64152a );
 a64157a <=( (not A201)  and  (not A200) );
 a64158a <=( A199  and  a64157a );
 a64159a <=( a64158a  and  a64153a );
 a64163a <=( A267  and  A265 );
 a64164a <=( (not A203)  and  a64163a );
 a64167a <=( A299  and  A298 );
 a64170a <=( (not A301)  and  (not A300) );
 a64171a <=( a64170a  and  a64167a );
 a64172a <=( a64171a  and  a64164a );
 a64176a <=( (not A167)  and  (not A169) );
 a64177a <=( (not A170)  and  a64176a );
 a64181a <=( (not A201)  and  (not A200) );
 a64182a <=( A199  and  a64181a );
 a64183a <=( a64182a  and  a64177a );
 a64187a <=( A267  and  A265 );
 a64188a <=( (not A203)  and  a64187a );
 a64191a <=( A299  and  A298 );
 a64194a <=( A302  and  (not A300) );
 a64195a <=( a64194a  and  a64191a );
 a64196a <=( a64195a  and  a64188a );
 a64200a <=( (not A167)  and  (not A169) );
 a64201a <=( (not A170)  and  a64200a );
 a64205a <=( (not A201)  and  (not A200) );
 a64206a <=( A199  and  a64205a );
 a64207a <=( a64206a  and  a64201a );
 a64211a <=( A267  and  A265 );
 a64212a <=( (not A203)  and  a64211a );
 a64215a <=( (not A299)  and  A298 );
 a64218a <=( A301  and  (not A300) );
 a64219a <=( a64218a  and  a64215a );
 a64220a <=( a64219a  and  a64212a );
 a64224a <=( (not A167)  and  (not A169) );
 a64225a <=( (not A170)  and  a64224a );
 a64229a <=( (not A201)  and  (not A200) );
 a64230a <=( A199  and  a64229a );
 a64231a <=( a64230a  and  a64225a );
 a64235a <=( A267  and  A265 );
 a64236a <=( (not A203)  and  a64235a );
 a64239a <=( (not A299)  and  A298 );
 a64242a <=( (not A302)  and  (not A300) );
 a64243a <=( a64242a  and  a64239a );
 a64244a <=( a64243a  and  a64236a );
 a64248a <=( (not A167)  and  (not A169) );
 a64249a <=( (not A170)  and  a64248a );
 a64253a <=( (not A201)  and  (not A200) );
 a64254a <=( A199  and  a64253a );
 a64255a <=( a64254a  and  a64249a );
 a64259a <=( A267  and  A265 );
 a64260a <=( (not A203)  and  a64259a );
 a64263a <=( A299  and  (not A298) );
 a64266a <=( A301  and  (not A300) );
 a64267a <=( a64266a  and  a64263a );
 a64268a <=( a64267a  and  a64260a );
 a64272a <=( (not A167)  and  (not A169) );
 a64273a <=( (not A170)  and  a64272a );
 a64277a <=( (not A201)  and  (not A200) );
 a64278a <=( A199  and  a64277a );
 a64279a <=( a64278a  and  a64273a );
 a64283a <=( A267  and  A265 );
 a64284a <=( (not A203)  and  a64283a );
 a64287a <=( A299  and  (not A298) );
 a64290a <=( (not A302)  and  (not A300) );
 a64291a <=( a64290a  and  a64287a );
 a64292a <=( a64291a  and  a64284a );
 a64296a <=( (not A167)  and  (not A169) );
 a64297a <=( (not A170)  and  a64296a );
 a64301a <=( (not A201)  and  (not A200) );
 a64302a <=( A199  and  a64301a );
 a64303a <=( a64302a  and  a64297a );
 a64307a <=( A267  and  A266 );
 a64308a <=( (not A203)  and  a64307a );
 a64311a <=( A299  and  A298 );
 a64314a <=( (not A301)  and  (not A300) );
 a64315a <=( a64314a  and  a64311a );
 a64316a <=( a64315a  and  a64308a );
 a64320a <=( (not A167)  and  (not A169) );
 a64321a <=( (not A170)  and  a64320a );
 a64325a <=( (not A201)  and  (not A200) );
 a64326a <=( A199  and  a64325a );
 a64327a <=( a64326a  and  a64321a );
 a64331a <=( A267  and  A266 );
 a64332a <=( (not A203)  and  a64331a );
 a64335a <=( A299  and  A298 );
 a64338a <=( A302  and  (not A300) );
 a64339a <=( a64338a  and  a64335a );
 a64340a <=( a64339a  and  a64332a );
 a64344a <=( (not A167)  and  (not A169) );
 a64345a <=( (not A170)  and  a64344a );
 a64349a <=( (not A201)  and  (not A200) );
 a64350a <=( A199  and  a64349a );
 a64351a <=( a64350a  and  a64345a );
 a64355a <=( A267  and  A266 );
 a64356a <=( (not A203)  and  a64355a );
 a64359a <=( (not A299)  and  A298 );
 a64362a <=( A301  and  (not A300) );
 a64363a <=( a64362a  and  a64359a );
 a64364a <=( a64363a  and  a64356a );
 a64368a <=( (not A167)  and  (not A169) );
 a64369a <=( (not A170)  and  a64368a );
 a64373a <=( (not A201)  and  (not A200) );
 a64374a <=( A199  and  a64373a );
 a64375a <=( a64374a  and  a64369a );
 a64379a <=( A267  and  A266 );
 a64380a <=( (not A203)  and  a64379a );
 a64383a <=( (not A299)  and  A298 );
 a64386a <=( (not A302)  and  (not A300) );
 a64387a <=( a64386a  and  a64383a );
 a64388a <=( a64387a  and  a64380a );
 a64392a <=( (not A167)  and  (not A169) );
 a64393a <=( (not A170)  and  a64392a );
 a64397a <=( (not A201)  and  (not A200) );
 a64398a <=( A199  and  a64397a );
 a64399a <=( a64398a  and  a64393a );
 a64403a <=( A267  and  A266 );
 a64404a <=( (not A203)  and  a64403a );
 a64407a <=( A299  and  (not A298) );
 a64410a <=( A301  and  (not A300) );
 a64411a <=( a64410a  and  a64407a );
 a64412a <=( a64411a  and  a64404a );
 a64416a <=( (not A167)  and  (not A169) );
 a64417a <=( (not A170)  and  a64416a );
 a64421a <=( (not A201)  and  (not A200) );
 a64422a <=( A199  and  a64421a );
 a64423a <=( a64422a  and  a64417a );
 a64427a <=( A267  and  A266 );
 a64428a <=( (not A203)  and  a64427a );
 a64431a <=( A299  and  (not A298) );
 a64434a <=( (not A302)  and  (not A300) );
 a64435a <=( a64434a  and  a64431a );
 a64436a <=( a64435a  and  a64428a );
 a64440a <=( (not A167)  and  (not A169) );
 a64441a <=( (not A170)  and  a64440a );
 a64445a <=( (not A202)  and  (not A200) );
 a64446a <=( (not A199)  and  a64445a );
 a64447a <=( a64446a  and  a64441a );
 a64451a <=( A268  and  A266 );
 a64452a <=( A265  and  a64451a );
 a64455a <=( (not A298)  and  (not A269) );
 a64458a <=( (not A301)  and  (not A299) );
 a64459a <=( a64458a  and  a64455a );
 a64460a <=( a64459a  and  a64452a );
 a64464a <=( (not A167)  and  (not A169) );
 a64465a <=( (not A170)  and  a64464a );
 a64469a <=( (not A202)  and  (not A200) );
 a64470a <=( (not A199)  and  a64469a );
 a64471a <=( a64470a  and  a64465a );
 a64475a <=( A268  and  A266 );
 a64476a <=( A265  and  a64475a );
 a64479a <=( (not A298)  and  (not A269) );
 a64482a <=( A302  and  (not A299) );
 a64483a <=( a64482a  and  a64479a );
 a64484a <=( a64483a  and  a64476a );
 a64488a <=( (not A167)  and  (not A169) );
 a64489a <=( (not A170)  and  a64488a );
 a64493a <=( (not A202)  and  (not A200) );
 a64494a <=( (not A199)  and  a64493a );
 a64495a <=( a64494a  and  a64489a );
 a64499a <=( (not A268)  and  A266 );
 a64500a <=( (not A265)  and  a64499a );
 a64503a <=( (not A298)  and  A269 );
 a64506a <=( (not A301)  and  (not A299) );
 a64507a <=( a64506a  and  a64503a );
 a64508a <=( a64507a  and  a64500a );
 a64512a <=( (not A167)  and  (not A169) );
 a64513a <=( (not A170)  and  a64512a );
 a64517a <=( (not A202)  and  (not A200) );
 a64518a <=( (not A199)  and  a64517a );
 a64519a <=( a64518a  and  a64513a );
 a64523a <=( (not A268)  and  A266 );
 a64524a <=( (not A265)  and  a64523a );
 a64527a <=( (not A298)  and  A269 );
 a64530a <=( A302  and  (not A299) );
 a64531a <=( a64530a  and  a64527a );
 a64532a <=( a64531a  and  a64524a );
 a64536a <=( (not A167)  and  (not A169) );
 a64537a <=( (not A170)  and  a64536a );
 a64541a <=( (not A202)  and  (not A200) );
 a64542a <=( (not A199)  and  a64541a );
 a64543a <=( a64542a  and  a64537a );
 a64547a <=( (not A268)  and  (not A266) );
 a64548a <=( A265  and  a64547a );
 a64551a <=( (not A298)  and  A269 );
 a64554a <=( (not A301)  and  (not A299) );
 a64555a <=( a64554a  and  a64551a );
 a64556a <=( a64555a  and  a64548a );
 a64560a <=( (not A167)  and  (not A169) );
 a64561a <=( (not A170)  and  a64560a );
 a64565a <=( (not A202)  and  (not A200) );
 a64566a <=( (not A199)  and  a64565a );
 a64567a <=( a64566a  and  a64561a );
 a64571a <=( (not A268)  and  (not A266) );
 a64572a <=( A265  and  a64571a );
 a64575a <=( (not A298)  and  A269 );
 a64578a <=( A302  and  (not A299) );
 a64579a <=( a64578a  and  a64575a );
 a64580a <=( a64579a  and  a64572a );
 a64584a <=( (not A167)  and  (not A169) );
 a64585a <=( (not A170)  and  a64584a );
 a64589a <=( (not A202)  and  (not A200) );
 a64590a <=( (not A199)  and  a64589a );
 a64591a <=( a64590a  and  a64585a );
 a64595a <=( A268  and  (not A266) );
 a64596a <=( (not A265)  and  a64595a );
 a64599a <=( (not A298)  and  (not A269) );
 a64602a <=( (not A301)  and  (not A299) );
 a64603a <=( a64602a  and  a64599a );
 a64604a <=( a64603a  and  a64596a );
 a64608a <=( (not A167)  and  (not A169) );
 a64609a <=( (not A170)  and  a64608a );
 a64613a <=( (not A202)  and  (not A200) );
 a64614a <=( (not A199)  and  a64613a );
 a64615a <=( a64614a  and  a64609a );
 a64619a <=( A268  and  (not A266) );
 a64620a <=( (not A265)  and  a64619a );
 a64623a <=( (not A298)  and  (not A269) );
 a64626a <=( A302  and  (not A299) );
 a64627a <=( a64626a  and  a64623a );
 a64628a <=( a64627a  and  a64620a );
 a64632a <=( (not A167)  and  (not A169) );
 a64633a <=( (not A170)  and  a64632a );
 a64637a <=( A203  and  (not A200) );
 a64638a <=( (not A199)  and  a64637a );
 a64639a <=( a64638a  and  a64633a );
 a64643a <=( A268  and  A266 );
 a64644a <=( A265  and  a64643a );
 a64647a <=( (not A298)  and  (not A269) );
 a64650a <=( (not A301)  and  (not A299) );
 a64651a <=( a64650a  and  a64647a );
 a64652a <=( a64651a  and  a64644a );
 a64656a <=( (not A167)  and  (not A169) );
 a64657a <=( (not A170)  and  a64656a );
 a64661a <=( A203  and  (not A200) );
 a64662a <=( (not A199)  and  a64661a );
 a64663a <=( a64662a  and  a64657a );
 a64667a <=( A268  and  A266 );
 a64668a <=( A265  and  a64667a );
 a64671a <=( (not A298)  and  (not A269) );
 a64674a <=( A302  and  (not A299) );
 a64675a <=( a64674a  and  a64671a );
 a64676a <=( a64675a  and  a64668a );
 a64680a <=( (not A167)  and  (not A169) );
 a64681a <=( (not A170)  and  a64680a );
 a64685a <=( A203  and  (not A200) );
 a64686a <=( (not A199)  and  a64685a );
 a64687a <=( a64686a  and  a64681a );
 a64691a <=( (not A268)  and  A266 );
 a64692a <=( (not A265)  and  a64691a );
 a64695a <=( (not A298)  and  A269 );
 a64698a <=( (not A301)  and  (not A299) );
 a64699a <=( a64698a  and  a64695a );
 a64700a <=( a64699a  and  a64692a );
 a64704a <=( (not A167)  and  (not A169) );
 a64705a <=( (not A170)  and  a64704a );
 a64709a <=( A203  and  (not A200) );
 a64710a <=( (not A199)  and  a64709a );
 a64711a <=( a64710a  and  a64705a );
 a64715a <=( (not A268)  and  A266 );
 a64716a <=( (not A265)  and  a64715a );
 a64719a <=( (not A298)  and  A269 );
 a64722a <=( A302  and  (not A299) );
 a64723a <=( a64722a  and  a64719a );
 a64724a <=( a64723a  and  a64716a );
 a64728a <=( (not A167)  and  (not A169) );
 a64729a <=( (not A170)  and  a64728a );
 a64733a <=( A203  and  (not A200) );
 a64734a <=( (not A199)  and  a64733a );
 a64735a <=( a64734a  and  a64729a );
 a64739a <=( (not A268)  and  (not A266) );
 a64740a <=( A265  and  a64739a );
 a64743a <=( (not A298)  and  A269 );
 a64746a <=( (not A301)  and  (not A299) );
 a64747a <=( a64746a  and  a64743a );
 a64748a <=( a64747a  and  a64740a );
 a64752a <=( (not A167)  and  (not A169) );
 a64753a <=( (not A170)  and  a64752a );
 a64757a <=( A203  and  (not A200) );
 a64758a <=( (not A199)  and  a64757a );
 a64759a <=( a64758a  and  a64753a );
 a64763a <=( (not A268)  and  (not A266) );
 a64764a <=( A265  and  a64763a );
 a64767a <=( (not A298)  and  A269 );
 a64770a <=( A302  and  (not A299) );
 a64771a <=( a64770a  and  a64767a );
 a64772a <=( a64771a  and  a64764a );
 a64776a <=( (not A167)  and  (not A169) );
 a64777a <=( (not A170)  and  a64776a );
 a64781a <=( A203  and  (not A200) );
 a64782a <=( (not A199)  and  a64781a );
 a64783a <=( a64782a  and  a64777a );
 a64787a <=( A268  and  (not A266) );
 a64788a <=( (not A265)  and  a64787a );
 a64791a <=( (not A298)  and  (not A269) );
 a64794a <=( (not A301)  and  (not A299) );
 a64795a <=( a64794a  and  a64791a );
 a64796a <=( a64795a  and  a64788a );
 a64800a <=( (not A167)  and  (not A169) );
 a64801a <=( (not A170)  and  a64800a );
 a64805a <=( A203  and  (not A200) );
 a64806a <=( (not A199)  and  a64805a );
 a64807a <=( a64806a  and  a64801a );
 a64811a <=( A268  and  (not A266) );
 a64812a <=( (not A265)  and  a64811a );
 a64815a <=( (not A298)  and  (not A269) );
 a64818a <=( A302  and  (not A299) );
 a64819a <=( a64818a  and  a64815a );
 a64820a <=( a64819a  and  a64812a );
 a64824a <=( (not A167)  and  (not A169) );
 a64825a <=( (not A170)  and  a64824a );
 a64829a <=( A202  and  (not A200) );
 a64830a <=( (not A199)  and  a64829a );
 a64831a <=( a64830a  and  a64825a );
 a64835a <=( A266  and  A265 );
 a64836a <=( (not A203)  and  a64835a );
 a64839a <=( (not A268)  and  (not A267) );
 a64842a <=( A300  and  A299 );
 a64843a <=( a64842a  and  a64839a );
 a64844a <=( a64843a  and  a64836a );
 a64848a <=( (not A167)  and  (not A169) );
 a64849a <=( (not A170)  and  a64848a );
 a64853a <=( A202  and  (not A200) );
 a64854a <=( (not A199)  and  a64853a );
 a64855a <=( a64854a  and  a64849a );
 a64859a <=( A266  and  A265 );
 a64860a <=( (not A203)  and  a64859a );
 a64863a <=( (not A268)  and  (not A267) );
 a64866a <=( A300  and  A298 );
 a64867a <=( a64866a  and  a64863a );
 a64868a <=( a64867a  and  a64860a );
 a64872a <=( (not A167)  and  (not A169) );
 a64873a <=( (not A170)  and  a64872a );
 a64877a <=( A202  and  (not A200) );
 a64878a <=( (not A199)  and  a64877a );
 a64879a <=( a64878a  and  a64873a );
 a64883a <=( A266  and  A265 );
 a64884a <=( (not A203)  and  a64883a );
 a64887a <=( A269  and  (not A267) );
 a64890a <=( A300  and  A299 );
 a64891a <=( a64890a  and  a64887a );
 a64892a <=( a64891a  and  a64884a );
 a64896a <=( (not A167)  and  (not A169) );
 a64897a <=( (not A170)  and  a64896a );
 a64901a <=( A202  and  (not A200) );
 a64902a <=( (not A199)  and  a64901a );
 a64903a <=( a64902a  and  a64897a );
 a64907a <=( A266  and  A265 );
 a64908a <=( (not A203)  and  a64907a );
 a64911a <=( A269  and  (not A267) );
 a64914a <=( A300  and  A298 );
 a64915a <=( a64914a  and  a64911a );
 a64916a <=( a64915a  and  a64908a );
 a64920a <=( (not A167)  and  (not A169) );
 a64921a <=( (not A170)  and  a64920a );
 a64925a <=( A202  and  (not A200) );
 a64926a <=( (not A199)  and  a64925a );
 a64927a <=( a64926a  and  a64921a );
 a64931a <=( A266  and  (not A265) );
 a64932a <=( (not A203)  and  a64931a );
 a64935a <=( A268  and  (not A267) );
 a64938a <=( A300  and  A299 );
 a64939a <=( a64938a  and  a64935a );
 a64940a <=( a64939a  and  a64932a );
 a64944a <=( (not A167)  and  (not A169) );
 a64945a <=( (not A170)  and  a64944a );
 a64949a <=( A202  and  (not A200) );
 a64950a <=( (not A199)  and  a64949a );
 a64951a <=( a64950a  and  a64945a );
 a64955a <=( A266  and  (not A265) );
 a64956a <=( (not A203)  and  a64955a );
 a64959a <=( A268  and  (not A267) );
 a64962a <=( A300  and  A298 );
 a64963a <=( a64962a  and  a64959a );
 a64964a <=( a64963a  and  a64956a );
 a64968a <=( (not A167)  and  (not A169) );
 a64969a <=( (not A170)  and  a64968a );
 a64973a <=( A202  and  (not A200) );
 a64974a <=( (not A199)  and  a64973a );
 a64975a <=( a64974a  and  a64969a );
 a64979a <=( A266  and  (not A265) );
 a64980a <=( (not A203)  and  a64979a );
 a64983a <=( (not A269)  and  (not A267) );
 a64986a <=( A300  and  A299 );
 a64987a <=( a64986a  and  a64983a );
 a64988a <=( a64987a  and  a64980a );
 a64992a <=( (not A167)  and  (not A169) );
 a64993a <=( (not A170)  and  a64992a );
 a64997a <=( A202  and  (not A200) );
 a64998a <=( (not A199)  and  a64997a );
 a64999a <=( a64998a  and  a64993a );
 a65003a <=( A266  and  (not A265) );
 a65004a <=( (not A203)  and  a65003a );
 a65007a <=( (not A269)  and  (not A267) );
 a65010a <=( A300  and  A298 );
 a65011a <=( a65010a  and  a65007a );
 a65012a <=( a65011a  and  a65004a );
 a65016a <=( (not A167)  and  (not A169) );
 a65017a <=( (not A170)  and  a65016a );
 a65021a <=( A202  and  (not A200) );
 a65022a <=( (not A199)  and  a65021a );
 a65023a <=( a65022a  and  a65017a );
 a65027a <=( (not A266)  and  A265 );
 a65028a <=( (not A203)  and  a65027a );
 a65031a <=( A268  and  (not A267) );
 a65034a <=( A300  and  A299 );
 a65035a <=( a65034a  and  a65031a );
 a65036a <=( a65035a  and  a65028a );
 a65040a <=( (not A167)  and  (not A169) );
 a65041a <=( (not A170)  and  a65040a );
 a65045a <=( A202  and  (not A200) );
 a65046a <=( (not A199)  and  a65045a );
 a65047a <=( a65046a  and  a65041a );
 a65051a <=( (not A266)  and  A265 );
 a65052a <=( (not A203)  and  a65051a );
 a65055a <=( A268  and  (not A267) );
 a65058a <=( A300  and  A298 );
 a65059a <=( a65058a  and  a65055a );
 a65060a <=( a65059a  and  a65052a );
 a65064a <=( (not A167)  and  (not A169) );
 a65065a <=( (not A170)  and  a65064a );
 a65069a <=( A202  and  (not A200) );
 a65070a <=( (not A199)  and  a65069a );
 a65071a <=( a65070a  and  a65065a );
 a65075a <=( (not A266)  and  A265 );
 a65076a <=( (not A203)  and  a65075a );
 a65079a <=( (not A269)  and  (not A267) );
 a65082a <=( A300  and  A299 );
 a65083a <=( a65082a  and  a65079a );
 a65084a <=( a65083a  and  a65076a );
 a65088a <=( (not A167)  and  (not A169) );
 a65089a <=( (not A170)  and  a65088a );
 a65093a <=( A202  and  (not A200) );
 a65094a <=( (not A199)  and  a65093a );
 a65095a <=( a65094a  and  a65089a );
 a65099a <=( (not A266)  and  A265 );
 a65100a <=( (not A203)  and  a65099a );
 a65103a <=( (not A269)  and  (not A267) );
 a65106a <=( A300  and  A298 );
 a65107a <=( a65106a  and  a65103a );
 a65108a <=( a65107a  and  a65100a );
 a65112a <=( A199  and  A166 );
 a65113a <=( A167  and  a65112a );
 a65116a <=( A202  and  A200 );
 a65119a <=( A265  and  (not A203) );
 a65120a <=( a65119a  and  a65116a );
 a65121a <=( a65120a  and  a65113a );
 a65125a <=( (not A268)  and  (not A267) );
 a65126a <=( A266  and  a65125a );
 a65129a <=( A299  and  A298 );
 a65132a <=( (not A302)  and  A301 );
 a65133a <=( a65132a  and  a65129a );
 a65134a <=( a65133a  and  a65126a );
 a65138a <=( A199  and  A166 );
 a65139a <=( A167  and  a65138a );
 a65142a <=( A202  and  A200 );
 a65145a <=( A265  and  (not A203) );
 a65146a <=( a65145a  and  a65142a );
 a65147a <=( a65146a  and  a65139a );
 a65151a <=( (not A268)  and  (not A267) );
 a65152a <=( A266  and  a65151a );
 a65155a <=( (not A299)  and  A298 );
 a65158a <=( A302  and  (not A301) );
 a65159a <=( a65158a  and  a65155a );
 a65160a <=( a65159a  and  a65152a );
 a65164a <=( A199  and  A166 );
 a65165a <=( A167  and  a65164a );
 a65168a <=( A202  and  A200 );
 a65171a <=( A265  and  (not A203) );
 a65172a <=( a65171a  and  a65168a );
 a65173a <=( a65172a  and  a65165a );
 a65177a <=( (not A268)  and  (not A267) );
 a65178a <=( A266  and  a65177a );
 a65181a <=( A299  and  (not A298) );
 a65184a <=( A302  and  (not A301) );
 a65185a <=( a65184a  and  a65181a );
 a65186a <=( a65185a  and  a65178a );
 a65190a <=( A199  and  A166 );
 a65191a <=( A167  and  a65190a );
 a65194a <=( A202  and  A200 );
 a65197a <=( A265  and  (not A203) );
 a65198a <=( a65197a  and  a65194a );
 a65199a <=( a65198a  and  a65191a );
 a65203a <=( (not A268)  and  (not A267) );
 a65204a <=( A266  and  a65203a );
 a65207a <=( (not A299)  and  (not A298) );
 a65210a <=( (not A302)  and  A301 );
 a65211a <=( a65210a  and  a65207a );
 a65212a <=( a65211a  and  a65204a );
 a65216a <=( A199  and  A166 );
 a65217a <=( A167  and  a65216a );
 a65220a <=( A202  and  A200 );
 a65223a <=( A265  and  (not A203) );
 a65224a <=( a65223a  and  a65220a );
 a65225a <=( a65224a  and  a65217a );
 a65229a <=( A269  and  (not A267) );
 a65230a <=( A266  and  a65229a );
 a65233a <=( A299  and  A298 );
 a65236a <=( (not A302)  and  A301 );
 a65237a <=( a65236a  and  a65233a );
 a65238a <=( a65237a  and  a65230a );
 a65242a <=( A199  and  A166 );
 a65243a <=( A167  and  a65242a );
 a65246a <=( A202  and  A200 );
 a65249a <=( A265  and  (not A203) );
 a65250a <=( a65249a  and  a65246a );
 a65251a <=( a65250a  and  a65243a );
 a65255a <=( A269  and  (not A267) );
 a65256a <=( A266  and  a65255a );
 a65259a <=( (not A299)  and  A298 );
 a65262a <=( A302  and  (not A301) );
 a65263a <=( a65262a  and  a65259a );
 a65264a <=( a65263a  and  a65256a );
 a65268a <=( A199  and  A166 );
 a65269a <=( A167  and  a65268a );
 a65272a <=( A202  and  A200 );
 a65275a <=( A265  and  (not A203) );
 a65276a <=( a65275a  and  a65272a );
 a65277a <=( a65276a  and  a65269a );
 a65281a <=( A269  and  (not A267) );
 a65282a <=( A266  and  a65281a );
 a65285a <=( A299  and  (not A298) );
 a65288a <=( A302  and  (not A301) );
 a65289a <=( a65288a  and  a65285a );
 a65290a <=( a65289a  and  a65282a );
 a65294a <=( A199  and  A166 );
 a65295a <=( A167  and  a65294a );
 a65298a <=( A202  and  A200 );
 a65301a <=( A265  and  (not A203) );
 a65302a <=( a65301a  and  a65298a );
 a65303a <=( a65302a  and  a65295a );
 a65307a <=( A269  and  (not A267) );
 a65308a <=( A266  and  a65307a );
 a65311a <=( (not A299)  and  (not A298) );
 a65314a <=( (not A302)  and  A301 );
 a65315a <=( a65314a  and  a65311a );
 a65316a <=( a65315a  and  a65308a );
 a65320a <=( A199  and  A166 );
 a65321a <=( A167  and  a65320a );
 a65324a <=( A202  and  A200 );
 a65327a <=( (not A265)  and  (not A203) );
 a65328a <=( a65327a  and  a65324a );
 a65329a <=( a65328a  and  a65321a );
 a65333a <=( A268  and  (not A267) );
 a65334a <=( A266  and  a65333a );
 a65337a <=( A299  and  A298 );
 a65340a <=( (not A302)  and  A301 );
 a65341a <=( a65340a  and  a65337a );
 a65342a <=( a65341a  and  a65334a );
 a65346a <=( A199  and  A166 );
 a65347a <=( A167  and  a65346a );
 a65350a <=( A202  and  A200 );
 a65353a <=( (not A265)  and  (not A203) );
 a65354a <=( a65353a  and  a65350a );
 a65355a <=( a65354a  and  a65347a );
 a65359a <=( A268  and  (not A267) );
 a65360a <=( A266  and  a65359a );
 a65363a <=( (not A299)  and  A298 );
 a65366a <=( A302  and  (not A301) );
 a65367a <=( a65366a  and  a65363a );
 a65368a <=( a65367a  and  a65360a );
 a65372a <=( A199  and  A166 );
 a65373a <=( A167  and  a65372a );
 a65376a <=( A202  and  A200 );
 a65379a <=( (not A265)  and  (not A203) );
 a65380a <=( a65379a  and  a65376a );
 a65381a <=( a65380a  and  a65373a );
 a65385a <=( A268  and  (not A267) );
 a65386a <=( A266  and  a65385a );
 a65389a <=( A299  and  (not A298) );
 a65392a <=( A302  and  (not A301) );
 a65393a <=( a65392a  and  a65389a );
 a65394a <=( a65393a  and  a65386a );
 a65398a <=( A199  and  A166 );
 a65399a <=( A167  and  a65398a );
 a65402a <=( A202  and  A200 );
 a65405a <=( (not A265)  and  (not A203) );
 a65406a <=( a65405a  and  a65402a );
 a65407a <=( a65406a  and  a65399a );
 a65411a <=( A268  and  (not A267) );
 a65412a <=( A266  and  a65411a );
 a65415a <=( (not A299)  and  (not A298) );
 a65418a <=( (not A302)  and  A301 );
 a65419a <=( a65418a  and  a65415a );
 a65420a <=( a65419a  and  a65412a );
 a65424a <=( A199  and  A166 );
 a65425a <=( A167  and  a65424a );
 a65428a <=( A202  and  A200 );
 a65431a <=( (not A265)  and  (not A203) );
 a65432a <=( a65431a  and  a65428a );
 a65433a <=( a65432a  and  a65425a );
 a65437a <=( (not A269)  and  (not A267) );
 a65438a <=( A266  and  a65437a );
 a65441a <=( A299  and  A298 );
 a65444a <=( (not A302)  and  A301 );
 a65445a <=( a65444a  and  a65441a );
 a65446a <=( a65445a  and  a65438a );
 a65450a <=( A199  and  A166 );
 a65451a <=( A167  and  a65450a );
 a65454a <=( A202  and  A200 );
 a65457a <=( (not A265)  and  (not A203) );
 a65458a <=( a65457a  and  a65454a );
 a65459a <=( a65458a  and  a65451a );
 a65463a <=( (not A269)  and  (not A267) );
 a65464a <=( A266  and  a65463a );
 a65467a <=( (not A299)  and  A298 );
 a65470a <=( A302  and  (not A301) );
 a65471a <=( a65470a  and  a65467a );
 a65472a <=( a65471a  and  a65464a );
 a65476a <=( A199  and  A166 );
 a65477a <=( A167  and  a65476a );
 a65480a <=( A202  and  A200 );
 a65483a <=( (not A265)  and  (not A203) );
 a65484a <=( a65483a  and  a65480a );
 a65485a <=( a65484a  and  a65477a );
 a65489a <=( (not A269)  and  (not A267) );
 a65490a <=( A266  and  a65489a );
 a65493a <=( A299  and  (not A298) );
 a65496a <=( A302  and  (not A301) );
 a65497a <=( a65496a  and  a65493a );
 a65498a <=( a65497a  and  a65490a );
 a65502a <=( A199  and  A166 );
 a65503a <=( A167  and  a65502a );
 a65506a <=( A202  and  A200 );
 a65509a <=( (not A265)  and  (not A203) );
 a65510a <=( a65509a  and  a65506a );
 a65511a <=( a65510a  and  a65503a );
 a65515a <=( (not A269)  and  (not A267) );
 a65516a <=( A266  and  a65515a );
 a65519a <=( (not A299)  and  (not A298) );
 a65522a <=( (not A302)  and  A301 );
 a65523a <=( a65522a  and  a65519a );
 a65524a <=( a65523a  and  a65516a );
 a65528a <=( A199  and  A166 );
 a65529a <=( A167  and  a65528a );
 a65532a <=( A202  and  A200 );
 a65535a <=( A265  and  (not A203) );
 a65536a <=( a65535a  and  a65532a );
 a65537a <=( a65536a  and  a65529a );
 a65541a <=( A268  and  (not A267) );
 a65542a <=( (not A266)  and  a65541a );
 a65545a <=( A299  and  A298 );
 a65548a <=( (not A302)  and  A301 );
 a65549a <=( a65548a  and  a65545a );
 a65550a <=( a65549a  and  a65542a );
 a65554a <=( A199  and  A166 );
 a65555a <=( A167  and  a65554a );
 a65558a <=( A202  and  A200 );
 a65561a <=( A265  and  (not A203) );
 a65562a <=( a65561a  and  a65558a );
 a65563a <=( a65562a  and  a65555a );
 a65567a <=( A268  and  (not A267) );
 a65568a <=( (not A266)  and  a65567a );
 a65571a <=( (not A299)  and  A298 );
 a65574a <=( A302  and  (not A301) );
 a65575a <=( a65574a  and  a65571a );
 a65576a <=( a65575a  and  a65568a );
 a65580a <=( A199  and  A166 );
 a65581a <=( A167  and  a65580a );
 a65584a <=( A202  and  A200 );
 a65587a <=( A265  and  (not A203) );
 a65588a <=( a65587a  and  a65584a );
 a65589a <=( a65588a  and  a65581a );
 a65593a <=( A268  and  (not A267) );
 a65594a <=( (not A266)  and  a65593a );
 a65597a <=( A299  and  (not A298) );
 a65600a <=( A302  and  (not A301) );
 a65601a <=( a65600a  and  a65597a );
 a65602a <=( a65601a  and  a65594a );
 a65606a <=( A199  and  A166 );
 a65607a <=( A167  and  a65606a );
 a65610a <=( A202  and  A200 );
 a65613a <=( A265  and  (not A203) );
 a65614a <=( a65613a  and  a65610a );
 a65615a <=( a65614a  and  a65607a );
 a65619a <=( A268  and  (not A267) );
 a65620a <=( (not A266)  and  a65619a );
 a65623a <=( (not A299)  and  (not A298) );
 a65626a <=( (not A302)  and  A301 );
 a65627a <=( a65626a  and  a65623a );
 a65628a <=( a65627a  and  a65620a );
 a65632a <=( A199  and  A166 );
 a65633a <=( A167  and  a65632a );
 a65636a <=( A202  and  A200 );
 a65639a <=( A265  and  (not A203) );
 a65640a <=( a65639a  and  a65636a );
 a65641a <=( a65640a  and  a65633a );
 a65645a <=( (not A269)  and  (not A267) );
 a65646a <=( (not A266)  and  a65645a );
 a65649a <=( A299  and  A298 );
 a65652a <=( (not A302)  and  A301 );
 a65653a <=( a65652a  and  a65649a );
 a65654a <=( a65653a  and  a65646a );
 a65658a <=( A199  and  A166 );
 a65659a <=( A167  and  a65658a );
 a65662a <=( A202  and  A200 );
 a65665a <=( A265  and  (not A203) );
 a65666a <=( a65665a  and  a65662a );
 a65667a <=( a65666a  and  a65659a );
 a65671a <=( (not A269)  and  (not A267) );
 a65672a <=( (not A266)  and  a65671a );
 a65675a <=( (not A299)  and  A298 );
 a65678a <=( A302  and  (not A301) );
 a65679a <=( a65678a  and  a65675a );
 a65680a <=( a65679a  and  a65672a );
 a65684a <=( A199  and  A166 );
 a65685a <=( A167  and  a65684a );
 a65688a <=( A202  and  A200 );
 a65691a <=( A265  and  (not A203) );
 a65692a <=( a65691a  and  a65688a );
 a65693a <=( a65692a  and  a65685a );
 a65697a <=( (not A269)  and  (not A267) );
 a65698a <=( (not A266)  and  a65697a );
 a65701a <=( A299  and  (not A298) );
 a65704a <=( A302  and  (not A301) );
 a65705a <=( a65704a  and  a65701a );
 a65706a <=( a65705a  and  a65698a );
 a65710a <=( A199  and  A166 );
 a65711a <=( A167  and  a65710a );
 a65714a <=( A202  and  A200 );
 a65717a <=( A265  and  (not A203) );
 a65718a <=( a65717a  and  a65714a );
 a65719a <=( a65718a  and  a65711a );
 a65723a <=( (not A269)  and  (not A267) );
 a65724a <=( (not A266)  and  a65723a );
 a65727a <=( (not A299)  and  (not A298) );
 a65730a <=( (not A302)  and  A301 );
 a65731a <=( a65730a  and  a65727a );
 a65732a <=( a65731a  and  a65724a );
 a65736a <=( A199  and  A166 );
 a65737a <=( A167  and  a65736a );
 a65740a <=( (not A201)  and  A200 );
 a65743a <=( A265  and  (not A202) );
 a65744a <=( a65743a  and  a65740a );
 a65745a <=( a65744a  and  a65737a );
 a65749a <=( (not A269)  and  A268 );
 a65750a <=( A266  and  a65749a );
 a65753a <=( A299  and  A298 );
 a65756a <=( (not A301)  and  (not A300) );
 a65757a <=( a65756a  and  a65753a );
 a65758a <=( a65757a  and  a65750a );
 a65762a <=( A199  and  A166 );
 a65763a <=( A167  and  a65762a );
 a65766a <=( (not A201)  and  A200 );
 a65769a <=( A265  and  (not A202) );
 a65770a <=( a65769a  and  a65766a );
 a65771a <=( a65770a  and  a65763a );
 a65775a <=( (not A269)  and  A268 );
 a65776a <=( A266  and  a65775a );
 a65779a <=( A299  and  A298 );
 a65782a <=( A302  and  (not A300) );
 a65783a <=( a65782a  and  a65779a );
 a65784a <=( a65783a  and  a65776a );
 a65788a <=( A199  and  A166 );
 a65789a <=( A167  and  a65788a );
 a65792a <=( (not A201)  and  A200 );
 a65795a <=( A265  and  (not A202) );
 a65796a <=( a65795a  and  a65792a );
 a65797a <=( a65796a  and  a65789a );
 a65801a <=( (not A269)  and  A268 );
 a65802a <=( A266  and  a65801a );
 a65805a <=( (not A299)  and  A298 );
 a65808a <=( A301  and  (not A300) );
 a65809a <=( a65808a  and  a65805a );
 a65810a <=( a65809a  and  a65802a );
 a65814a <=( A199  and  A166 );
 a65815a <=( A167  and  a65814a );
 a65818a <=( (not A201)  and  A200 );
 a65821a <=( A265  and  (not A202) );
 a65822a <=( a65821a  and  a65818a );
 a65823a <=( a65822a  and  a65815a );
 a65827a <=( (not A269)  and  A268 );
 a65828a <=( A266  and  a65827a );
 a65831a <=( (not A299)  and  A298 );
 a65834a <=( (not A302)  and  (not A300) );
 a65835a <=( a65834a  and  a65831a );
 a65836a <=( a65835a  and  a65828a );
 a65840a <=( A199  and  A166 );
 a65841a <=( A167  and  a65840a );
 a65844a <=( (not A201)  and  A200 );
 a65847a <=( A265  and  (not A202) );
 a65848a <=( a65847a  and  a65844a );
 a65849a <=( a65848a  and  a65841a );
 a65853a <=( (not A269)  and  A268 );
 a65854a <=( A266  and  a65853a );
 a65857a <=( A299  and  (not A298) );
 a65860a <=( A301  and  (not A300) );
 a65861a <=( a65860a  and  a65857a );
 a65862a <=( a65861a  and  a65854a );
 a65866a <=( A199  and  A166 );
 a65867a <=( A167  and  a65866a );
 a65870a <=( (not A201)  and  A200 );
 a65873a <=( A265  and  (not A202) );
 a65874a <=( a65873a  and  a65870a );
 a65875a <=( a65874a  and  a65867a );
 a65879a <=( (not A269)  and  A268 );
 a65880a <=( A266  and  a65879a );
 a65883a <=( A299  and  (not A298) );
 a65886a <=( (not A302)  and  (not A300) );
 a65887a <=( a65886a  and  a65883a );
 a65888a <=( a65887a  and  a65880a );
 a65892a <=( A199  and  A166 );
 a65893a <=( A167  and  a65892a );
 a65896a <=( (not A201)  and  A200 );
 a65899a <=( (not A265)  and  (not A202) );
 a65900a <=( a65899a  and  a65896a );
 a65901a <=( a65900a  and  a65893a );
 a65905a <=( A269  and  (not A268) );
 a65906a <=( A266  and  a65905a );
 a65909a <=( A299  and  A298 );
 a65912a <=( (not A301)  and  (not A300) );
 a65913a <=( a65912a  and  a65909a );
 a65914a <=( a65913a  and  a65906a );
 a65918a <=( A199  and  A166 );
 a65919a <=( A167  and  a65918a );
 a65922a <=( (not A201)  and  A200 );
 a65925a <=( (not A265)  and  (not A202) );
 a65926a <=( a65925a  and  a65922a );
 a65927a <=( a65926a  and  a65919a );
 a65931a <=( A269  and  (not A268) );
 a65932a <=( A266  and  a65931a );
 a65935a <=( A299  and  A298 );
 a65938a <=( A302  and  (not A300) );
 a65939a <=( a65938a  and  a65935a );
 a65940a <=( a65939a  and  a65932a );
 a65944a <=( A199  and  A166 );
 a65945a <=( A167  and  a65944a );
 a65948a <=( (not A201)  and  A200 );
 a65951a <=( (not A265)  and  (not A202) );
 a65952a <=( a65951a  and  a65948a );
 a65953a <=( a65952a  and  a65945a );
 a65957a <=( A269  and  (not A268) );
 a65958a <=( A266  and  a65957a );
 a65961a <=( (not A299)  and  A298 );
 a65964a <=( A301  and  (not A300) );
 a65965a <=( a65964a  and  a65961a );
 a65966a <=( a65965a  and  a65958a );
 a65970a <=( A199  and  A166 );
 a65971a <=( A167  and  a65970a );
 a65974a <=( (not A201)  and  A200 );
 a65977a <=( (not A265)  and  (not A202) );
 a65978a <=( a65977a  and  a65974a );
 a65979a <=( a65978a  and  a65971a );
 a65983a <=( A269  and  (not A268) );
 a65984a <=( A266  and  a65983a );
 a65987a <=( (not A299)  and  A298 );
 a65990a <=( (not A302)  and  (not A300) );
 a65991a <=( a65990a  and  a65987a );
 a65992a <=( a65991a  and  a65984a );
 a65996a <=( A199  and  A166 );
 a65997a <=( A167  and  a65996a );
 a66000a <=( (not A201)  and  A200 );
 a66003a <=( (not A265)  and  (not A202) );
 a66004a <=( a66003a  and  a66000a );
 a66005a <=( a66004a  and  a65997a );
 a66009a <=( A269  and  (not A268) );
 a66010a <=( A266  and  a66009a );
 a66013a <=( A299  and  (not A298) );
 a66016a <=( A301  and  (not A300) );
 a66017a <=( a66016a  and  a66013a );
 a66018a <=( a66017a  and  a66010a );
 a66022a <=( A199  and  A166 );
 a66023a <=( A167  and  a66022a );
 a66026a <=( (not A201)  and  A200 );
 a66029a <=( (not A265)  and  (not A202) );
 a66030a <=( a66029a  and  a66026a );
 a66031a <=( a66030a  and  a66023a );
 a66035a <=( A269  and  (not A268) );
 a66036a <=( A266  and  a66035a );
 a66039a <=( A299  and  (not A298) );
 a66042a <=( (not A302)  and  (not A300) );
 a66043a <=( a66042a  and  a66039a );
 a66044a <=( a66043a  and  a66036a );
 a66048a <=( A199  and  A166 );
 a66049a <=( A167  and  a66048a );
 a66052a <=( (not A201)  and  A200 );
 a66055a <=( A265  and  (not A202) );
 a66056a <=( a66055a  and  a66052a );
 a66057a <=( a66056a  and  a66049a );
 a66061a <=( A269  and  (not A268) );
 a66062a <=( (not A266)  and  a66061a );
 a66065a <=( A299  and  A298 );
 a66068a <=( (not A301)  and  (not A300) );
 a66069a <=( a66068a  and  a66065a );
 a66070a <=( a66069a  and  a66062a );
 a66074a <=( A199  and  A166 );
 a66075a <=( A167  and  a66074a );
 a66078a <=( (not A201)  and  A200 );
 a66081a <=( A265  and  (not A202) );
 a66082a <=( a66081a  and  a66078a );
 a66083a <=( a66082a  and  a66075a );
 a66087a <=( A269  and  (not A268) );
 a66088a <=( (not A266)  and  a66087a );
 a66091a <=( A299  and  A298 );
 a66094a <=( A302  and  (not A300) );
 a66095a <=( a66094a  and  a66091a );
 a66096a <=( a66095a  and  a66088a );
 a66100a <=( A199  and  A166 );
 a66101a <=( A167  and  a66100a );
 a66104a <=( (not A201)  and  A200 );
 a66107a <=( A265  and  (not A202) );
 a66108a <=( a66107a  and  a66104a );
 a66109a <=( a66108a  and  a66101a );
 a66113a <=( A269  and  (not A268) );
 a66114a <=( (not A266)  and  a66113a );
 a66117a <=( (not A299)  and  A298 );
 a66120a <=( A301  and  (not A300) );
 a66121a <=( a66120a  and  a66117a );
 a66122a <=( a66121a  and  a66114a );
 a66126a <=( A199  and  A166 );
 a66127a <=( A167  and  a66126a );
 a66130a <=( (not A201)  and  A200 );
 a66133a <=( A265  and  (not A202) );
 a66134a <=( a66133a  and  a66130a );
 a66135a <=( a66134a  and  a66127a );
 a66139a <=( A269  and  (not A268) );
 a66140a <=( (not A266)  and  a66139a );
 a66143a <=( (not A299)  and  A298 );
 a66146a <=( (not A302)  and  (not A300) );
 a66147a <=( a66146a  and  a66143a );
 a66148a <=( a66147a  and  a66140a );
 a66152a <=( A199  and  A166 );
 a66153a <=( A167  and  a66152a );
 a66156a <=( (not A201)  and  A200 );
 a66159a <=( A265  and  (not A202) );
 a66160a <=( a66159a  and  a66156a );
 a66161a <=( a66160a  and  a66153a );
 a66165a <=( A269  and  (not A268) );
 a66166a <=( (not A266)  and  a66165a );
 a66169a <=( A299  and  (not A298) );
 a66172a <=( A301  and  (not A300) );
 a66173a <=( a66172a  and  a66169a );
 a66174a <=( a66173a  and  a66166a );
 a66178a <=( A199  and  A166 );
 a66179a <=( A167  and  a66178a );
 a66182a <=( (not A201)  and  A200 );
 a66185a <=( A265  and  (not A202) );
 a66186a <=( a66185a  and  a66182a );
 a66187a <=( a66186a  and  a66179a );
 a66191a <=( A269  and  (not A268) );
 a66192a <=( (not A266)  and  a66191a );
 a66195a <=( A299  and  (not A298) );
 a66198a <=( (not A302)  and  (not A300) );
 a66199a <=( a66198a  and  a66195a );
 a66200a <=( a66199a  and  a66192a );
 a66204a <=( A199  and  A166 );
 a66205a <=( A167  and  a66204a );
 a66208a <=( (not A201)  and  A200 );
 a66211a <=( (not A265)  and  (not A202) );
 a66212a <=( a66211a  and  a66208a );
 a66213a <=( a66212a  and  a66205a );
 a66217a <=( (not A269)  and  A268 );
 a66218a <=( (not A266)  and  a66217a );
 a66221a <=( A299  and  A298 );
 a66224a <=( (not A301)  and  (not A300) );
 a66225a <=( a66224a  and  a66221a );
 a66226a <=( a66225a  and  a66218a );
 a66230a <=( A199  and  A166 );
 a66231a <=( A167  and  a66230a );
 a66234a <=( (not A201)  and  A200 );
 a66237a <=( (not A265)  and  (not A202) );
 a66238a <=( a66237a  and  a66234a );
 a66239a <=( a66238a  and  a66231a );
 a66243a <=( (not A269)  and  A268 );
 a66244a <=( (not A266)  and  a66243a );
 a66247a <=( A299  and  A298 );
 a66250a <=( A302  and  (not A300) );
 a66251a <=( a66250a  and  a66247a );
 a66252a <=( a66251a  and  a66244a );
 a66256a <=( A199  and  A166 );
 a66257a <=( A167  and  a66256a );
 a66260a <=( (not A201)  and  A200 );
 a66263a <=( (not A265)  and  (not A202) );
 a66264a <=( a66263a  and  a66260a );
 a66265a <=( a66264a  and  a66257a );
 a66269a <=( (not A269)  and  A268 );
 a66270a <=( (not A266)  and  a66269a );
 a66273a <=( (not A299)  and  A298 );
 a66276a <=( A301  and  (not A300) );
 a66277a <=( a66276a  and  a66273a );
 a66278a <=( a66277a  and  a66270a );
 a66282a <=( A199  and  A166 );
 a66283a <=( A167  and  a66282a );
 a66286a <=( (not A201)  and  A200 );
 a66289a <=( (not A265)  and  (not A202) );
 a66290a <=( a66289a  and  a66286a );
 a66291a <=( a66290a  and  a66283a );
 a66295a <=( (not A269)  and  A268 );
 a66296a <=( (not A266)  and  a66295a );
 a66299a <=( (not A299)  and  A298 );
 a66302a <=( (not A302)  and  (not A300) );
 a66303a <=( a66302a  and  a66299a );
 a66304a <=( a66303a  and  a66296a );
 a66308a <=( A199  and  A166 );
 a66309a <=( A167  and  a66308a );
 a66312a <=( (not A201)  and  A200 );
 a66315a <=( (not A265)  and  (not A202) );
 a66316a <=( a66315a  and  a66312a );
 a66317a <=( a66316a  and  a66309a );
 a66321a <=( (not A269)  and  A268 );
 a66322a <=( (not A266)  and  a66321a );
 a66325a <=( A299  and  (not A298) );
 a66328a <=( A301  and  (not A300) );
 a66329a <=( a66328a  and  a66325a );
 a66330a <=( a66329a  and  a66322a );
 a66334a <=( A199  and  A166 );
 a66335a <=( A167  and  a66334a );
 a66338a <=( (not A201)  and  A200 );
 a66341a <=( (not A265)  and  (not A202) );
 a66342a <=( a66341a  and  a66338a );
 a66343a <=( a66342a  and  a66335a );
 a66347a <=( (not A269)  and  A268 );
 a66348a <=( (not A266)  and  a66347a );
 a66351a <=( A299  and  (not A298) );
 a66354a <=( (not A302)  and  (not A300) );
 a66355a <=( a66354a  and  a66351a );
 a66356a <=( a66355a  and  a66348a );
 a66360a <=( A199  and  A166 );
 a66361a <=( A167  and  a66360a );
 a66364a <=( (not A201)  and  A200 );
 a66367a <=( A265  and  A203 );
 a66368a <=( a66367a  and  a66364a );
 a66369a <=( a66368a  and  a66361a );
 a66373a <=( (not A269)  and  A268 );
 a66374a <=( A266  and  a66373a );
 a66377a <=( A299  and  A298 );
 a66380a <=( (not A301)  and  (not A300) );
 a66381a <=( a66380a  and  a66377a );
 a66382a <=( a66381a  and  a66374a );
 a66386a <=( A199  and  A166 );
 a66387a <=( A167  and  a66386a );
 a66390a <=( (not A201)  and  A200 );
 a66393a <=( A265  and  A203 );
 a66394a <=( a66393a  and  a66390a );
 a66395a <=( a66394a  and  a66387a );
 a66399a <=( (not A269)  and  A268 );
 a66400a <=( A266  and  a66399a );
 a66403a <=( A299  and  A298 );
 a66406a <=( A302  and  (not A300) );
 a66407a <=( a66406a  and  a66403a );
 a66408a <=( a66407a  and  a66400a );
 a66412a <=( A199  and  A166 );
 a66413a <=( A167  and  a66412a );
 a66416a <=( (not A201)  and  A200 );
 a66419a <=( A265  and  A203 );
 a66420a <=( a66419a  and  a66416a );
 a66421a <=( a66420a  and  a66413a );
 a66425a <=( (not A269)  and  A268 );
 a66426a <=( A266  and  a66425a );
 a66429a <=( (not A299)  and  A298 );
 a66432a <=( A301  and  (not A300) );
 a66433a <=( a66432a  and  a66429a );
 a66434a <=( a66433a  and  a66426a );
 a66438a <=( A199  and  A166 );
 a66439a <=( A167  and  a66438a );
 a66442a <=( (not A201)  and  A200 );
 a66445a <=( A265  and  A203 );
 a66446a <=( a66445a  and  a66442a );
 a66447a <=( a66446a  and  a66439a );
 a66451a <=( (not A269)  and  A268 );
 a66452a <=( A266  and  a66451a );
 a66455a <=( (not A299)  and  A298 );
 a66458a <=( (not A302)  and  (not A300) );
 a66459a <=( a66458a  and  a66455a );
 a66460a <=( a66459a  and  a66452a );
 a66464a <=( A199  and  A166 );
 a66465a <=( A167  and  a66464a );
 a66468a <=( (not A201)  and  A200 );
 a66471a <=( A265  and  A203 );
 a66472a <=( a66471a  and  a66468a );
 a66473a <=( a66472a  and  a66465a );
 a66477a <=( (not A269)  and  A268 );
 a66478a <=( A266  and  a66477a );
 a66481a <=( A299  and  (not A298) );
 a66484a <=( A301  and  (not A300) );
 a66485a <=( a66484a  and  a66481a );
 a66486a <=( a66485a  and  a66478a );
 a66490a <=( A199  and  A166 );
 a66491a <=( A167  and  a66490a );
 a66494a <=( (not A201)  and  A200 );
 a66497a <=( A265  and  A203 );
 a66498a <=( a66497a  and  a66494a );
 a66499a <=( a66498a  and  a66491a );
 a66503a <=( (not A269)  and  A268 );
 a66504a <=( A266  and  a66503a );
 a66507a <=( A299  and  (not A298) );
 a66510a <=( (not A302)  and  (not A300) );
 a66511a <=( a66510a  and  a66507a );
 a66512a <=( a66511a  and  a66504a );
 a66516a <=( A199  and  A166 );
 a66517a <=( A167  and  a66516a );
 a66520a <=( (not A201)  and  A200 );
 a66523a <=( (not A265)  and  A203 );
 a66524a <=( a66523a  and  a66520a );
 a66525a <=( a66524a  and  a66517a );
 a66529a <=( A269  and  (not A268) );
 a66530a <=( A266  and  a66529a );
 a66533a <=( A299  and  A298 );
 a66536a <=( (not A301)  and  (not A300) );
 a66537a <=( a66536a  and  a66533a );
 a66538a <=( a66537a  and  a66530a );
 a66542a <=( A199  and  A166 );
 a66543a <=( A167  and  a66542a );
 a66546a <=( (not A201)  and  A200 );
 a66549a <=( (not A265)  and  A203 );
 a66550a <=( a66549a  and  a66546a );
 a66551a <=( a66550a  and  a66543a );
 a66555a <=( A269  and  (not A268) );
 a66556a <=( A266  and  a66555a );
 a66559a <=( A299  and  A298 );
 a66562a <=( A302  and  (not A300) );
 a66563a <=( a66562a  and  a66559a );
 a66564a <=( a66563a  and  a66556a );
 a66568a <=( A199  and  A166 );
 a66569a <=( A167  and  a66568a );
 a66572a <=( (not A201)  and  A200 );
 a66575a <=( (not A265)  and  A203 );
 a66576a <=( a66575a  and  a66572a );
 a66577a <=( a66576a  and  a66569a );
 a66581a <=( A269  and  (not A268) );
 a66582a <=( A266  and  a66581a );
 a66585a <=( (not A299)  and  A298 );
 a66588a <=( A301  and  (not A300) );
 a66589a <=( a66588a  and  a66585a );
 a66590a <=( a66589a  and  a66582a );
 a66594a <=( A199  and  A166 );
 a66595a <=( A167  and  a66594a );
 a66598a <=( (not A201)  and  A200 );
 a66601a <=( (not A265)  and  A203 );
 a66602a <=( a66601a  and  a66598a );
 a66603a <=( a66602a  and  a66595a );
 a66607a <=( A269  and  (not A268) );
 a66608a <=( A266  and  a66607a );
 a66611a <=( (not A299)  and  A298 );
 a66614a <=( (not A302)  and  (not A300) );
 a66615a <=( a66614a  and  a66611a );
 a66616a <=( a66615a  and  a66608a );
 a66620a <=( A199  and  A166 );
 a66621a <=( A167  and  a66620a );
 a66624a <=( (not A201)  and  A200 );
 a66627a <=( (not A265)  and  A203 );
 a66628a <=( a66627a  and  a66624a );
 a66629a <=( a66628a  and  a66621a );
 a66633a <=( A269  and  (not A268) );
 a66634a <=( A266  and  a66633a );
 a66637a <=( A299  and  (not A298) );
 a66640a <=( A301  and  (not A300) );
 a66641a <=( a66640a  and  a66637a );
 a66642a <=( a66641a  and  a66634a );
 a66646a <=( A199  and  A166 );
 a66647a <=( A167  and  a66646a );
 a66650a <=( (not A201)  and  A200 );
 a66653a <=( (not A265)  and  A203 );
 a66654a <=( a66653a  and  a66650a );
 a66655a <=( a66654a  and  a66647a );
 a66659a <=( A269  and  (not A268) );
 a66660a <=( A266  and  a66659a );
 a66663a <=( A299  and  (not A298) );
 a66666a <=( (not A302)  and  (not A300) );
 a66667a <=( a66666a  and  a66663a );
 a66668a <=( a66667a  and  a66660a );
 a66672a <=( A199  and  A166 );
 a66673a <=( A167  and  a66672a );
 a66676a <=( (not A201)  and  A200 );
 a66679a <=( A265  and  A203 );
 a66680a <=( a66679a  and  a66676a );
 a66681a <=( a66680a  and  a66673a );
 a66685a <=( A269  and  (not A268) );
 a66686a <=( (not A266)  and  a66685a );
 a66689a <=( A299  and  A298 );
 a66692a <=( (not A301)  and  (not A300) );
 a66693a <=( a66692a  and  a66689a );
 a66694a <=( a66693a  and  a66686a );
 a66698a <=( A199  and  A166 );
 a66699a <=( A167  and  a66698a );
 a66702a <=( (not A201)  and  A200 );
 a66705a <=( A265  and  A203 );
 a66706a <=( a66705a  and  a66702a );
 a66707a <=( a66706a  and  a66699a );
 a66711a <=( A269  and  (not A268) );
 a66712a <=( (not A266)  and  a66711a );
 a66715a <=( A299  and  A298 );
 a66718a <=( A302  and  (not A300) );
 a66719a <=( a66718a  and  a66715a );
 a66720a <=( a66719a  and  a66712a );
 a66724a <=( A199  and  A166 );
 a66725a <=( A167  and  a66724a );
 a66728a <=( (not A201)  and  A200 );
 a66731a <=( A265  and  A203 );
 a66732a <=( a66731a  and  a66728a );
 a66733a <=( a66732a  and  a66725a );
 a66737a <=( A269  and  (not A268) );
 a66738a <=( (not A266)  and  a66737a );
 a66741a <=( (not A299)  and  A298 );
 a66744a <=( A301  and  (not A300) );
 a66745a <=( a66744a  and  a66741a );
 a66746a <=( a66745a  and  a66738a );
 a66750a <=( A199  and  A166 );
 a66751a <=( A167  and  a66750a );
 a66754a <=( (not A201)  and  A200 );
 a66757a <=( A265  and  A203 );
 a66758a <=( a66757a  and  a66754a );
 a66759a <=( a66758a  and  a66751a );
 a66763a <=( A269  and  (not A268) );
 a66764a <=( (not A266)  and  a66763a );
 a66767a <=( (not A299)  and  A298 );
 a66770a <=( (not A302)  and  (not A300) );
 a66771a <=( a66770a  and  a66767a );
 a66772a <=( a66771a  and  a66764a );
 a66776a <=( A199  and  A166 );
 a66777a <=( A167  and  a66776a );
 a66780a <=( (not A201)  and  A200 );
 a66783a <=( A265  and  A203 );
 a66784a <=( a66783a  and  a66780a );
 a66785a <=( a66784a  and  a66777a );
 a66789a <=( A269  and  (not A268) );
 a66790a <=( (not A266)  and  a66789a );
 a66793a <=( A299  and  (not A298) );
 a66796a <=( A301  and  (not A300) );
 a66797a <=( a66796a  and  a66793a );
 a66798a <=( a66797a  and  a66790a );
 a66802a <=( A199  and  A166 );
 a66803a <=( A167  and  a66802a );
 a66806a <=( (not A201)  and  A200 );
 a66809a <=( A265  and  A203 );
 a66810a <=( a66809a  and  a66806a );
 a66811a <=( a66810a  and  a66803a );
 a66815a <=( A269  and  (not A268) );
 a66816a <=( (not A266)  and  a66815a );
 a66819a <=( A299  and  (not A298) );
 a66822a <=( (not A302)  and  (not A300) );
 a66823a <=( a66822a  and  a66819a );
 a66824a <=( a66823a  and  a66816a );
 a66828a <=( A199  and  A166 );
 a66829a <=( A167  and  a66828a );
 a66832a <=( (not A201)  and  A200 );
 a66835a <=( (not A265)  and  A203 );
 a66836a <=( a66835a  and  a66832a );
 a66837a <=( a66836a  and  a66829a );
 a66841a <=( (not A269)  and  A268 );
 a66842a <=( (not A266)  and  a66841a );
 a66845a <=( A299  and  A298 );
 a66848a <=( (not A301)  and  (not A300) );
 a66849a <=( a66848a  and  a66845a );
 a66850a <=( a66849a  and  a66842a );
 a66854a <=( A199  and  A166 );
 a66855a <=( A167  and  a66854a );
 a66858a <=( (not A201)  and  A200 );
 a66861a <=( (not A265)  and  A203 );
 a66862a <=( a66861a  and  a66858a );
 a66863a <=( a66862a  and  a66855a );
 a66867a <=( (not A269)  and  A268 );
 a66868a <=( (not A266)  and  a66867a );
 a66871a <=( A299  and  A298 );
 a66874a <=( A302  and  (not A300) );
 a66875a <=( a66874a  and  a66871a );
 a66876a <=( a66875a  and  a66868a );
 a66880a <=( A199  and  A166 );
 a66881a <=( A167  and  a66880a );
 a66884a <=( (not A201)  and  A200 );
 a66887a <=( (not A265)  and  A203 );
 a66888a <=( a66887a  and  a66884a );
 a66889a <=( a66888a  and  a66881a );
 a66893a <=( (not A269)  and  A268 );
 a66894a <=( (not A266)  and  a66893a );
 a66897a <=( (not A299)  and  A298 );
 a66900a <=( A301  and  (not A300) );
 a66901a <=( a66900a  and  a66897a );
 a66902a <=( a66901a  and  a66894a );
 a66906a <=( A199  and  A166 );
 a66907a <=( A167  and  a66906a );
 a66910a <=( (not A201)  and  A200 );
 a66913a <=( (not A265)  and  A203 );
 a66914a <=( a66913a  and  a66910a );
 a66915a <=( a66914a  and  a66907a );
 a66919a <=( (not A269)  and  A268 );
 a66920a <=( (not A266)  and  a66919a );
 a66923a <=( (not A299)  and  A298 );
 a66926a <=( (not A302)  and  (not A300) );
 a66927a <=( a66926a  and  a66923a );
 a66928a <=( a66927a  and  a66920a );
 a66932a <=( A199  and  A166 );
 a66933a <=( A167  and  a66932a );
 a66936a <=( (not A201)  and  A200 );
 a66939a <=( (not A265)  and  A203 );
 a66940a <=( a66939a  and  a66936a );
 a66941a <=( a66940a  and  a66933a );
 a66945a <=( (not A269)  and  A268 );
 a66946a <=( (not A266)  and  a66945a );
 a66949a <=( A299  and  (not A298) );
 a66952a <=( A301  and  (not A300) );
 a66953a <=( a66952a  and  a66949a );
 a66954a <=( a66953a  and  a66946a );
 a66958a <=( A199  and  A166 );
 a66959a <=( A167  and  a66958a );
 a66962a <=( (not A201)  and  A200 );
 a66965a <=( (not A265)  and  A203 );
 a66966a <=( a66965a  and  a66962a );
 a66967a <=( a66966a  and  a66959a );
 a66971a <=( (not A269)  and  A268 );
 a66972a <=( (not A266)  and  a66971a );
 a66975a <=( A299  and  (not A298) );
 a66978a <=( (not A302)  and  (not A300) );
 a66979a <=( a66978a  and  a66975a );
 a66980a <=( a66979a  and  a66972a );
 a66984a <=( (not A199)  and  A166 );
 a66985a <=( A167  and  a66984a );
 a66988a <=( (not A202)  and  A200 );
 a66991a <=( A265  and  A203 );
 a66992a <=( a66991a  and  a66988a );
 a66993a <=( a66992a  and  a66985a );
 a66997a <=( (not A268)  and  (not A267) );
 a66998a <=( A266  and  a66997a );
 a67001a <=( A299  and  A298 );
 a67004a <=( (not A302)  and  A301 );
 a67005a <=( a67004a  and  a67001a );
 a67006a <=( a67005a  and  a66998a );
 a67010a <=( (not A199)  and  A166 );
 a67011a <=( A167  and  a67010a );
 a67014a <=( (not A202)  and  A200 );
 a67017a <=( A265  and  A203 );
 a67018a <=( a67017a  and  a67014a );
 a67019a <=( a67018a  and  a67011a );
 a67023a <=( (not A268)  and  (not A267) );
 a67024a <=( A266  and  a67023a );
 a67027a <=( (not A299)  and  A298 );
 a67030a <=( A302  and  (not A301) );
 a67031a <=( a67030a  and  a67027a );
 a67032a <=( a67031a  and  a67024a );
 a67036a <=( (not A199)  and  A166 );
 a67037a <=( A167  and  a67036a );
 a67040a <=( (not A202)  and  A200 );
 a67043a <=( A265  and  A203 );
 a67044a <=( a67043a  and  a67040a );
 a67045a <=( a67044a  and  a67037a );
 a67049a <=( (not A268)  and  (not A267) );
 a67050a <=( A266  and  a67049a );
 a67053a <=( A299  and  (not A298) );
 a67056a <=( A302  and  (not A301) );
 a67057a <=( a67056a  and  a67053a );
 a67058a <=( a67057a  and  a67050a );
 a67062a <=( (not A199)  and  A166 );
 a67063a <=( A167  and  a67062a );
 a67066a <=( (not A202)  and  A200 );
 a67069a <=( A265  and  A203 );
 a67070a <=( a67069a  and  a67066a );
 a67071a <=( a67070a  and  a67063a );
 a67075a <=( (not A268)  and  (not A267) );
 a67076a <=( A266  and  a67075a );
 a67079a <=( (not A299)  and  (not A298) );
 a67082a <=( (not A302)  and  A301 );
 a67083a <=( a67082a  and  a67079a );
 a67084a <=( a67083a  and  a67076a );
 a67088a <=( (not A199)  and  A166 );
 a67089a <=( A167  and  a67088a );
 a67092a <=( (not A202)  and  A200 );
 a67095a <=( A265  and  A203 );
 a67096a <=( a67095a  and  a67092a );
 a67097a <=( a67096a  and  a67089a );
 a67101a <=( A269  and  (not A267) );
 a67102a <=( A266  and  a67101a );
 a67105a <=( A299  and  A298 );
 a67108a <=( (not A302)  and  A301 );
 a67109a <=( a67108a  and  a67105a );
 a67110a <=( a67109a  and  a67102a );
 a67114a <=( (not A199)  and  A166 );
 a67115a <=( A167  and  a67114a );
 a67118a <=( (not A202)  and  A200 );
 a67121a <=( A265  and  A203 );
 a67122a <=( a67121a  and  a67118a );
 a67123a <=( a67122a  and  a67115a );
 a67127a <=( A269  and  (not A267) );
 a67128a <=( A266  and  a67127a );
 a67131a <=( (not A299)  and  A298 );
 a67134a <=( A302  and  (not A301) );
 a67135a <=( a67134a  and  a67131a );
 a67136a <=( a67135a  and  a67128a );
 a67140a <=( (not A199)  and  A166 );
 a67141a <=( A167  and  a67140a );
 a67144a <=( (not A202)  and  A200 );
 a67147a <=( A265  and  A203 );
 a67148a <=( a67147a  and  a67144a );
 a67149a <=( a67148a  and  a67141a );
 a67153a <=( A269  and  (not A267) );
 a67154a <=( A266  and  a67153a );
 a67157a <=( A299  and  (not A298) );
 a67160a <=( A302  and  (not A301) );
 a67161a <=( a67160a  and  a67157a );
 a67162a <=( a67161a  and  a67154a );
 a67166a <=( (not A199)  and  A166 );
 a67167a <=( A167  and  a67166a );
 a67170a <=( (not A202)  and  A200 );
 a67173a <=( A265  and  A203 );
 a67174a <=( a67173a  and  a67170a );
 a67175a <=( a67174a  and  a67167a );
 a67179a <=( A269  and  (not A267) );
 a67180a <=( A266  and  a67179a );
 a67183a <=( (not A299)  and  (not A298) );
 a67186a <=( (not A302)  and  A301 );
 a67187a <=( a67186a  and  a67183a );
 a67188a <=( a67187a  and  a67180a );
 a67192a <=( (not A199)  and  A166 );
 a67193a <=( A167  and  a67192a );
 a67196a <=( (not A202)  and  A200 );
 a67199a <=( (not A265)  and  A203 );
 a67200a <=( a67199a  and  a67196a );
 a67201a <=( a67200a  and  a67193a );
 a67205a <=( A268  and  (not A267) );
 a67206a <=( A266  and  a67205a );
 a67209a <=( A299  and  A298 );
 a67212a <=( (not A302)  and  A301 );
 a67213a <=( a67212a  and  a67209a );
 a67214a <=( a67213a  and  a67206a );
 a67218a <=( (not A199)  and  A166 );
 a67219a <=( A167  and  a67218a );
 a67222a <=( (not A202)  and  A200 );
 a67225a <=( (not A265)  and  A203 );
 a67226a <=( a67225a  and  a67222a );
 a67227a <=( a67226a  and  a67219a );
 a67231a <=( A268  and  (not A267) );
 a67232a <=( A266  and  a67231a );
 a67235a <=( (not A299)  and  A298 );
 a67238a <=( A302  and  (not A301) );
 a67239a <=( a67238a  and  a67235a );
 a67240a <=( a67239a  and  a67232a );
 a67244a <=( (not A199)  and  A166 );
 a67245a <=( A167  and  a67244a );
 a67248a <=( (not A202)  and  A200 );
 a67251a <=( (not A265)  and  A203 );
 a67252a <=( a67251a  and  a67248a );
 a67253a <=( a67252a  and  a67245a );
 a67257a <=( A268  and  (not A267) );
 a67258a <=( A266  and  a67257a );
 a67261a <=( A299  and  (not A298) );
 a67264a <=( A302  and  (not A301) );
 a67265a <=( a67264a  and  a67261a );
 a67266a <=( a67265a  and  a67258a );
 a67270a <=( (not A199)  and  A166 );
 a67271a <=( A167  and  a67270a );
 a67274a <=( (not A202)  and  A200 );
 a67277a <=( (not A265)  and  A203 );
 a67278a <=( a67277a  and  a67274a );
 a67279a <=( a67278a  and  a67271a );
 a67283a <=( A268  and  (not A267) );
 a67284a <=( A266  and  a67283a );
 a67287a <=( (not A299)  and  (not A298) );
 a67290a <=( (not A302)  and  A301 );
 a67291a <=( a67290a  and  a67287a );
 a67292a <=( a67291a  and  a67284a );
 a67296a <=( (not A199)  and  A166 );
 a67297a <=( A167  and  a67296a );
 a67300a <=( (not A202)  and  A200 );
 a67303a <=( (not A265)  and  A203 );
 a67304a <=( a67303a  and  a67300a );
 a67305a <=( a67304a  and  a67297a );
 a67309a <=( (not A269)  and  (not A267) );
 a67310a <=( A266  and  a67309a );
 a67313a <=( A299  and  A298 );
 a67316a <=( (not A302)  and  A301 );
 a67317a <=( a67316a  and  a67313a );
 a67318a <=( a67317a  and  a67310a );
 a67322a <=( (not A199)  and  A166 );
 a67323a <=( A167  and  a67322a );
 a67326a <=( (not A202)  and  A200 );
 a67329a <=( (not A265)  and  A203 );
 a67330a <=( a67329a  and  a67326a );
 a67331a <=( a67330a  and  a67323a );
 a67335a <=( (not A269)  and  (not A267) );
 a67336a <=( A266  and  a67335a );
 a67339a <=( (not A299)  and  A298 );
 a67342a <=( A302  and  (not A301) );
 a67343a <=( a67342a  and  a67339a );
 a67344a <=( a67343a  and  a67336a );
 a67348a <=( (not A199)  and  A166 );
 a67349a <=( A167  and  a67348a );
 a67352a <=( (not A202)  and  A200 );
 a67355a <=( (not A265)  and  A203 );
 a67356a <=( a67355a  and  a67352a );
 a67357a <=( a67356a  and  a67349a );
 a67361a <=( (not A269)  and  (not A267) );
 a67362a <=( A266  and  a67361a );
 a67365a <=( A299  and  (not A298) );
 a67368a <=( A302  and  (not A301) );
 a67369a <=( a67368a  and  a67365a );
 a67370a <=( a67369a  and  a67362a );
 a67374a <=( (not A199)  and  A166 );
 a67375a <=( A167  and  a67374a );
 a67378a <=( (not A202)  and  A200 );
 a67381a <=( (not A265)  and  A203 );
 a67382a <=( a67381a  and  a67378a );
 a67383a <=( a67382a  and  a67375a );
 a67387a <=( (not A269)  and  (not A267) );
 a67388a <=( A266  and  a67387a );
 a67391a <=( (not A299)  and  (not A298) );
 a67394a <=( (not A302)  and  A301 );
 a67395a <=( a67394a  and  a67391a );
 a67396a <=( a67395a  and  a67388a );
 a67400a <=( (not A199)  and  A166 );
 a67401a <=( A167  and  a67400a );
 a67404a <=( (not A202)  and  A200 );
 a67407a <=( A265  and  A203 );
 a67408a <=( a67407a  and  a67404a );
 a67409a <=( a67408a  and  a67401a );
 a67413a <=( A268  and  (not A267) );
 a67414a <=( (not A266)  and  a67413a );
 a67417a <=( A299  and  A298 );
 a67420a <=( (not A302)  and  A301 );
 a67421a <=( a67420a  and  a67417a );
 a67422a <=( a67421a  and  a67414a );
 a67426a <=( (not A199)  and  A166 );
 a67427a <=( A167  and  a67426a );
 a67430a <=( (not A202)  and  A200 );
 a67433a <=( A265  and  A203 );
 a67434a <=( a67433a  and  a67430a );
 a67435a <=( a67434a  and  a67427a );
 a67439a <=( A268  and  (not A267) );
 a67440a <=( (not A266)  and  a67439a );
 a67443a <=( (not A299)  and  A298 );
 a67446a <=( A302  and  (not A301) );
 a67447a <=( a67446a  and  a67443a );
 a67448a <=( a67447a  and  a67440a );
 a67452a <=( (not A199)  and  A166 );
 a67453a <=( A167  and  a67452a );
 a67456a <=( (not A202)  and  A200 );
 a67459a <=( A265  and  A203 );
 a67460a <=( a67459a  and  a67456a );
 a67461a <=( a67460a  and  a67453a );
 a67465a <=( A268  and  (not A267) );
 a67466a <=( (not A266)  and  a67465a );
 a67469a <=( A299  and  (not A298) );
 a67472a <=( A302  and  (not A301) );
 a67473a <=( a67472a  and  a67469a );
 a67474a <=( a67473a  and  a67466a );
 a67478a <=( (not A199)  and  A166 );
 a67479a <=( A167  and  a67478a );
 a67482a <=( (not A202)  and  A200 );
 a67485a <=( A265  and  A203 );
 a67486a <=( a67485a  and  a67482a );
 a67487a <=( a67486a  and  a67479a );
 a67491a <=( A268  and  (not A267) );
 a67492a <=( (not A266)  and  a67491a );
 a67495a <=( (not A299)  and  (not A298) );
 a67498a <=( (not A302)  and  A301 );
 a67499a <=( a67498a  and  a67495a );
 a67500a <=( a67499a  and  a67492a );
 a67504a <=( (not A199)  and  A166 );
 a67505a <=( A167  and  a67504a );
 a67508a <=( (not A202)  and  A200 );
 a67511a <=( A265  and  A203 );
 a67512a <=( a67511a  and  a67508a );
 a67513a <=( a67512a  and  a67505a );
 a67517a <=( (not A269)  and  (not A267) );
 a67518a <=( (not A266)  and  a67517a );
 a67521a <=( A299  and  A298 );
 a67524a <=( (not A302)  and  A301 );
 a67525a <=( a67524a  and  a67521a );
 a67526a <=( a67525a  and  a67518a );
 a67530a <=( (not A199)  and  A166 );
 a67531a <=( A167  and  a67530a );
 a67534a <=( (not A202)  and  A200 );
 a67537a <=( A265  and  A203 );
 a67538a <=( a67537a  and  a67534a );
 a67539a <=( a67538a  and  a67531a );
 a67543a <=( (not A269)  and  (not A267) );
 a67544a <=( (not A266)  and  a67543a );
 a67547a <=( (not A299)  and  A298 );
 a67550a <=( A302  and  (not A301) );
 a67551a <=( a67550a  and  a67547a );
 a67552a <=( a67551a  and  a67544a );
 a67556a <=( (not A199)  and  A166 );
 a67557a <=( A167  and  a67556a );
 a67560a <=( (not A202)  and  A200 );
 a67563a <=( A265  and  A203 );
 a67564a <=( a67563a  and  a67560a );
 a67565a <=( a67564a  and  a67557a );
 a67569a <=( (not A269)  and  (not A267) );
 a67570a <=( (not A266)  and  a67569a );
 a67573a <=( A299  and  (not A298) );
 a67576a <=( A302  and  (not A301) );
 a67577a <=( a67576a  and  a67573a );
 a67578a <=( a67577a  and  a67570a );
 a67582a <=( (not A199)  and  A166 );
 a67583a <=( A167  and  a67582a );
 a67586a <=( (not A202)  and  A200 );
 a67589a <=( A265  and  A203 );
 a67590a <=( a67589a  and  a67586a );
 a67591a <=( a67590a  and  a67583a );
 a67595a <=( (not A269)  and  (not A267) );
 a67596a <=( (not A266)  and  a67595a );
 a67599a <=( (not A299)  and  (not A298) );
 a67602a <=( (not A302)  and  A301 );
 a67603a <=( a67602a  and  a67599a );
 a67604a <=( a67603a  and  a67596a );
 a67608a <=( (not A199)  and  A166 );
 a67609a <=( A167  and  a67608a );
 a67612a <=( (not A201)  and  A200 );
 a67615a <=( A265  and  A202 );
 a67616a <=( a67615a  and  a67612a );
 a67617a <=( a67616a  and  a67609a );
 a67621a <=( (not A269)  and  A268 );
 a67622a <=( A266  and  a67621a );
 a67625a <=( A299  and  A298 );
 a67628a <=( (not A301)  and  (not A300) );
 a67629a <=( a67628a  and  a67625a );
 a67630a <=( a67629a  and  a67622a );
 a67634a <=( (not A199)  and  A166 );
 a67635a <=( A167  and  a67634a );
 a67638a <=( (not A201)  and  A200 );
 a67641a <=( A265  and  A202 );
 a67642a <=( a67641a  and  a67638a );
 a67643a <=( a67642a  and  a67635a );
 a67647a <=( (not A269)  and  A268 );
 a67648a <=( A266  and  a67647a );
 a67651a <=( A299  and  A298 );
 a67654a <=( A302  and  (not A300) );
 a67655a <=( a67654a  and  a67651a );
 a67656a <=( a67655a  and  a67648a );
 a67660a <=( (not A199)  and  A166 );
 a67661a <=( A167  and  a67660a );
 a67664a <=( (not A201)  and  A200 );
 a67667a <=( A265  and  A202 );
 a67668a <=( a67667a  and  a67664a );
 a67669a <=( a67668a  and  a67661a );
 a67673a <=( (not A269)  and  A268 );
 a67674a <=( A266  and  a67673a );
 a67677a <=( (not A299)  and  A298 );
 a67680a <=( A301  and  (not A300) );
 a67681a <=( a67680a  and  a67677a );
 a67682a <=( a67681a  and  a67674a );
 a67686a <=( (not A199)  and  A166 );
 a67687a <=( A167  and  a67686a );
 a67690a <=( (not A201)  and  A200 );
 a67693a <=( A265  and  A202 );
 a67694a <=( a67693a  and  a67690a );
 a67695a <=( a67694a  and  a67687a );
 a67699a <=( (not A269)  and  A268 );
 a67700a <=( A266  and  a67699a );
 a67703a <=( (not A299)  and  A298 );
 a67706a <=( (not A302)  and  (not A300) );
 a67707a <=( a67706a  and  a67703a );
 a67708a <=( a67707a  and  a67700a );
 a67712a <=( (not A199)  and  A166 );
 a67713a <=( A167  and  a67712a );
 a67716a <=( (not A201)  and  A200 );
 a67719a <=( A265  and  A202 );
 a67720a <=( a67719a  and  a67716a );
 a67721a <=( a67720a  and  a67713a );
 a67725a <=( (not A269)  and  A268 );
 a67726a <=( A266  and  a67725a );
 a67729a <=( A299  and  (not A298) );
 a67732a <=( A301  and  (not A300) );
 a67733a <=( a67732a  and  a67729a );
 a67734a <=( a67733a  and  a67726a );
 a67738a <=( (not A199)  and  A166 );
 a67739a <=( A167  and  a67738a );
 a67742a <=( (not A201)  and  A200 );
 a67745a <=( A265  and  A202 );
 a67746a <=( a67745a  and  a67742a );
 a67747a <=( a67746a  and  a67739a );
 a67751a <=( (not A269)  and  A268 );
 a67752a <=( A266  and  a67751a );
 a67755a <=( A299  and  (not A298) );
 a67758a <=( (not A302)  and  (not A300) );
 a67759a <=( a67758a  and  a67755a );
 a67760a <=( a67759a  and  a67752a );
 a67764a <=( (not A199)  and  A166 );
 a67765a <=( A167  and  a67764a );
 a67768a <=( (not A201)  and  A200 );
 a67771a <=( (not A265)  and  A202 );
 a67772a <=( a67771a  and  a67768a );
 a67773a <=( a67772a  and  a67765a );
 a67777a <=( A269  and  (not A268) );
 a67778a <=( A266  and  a67777a );
 a67781a <=( A299  and  A298 );
 a67784a <=( (not A301)  and  (not A300) );
 a67785a <=( a67784a  and  a67781a );
 a67786a <=( a67785a  and  a67778a );
 a67790a <=( (not A199)  and  A166 );
 a67791a <=( A167  and  a67790a );
 a67794a <=( (not A201)  and  A200 );
 a67797a <=( (not A265)  and  A202 );
 a67798a <=( a67797a  and  a67794a );
 a67799a <=( a67798a  and  a67791a );
 a67803a <=( A269  and  (not A268) );
 a67804a <=( A266  and  a67803a );
 a67807a <=( A299  and  A298 );
 a67810a <=( A302  and  (not A300) );
 a67811a <=( a67810a  and  a67807a );
 a67812a <=( a67811a  and  a67804a );
 a67816a <=( (not A199)  and  A166 );
 a67817a <=( A167  and  a67816a );
 a67820a <=( (not A201)  and  A200 );
 a67823a <=( (not A265)  and  A202 );
 a67824a <=( a67823a  and  a67820a );
 a67825a <=( a67824a  and  a67817a );
 a67829a <=( A269  and  (not A268) );
 a67830a <=( A266  and  a67829a );
 a67833a <=( (not A299)  and  A298 );
 a67836a <=( A301  and  (not A300) );
 a67837a <=( a67836a  and  a67833a );
 a67838a <=( a67837a  and  a67830a );
 a67842a <=( (not A199)  and  A166 );
 a67843a <=( A167  and  a67842a );
 a67846a <=( (not A201)  and  A200 );
 a67849a <=( (not A265)  and  A202 );
 a67850a <=( a67849a  and  a67846a );
 a67851a <=( a67850a  and  a67843a );
 a67855a <=( A269  and  (not A268) );
 a67856a <=( A266  and  a67855a );
 a67859a <=( (not A299)  and  A298 );
 a67862a <=( (not A302)  and  (not A300) );
 a67863a <=( a67862a  and  a67859a );
 a67864a <=( a67863a  and  a67856a );
 a67868a <=( (not A199)  and  A166 );
 a67869a <=( A167  and  a67868a );
 a67872a <=( (not A201)  and  A200 );
 a67875a <=( (not A265)  and  A202 );
 a67876a <=( a67875a  and  a67872a );
 a67877a <=( a67876a  and  a67869a );
 a67881a <=( A269  and  (not A268) );
 a67882a <=( A266  and  a67881a );
 a67885a <=( A299  and  (not A298) );
 a67888a <=( A301  and  (not A300) );
 a67889a <=( a67888a  and  a67885a );
 a67890a <=( a67889a  and  a67882a );
 a67894a <=( (not A199)  and  A166 );
 a67895a <=( A167  and  a67894a );
 a67898a <=( (not A201)  and  A200 );
 a67901a <=( (not A265)  and  A202 );
 a67902a <=( a67901a  and  a67898a );
 a67903a <=( a67902a  and  a67895a );
 a67907a <=( A269  and  (not A268) );
 a67908a <=( A266  and  a67907a );
 a67911a <=( A299  and  (not A298) );
 a67914a <=( (not A302)  and  (not A300) );
 a67915a <=( a67914a  and  a67911a );
 a67916a <=( a67915a  and  a67908a );
 a67920a <=( (not A199)  and  A166 );
 a67921a <=( A167  and  a67920a );
 a67924a <=( (not A201)  and  A200 );
 a67927a <=( A265  and  A202 );
 a67928a <=( a67927a  and  a67924a );
 a67929a <=( a67928a  and  a67921a );
 a67933a <=( A269  and  (not A268) );
 a67934a <=( (not A266)  and  a67933a );
 a67937a <=( A299  and  A298 );
 a67940a <=( (not A301)  and  (not A300) );
 a67941a <=( a67940a  and  a67937a );
 a67942a <=( a67941a  and  a67934a );
 a67946a <=( (not A199)  and  A166 );
 a67947a <=( A167  and  a67946a );
 a67950a <=( (not A201)  and  A200 );
 a67953a <=( A265  and  A202 );
 a67954a <=( a67953a  and  a67950a );
 a67955a <=( a67954a  and  a67947a );
 a67959a <=( A269  and  (not A268) );
 a67960a <=( (not A266)  and  a67959a );
 a67963a <=( A299  and  A298 );
 a67966a <=( A302  and  (not A300) );
 a67967a <=( a67966a  and  a67963a );
 a67968a <=( a67967a  and  a67960a );
 a67972a <=( (not A199)  and  A166 );
 a67973a <=( A167  and  a67972a );
 a67976a <=( (not A201)  and  A200 );
 a67979a <=( A265  and  A202 );
 a67980a <=( a67979a  and  a67976a );
 a67981a <=( a67980a  and  a67973a );
 a67985a <=( A269  and  (not A268) );
 a67986a <=( (not A266)  and  a67985a );
 a67989a <=( (not A299)  and  A298 );
 a67992a <=( A301  and  (not A300) );
 a67993a <=( a67992a  and  a67989a );
 a67994a <=( a67993a  and  a67986a );
 a67998a <=( (not A199)  and  A166 );
 a67999a <=( A167  and  a67998a );
 a68002a <=( (not A201)  and  A200 );
 a68005a <=( A265  and  A202 );
 a68006a <=( a68005a  and  a68002a );
 a68007a <=( a68006a  and  a67999a );
 a68011a <=( A269  and  (not A268) );
 a68012a <=( (not A266)  and  a68011a );
 a68015a <=( (not A299)  and  A298 );
 a68018a <=( (not A302)  and  (not A300) );
 a68019a <=( a68018a  and  a68015a );
 a68020a <=( a68019a  and  a68012a );
 a68024a <=( (not A199)  and  A166 );
 a68025a <=( A167  and  a68024a );
 a68028a <=( (not A201)  and  A200 );
 a68031a <=( A265  and  A202 );
 a68032a <=( a68031a  and  a68028a );
 a68033a <=( a68032a  and  a68025a );
 a68037a <=( A269  and  (not A268) );
 a68038a <=( (not A266)  and  a68037a );
 a68041a <=( A299  and  (not A298) );
 a68044a <=( A301  and  (not A300) );
 a68045a <=( a68044a  and  a68041a );
 a68046a <=( a68045a  and  a68038a );
 a68050a <=( (not A199)  and  A166 );
 a68051a <=( A167  and  a68050a );
 a68054a <=( (not A201)  and  A200 );
 a68057a <=( A265  and  A202 );
 a68058a <=( a68057a  and  a68054a );
 a68059a <=( a68058a  and  a68051a );
 a68063a <=( A269  and  (not A268) );
 a68064a <=( (not A266)  and  a68063a );
 a68067a <=( A299  and  (not A298) );
 a68070a <=( (not A302)  and  (not A300) );
 a68071a <=( a68070a  and  a68067a );
 a68072a <=( a68071a  and  a68064a );
 a68076a <=( (not A199)  and  A166 );
 a68077a <=( A167  and  a68076a );
 a68080a <=( (not A201)  and  A200 );
 a68083a <=( (not A265)  and  A202 );
 a68084a <=( a68083a  and  a68080a );
 a68085a <=( a68084a  and  a68077a );
 a68089a <=( (not A269)  and  A268 );
 a68090a <=( (not A266)  and  a68089a );
 a68093a <=( A299  and  A298 );
 a68096a <=( (not A301)  and  (not A300) );
 a68097a <=( a68096a  and  a68093a );
 a68098a <=( a68097a  and  a68090a );
 a68102a <=( (not A199)  and  A166 );
 a68103a <=( A167  and  a68102a );
 a68106a <=( (not A201)  and  A200 );
 a68109a <=( (not A265)  and  A202 );
 a68110a <=( a68109a  and  a68106a );
 a68111a <=( a68110a  and  a68103a );
 a68115a <=( (not A269)  and  A268 );
 a68116a <=( (not A266)  and  a68115a );
 a68119a <=( A299  and  A298 );
 a68122a <=( A302  and  (not A300) );
 a68123a <=( a68122a  and  a68119a );
 a68124a <=( a68123a  and  a68116a );
 a68128a <=( (not A199)  and  A166 );
 a68129a <=( A167  and  a68128a );
 a68132a <=( (not A201)  and  A200 );
 a68135a <=( (not A265)  and  A202 );
 a68136a <=( a68135a  and  a68132a );
 a68137a <=( a68136a  and  a68129a );
 a68141a <=( (not A269)  and  A268 );
 a68142a <=( (not A266)  and  a68141a );
 a68145a <=( (not A299)  and  A298 );
 a68148a <=( A301  and  (not A300) );
 a68149a <=( a68148a  and  a68145a );
 a68150a <=( a68149a  and  a68142a );
 a68154a <=( (not A199)  and  A166 );
 a68155a <=( A167  and  a68154a );
 a68158a <=( (not A201)  and  A200 );
 a68161a <=( (not A265)  and  A202 );
 a68162a <=( a68161a  and  a68158a );
 a68163a <=( a68162a  and  a68155a );
 a68167a <=( (not A269)  and  A268 );
 a68168a <=( (not A266)  and  a68167a );
 a68171a <=( (not A299)  and  A298 );
 a68174a <=( (not A302)  and  (not A300) );
 a68175a <=( a68174a  and  a68171a );
 a68176a <=( a68175a  and  a68168a );
 a68180a <=( (not A199)  and  A166 );
 a68181a <=( A167  and  a68180a );
 a68184a <=( (not A201)  and  A200 );
 a68187a <=( (not A265)  and  A202 );
 a68188a <=( a68187a  and  a68184a );
 a68189a <=( a68188a  and  a68181a );
 a68193a <=( (not A269)  and  A268 );
 a68194a <=( (not A266)  and  a68193a );
 a68197a <=( A299  and  (not A298) );
 a68200a <=( A301  and  (not A300) );
 a68201a <=( a68200a  and  a68197a );
 a68202a <=( a68201a  and  a68194a );
 a68206a <=( (not A199)  and  A166 );
 a68207a <=( A167  and  a68206a );
 a68210a <=( (not A201)  and  A200 );
 a68213a <=( (not A265)  and  A202 );
 a68214a <=( a68213a  and  a68210a );
 a68215a <=( a68214a  and  a68207a );
 a68219a <=( (not A269)  and  A268 );
 a68220a <=( (not A266)  and  a68219a );
 a68223a <=( A299  and  (not A298) );
 a68226a <=( (not A302)  and  (not A300) );
 a68227a <=( a68226a  and  a68223a );
 a68228a <=( a68227a  and  a68220a );
 a68232a <=( (not A199)  and  A166 );
 a68233a <=( A167  and  a68232a );
 a68236a <=( (not A201)  and  A200 );
 a68239a <=( A265  and  (not A203) );
 a68240a <=( a68239a  and  a68236a );
 a68241a <=( a68240a  and  a68233a );
 a68245a <=( (not A269)  and  A268 );
 a68246a <=( A266  and  a68245a );
 a68249a <=( A299  and  A298 );
 a68252a <=( (not A301)  and  (not A300) );
 a68253a <=( a68252a  and  a68249a );
 a68254a <=( a68253a  and  a68246a );
 a68258a <=( (not A199)  and  A166 );
 a68259a <=( A167  and  a68258a );
 a68262a <=( (not A201)  and  A200 );
 a68265a <=( A265  and  (not A203) );
 a68266a <=( a68265a  and  a68262a );
 a68267a <=( a68266a  and  a68259a );
 a68271a <=( (not A269)  and  A268 );
 a68272a <=( A266  and  a68271a );
 a68275a <=( A299  and  A298 );
 a68278a <=( A302  and  (not A300) );
 a68279a <=( a68278a  and  a68275a );
 a68280a <=( a68279a  and  a68272a );
 a68284a <=( (not A199)  and  A166 );
 a68285a <=( A167  and  a68284a );
 a68288a <=( (not A201)  and  A200 );
 a68291a <=( A265  and  (not A203) );
 a68292a <=( a68291a  and  a68288a );
 a68293a <=( a68292a  and  a68285a );
 a68297a <=( (not A269)  and  A268 );
 a68298a <=( A266  and  a68297a );
 a68301a <=( (not A299)  and  A298 );
 a68304a <=( A301  and  (not A300) );
 a68305a <=( a68304a  and  a68301a );
 a68306a <=( a68305a  and  a68298a );
 a68310a <=( (not A199)  and  A166 );
 a68311a <=( A167  and  a68310a );
 a68314a <=( (not A201)  and  A200 );
 a68317a <=( A265  and  (not A203) );
 a68318a <=( a68317a  and  a68314a );
 a68319a <=( a68318a  and  a68311a );
 a68323a <=( (not A269)  and  A268 );
 a68324a <=( A266  and  a68323a );
 a68327a <=( (not A299)  and  A298 );
 a68330a <=( (not A302)  and  (not A300) );
 a68331a <=( a68330a  and  a68327a );
 a68332a <=( a68331a  and  a68324a );
 a68336a <=( (not A199)  and  A166 );
 a68337a <=( A167  and  a68336a );
 a68340a <=( (not A201)  and  A200 );
 a68343a <=( A265  and  (not A203) );
 a68344a <=( a68343a  and  a68340a );
 a68345a <=( a68344a  and  a68337a );
 a68349a <=( (not A269)  and  A268 );
 a68350a <=( A266  and  a68349a );
 a68353a <=( A299  and  (not A298) );
 a68356a <=( A301  and  (not A300) );
 a68357a <=( a68356a  and  a68353a );
 a68358a <=( a68357a  and  a68350a );
 a68362a <=( (not A199)  and  A166 );
 a68363a <=( A167  and  a68362a );
 a68366a <=( (not A201)  and  A200 );
 a68369a <=( A265  and  (not A203) );
 a68370a <=( a68369a  and  a68366a );
 a68371a <=( a68370a  and  a68363a );
 a68375a <=( (not A269)  and  A268 );
 a68376a <=( A266  and  a68375a );
 a68379a <=( A299  and  (not A298) );
 a68382a <=( (not A302)  and  (not A300) );
 a68383a <=( a68382a  and  a68379a );
 a68384a <=( a68383a  and  a68376a );
 a68388a <=( (not A199)  and  A166 );
 a68389a <=( A167  and  a68388a );
 a68392a <=( (not A201)  and  A200 );
 a68395a <=( (not A265)  and  (not A203) );
 a68396a <=( a68395a  and  a68392a );
 a68397a <=( a68396a  and  a68389a );
 a68401a <=( A269  and  (not A268) );
 a68402a <=( A266  and  a68401a );
 a68405a <=( A299  and  A298 );
 a68408a <=( (not A301)  and  (not A300) );
 a68409a <=( a68408a  and  a68405a );
 a68410a <=( a68409a  and  a68402a );
 a68414a <=( (not A199)  and  A166 );
 a68415a <=( A167  and  a68414a );
 a68418a <=( (not A201)  and  A200 );
 a68421a <=( (not A265)  and  (not A203) );
 a68422a <=( a68421a  and  a68418a );
 a68423a <=( a68422a  and  a68415a );
 a68427a <=( A269  and  (not A268) );
 a68428a <=( A266  and  a68427a );
 a68431a <=( A299  and  A298 );
 a68434a <=( A302  and  (not A300) );
 a68435a <=( a68434a  and  a68431a );
 a68436a <=( a68435a  and  a68428a );
 a68440a <=( (not A199)  and  A166 );
 a68441a <=( A167  and  a68440a );
 a68444a <=( (not A201)  and  A200 );
 a68447a <=( (not A265)  and  (not A203) );
 a68448a <=( a68447a  and  a68444a );
 a68449a <=( a68448a  and  a68441a );
 a68453a <=( A269  and  (not A268) );
 a68454a <=( A266  and  a68453a );
 a68457a <=( (not A299)  and  A298 );
 a68460a <=( A301  and  (not A300) );
 a68461a <=( a68460a  and  a68457a );
 a68462a <=( a68461a  and  a68454a );
 a68466a <=( (not A199)  and  A166 );
 a68467a <=( A167  and  a68466a );
 a68470a <=( (not A201)  and  A200 );
 a68473a <=( (not A265)  and  (not A203) );
 a68474a <=( a68473a  and  a68470a );
 a68475a <=( a68474a  and  a68467a );
 a68479a <=( A269  and  (not A268) );
 a68480a <=( A266  and  a68479a );
 a68483a <=( (not A299)  and  A298 );
 a68486a <=( (not A302)  and  (not A300) );
 a68487a <=( a68486a  and  a68483a );
 a68488a <=( a68487a  and  a68480a );
 a68492a <=( (not A199)  and  A166 );
 a68493a <=( A167  and  a68492a );
 a68496a <=( (not A201)  and  A200 );
 a68499a <=( (not A265)  and  (not A203) );
 a68500a <=( a68499a  and  a68496a );
 a68501a <=( a68500a  and  a68493a );
 a68505a <=( A269  and  (not A268) );
 a68506a <=( A266  and  a68505a );
 a68509a <=( A299  and  (not A298) );
 a68512a <=( A301  and  (not A300) );
 a68513a <=( a68512a  and  a68509a );
 a68514a <=( a68513a  and  a68506a );
 a68518a <=( (not A199)  and  A166 );
 a68519a <=( A167  and  a68518a );
 a68522a <=( (not A201)  and  A200 );
 a68525a <=( (not A265)  and  (not A203) );
 a68526a <=( a68525a  and  a68522a );
 a68527a <=( a68526a  and  a68519a );
 a68531a <=( A269  and  (not A268) );
 a68532a <=( A266  and  a68531a );
 a68535a <=( A299  and  (not A298) );
 a68538a <=( (not A302)  and  (not A300) );
 a68539a <=( a68538a  and  a68535a );
 a68540a <=( a68539a  and  a68532a );
 a68544a <=( (not A199)  and  A166 );
 a68545a <=( A167  and  a68544a );
 a68548a <=( (not A201)  and  A200 );
 a68551a <=( A265  and  (not A203) );
 a68552a <=( a68551a  and  a68548a );
 a68553a <=( a68552a  and  a68545a );
 a68557a <=( A269  and  (not A268) );
 a68558a <=( (not A266)  and  a68557a );
 a68561a <=( A299  and  A298 );
 a68564a <=( (not A301)  and  (not A300) );
 a68565a <=( a68564a  and  a68561a );
 a68566a <=( a68565a  and  a68558a );
 a68570a <=( (not A199)  and  A166 );
 a68571a <=( A167  and  a68570a );
 a68574a <=( (not A201)  and  A200 );
 a68577a <=( A265  and  (not A203) );
 a68578a <=( a68577a  and  a68574a );
 a68579a <=( a68578a  and  a68571a );
 a68583a <=( A269  and  (not A268) );
 a68584a <=( (not A266)  and  a68583a );
 a68587a <=( A299  and  A298 );
 a68590a <=( A302  and  (not A300) );
 a68591a <=( a68590a  and  a68587a );
 a68592a <=( a68591a  and  a68584a );
 a68596a <=( (not A199)  and  A166 );
 a68597a <=( A167  and  a68596a );
 a68600a <=( (not A201)  and  A200 );
 a68603a <=( A265  and  (not A203) );
 a68604a <=( a68603a  and  a68600a );
 a68605a <=( a68604a  and  a68597a );
 a68609a <=( A269  and  (not A268) );
 a68610a <=( (not A266)  and  a68609a );
 a68613a <=( (not A299)  and  A298 );
 a68616a <=( A301  and  (not A300) );
 a68617a <=( a68616a  and  a68613a );
 a68618a <=( a68617a  and  a68610a );
 a68622a <=( (not A199)  and  A166 );
 a68623a <=( A167  and  a68622a );
 a68626a <=( (not A201)  and  A200 );
 a68629a <=( A265  and  (not A203) );
 a68630a <=( a68629a  and  a68626a );
 a68631a <=( a68630a  and  a68623a );
 a68635a <=( A269  and  (not A268) );
 a68636a <=( (not A266)  and  a68635a );
 a68639a <=( (not A299)  and  A298 );
 a68642a <=( (not A302)  and  (not A300) );
 a68643a <=( a68642a  and  a68639a );
 a68644a <=( a68643a  and  a68636a );
 a68648a <=( (not A199)  and  A166 );
 a68649a <=( A167  and  a68648a );
 a68652a <=( (not A201)  and  A200 );
 a68655a <=( A265  and  (not A203) );
 a68656a <=( a68655a  and  a68652a );
 a68657a <=( a68656a  and  a68649a );
 a68661a <=( A269  and  (not A268) );
 a68662a <=( (not A266)  and  a68661a );
 a68665a <=( A299  and  (not A298) );
 a68668a <=( A301  and  (not A300) );
 a68669a <=( a68668a  and  a68665a );
 a68670a <=( a68669a  and  a68662a );
 a68674a <=( (not A199)  and  A166 );
 a68675a <=( A167  and  a68674a );
 a68678a <=( (not A201)  and  A200 );
 a68681a <=( A265  and  (not A203) );
 a68682a <=( a68681a  and  a68678a );
 a68683a <=( a68682a  and  a68675a );
 a68687a <=( A269  and  (not A268) );
 a68688a <=( (not A266)  and  a68687a );
 a68691a <=( A299  and  (not A298) );
 a68694a <=( (not A302)  and  (not A300) );
 a68695a <=( a68694a  and  a68691a );
 a68696a <=( a68695a  and  a68688a );
 a68700a <=( (not A199)  and  A166 );
 a68701a <=( A167  and  a68700a );
 a68704a <=( (not A201)  and  A200 );
 a68707a <=( (not A265)  and  (not A203) );
 a68708a <=( a68707a  and  a68704a );
 a68709a <=( a68708a  and  a68701a );
 a68713a <=( (not A269)  and  A268 );
 a68714a <=( (not A266)  and  a68713a );
 a68717a <=( A299  and  A298 );
 a68720a <=( (not A301)  and  (not A300) );
 a68721a <=( a68720a  and  a68717a );
 a68722a <=( a68721a  and  a68714a );
 a68726a <=( (not A199)  and  A166 );
 a68727a <=( A167  and  a68726a );
 a68730a <=( (not A201)  and  A200 );
 a68733a <=( (not A265)  and  (not A203) );
 a68734a <=( a68733a  and  a68730a );
 a68735a <=( a68734a  and  a68727a );
 a68739a <=( (not A269)  and  A268 );
 a68740a <=( (not A266)  and  a68739a );
 a68743a <=( A299  and  A298 );
 a68746a <=( A302  and  (not A300) );
 a68747a <=( a68746a  and  a68743a );
 a68748a <=( a68747a  and  a68740a );
 a68752a <=( (not A199)  and  A166 );
 a68753a <=( A167  and  a68752a );
 a68756a <=( (not A201)  and  A200 );
 a68759a <=( (not A265)  and  (not A203) );
 a68760a <=( a68759a  and  a68756a );
 a68761a <=( a68760a  and  a68753a );
 a68765a <=( (not A269)  and  A268 );
 a68766a <=( (not A266)  and  a68765a );
 a68769a <=( (not A299)  and  A298 );
 a68772a <=( A301  and  (not A300) );
 a68773a <=( a68772a  and  a68769a );
 a68774a <=( a68773a  and  a68766a );
 a68778a <=( (not A199)  and  A166 );
 a68779a <=( A167  and  a68778a );
 a68782a <=( (not A201)  and  A200 );
 a68785a <=( (not A265)  and  (not A203) );
 a68786a <=( a68785a  and  a68782a );
 a68787a <=( a68786a  and  a68779a );
 a68791a <=( (not A269)  and  A268 );
 a68792a <=( (not A266)  and  a68791a );
 a68795a <=( (not A299)  and  A298 );
 a68798a <=( (not A302)  and  (not A300) );
 a68799a <=( a68798a  and  a68795a );
 a68800a <=( a68799a  and  a68792a );
 a68804a <=( (not A199)  and  A166 );
 a68805a <=( A167  and  a68804a );
 a68808a <=( (not A201)  and  A200 );
 a68811a <=( (not A265)  and  (not A203) );
 a68812a <=( a68811a  and  a68808a );
 a68813a <=( a68812a  and  a68805a );
 a68817a <=( (not A269)  and  A268 );
 a68818a <=( (not A266)  and  a68817a );
 a68821a <=( A299  and  (not A298) );
 a68824a <=( A301  and  (not A300) );
 a68825a <=( a68824a  and  a68821a );
 a68826a <=( a68825a  and  a68818a );
 a68830a <=( (not A199)  and  A166 );
 a68831a <=( A167  and  a68830a );
 a68834a <=( (not A201)  and  A200 );
 a68837a <=( (not A265)  and  (not A203) );
 a68838a <=( a68837a  and  a68834a );
 a68839a <=( a68838a  and  a68831a );
 a68843a <=( (not A269)  and  A268 );
 a68844a <=( (not A266)  and  a68843a );
 a68847a <=( A299  and  (not A298) );
 a68850a <=( (not A302)  and  (not A300) );
 a68851a <=( a68850a  and  a68847a );
 a68852a <=( a68851a  and  a68844a );
 a68856a <=( A199  and  A166 );
 a68857a <=( A167  and  a68856a );
 a68860a <=( (not A202)  and  (not A200) );
 a68863a <=( A265  and  A203 );
 a68864a <=( a68863a  and  a68860a );
 a68865a <=( a68864a  and  a68857a );
 a68869a <=( (not A268)  and  (not A267) );
 a68870a <=( A266  and  a68869a );
 a68873a <=( A299  and  A298 );
 a68876a <=( (not A302)  and  A301 );
 a68877a <=( a68876a  and  a68873a );
 a68878a <=( a68877a  and  a68870a );
 a68882a <=( A199  and  A166 );
 a68883a <=( A167  and  a68882a );
 a68886a <=( (not A202)  and  (not A200) );
 a68889a <=( A265  and  A203 );
 a68890a <=( a68889a  and  a68886a );
 a68891a <=( a68890a  and  a68883a );
 a68895a <=( (not A268)  and  (not A267) );
 a68896a <=( A266  and  a68895a );
 a68899a <=( (not A299)  and  A298 );
 a68902a <=( A302  and  (not A301) );
 a68903a <=( a68902a  and  a68899a );
 a68904a <=( a68903a  and  a68896a );
 a68908a <=( A199  and  A166 );
 a68909a <=( A167  and  a68908a );
 a68912a <=( (not A202)  and  (not A200) );
 a68915a <=( A265  and  A203 );
 a68916a <=( a68915a  and  a68912a );
 a68917a <=( a68916a  and  a68909a );
 a68921a <=( (not A268)  and  (not A267) );
 a68922a <=( A266  and  a68921a );
 a68925a <=( A299  and  (not A298) );
 a68928a <=( A302  and  (not A301) );
 a68929a <=( a68928a  and  a68925a );
 a68930a <=( a68929a  and  a68922a );
 a68934a <=( A199  and  A166 );
 a68935a <=( A167  and  a68934a );
 a68938a <=( (not A202)  and  (not A200) );
 a68941a <=( A265  and  A203 );
 a68942a <=( a68941a  and  a68938a );
 a68943a <=( a68942a  and  a68935a );
 a68947a <=( (not A268)  and  (not A267) );
 a68948a <=( A266  and  a68947a );
 a68951a <=( (not A299)  and  (not A298) );
 a68954a <=( (not A302)  and  A301 );
 a68955a <=( a68954a  and  a68951a );
 a68956a <=( a68955a  and  a68948a );
 a68960a <=( A199  and  A166 );
 a68961a <=( A167  and  a68960a );
 a68964a <=( (not A202)  and  (not A200) );
 a68967a <=( A265  and  A203 );
 a68968a <=( a68967a  and  a68964a );
 a68969a <=( a68968a  and  a68961a );
 a68973a <=( A269  and  (not A267) );
 a68974a <=( A266  and  a68973a );
 a68977a <=( A299  and  A298 );
 a68980a <=( (not A302)  and  A301 );
 a68981a <=( a68980a  and  a68977a );
 a68982a <=( a68981a  and  a68974a );
 a68986a <=( A199  and  A166 );
 a68987a <=( A167  and  a68986a );
 a68990a <=( (not A202)  and  (not A200) );
 a68993a <=( A265  and  A203 );
 a68994a <=( a68993a  and  a68990a );
 a68995a <=( a68994a  and  a68987a );
 a68999a <=( A269  and  (not A267) );
 a69000a <=( A266  and  a68999a );
 a69003a <=( (not A299)  and  A298 );
 a69006a <=( A302  and  (not A301) );
 a69007a <=( a69006a  and  a69003a );
 a69008a <=( a69007a  and  a69000a );
 a69012a <=( A199  and  A166 );
 a69013a <=( A167  and  a69012a );
 a69016a <=( (not A202)  and  (not A200) );
 a69019a <=( A265  and  A203 );
 a69020a <=( a69019a  and  a69016a );
 a69021a <=( a69020a  and  a69013a );
 a69025a <=( A269  and  (not A267) );
 a69026a <=( A266  and  a69025a );
 a69029a <=( A299  and  (not A298) );
 a69032a <=( A302  and  (not A301) );
 a69033a <=( a69032a  and  a69029a );
 a69034a <=( a69033a  and  a69026a );
 a69038a <=( A199  and  A166 );
 a69039a <=( A167  and  a69038a );
 a69042a <=( (not A202)  and  (not A200) );
 a69045a <=( A265  and  A203 );
 a69046a <=( a69045a  and  a69042a );
 a69047a <=( a69046a  and  a69039a );
 a69051a <=( A269  and  (not A267) );
 a69052a <=( A266  and  a69051a );
 a69055a <=( (not A299)  and  (not A298) );
 a69058a <=( (not A302)  and  A301 );
 a69059a <=( a69058a  and  a69055a );
 a69060a <=( a69059a  and  a69052a );
 a69064a <=( A199  and  A166 );
 a69065a <=( A167  and  a69064a );
 a69068a <=( (not A202)  and  (not A200) );
 a69071a <=( (not A265)  and  A203 );
 a69072a <=( a69071a  and  a69068a );
 a69073a <=( a69072a  and  a69065a );
 a69077a <=( A268  and  (not A267) );
 a69078a <=( A266  and  a69077a );
 a69081a <=( A299  and  A298 );
 a69084a <=( (not A302)  and  A301 );
 a69085a <=( a69084a  and  a69081a );
 a69086a <=( a69085a  and  a69078a );
 a69090a <=( A199  and  A166 );
 a69091a <=( A167  and  a69090a );
 a69094a <=( (not A202)  and  (not A200) );
 a69097a <=( (not A265)  and  A203 );
 a69098a <=( a69097a  and  a69094a );
 a69099a <=( a69098a  and  a69091a );
 a69103a <=( A268  and  (not A267) );
 a69104a <=( A266  and  a69103a );
 a69107a <=( (not A299)  and  A298 );
 a69110a <=( A302  and  (not A301) );
 a69111a <=( a69110a  and  a69107a );
 a69112a <=( a69111a  and  a69104a );
 a69116a <=( A199  and  A166 );
 a69117a <=( A167  and  a69116a );
 a69120a <=( (not A202)  and  (not A200) );
 a69123a <=( (not A265)  and  A203 );
 a69124a <=( a69123a  and  a69120a );
 a69125a <=( a69124a  and  a69117a );
 a69129a <=( A268  and  (not A267) );
 a69130a <=( A266  and  a69129a );
 a69133a <=( A299  and  (not A298) );
 a69136a <=( A302  and  (not A301) );
 a69137a <=( a69136a  and  a69133a );
 a69138a <=( a69137a  and  a69130a );
 a69142a <=( A199  and  A166 );
 a69143a <=( A167  and  a69142a );
 a69146a <=( (not A202)  and  (not A200) );
 a69149a <=( (not A265)  and  A203 );
 a69150a <=( a69149a  and  a69146a );
 a69151a <=( a69150a  and  a69143a );
 a69155a <=( A268  and  (not A267) );
 a69156a <=( A266  and  a69155a );
 a69159a <=( (not A299)  and  (not A298) );
 a69162a <=( (not A302)  and  A301 );
 a69163a <=( a69162a  and  a69159a );
 a69164a <=( a69163a  and  a69156a );
 a69168a <=( A199  and  A166 );
 a69169a <=( A167  and  a69168a );
 a69172a <=( (not A202)  and  (not A200) );
 a69175a <=( (not A265)  and  A203 );
 a69176a <=( a69175a  and  a69172a );
 a69177a <=( a69176a  and  a69169a );
 a69181a <=( (not A269)  and  (not A267) );
 a69182a <=( A266  and  a69181a );
 a69185a <=( A299  and  A298 );
 a69188a <=( (not A302)  and  A301 );
 a69189a <=( a69188a  and  a69185a );
 a69190a <=( a69189a  and  a69182a );
 a69194a <=( A199  and  A166 );
 a69195a <=( A167  and  a69194a );
 a69198a <=( (not A202)  and  (not A200) );
 a69201a <=( (not A265)  and  A203 );
 a69202a <=( a69201a  and  a69198a );
 a69203a <=( a69202a  and  a69195a );
 a69207a <=( (not A269)  and  (not A267) );
 a69208a <=( A266  and  a69207a );
 a69211a <=( (not A299)  and  A298 );
 a69214a <=( A302  and  (not A301) );
 a69215a <=( a69214a  and  a69211a );
 a69216a <=( a69215a  and  a69208a );
 a69220a <=( A199  and  A166 );
 a69221a <=( A167  and  a69220a );
 a69224a <=( (not A202)  and  (not A200) );
 a69227a <=( (not A265)  and  A203 );
 a69228a <=( a69227a  and  a69224a );
 a69229a <=( a69228a  and  a69221a );
 a69233a <=( (not A269)  and  (not A267) );
 a69234a <=( A266  and  a69233a );
 a69237a <=( A299  and  (not A298) );
 a69240a <=( A302  and  (not A301) );
 a69241a <=( a69240a  and  a69237a );
 a69242a <=( a69241a  and  a69234a );
 a69246a <=( A199  and  A166 );
 a69247a <=( A167  and  a69246a );
 a69250a <=( (not A202)  and  (not A200) );
 a69253a <=( (not A265)  and  A203 );
 a69254a <=( a69253a  and  a69250a );
 a69255a <=( a69254a  and  a69247a );
 a69259a <=( (not A269)  and  (not A267) );
 a69260a <=( A266  and  a69259a );
 a69263a <=( (not A299)  and  (not A298) );
 a69266a <=( (not A302)  and  A301 );
 a69267a <=( a69266a  and  a69263a );
 a69268a <=( a69267a  and  a69260a );
 a69272a <=( A199  and  A166 );
 a69273a <=( A167  and  a69272a );
 a69276a <=( (not A202)  and  (not A200) );
 a69279a <=( A265  and  A203 );
 a69280a <=( a69279a  and  a69276a );
 a69281a <=( a69280a  and  a69273a );
 a69285a <=( A268  and  (not A267) );
 a69286a <=( (not A266)  and  a69285a );
 a69289a <=( A299  and  A298 );
 a69292a <=( (not A302)  and  A301 );
 a69293a <=( a69292a  and  a69289a );
 a69294a <=( a69293a  and  a69286a );
 a69298a <=( A199  and  A166 );
 a69299a <=( A167  and  a69298a );
 a69302a <=( (not A202)  and  (not A200) );
 a69305a <=( A265  and  A203 );
 a69306a <=( a69305a  and  a69302a );
 a69307a <=( a69306a  and  a69299a );
 a69311a <=( A268  and  (not A267) );
 a69312a <=( (not A266)  and  a69311a );
 a69315a <=( (not A299)  and  A298 );
 a69318a <=( A302  and  (not A301) );
 a69319a <=( a69318a  and  a69315a );
 a69320a <=( a69319a  and  a69312a );
 a69324a <=( A199  and  A166 );
 a69325a <=( A167  and  a69324a );
 a69328a <=( (not A202)  and  (not A200) );
 a69331a <=( A265  and  A203 );
 a69332a <=( a69331a  and  a69328a );
 a69333a <=( a69332a  and  a69325a );
 a69337a <=( A268  and  (not A267) );
 a69338a <=( (not A266)  and  a69337a );
 a69341a <=( A299  and  (not A298) );
 a69344a <=( A302  and  (not A301) );
 a69345a <=( a69344a  and  a69341a );
 a69346a <=( a69345a  and  a69338a );
 a69350a <=( A199  and  A166 );
 a69351a <=( A167  and  a69350a );
 a69354a <=( (not A202)  and  (not A200) );
 a69357a <=( A265  and  A203 );
 a69358a <=( a69357a  and  a69354a );
 a69359a <=( a69358a  and  a69351a );
 a69363a <=( A268  and  (not A267) );
 a69364a <=( (not A266)  and  a69363a );
 a69367a <=( (not A299)  and  (not A298) );
 a69370a <=( (not A302)  and  A301 );
 a69371a <=( a69370a  and  a69367a );
 a69372a <=( a69371a  and  a69364a );
 a69376a <=( A199  and  A166 );
 a69377a <=( A167  and  a69376a );
 a69380a <=( (not A202)  and  (not A200) );
 a69383a <=( A265  and  A203 );
 a69384a <=( a69383a  and  a69380a );
 a69385a <=( a69384a  and  a69377a );
 a69389a <=( (not A269)  and  (not A267) );
 a69390a <=( (not A266)  and  a69389a );
 a69393a <=( A299  and  A298 );
 a69396a <=( (not A302)  and  A301 );
 a69397a <=( a69396a  and  a69393a );
 a69398a <=( a69397a  and  a69390a );
 a69402a <=( A199  and  A166 );
 a69403a <=( A167  and  a69402a );
 a69406a <=( (not A202)  and  (not A200) );
 a69409a <=( A265  and  A203 );
 a69410a <=( a69409a  and  a69406a );
 a69411a <=( a69410a  and  a69403a );
 a69415a <=( (not A269)  and  (not A267) );
 a69416a <=( (not A266)  and  a69415a );
 a69419a <=( (not A299)  and  A298 );
 a69422a <=( A302  and  (not A301) );
 a69423a <=( a69422a  and  a69419a );
 a69424a <=( a69423a  and  a69416a );
 a69428a <=( A199  and  A166 );
 a69429a <=( A167  and  a69428a );
 a69432a <=( (not A202)  and  (not A200) );
 a69435a <=( A265  and  A203 );
 a69436a <=( a69435a  and  a69432a );
 a69437a <=( a69436a  and  a69429a );
 a69441a <=( (not A269)  and  (not A267) );
 a69442a <=( (not A266)  and  a69441a );
 a69445a <=( A299  and  (not A298) );
 a69448a <=( A302  and  (not A301) );
 a69449a <=( a69448a  and  a69445a );
 a69450a <=( a69449a  and  a69442a );
 a69454a <=( A199  and  A166 );
 a69455a <=( A167  and  a69454a );
 a69458a <=( (not A202)  and  (not A200) );
 a69461a <=( A265  and  A203 );
 a69462a <=( a69461a  and  a69458a );
 a69463a <=( a69462a  and  a69455a );
 a69467a <=( (not A269)  and  (not A267) );
 a69468a <=( (not A266)  and  a69467a );
 a69471a <=( (not A299)  and  (not A298) );
 a69474a <=( (not A302)  and  A301 );
 a69475a <=( a69474a  and  a69471a );
 a69476a <=( a69475a  and  a69468a );
 a69480a <=( A199  and  A166 );
 a69481a <=( A167  and  a69480a );
 a69484a <=( (not A201)  and  (not A200) );
 a69487a <=( A265  and  A202 );
 a69488a <=( a69487a  and  a69484a );
 a69489a <=( a69488a  and  a69481a );
 a69493a <=( (not A269)  and  A268 );
 a69494a <=( A266  and  a69493a );
 a69497a <=( A299  and  A298 );
 a69500a <=( (not A301)  and  (not A300) );
 a69501a <=( a69500a  and  a69497a );
 a69502a <=( a69501a  and  a69494a );
 a69506a <=( A199  and  A166 );
 a69507a <=( A167  and  a69506a );
 a69510a <=( (not A201)  and  (not A200) );
 a69513a <=( A265  and  A202 );
 a69514a <=( a69513a  and  a69510a );
 a69515a <=( a69514a  and  a69507a );
 a69519a <=( (not A269)  and  A268 );
 a69520a <=( A266  and  a69519a );
 a69523a <=( A299  and  A298 );
 a69526a <=( A302  and  (not A300) );
 a69527a <=( a69526a  and  a69523a );
 a69528a <=( a69527a  and  a69520a );
 a69532a <=( A199  and  A166 );
 a69533a <=( A167  and  a69532a );
 a69536a <=( (not A201)  and  (not A200) );
 a69539a <=( A265  and  A202 );
 a69540a <=( a69539a  and  a69536a );
 a69541a <=( a69540a  and  a69533a );
 a69545a <=( (not A269)  and  A268 );
 a69546a <=( A266  and  a69545a );
 a69549a <=( (not A299)  and  A298 );
 a69552a <=( A301  and  (not A300) );
 a69553a <=( a69552a  and  a69549a );
 a69554a <=( a69553a  and  a69546a );
 a69558a <=( A199  and  A166 );
 a69559a <=( A167  and  a69558a );
 a69562a <=( (not A201)  and  (not A200) );
 a69565a <=( A265  and  A202 );
 a69566a <=( a69565a  and  a69562a );
 a69567a <=( a69566a  and  a69559a );
 a69571a <=( (not A269)  and  A268 );
 a69572a <=( A266  and  a69571a );
 a69575a <=( (not A299)  and  A298 );
 a69578a <=( (not A302)  and  (not A300) );
 a69579a <=( a69578a  and  a69575a );
 a69580a <=( a69579a  and  a69572a );
 a69584a <=( A199  and  A166 );
 a69585a <=( A167  and  a69584a );
 a69588a <=( (not A201)  and  (not A200) );
 a69591a <=( A265  and  A202 );
 a69592a <=( a69591a  and  a69588a );
 a69593a <=( a69592a  and  a69585a );
 a69597a <=( (not A269)  and  A268 );
 a69598a <=( A266  and  a69597a );
 a69601a <=( A299  and  (not A298) );
 a69604a <=( A301  and  (not A300) );
 a69605a <=( a69604a  and  a69601a );
 a69606a <=( a69605a  and  a69598a );
 a69610a <=( A199  and  A166 );
 a69611a <=( A167  and  a69610a );
 a69614a <=( (not A201)  and  (not A200) );
 a69617a <=( A265  and  A202 );
 a69618a <=( a69617a  and  a69614a );
 a69619a <=( a69618a  and  a69611a );
 a69623a <=( (not A269)  and  A268 );
 a69624a <=( A266  and  a69623a );
 a69627a <=( A299  and  (not A298) );
 a69630a <=( (not A302)  and  (not A300) );
 a69631a <=( a69630a  and  a69627a );
 a69632a <=( a69631a  and  a69624a );
 a69636a <=( A199  and  A166 );
 a69637a <=( A167  and  a69636a );
 a69640a <=( (not A201)  and  (not A200) );
 a69643a <=( (not A265)  and  A202 );
 a69644a <=( a69643a  and  a69640a );
 a69645a <=( a69644a  and  a69637a );
 a69649a <=( A269  and  (not A268) );
 a69650a <=( A266  and  a69649a );
 a69653a <=( A299  and  A298 );
 a69656a <=( (not A301)  and  (not A300) );
 a69657a <=( a69656a  and  a69653a );
 a69658a <=( a69657a  and  a69650a );
 a69662a <=( A199  and  A166 );
 a69663a <=( A167  and  a69662a );
 a69666a <=( (not A201)  and  (not A200) );
 a69669a <=( (not A265)  and  A202 );
 a69670a <=( a69669a  and  a69666a );
 a69671a <=( a69670a  and  a69663a );
 a69675a <=( A269  and  (not A268) );
 a69676a <=( A266  and  a69675a );
 a69679a <=( A299  and  A298 );
 a69682a <=( A302  and  (not A300) );
 a69683a <=( a69682a  and  a69679a );
 a69684a <=( a69683a  and  a69676a );
 a69688a <=( A199  and  A166 );
 a69689a <=( A167  and  a69688a );
 a69692a <=( (not A201)  and  (not A200) );
 a69695a <=( (not A265)  and  A202 );
 a69696a <=( a69695a  and  a69692a );
 a69697a <=( a69696a  and  a69689a );
 a69701a <=( A269  and  (not A268) );
 a69702a <=( A266  and  a69701a );
 a69705a <=( (not A299)  and  A298 );
 a69708a <=( A301  and  (not A300) );
 a69709a <=( a69708a  and  a69705a );
 a69710a <=( a69709a  and  a69702a );
 a69714a <=( A199  and  A166 );
 a69715a <=( A167  and  a69714a );
 a69718a <=( (not A201)  and  (not A200) );
 a69721a <=( (not A265)  and  A202 );
 a69722a <=( a69721a  and  a69718a );
 a69723a <=( a69722a  and  a69715a );
 a69727a <=( A269  and  (not A268) );
 a69728a <=( A266  and  a69727a );
 a69731a <=( (not A299)  and  A298 );
 a69734a <=( (not A302)  and  (not A300) );
 a69735a <=( a69734a  and  a69731a );
 a69736a <=( a69735a  and  a69728a );
 a69740a <=( A199  and  A166 );
 a69741a <=( A167  and  a69740a );
 a69744a <=( (not A201)  and  (not A200) );
 a69747a <=( (not A265)  and  A202 );
 a69748a <=( a69747a  and  a69744a );
 a69749a <=( a69748a  and  a69741a );
 a69753a <=( A269  and  (not A268) );
 a69754a <=( A266  and  a69753a );
 a69757a <=( A299  and  (not A298) );
 a69760a <=( A301  and  (not A300) );
 a69761a <=( a69760a  and  a69757a );
 a69762a <=( a69761a  and  a69754a );
 a69766a <=( A199  and  A166 );
 a69767a <=( A167  and  a69766a );
 a69770a <=( (not A201)  and  (not A200) );
 a69773a <=( (not A265)  and  A202 );
 a69774a <=( a69773a  and  a69770a );
 a69775a <=( a69774a  and  a69767a );
 a69779a <=( A269  and  (not A268) );
 a69780a <=( A266  and  a69779a );
 a69783a <=( A299  and  (not A298) );
 a69786a <=( (not A302)  and  (not A300) );
 a69787a <=( a69786a  and  a69783a );
 a69788a <=( a69787a  and  a69780a );
 a69792a <=( A199  and  A166 );
 a69793a <=( A167  and  a69792a );
 a69796a <=( (not A201)  and  (not A200) );
 a69799a <=( A265  and  A202 );
 a69800a <=( a69799a  and  a69796a );
 a69801a <=( a69800a  and  a69793a );
 a69805a <=( A269  and  (not A268) );
 a69806a <=( (not A266)  and  a69805a );
 a69809a <=( A299  and  A298 );
 a69812a <=( (not A301)  and  (not A300) );
 a69813a <=( a69812a  and  a69809a );
 a69814a <=( a69813a  and  a69806a );
 a69818a <=( A199  and  A166 );
 a69819a <=( A167  and  a69818a );
 a69822a <=( (not A201)  and  (not A200) );
 a69825a <=( A265  and  A202 );
 a69826a <=( a69825a  and  a69822a );
 a69827a <=( a69826a  and  a69819a );
 a69831a <=( A269  and  (not A268) );
 a69832a <=( (not A266)  and  a69831a );
 a69835a <=( A299  and  A298 );
 a69838a <=( A302  and  (not A300) );
 a69839a <=( a69838a  and  a69835a );
 a69840a <=( a69839a  and  a69832a );
 a69844a <=( A199  and  A166 );
 a69845a <=( A167  and  a69844a );
 a69848a <=( (not A201)  and  (not A200) );
 a69851a <=( A265  and  A202 );
 a69852a <=( a69851a  and  a69848a );
 a69853a <=( a69852a  and  a69845a );
 a69857a <=( A269  and  (not A268) );
 a69858a <=( (not A266)  and  a69857a );
 a69861a <=( (not A299)  and  A298 );
 a69864a <=( A301  and  (not A300) );
 a69865a <=( a69864a  and  a69861a );
 a69866a <=( a69865a  and  a69858a );
 a69870a <=( A199  and  A166 );
 a69871a <=( A167  and  a69870a );
 a69874a <=( (not A201)  and  (not A200) );
 a69877a <=( A265  and  A202 );
 a69878a <=( a69877a  and  a69874a );
 a69879a <=( a69878a  and  a69871a );
 a69883a <=( A269  and  (not A268) );
 a69884a <=( (not A266)  and  a69883a );
 a69887a <=( (not A299)  and  A298 );
 a69890a <=( (not A302)  and  (not A300) );
 a69891a <=( a69890a  and  a69887a );
 a69892a <=( a69891a  and  a69884a );
 a69896a <=( A199  and  A166 );
 a69897a <=( A167  and  a69896a );
 a69900a <=( (not A201)  and  (not A200) );
 a69903a <=( A265  and  A202 );
 a69904a <=( a69903a  and  a69900a );
 a69905a <=( a69904a  and  a69897a );
 a69909a <=( A269  and  (not A268) );
 a69910a <=( (not A266)  and  a69909a );
 a69913a <=( A299  and  (not A298) );
 a69916a <=( A301  and  (not A300) );
 a69917a <=( a69916a  and  a69913a );
 a69918a <=( a69917a  and  a69910a );
 a69922a <=( A199  and  A166 );
 a69923a <=( A167  and  a69922a );
 a69926a <=( (not A201)  and  (not A200) );
 a69929a <=( A265  and  A202 );
 a69930a <=( a69929a  and  a69926a );
 a69931a <=( a69930a  and  a69923a );
 a69935a <=( A269  and  (not A268) );
 a69936a <=( (not A266)  and  a69935a );
 a69939a <=( A299  and  (not A298) );
 a69942a <=( (not A302)  and  (not A300) );
 a69943a <=( a69942a  and  a69939a );
 a69944a <=( a69943a  and  a69936a );
 a69948a <=( A199  and  A166 );
 a69949a <=( A167  and  a69948a );
 a69952a <=( (not A201)  and  (not A200) );
 a69955a <=( (not A265)  and  A202 );
 a69956a <=( a69955a  and  a69952a );
 a69957a <=( a69956a  and  a69949a );
 a69961a <=( (not A269)  and  A268 );
 a69962a <=( (not A266)  and  a69961a );
 a69965a <=( A299  and  A298 );
 a69968a <=( (not A301)  and  (not A300) );
 a69969a <=( a69968a  and  a69965a );
 a69970a <=( a69969a  and  a69962a );
 a69974a <=( A199  and  A166 );
 a69975a <=( A167  and  a69974a );
 a69978a <=( (not A201)  and  (not A200) );
 a69981a <=( (not A265)  and  A202 );
 a69982a <=( a69981a  and  a69978a );
 a69983a <=( a69982a  and  a69975a );
 a69987a <=( (not A269)  and  A268 );
 a69988a <=( (not A266)  and  a69987a );
 a69991a <=( A299  and  A298 );
 a69994a <=( A302  and  (not A300) );
 a69995a <=( a69994a  and  a69991a );
 a69996a <=( a69995a  and  a69988a );
 a70000a <=( A199  and  A166 );
 a70001a <=( A167  and  a70000a );
 a70004a <=( (not A201)  and  (not A200) );
 a70007a <=( (not A265)  and  A202 );
 a70008a <=( a70007a  and  a70004a );
 a70009a <=( a70008a  and  a70001a );
 a70013a <=( (not A269)  and  A268 );
 a70014a <=( (not A266)  and  a70013a );
 a70017a <=( (not A299)  and  A298 );
 a70020a <=( A301  and  (not A300) );
 a70021a <=( a70020a  and  a70017a );
 a70022a <=( a70021a  and  a70014a );
 a70026a <=( A199  and  A166 );
 a70027a <=( A167  and  a70026a );
 a70030a <=( (not A201)  and  (not A200) );
 a70033a <=( (not A265)  and  A202 );
 a70034a <=( a70033a  and  a70030a );
 a70035a <=( a70034a  and  a70027a );
 a70039a <=( (not A269)  and  A268 );
 a70040a <=( (not A266)  and  a70039a );
 a70043a <=( (not A299)  and  A298 );
 a70046a <=( (not A302)  and  (not A300) );
 a70047a <=( a70046a  and  a70043a );
 a70048a <=( a70047a  and  a70040a );
 a70052a <=( A199  and  A166 );
 a70053a <=( A167  and  a70052a );
 a70056a <=( (not A201)  and  (not A200) );
 a70059a <=( (not A265)  and  A202 );
 a70060a <=( a70059a  and  a70056a );
 a70061a <=( a70060a  and  a70053a );
 a70065a <=( (not A269)  and  A268 );
 a70066a <=( (not A266)  and  a70065a );
 a70069a <=( A299  and  (not A298) );
 a70072a <=( A301  and  (not A300) );
 a70073a <=( a70072a  and  a70069a );
 a70074a <=( a70073a  and  a70066a );
 a70078a <=( A199  and  A166 );
 a70079a <=( A167  and  a70078a );
 a70082a <=( (not A201)  and  (not A200) );
 a70085a <=( (not A265)  and  A202 );
 a70086a <=( a70085a  and  a70082a );
 a70087a <=( a70086a  and  a70079a );
 a70091a <=( (not A269)  and  A268 );
 a70092a <=( (not A266)  and  a70091a );
 a70095a <=( A299  and  (not A298) );
 a70098a <=( (not A302)  and  (not A300) );
 a70099a <=( a70098a  and  a70095a );
 a70100a <=( a70099a  and  a70092a );
 a70104a <=( A199  and  A166 );
 a70105a <=( A167  and  a70104a );
 a70108a <=( (not A201)  and  (not A200) );
 a70111a <=( A265  and  (not A203) );
 a70112a <=( a70111a  and  a70108a );
 a70113a <=( a70112a  and  a70105a );
 a70117a <=( (not A269)  and  A268 );
 a70118a <=( A266  and  a70117a );
 a70121a <=( A299  and  A298 );
 a70124a <=( (not A301)  and  (not A300) );
 a70125a <=( a70124a  and  a70121a );
 a70126a <=( a70125a  and  a70118a );
 a70130a <=( A199  and  A166 );
 a70131a <=( A167  and  a70130a );
 a70134a <=( (not A201)  and  (not A200) );
 a70137a <=( A265  and  (not A203) );
 a70138a <=( a70137a  and  a70134a );
 a70139a <=( a70138a  and  a70131a );
 a70143a <=( (not A269)  and  A268 );
 a70144a <=( A266  and  a70143a );
 a70147a <=( A299  and  A298 );
 a70150a <=( A302  and  (not A300) );
 a70151a <=( a70150a  and  a70147a );
 a70152a <=( a70151a  and  a70144a );
 a70156a <=( A199  and  A166 );
 a70157a <=( A167  and  a70156a );
 a70160a <=( (not A201)  and  (not A200) );
 a70163a <=( A265  and  (not A203) );
 a70164a <=( a70163a  and  a70160a );
 a70165a <=( a70164a  and  a70157a );
 a70169a <=( (not A269)  and  A268 );
 a70170a <=( A266  and  a70169a );
 a70173a <=( (not A299)  and  A298 );
 a70176a <=( A301  and  (not A300) );
 a70177a <=( a70176a  and  a70173a );
 a70178a <=( a70177a  and  a70170a );
 a70182a <=( A199  and  A166 );
 a70183a <=( A167  and  a70182a );
 a70186a <=( (not A201)  and  (not A200) );
 a70189a <=( A265  and  (not A203) );
 a70190a <=( a70189a  and  a70186a );
 a70191a <=( a70190a  and  a70183a );
 a70195a <=( (not A269)  and  A268 );
 a70196a <=( A266  and  a70195a );
 a70199a <=( (not A299)  and  A298 );
 a70202a <=( (not A302)  and  (not A300) );
 a70203a <=( a70202a  and  a70199a );
 a70204a <=( a70203a  and  a70196a );
 a70208a <=( A199  and  A166 );
 a70209a <=( A167  and  a70208a );
 a70212a <=( (not A201)  and  (not A200) );
 a70215a <=( A265  and  (not A203) );
 a70216a <=( a70215a  and  a70212a );
 a70217a <=( a70216a  and  a70209a );
 a70221a <=( (not A269)  and  A268 );
 a70222a <=( A266  and  a70221a );
 a70225a <=( A299  and  (not A298) );
 a70228a <=( A301  and  (not A300) );
 a70229a <=( a70228a  and  a70225a );
 a70230a <=( a70229a  and  a70222a );
 a70234a <=( A199  and  A166 );
 a70235a <=( A167  and  a70234a );
 a70238a <=( (not A201)  and  (not A200) );
 a70241a <=( A265  and  (not A203) );
 a70242a <=( a70241a  and  a70238a );
 a70243a <=( a70242a  and  a70235a );
 a70247a <=( (not A269)  and  A268 );
 a70248a <=( A266  and  a70247a );
 a70251a <=( A299  and  (not A298) );
 a70254a <=( (not A302)  and  (not A300) );
 a70255a <=( a70254a  and  a70251a );
 a70256a <=( a70255a  and  a70248a );
 a70260a <=( A199  and  A166 );
 a70261a <=( A167  and  a70260a );
 a70264a <=( (not A201)  and  (not A200) );
 a70267a <=( (not A265)  and  (not A203) );
 a70268a <=( a70267a  and  a70264a );
 a70269a <=( a70268a  and  a70261a );
 a70273a <=( A269  and  (not A268) );
 a70274a <=( A266  and  a70273a );
 a70277a <=( A299  and  A298 );
 a70280a <=( (not A301)  and  (not A300) );
 a70281a <=( a70280a  and  a70277a );
 a70282a <=( a70281a  and  a70274a );
 a70286a <=( A199  and  A166 );
 a70287a <=( A167  and  a70286a );
 a70290a <=( (not A201)  and  (not A200) );
 a70293a <=( (not A265)  and  (not A203) );
 a70294a <=( a70293a  and  a70290a );
 a70295a <=( a70294a  and  a70287a );
 a70299a <=( A269  and  (not A268) );
 a70300a <=( A266  and  a70299a );
 a70303a <=( A299  and  A298 );
 a70306a <=( A302  and  (not A300) );
 a70307a <=( a70306a  and  a70303a );
 a70308a <=( a70307a  and  a70300a );
 a70312a <=( A199  and  A166 );
 a70313a <=( A167  and  a70312a );
 a70316a <=( (not A201)  and  (not A200) );
 a70319a <=( (not A265)  and  (not A203) );
 a70320a <=( a70319a  and  a70316a );
 a70321a <=( a70320a  and  a70313a );
 a70325a <=( A269  and  (not A268) );
 a70326a <=( A266  and  a70325a );
 a70329a <=( (not A299)  and  A298 );
 a70332a <=( A301  and  (not A300) );
 a70333a <=( a70332a  and  a70329a );
 a70334a <=( a70333a  and  a70326a );
 a70338a <=( A199  and  A166 );
 a70339a <=( A167  and  a70338a );
 a70342a <=( (not A201)  and  (not A200) );
 a70345a <=( (not A265)  and  (not A203) );
 a70346a <=( a70345a  and  a70342a );
 a70347a <=( a70346a  and  a70339a );
 a70351a <=( A269  and  (not A268) );
 a70352a <=( A266  and  a70351a );
 a70355a <=( (not A299)  and  A298 );
 a70358a <=( (not A302)  and  (not A300) );
 a70359a <=( a70358a  and  a70355a );
 a70360a <=( a70359a  and  a70352a );
 a70364a <=( A199  and  A166 );
 a70365a <=( A167  and  a70364a );
 a70368a <=( (not A201)  and  (not A200) );
 a70371a <=( (not A265)  and  (not A203) );
 a70372a <=( a70371a  and  a70368a );
 a70373a <=( a70372a  and  a70365a );
 a70377a <=( A269  and  (not A268) );
 a70378a <=( A266  and  a70377a );
 a70381a <=( A299  and  (not A298) );
 a70384a <=( A301  and  (not A300) );
 a70385a <=( a70384a  and  a70381a );
 a70386a <=( a70385a  and  a70378a );
 a70390a <=( A199  and  A166 );
 a70391a <=( A167  and  a70390a );
 a70394a <=( (not A201)  and  (not A200) );
 a70397a <=( (not A265)  and  (not A203) );
 a70398a <=( a70397a  and  a70394a );
 a70399a <=( a70398a  and  a70391a );
 a70403a <=( A269  and  (not A268) );
 a70404a <=( A266  and  a70403a );
 a70407a <=( A299  and  (not A298) );
 a70410a <=( (not A302)  and  (not A300) );
 a70411a <=( a70410a  and  a70407a );
 a70412a <=( a70411a  and  a70404a );
 a70416a <=( A199  and  A166 );
 a70417a <=( A167  and  a70416a );
 a70420a <=( (not A201)  and  (not A200) );
 a70423a <=( A265  and  (not A203) );
 a70424a <=( a70423a  and  a70420a );
 a70425a <=( a70424a  and  a70417a );
 a70429a <=( A269  and  (not A268) );
 a70430a <=( (not A266)  and  a70429a );
 a70433a <=( A299  and  A298 );
 a70436a <=( (not A301)  and  (not A300) );
 a70437a <=( a70436a  and  a70433a );
 a70438a <=( a70437a  and  a70430a );
 a70442a <=( A199  and  A166 );
 a70443a <=( A167  and  a70442a );
 a70446a <=( (not A201)  and  (not A200) );
 a70449a <=( A265  and  (not A203) );
 a70450a <=( a70449a  and  a70446a );
 a70451a <=( a70450a  and  a70443a );
 a70455a <=( A269  and  (not A268) );
 a70456a <=( (not A266)  and  a70455a );
 a70459a <=( A299  and  A298 );
 a70462a <=( A302  and  (not A300) );
 a70463a <=( a70462a  and  a70459a );
 a70464a <=( a70463a  and  a70456a );
 a70468a <=( A199  and  A166 );
 a70469a <=( A167  and  a70468a );
 a70472a <=( (not A201)  and  (not A200) );
 a70475a <=( A265  and  (not A203) );
 a70476a <=( a70475a  and  a70472a );
 a70477a <=( a70476a  and  a70469a );
 a70481a <=( A269  and  (not A268) );
 a70482a <=( (not A266)  and  a70481a );
 a70485a <=( (not A299)  and  A298 );
 a70488a <=( A301  and  (not A300) );
 a70489a <=( a70488a  and  a70485a );
 a70490a <=( a70489a  and  a70482a );
 a70494a <=( A199  and  A166 );
 a70495a <=( A167  and  a70494a );
 a70498a <=( (not A201)  and  (not A200) );
 a70501a <=( A265  and  (not A203) );
 a70502a <=( a70501a  and  a70498a );
 a70503a <=( a70502a  and  a70495a );
 a70507a <=( A269  and  (not A268) );
 a70508a <=( (not A266)  and  a70507a );
 a70511a <=( (not A299)  and  A298 );
 a70514a <=( (not A302)  and  (not A300) );
 a70515a <=( a70514a  and  a70511a );
 a70516a <=( a70515a  and  a70508a );
 a70520a <=( A199  and  A166 );
 a70521a <=( A167  and  a70520a );
 a70524a <=( (not A201)  and  (not A200) );
 a70527a <=( A265  and  (not A203) );
 a70528a <=( a70527a  and  a70524a );
 a70529a <=( a70528a  and  a70521a );
 a70533a <=( A269  and  (not A268) );
 a70534a <=( (not A266)  and  a70533a );
 a70537a <=( A299  and  (not A298) );
 a70540a <=( A301  and  (not A300) );
 a70541a <=( a70540a  and  a70537a );
 a70542a <=( a70541a  and  a70534a );
 a70546a <=( A199  and  A166 );
 a70547a <=( A167  and  a70546a );
 a70550a <=( (not A201)  and  (not A200) );
 a70553a <=( A265  and  (not A203) );
 a70554a <=( a70553a  and  a70550a );
 a70555a <=( a70554a  and  a70547a );
 a70559a <=( A269  and  (not A268) );
 a70560a <=( (not A266)  and  a70559a );
 a70563a <=( A299  and  (not A298) );
 a70566a <=( (not A302)  and  (not A300) );
 a70567a <=( a70566a  and  a70563a );
 a70568a <=( a70567a  and  a70560a );
 a70572a <=( A199  and  A166 );
 a70573a <=( A167  and  a70572a );
 a70576a <=( (not A201)  and  (not A200) );
 a70579a <=( (not A265)  and  (not A203) );
 a70580a <=( a70579a  and  a70576a );
 a70581a <=( a70580a  and  a70573a );
 a70585a <=( (not A269)  and  A268 );
 a70586a <=( (not A266)  and  a70585a );
 a70589a <=( A299  and  A298 );
 a70592a <=( (not A301)  and  (not A300) );
 a70593a <=( a70592a  and  a70589a );
 a70594a <=( a70593a  and  a70586a );
 a70598a <=( A199  and  A166 );
 a70599a <=( A167  and  a70598a );
 a70602a <=( (not A201)  and  (not A200) );
 a70605a <=( (not A265)  and  (not A203) );
 a70606a <=( a70605a  and  a70602a );
 a70607a <=( a70606a  and  a70599a );
 a70611a <=( (not A269)  and  A268 );
 a70612a <=( (not A266)  and  a70611a );
 a70615a <=( A299  and  A298 );
 a70618a <=( A302  and  (not A300) );
 a70619a <=( a70618a  and  a70615a );
 a70620a <=( a70619a  and  a70612a );
 a70624a <=( A199  and  A166 );
 a70625a <=( A167  and  a70624a );
 a70628a <=( (not A201)  and  (not A200) );
 a70631a <=( (not A265)  and  (not A203) );
 a70632a <=( a70631a  and  a70628a );
 a70633a <=( a70632a  and  a70625a );
 a70637a <=( (not A269)  and  A268 );
 a70638a <=( (not A266)  and  a70637a );
 a70641a <=( (not A299)  and  A298 );
 a70644a <=( A301  and  (not A300) );
 a70645a <=( a70644a  and  a70641a );
 a70646a <=( a70645a  and  a70638a );
 a70650a <=( A199  and  A166 );
 a70651a <=( A167  and  a70650a );
 a70654a <=( (not A201)  and  (not A200) );
 a70657a <=( (not A265)  and  (not A203) );
 a70658a <=( a70657a  and  a70654a );
 a70659a <=( a70658a  and  a70651a );
 a70663a <=( (not A269)  and  A268 );
 a70664a <=( (not A266)  and  a70663a );
 a70667a <=( (not A299)  and  A298 );
 a70670a <=( (not A302)  and  (not A300) );
 a70671a <=( a70670a  and  a70667a );
 a70672a <=( a70671a  and  a70664a );
 a70676a <=( A199  and  A166 );
 a70677a <=( A167  and  a70676a );
 a70680a <=( (not A201)  and  (not A200) );
 a70683a <=( (not A265)  and  (not A203) );
 a70684a <=( a70683a  and  a70680a );
 a70685a <=( a70684a  and  a70677a );
 a70689a <=( (not A269)  and  A268 );
 a70690a <=( (not A266)  and  a70689a );
 a70693a <=( A299  and  (not A298) );
 a70696a <=( A301  and  (not A300) );
 a70697a <=( a70696a  and  a70693a );
 a70698a <=( a70697a  and  a70690a );
 a70702a <=( A199  and  A166 );
 a70703a <=( A167  and  a70702a );
 a70706a <=( (not A201)  and  (not A200) );
 a70709a <=( (not A265)  and  (not A203) );
 a70710a <=( a70709a  and  a70706a );
 a70711a <=( a70710a  and  a70703a );
 a70715a <=( (not A269)  and  A268 );
 a70716a <=( (not A266)  and  a70715a );
 a70719a <=( A299  and  (not A298) );
 a70722a <=( (not A302)  and  (not A300) );
 a70723a <=( a70722a  and  a70719a );
 a70724a <=( a70723a  and  a70716a );
 a70728a <=( (not A199)  and  A166 );
 a70729a <=( A167  and  a70728a );
 a70732a <=( A202  and  (not A200) );
 a70735a <=( A265  and  (not A203) );
 a70736a <=( a70735a  and  a70732a );
 a70737a <=( a70736a  and  a70729a );
 a70741a <=( (not A268)  and  (not A267) );
 a70742a <=( A266  and  a70741a );
 a70745a <=( A299  and  A298 );
 a70748a <=( (not A302)  and  A301 );
 a70749a <=( a70748a  and  a70745a );
 a70750a <=( a70749a  and  a70742a );
 a70754a <=( (not A199)  and  A166 );
 a70755a <=( A167  and  a70754a );
 a70758a <=( A202  and  (not A200) );
 a70761a <=( A265  and  (not A203) );
 a70762a <=( a70761a  and  a70758a );
 a70763a <=( a70762a  and  a70755a );
 a70767a <=( (not A268)  and  (not A267) );
 a70768a <=( A266  and  a70767a );
 a70771a <=( (not A299)  and  A298 );
 a70774a <=( A302  and  (not A301) );
 a70775a <=( a70774a  and  a70771a );
 a70776a <=( a70775a  and  a70768a );
 a70780a <=( (not A199)  and  A166 );
 a70781a <=( A167  and  a70780a );
 a70784a <=( A202  and  (not A200) );
 a70787a <=( A265  and  (not A203) );
 a70788a <=( a70787a  and  a70784a );
 a70789a <=( a70788a  and  a70781a );
 a70793a <=( (not A268)  and  (not A267) );
 a70794a <=( A266  and  a70793a );
 a70797a <=( A299  and  (not A298) );
 a70800a <=( A302  and  (not A301) );
 a70801a <=( a70800a  and  a70797a );
 a70802a <=( a70801a  and  a70794a );
 a70806a <=( (not A199)  and  A166 );
 a70807a <=( A167  and  a70806a );
 a70810a <=( A202  and  (not A200) );
 a70813a <=( A265  and  (not A203) );
 a70814a <=( a70813a  and  a70810a );
 a70815a <=( a70814a  and  a70807a );
 a70819a <=( (not A268)  and  (not A267) );
 a70820a <=( A266  and  a70819a );
 a70823a <=( (not A299)  and  (not A298) );
 a70826a <=( (not A302)  and  A301 );
 a70827a <=( a70826a  and  a70823a );
 a70828a <=( a70827a  and  a70820a );
 a70832a <=( (not A199)  and  A166 );
 a70833a <=( A167  and  a70832a );
 a70836a <=( A202  and  (not A200) );
 a70839a <=( A265  and  (not A203) );
 a70840a <=( a70839a  and  a70836a );
 a70841a <=( a70840a  and  a70833a );
 a70845a <=( A269  and  (not A267) );
 a70846a <=( A266  and  a70845a );
 a70849a <=( A299  and  A298 );
 a70852a <=( (not A302)  and  A301 );
 a70853a <=( a70852a  and  a70849a );
 a70854a <=( a70853a  and  a70846a );
 a70858a <=( (not A199)  and  A166 );
 a70859a <=( A167  and  a70858a );
 a70862a <=( A202  and  (not A200) );
 a70865a <=( A265  and  (not A203) );
 a70866a <=( a70865a  and  a70862a );
 a70867a <=( a70866a  and  a70859a );
 a70871a <=( A269  and  (not A267) );
 a70872a <=( A266  and  a70871a );
 a70875a <=( (not A299)  and  A298 );
 a70878a <=( A302  and  (not A301) );
 a70879a <=( a70878a  and  a70875a );
 a70880a <=( a70879a  and  a70872a );
 a70884a <=( (not A199)  and  A166 );
 a70885a <=( A167  and  a70884a );
 a70888a <=( A202  and  (not A200) );
 a70891a <=( A265  and  (not A203) );
 a70892a <=( a70891a  and  a70888a );
 a70893a <=( a70892a  and  a70885a );
 a70897a <=( A269  and  (not A267) );
 a70898a <=( A266  and  a70897a );
 a70901a <=( A299  and  (not A298) );
 a70904a <=( A302  and  (not A301) );
 a70905a <=( a70904a  and  a70901a );
 a70906a <=( a70905a  and  a70898a );
 a70910a <=( (not A199)  and  A166 );
 a70911a <=( A167  and  a70910a );
 a70914a <=( A202  and  (not A200) );
 a70917a <=( A265  and  (not A203) );
 a70918a <=( a70917a  and  a70914a );
 a70919a <=( a70918a  and  a70911a );
 a70923a <=( A269  and  (not A267) );
 a70924a <=( A266  and  a70923a );
 a70927a <=( (not A299)  and  (not A298) );
 a70930a <=( (not A302)  and  A301 );
 a70931a <=( a70930a  and  a70927a );
 a70932a <=( a70931a  and  a70924a );
 a70936a <=( (not A199)  and  A166 );
 a70937a <=( A167  and  a70936a );
 a70940a <=( A202  and  (not A200) );
 a70943a <=( (not A265)  and  (not A203) );
 a70944a <=( a70943a  and  a70940a );
 a70945a <=( a70944a  and  a70937a );
 a70949a <=( A268  and  (not A267) );
 a70950a <=( A266  and  a70949a );
 a70953a <=( A299  and  A298 );
 a70956a <=( (not A302)  and  A301 );
 a70957a <=( a70956a  and  a70953a );
 a70958a <=( a70957a  and  a70950a );
 a70962a <=( (not A199)  and  A166 );
 a70963a <=( A167  and  a70962a );
 a70966a <=( A202  and  (not A200) );
 a70969a <=( (not A265)  and  (not A203) );
 a70970a <=( a70969a  and  a70966a );
 a70971a <=( a70970a  and  a70963a );
 a70975a <=( A268  and  (not A267) );
 a70976a <=( A266  and  a70975a );
 a70979a <=( (not A299)  and  A298 );
 a70982a <=( A302  and  (not A301) );
 a70983a <=( a70982a  and  a70979a );
 a70984a <=( a70983a  and  a70976a );
 a70988a <=( (not A199)  and  A166 );
 a70989a <=( A167  and  a70988a );
 a70992a <=( A202  and  (not A200) );
 a70995a <=( (not A265)  and  (not A203) );
 a70996a <=( a70995a  and  a70992a );
 a70997a <=( a70996a  and  a70989a );
 a71001a <=( A268  and  (not A267) );
 a71002a <=( A266  and  a71001a );
 a71005a <=( A299  and  (not A298) );
 a71008a <=( A302  and  (not A301) );
 a71009a <=( a71008a  and  a71005a );
 a71010a <=( a71009a  and  a71002a );
 a71014a <=( (not A199)  and  A166 );
 a71015a <=( A167  and  a71014a );
 a71018a <=( A202  and  (not A200) );
 a71021a <=( (not A265)  and  (not A203) );
 a71022a <=( a71021a  and  a71018a );
 a71023a <=( a71022a  and  a71015a );
 a71027a <=( A268  and  (not A267) );
 a71028a <=( A266  and  a71027a );
 a71031a <=( (not A299)  and  (not A298) );
 a71034a <=( (not A302)  and  A301 );
 a71035a <=( a71034a  and  a71031a );
 a71036a <=( a71035a  and  a71028a );
 a71040a <=( (not A199)  and  A166 );
 a71041a <=( A167  and  a71040a );
 a71044a <=( A202  and  (not A200) );
 a71047a <=( (not A265)  and  (not A203) );
 a71048a <=( a71047a  and  a71044a );
 a71049a <=( a71048a  and  a71041a );
 a71053a <=( (not A269)  and  (not A267) );
 a71054a <=( A266  and  a71053a );
 a71057a <=( A299  and  A298 );
 a71060a <=( (not A302)  and  A301 );
 a71061a <=( a71060a  and  a71057a );
 a71062a <=( a71061a  and  a71054a );
 a71066a <=( (not A199)  and  A166 );
 a71067a <=( A167  and  a71066a );
 a71070a <=( A202  and  (not A200) );
 a71073a <=( (not A265)  and  (not A203) );
 a71074a <=( a71073a  and  a71070a );
 a71075a <=( a71074a  and  a71067a );
 a71079a <=( (not A269)  and  (not A267) );
 a71080a <=( A266  and  a71079a );
 a71083a <=( (not A299)  and  A298 );
 a71086a <=( A302  and  (not A301) );
 a71087a <=( a71086a  and  a71083a );
 a71088a <=( a71087a  and  a71080a );
 a71092a <=( (not A199)  and  A166 );
 a71093a <=( A167  and  a71092a );
 a71096a <=( A202  and  (not A200) );
 a71099a <=( (not A265)  and  (not A203) );
 a71100a <=( a71099a  and  a71096a );
 a71101a <=( a71100a  and  a71093a );
 a71105a <=( (not A269)  and  (not A267) );
 a71106a <=( A266  and  a71105a );
 a71109a <=( A299  and  (not A298) );
 a71112a <=( A302  and  (not A301) );
 a71113a <=( a71112a  and  a71109a );
 a71114a <=( a71113a  and  a71106a );
 a71118a <=( (not A199)  and  A166 );
 a71119a <=( A167  and  a71118a );
 a71122a <=( A202  and  (not A200) );
 a71125a <=( (not A265)  and  (not A203) );
 a71126a <=( a71125a  and  a71122a );
 a71127a <=( a71126a  and  a71119a );
 a71131a <=( (not A269)  and  (not A267) );
 a71132a <=( A266  and  a71131a );
 a71135a <=( (not A299)  and  (not A298) );
 a71138a <=( (not A302)  and  A301 );
 a71139a <=( a71138a  and  a71135a );
 a71140a <=( a71139a  and  a71132a );
 a71144a <=( (not A199)  and  A166 );
 a71145a <=( A167  and  a71144a );
 a71148a <=( A202  and  (not A200) );
 a71151a <=( A265  and  (not A203) );
 a71152a <=( a71151a  and  a71148a );
 a71153a <=( a71152a  and  a71145a );
 a71157a <=( A268  and  (not A267) );
 a71158a <=( (not A266)  and  a71157a );
 a71161a <=( A299  and  A298 );
 a71164a <=( (not A302)  and  A301 );
 a71165a <=( a71164a  and  a71161a );
 a71166a <=( a71165a  and  a71158a );
 a71170a <=( (not A199)  and  A166 );
 a71171a <=( A167  and  a71170a );
 a71174a <=( A202  and  (not A200) );
 a71177a <=( A265  and  (not A203) );
 a71178a <=( a71177a  and  a71174a );
 a71179a <=( a71178a  and  a71171a );
 a71183a <=( A268  and  (not A267) );
 a71184a <=( (not A266)  and  a71183a );
 a71187a <=( (not A299)  and  A298 );
 a71190a <=( A302  and  (not A301) );
 a71191a <=( a71190a  and  a71187a );
 a71192a <=( a71191a  and  a71184a );
 a71196a <=( (not A199)  and  A166 );
 a71197a <=( A167  and  a71196a );
 a71200a <=( A202  and  (not A200) );
 a71203a <=( A265  and  (not A203) );
 a71204a <=( a71203a  and  a71200a );
 a71205a <=( a71204a  and  a71197a );
 a71209a <=( A268  and  (not A267) );
 a71210a <=( (not A266)  and  a71209a );
 a71213a <=( A299  and  (not A298) );
 a71216a <=( A302  and  (not A301) );
 a71217a <=( a71216a  and  a71213a );
 a71218a <=( a71217a  and  a71210a );
 a71222a <=( (not A199)  and  A166 );
 a71223a <=( A167  and  a71222a );
 a71226a <=( A202  and  (not A200) );
 a71229a <=( A265  and  (not A203) );
 a71230a <=( a71229a  and  a71226a );
 a71231a <=( a71230a  and  a71223a );
 a71235a <=( A268  and  (not A267) );
 a71236a <=( (not A266)  and  a71235a );
 a71239a <=( (not A299)  and  (not A298) );
 a71242a <=( (not A302)  and  A301 );
 a71243a <=( a71242a  and  a71239a );
 a71244a <=( a71243a  and  a71236a );
 a71248a <=( (not A199)  and  A166 );
 a71249a <=( A167  and  a71248a );
 a71252a <=( A202  and  (not A200) );
 a71255a <=( A265  and  (not A203) );
 a71256a <=( a71255a  and  a71252a );
 a71257a <=( a71256a  and  a71249a );
 a71261a <=( (not A269)  and  (not A267) );
 a71262a <=( (not A266)  and  a71261a );
 a71265a <=( A299  and  A298 );
 a71268a <=( (not A302)  and  A301 );
 a71269a <=( a71268a  and  a71265a );
 a71270a <=( a71269a  and  a71262a );
 a71274a <=( (not A199)  and  A166 );
 a71275a <=( A167  and  a71274a );
 a71278a <=( A202  and  (not A200) );
 a71281a <=( A265  and  (not A203) );
 a71282a <=( a71281a  and  a71278a );
 a71283a <=( a71282a  and  a71275a );
 a71287a <=( (not A269)  and  (not A267) );
 a71288a <=( (not A266)  and  a71287a );
 a71291a <=( (not A299)  and  A298 );
 a71294a <=( A302  and  (not A301) );
 a71295a <=( a71294a  and  a71291a );
 a71296a <=( a71295a  and  a71288a );
 a71300a <=( (not A199)  and  A166 );
 a71301a <=( A167  and  a71300a );
 a71304a <=( A202  and  (not A200) );
 a71307a <=( A265  and  (not A203) );
 a71308a <=( a71307a  and  a71304a );
 a71309a <=( a71308a  and  a71301a );
 a71313a <=( (not A269)  and  (not A267) );
 a71314a <=( (not A266)  and  a71313a );
 a71317a <=( A299  and  (not A298) );
 a71320a <=( A302  and  (not A301) );
 a71321a <=( a71320a  and  a71317a );
 a71322a <=( a71321a  and  a71314a );
 a71326a <=( (not A199)  and  A166 );
 a71327a <=( A167  and  a71326a );
 a71330a <=( A202  and  (not A200) );
 a71333a <=( A265  and  (not A203) );
 a71334a <=( a71333a  and  a71330a );
 a71335a <=( a71334a  and  a71327a );
 a71339a <=( (not A269)  and  (not A267) );
 a71340a <=( (not A266)  and  a71339a );
 a71343a <=( (not A299)  and  (not A298) );
 a71346a <=( (not A302)  and  A301 );
 a71347a <=( a71346a  and  a71343a );
 a71348a <=( a71347a  and  a71340a );
 a71352a <=( A199  and  (not A166) );
 a71353a <=( A167  and  a71352a );
 a71356a <=( A202  and  A200 );
 a71359a <=( A265  and  (not A203) );
 a71360a <=( a71359a  and  a71356a );
 a71361a <=( a71360a  and  a71353a );
 a71365a <=( (not A269)  and  A268 );
 a71366a <=( A266  and  a71365a );
 a71369a <=( A299  and  A298 );
 a71372a <=( (not A301)  and  (not A300) );
 a71373a <=( a71372a  and  a71369a );
 a71374a <=( a71373a  and  a71366a );
 a71378a <=( A199  and  (not A166) );
 a71379a <=( A167  and  a71378a );
 a71382a <=( A202  and  A200 );
 a71385a <=( A265  and  (not A203) );
 a71386a <=( a71385a  and  a71382a );
 a71387a <=( a71386a  and  a71379a );
 a71391a <=( (not A269)  and  A268 );
 a71392a <=( A266  and  a71391a );
 a71395a <=( A299  and  A298 );
 a71398a <=( A302  and  (not A300) );
 a71399a <=( a71398a  and  a71395a );
 a71400a <=( a71399a  and  a71392a );
 a71404a <=( A199  and  (not A166) );
 a71405a <=( A167  and  a71404a );
 a71408a <=( A202  and  A200 );
 a71411a <=( A265  and  (not A203) );
 a71412a <=( a71411a  and  a71408a );
 a71413a <=( a71412a  and  a71405a );
 a71417a <=( (not A269)  and  A268 );
 a71418a <=( A266  and  a71417a );
 a71421a <=( (not A299)  and  A298 );
 a71424a <=( A301  and  (not A300) );
 a71425a <=( a71424a  and  a71421a );
 a71426a <=( a71425a  and  a71418a );
 a71430a <=( A199  and  (not A166) );
 a71431a <=( A167  and  a71430a );
 a71434a <=( A202  and  A200 );
 a71437a <=( A265  and  (not A203) );
 a71438a <=( a71437a  and  a71434a );
 a71439a <=( a71438a  and  a71431a );
 a71443a <=( (not A269)  and  A268 );
 a71444a <=( A266  and  a71443a );
 a71447a <=( (not A299)  and  A298 );
 a71450a <=( (not A302)  and  (not A300) );
 a71451a <=( a71450a  and  a71447a );
 a71452a <=( a71451a  and  a71444a );
 a71456a <=( A199  and  (not A166) );
 a71457a <=( A167  and  a71456a );
 a71460a <=( A202  and  A200 );
 a71463a <=( A265  and  (not A203) );
 a71464a <=( a71463a  and  a71460a );
 a71465a <=( a71464a  and  a71457a );
 a71469a <=( (not A269)  and  A268 );
 a71470a <=( A266  and  a71469a );
 a71473a <=( A299  and  (not A298) );
 a71476a <=( A301  and  (not A300) );
 a71477a <=( a71476a  and  a71473a );
 a71478a <=( a71477a  and  a71470a );
 a71482a <=( A199  and  (not A166) );
 a71483a <=( A167  and  a71482a );
 a71486a <=( A202  and  A200 );
 a71489a <=( A265  and  (not A203) );
 a71490a <=( a71489a  and  a71486a );
 a71491a <=( a71490a  and  a71483a );
 a71495a <=( (not A269)  and  A268 );
 a71496a <=( A266  and  a71495a );
 a71499a <=( A299  and  (not A298) );
 a71502a <=( (not A302)  and  (not A300) );
 a71503a <=( a71502a  and  a71499a );
 a71504a <=( a71503a  and  a71496a );
 a71508a <=( A199  and  (not A166) );
 a71509a <=( A167  and  a71508a );
 a71512a <=( A202  and  A200 );
 a71515a <=( (not A265)  and  (not A203) );
 a71516a <=( a71515a  and  a71512a );
 a71517a <=( a71516a  and  a71509a );
 a71521a <=( A269  and  (not A268) );
 a71522a <=( A266  and  a71521a );
 a71525a <=( A299  and  A298 );
 a71528a <=( (not A301)  and  (not A300) );
 a71529a <=( a71528a  and  a71525a );
 a71530a <=( a71529a  and  a71522a );
 a71534a <=( A199  and  (not A166) );
 a71535a <=( A167  and  a71534a );
 a71538a <=( A202  and  A200 );
 a71541a <=( (not A265)  and  (not A203) );
 a71542a <=( a71541a  and  a71538a );
 a71543a <=( a71542a  and  a71535a );
 a71547a <=( A269  and  (not A268) );
 a71548a <=( A266  and  a71547a );
 a71551a <=( A299  and  A298 );
 a71554a <=( A302  and  (not A300) );
 a71555a <=( a71554a  and  a71551a );
 a71556a <=( a71555a  and  a71548a );
 a71560a <=( A199  and  (not A166) );
 a71561a <=( A167  and  a71560a );
 a71564a <=( A202  and  A200 );
 a71567a <=( (not A265)  and  (not A203) );
 a71568a <=( a71567a  and  a71564a );
 a71569a <=( a71568a  and  a71561a );
 a71573a <=( A269  and  (not A268) );
 a71574a <=( A266  and  a71573a );
 a71577a <=( (not A299)  and  A298 );
 a71580a <=( A301  and  (not A300) );
 a71581a <=( a71580a  and  a71577a );
 a71582a <=( a71581a  and  a71574a );
 a71586a <=( A199  and  (not A166) );
 a71587a <=( A167  and  a71586a );
 a71590a <=( A202  and  A200 );
 a71593a <=( (not A265)  and  (not A203) );
 a71594a <=( a71593a  and  a71590a );
 a71595a <=( a71594a  and  a71587a );
 a71599a <=( A269  and  (not A268) );
 a71600a <=( A266  and  a71599a );
 a71603a <=( (not A299)  and  A298 );
 a71606a <=( (not A302)  and  (not A300) );
 a71607a <=( a71606a  and  a71603a );
 a71608a <=( a71607a  and  a71600a );
 a71612a <=( A199  and  (not A166) );
 a71613a <=( A167  and  a71612a );
 a71616a <=( A202  and  A200 );
 a71619a <=( (not A265)  and  (not A203) );
 a71620a <=( a71619a  and  a71616a );
 a71621a <=( a71620a  and  a71613a );
 a71625a <=( A269  and  (not A268) );
 a71626a <=( A266  and  a71625a );
 a71629a <=( A299  and  (not A298) );
 a71632a <=( A301  and  (not A300) );
 a71633a <=( a71632a  and  a71629a );
 a71634a <=( a71633a  and  a71626a );
 a71638a <=( A199  and  (not A166) );
 a71639a <=( A167  and  a71638a );
 a71642a <=( A202  and  A200 );
 a71645a <=( (not A265)  and  (not A203) );
 a71646a <=( a71645a  and  a71642a );
 a71647a <=( a71646a  and  a71639a );
 a71651a <=( A269  and  (not A268) );
 a71652a <=( A266  and  a71651a );
 a71655a <=( A299  and  (not A298) );
 a71658a <=( (not A302)  and  (not A300) );
 a71659a <=( a71658a  and  a71655a );
 a71660a <=( a71659a  and  a71652a );
 a71664a <=( A199  and  (not A166) );
 a71665a <=( A167  and  a71664a );
 a71668a <=( A202  and  A200 );
 a71671a <=( A265  and  (not A203) );
 a71672a <=( a71671a  and  a71668a );
 a71673a <=( a71672a  and  a71665a );
 a71677a <=( A269  and  (not A268) );
 a71678a <=( (not A266)  and  a71677a );
 a71681a <=( A299  and  A298 );
 a71684a <=( (not A301)  and  (not A300) );
 a71685a <=( a71684a  and  a71681a );
 a71686a <=( a71685a  and  a71678a );
 a71690a <=( A199  and  (not A166) );
 a71691a <=( A167  and  a71690a );
 a71694a <=( A202  and  A200 );
 a71697a <=( A265  and  (not A203) );
 a71698a <=( a71697a  and  a71694a );
 a71699a <=( a71698a  and  a71691a );
 a71703a <=( A269  and  (not A268) );
 a71704a <=( (not A266)  and  a71703a );
 a71707a <=( A299  and  A298 );
 a71710a <=( A302  and  (not A300) );
 a71711a <=( a71710a  and  a71707a );
 a71712a <=( a71711a  and  a71704a );
 a71716a <=( A199  and  (not A166) );
 a71717a <=( A167  and  a71716a );
 a71720a <=( A202  and  A200 );
 a71723a <=( A265  and  (not A203) );
 a71724a <=( a71723a  and  a71720a );
 a71725a <=( a71724a  and  a71717a );
 a71729a <=( A269  and  (not A268) );
 a71730a <=( (not A266)  and  a71729a );
 a71733a <=( (not A299)  and  A298 );
 a71736a <=( A301  and  (not A300) );
 a71737a <=( a71736a  and  a71733a );
 a71738a <=( a71737a  and  a71730a );
 a71742a <=( A199  and  (not A166) );
 a71743a <=( A167  and  a71742a );
 a71746a <=( A202  and  A200 );
 a71749a <=( A265  and  (not A203) );
 a71750a <=( a71749a  and  a71746a );
 a71751a <=( a71750a  and  a71743a );
 a71755a <=( A269  and  (not A268) );
 a71756a <=( (not A266)  and  a71755a );
 a71759a <=( (not A299)  and  A298 );
 a71762a <=( (not A302)  and  (not A300) );
 a71763a <=( a71762a  and  a71759a );
 a71764a <=( a71763a  and  a71756a );
 a71768a <=( A199  and  (not A166) );
 a71769a <=( A167  and  a71768a );
 a71772a <=( A202  and  A200 );
 a71775a <=( A265  and  (not A203) );
 a71776a <=( a71775a  and  a71772a );
 a71777a <=( a71776a  and  a71769a );
 a71781a <=( A269  and  (not A268) );
 a71782a <=( (not A266)  and  a71781a );
 a71785a <=( A299  and  (not A298) );
 a71788a <=( A301  and  (not A300) );
 a71789a <=( a71788a  and  a71785a );
 a71790a <=( a71789a  and  a71782a );
 a71794a <=( A199  and  (not A166) );
 a71795a <=( A167  and  a71794a );
 a71798a <=( A202  and  A200 );
 a71801a <=( A265  and  (not A203) );
 a71802a <=( a71801a  and  a71798a );
 a71803a <=( a71802a  and  a71795a );
 a71807a <=( A269  and  (not A268) );
 a71808a <=( (not A266)  and  a71807a );
 a71811a <=( A299  and  (not A298) );
 a71814a <=( (not A302)  and  (not A300) );
 a71815a <=( a71814a  and  a71811a );
 a71816a <=( a71815a  and  a71808a );
 a71820a <=( A199  and  (not A166) );
 a71821a <=( A167  and  a71820a );
 a71824a <=( A202  and  A200 );
 a71827a <=( (not A265)  and  (not A203) );
 a71828a <=( a71827a  and  a71824a );
 a71829a <=( a71828a  and  a71821a );
 a71833a <=( (not A269)  and  A268 );
 a71834a <=( (not A266)  and  a71833a );
 a71837a <=( A299  and  A298 );
 a71840a <=( (not A301)  and  (not A300) );
 a71841a <=( a71840a  and  a71837a );
 a71842a <=( a71841a  and  a71834a );
 a71846a <=( A199  and  (not A166) );
 a71847a <=( A167  and  a71846a );
 a71850a <=( A202  and  A200 );
 a71853a <=( (not A265)  and  (not A203) );
 a71854a <=( a71853a  and  a71850a );
 a71855a <=( a71854a  and  a71847a );
 a71859a <=( (not A269)  and  A268 );
 a71860a <=( (not A266)  and  a71859a );
 a71863a <=( A299  and  A298 );
 a71866a <=( A302  and  (not A300) );
 a71867a <=( a71866a  and  a71863a );
 a71868a <=( a71867a  and  a71860a );
 a71872a <=( A199  and  (not A166) );
 a71873a <=( A167  and  a71872a );
 a71876a <=( A202  and  A200 );
 a71879a <=( (not A265)  and  (not A203) );
 a71880a <=( a71879a  and  a71876a );
 a71881a <=( a71880a  and  a71873a );
 a71885a <=( (not A269)  and  A268 );
 a71886a <=( (not A266)  and  a71885a );
 a71889a <=( (not A299)  and  A298 );
 a71892a <=( A301  and  (not A300) );
 a71893a <=( a71892a  and  a71889a );
 a71894a <=( a71893a  and  a71886a );
 a71898a <=( A199  and  (not A166) );
 a71899a <=( A167  and  a71898a );
 a71902a <=( A202  and  A200 );
 a71905a <=( (not A265)  and  (not A203) );
 a71906a <=( a71905a  and  a71902a );
 a71907a <=( a71906a  and  a71899a );
 a71911a <=( (not A269)  and  A268 );
 a71912a <=( (not A266)  and  a71911a );
 a71915a <=( (not A299)  and  A298 );
 a71918a <=( (not A302)  and  (not A300) );
 a71919a <=( a71918a  and  a71915a );
 a71920a <=( a71919a  and  a71912a );
 a71924a <=( A199  and  (not A166) );
 a71925a <=( A167  and  a71924a );
 a71928a <=( A202  and  A200 );
 a71931a <=( (not A265)  and  (not A203) );
 a71932a <=( a71931a  and  a71928a );
 a71933a <=( a71932a  and  a71925a );
 a71937a <=( (not A269)  and  A268 );
 a71938a <=( (not A266)  and  a71937a );
 a71941a <=( A299  and  (not A298) );
 a71944a <=( A301  and  (not A300) );
 a71945a <=( a71944a  and  a71941a );
 a71946a <=( a71945a  and  a71938a );
 a71950a <=( A199  and  (not A166) );
 a71951a <=( A167  and  a71950a );
 a71954a <=( A202  and  A200 );
 a71957a <=( (not A265)  and  (not A203) );
 a71958a <=( a71957a  and  a71954a );
 a71959a <=( a71958a  and  a71951a );
 a71963a <=( (not A269)  and  A268 );
 a71964a <=( (not A266)  and  a71963a );
 a71967a <=( A299  and  (not A298) );
 a71970a <=( (not A302)  and  (not A300) );
 a71971a <=( a71970a  and  a71967a );
 a71972a <=( a71971a  and  a71964a );
 a71976a <=( A199  and  (not A166) );
 a71977a <=( A167  and  a71976a );
 a71980a <=( (not A201)  and  A200 );
 a71983a <=( A265  and  (not A202) );
 a71984a <=( a71983a  and  a71980a );
 a71985a <=( a71984a  and  a71977a );
 a71989a <=( (not A268)  and  (not A267) );
 a71990a <=( A266  and  a71989a );
 a71993a <=( A299  and  A298 );
 a71996a <=( (not A302)  and  A301 );
 a71997a <=( a71996a  and  a71993a );
 a71998a <=( a71997a  and  a71990a );
 a72002a <=( A199  and  (not A166) );
 a72003a <=( A167  and  a72002a );
 a72006a <=( (not A201)  and  A200 );
 a72009a <=( A265  and  (not A202) );
 a72010a <=( a72009a  and  a72006a );
 a72011a <=( a72010a  and  a72003a );
 a72015a <=( (not A268)  and  (not A267) );
 a72016a <=( A266  and  a72015a );
 a72019a <=( (not A299)  and  A298 );
 a72022a <=( A302  and  (not A301) );
 a72023a <=( a72022a  and  a72019a );
 a72024a <=( a72023a  and  a72016a );
 a72028a <=( A199  and  (not A166) );
 a72029a <=( A167  and  a72028a );
 a72032a <=( (not A201)  and  A200 );
 a72035a <=( A265  and  (not A202) );
 a72036a <=( a72035a  and  a72032a );
 a72037a <=( a72036a  and  a72029a );
 a72041a <=( (not A268)  and  (not A267) );
 a72042a <=( A266  and  a72041a );
 a72045a <=( A299  and  (not A298) );
 a72048a <=( A302  and  (not A301) );
 a72049a <=( a72048a  and  a72045a );
 a72050a <=( a72049a  and  a72042a );
 a72054a <=( A199  and  (not A166) );
 a72055a <=( A167  and  a72054a );
 a72058a <=( (not A201)  and  A200 );
 a72061a <=( A265  and  (not A202) );
 a72062a <=( a72061a  and  a72058a );
 a72063a <=( a72062a  and  a72055a );
 a72067a <=( (not A268)  and  (not A267) );
 a72068a <=( A266  and  a72067a );
 a72071a <=( (not A299)  and  (not A298) );
 a72074a <=( (not A302)  and  A301 );
 a72075a <=( a72074a  and  a72071a );
 a72076a <=( a72075a  and  a72068a );
 a72080a <=( A199  and  (not A166) );
 a72081a <=( A167  and  a72080a );
 a72084a <=( (not A201)  and  A200 );
 a72087a <=( A265  and  (not A202) );
 a72088a <=( a72087a  and  a72084a );
 a72089a <=( a72088a  and  a72081a );
 a72093a <=( A269  and  (not A267) );
 a72094a <=( A266  and  a72093a );
 a72097a <=( A299  and  A298 );
 a72100a <=( (not A302)  and  A301 );
 a72101a <=( a72100a  and  a72097a );
 a72102a <=( a72101a  and  a72094a );
 a72106a <=( A199  and  (not A166) );
 a72107a <=( A167  and  a72106a );
 a72110a <=( (not A201)  and  A200 );
 a72113a <=( A265  and  (not A202) );
 a72114a <=( a72113a  and  a72110a );
 a72115a <=( a72114a  and  a72107a );
 a72119a <=( A269  and  (not A267) );
 a72120a <=( A266  and  a72119a );
 a72123a <=( (not A299)  and  A298 );
 a72126a <=( A302  and  (not A301) );
 a72127a <=( a72126a  and  a72123a );
 a72128a <=( a72127a  and  a72120a );
 a72132a <=( A199  and  (not A166) );
 a72133a <=( A167  and  a72132a );
 a72136a <=( (not A201)  and  A200 );
 a72139a <=( A265  and  (not A202) );
 a72140a <=( a72139a  and  a72136a );
 a72141a <=( a72140a  and  a72133a );
 a72145a <=( A269  and  (not A267) );
 a72146a <=( A266  and  a72145a );
 a72149a <=( A299  and  (not A298) );
 a72152a <=( A302  and  (not A301) );
 a72153a <=( a72152a  and  a72149a );
 a72154a <=( a72153a  and  a72146a );
 a72158a <=( A199  and  (not A166) );
 a72159a <=( A167  and  a72158a );
 a72162a <=( (not A201)  and  A200 );
 a72165a <=( A265  and  (not A202) );
 a72166a <=( a72165a  and  a72162a );
 a72167a <=( a72166a  and  a72159a );
 a72171a <=( A269  and  (not A267) );
 a72172a <=( A266  and  a72171a );
 a72175a <=( (not A299)  and  (not A298) );
 a72178a <=( (not A302)  and  A301 );
 a72179a <=( a72178a  and  a72175a );
 a72180a <=( a72179a  and  a72172a );
 a72184a <=( A199  and  (not A166) );
 a72185a <=( A167  and  a72184a );
 a72188a <=( (not A201)  and  A200 );
 a72191a <=( (not A265)  and  (not A202) );
 a72192a <=( a72191a  and  a72188a );
 a72193a <=( a72192a  and  a72185a );
 a72197a <=( A268  and  (not A267) );
 a72198a <=( A266  and  a72197a );
 a72201a <=( A299  and  A298 );
 a72204a <=( (not A302)  and  A301 );
 a72205a <=( a72204a  and  a72201a );
 a72206a <=( a72205a  and  a72198a );
 a72210a <=( A199  and  (not A166) );
 a72211a <=( A167  and  a72210a );
 a72214a <=( (not A201)  and  A200 );
 a72217a <=( (not A265)  and  (not A202) );
 a72218a <=( a72217a  and  a72214a );
 a72219a <=( a72218a  and  a72211a );
 a72223a <=( A268  and  (not A267) );
 a72224a <=( A266  and  a72223a );
 a72227a <=( (not A299)  and  A298 );
 a72230a <=( A302  and  (not A301) );
 a72231a <=( a72230a  and  a72227a );
 a72232a <=( a72231a  and  a72224a );
 a72236a <=( A199  and  (not A166) );
 a72237a <=( A167  and  a72236a );
 a72240a <=( (not A201)  and  A200 );
 a72243a <=( (not A265)  and  (not A202) );
 a72244a <=( a72243a  and  a72240a );
 a72245a <=( a72244a  and  a72237a );
 a72249a <=( A268  and  (not A267) );
 a72250a <=( A266  and  a72249a );
 a72253a <=( A299  and  (not A298) );
 a72256a <=( A302  and  (not A301) );
 a72257a <=( a72256a  and  a72253a );
 a72258a <=( a72257a  and  a72250a );
 a72262a <=( A199  and  (not A166) );
 a72263a <=( A167  and  a72262a );
 a72266a <=( (not A201)  and  A200 );
 a72269a <=( (not A265)  and  (not A202) );
 a72270a <=( a72269a  and  a72266a );
 a72271a <=( a72270a  and  a72263a );
 a72275a <=( A268  and  (not A267) );
 a72276a <=( A266  and  a72275a );
 a72279a <=( (not A299)  and  (not A298) );
 a72282a <=( (not A302)  and  A301 );
 a72283a <=( a72282a  and  a72279a );
 a72284a <=( a72283a  and  a72276a );
 a72288a <=( A199  and  (not A166) );
 a72289a <=( A167  and  a72288a );
 a72292a <=( (not A201)  and  A200 );
 a72295a <=( (not A265)  and  (not A202) );
 a72296a <=( a72295a  and  a72292a );
 a72297a <=( a72296a  and  a72289a );
 a72301a <=( (not A269)  and  (not A267) );
 a72302a <=( A266  and  a72301a );
 a72305a <=( A299  and  A298 );
 a72308a <=( (not A302)  and  A301 );
 a72309a <=( a72308a  and  a72305a );
 a72310a <=( a72309a  and  a72302a );
 a72314a <=( A199  and  (not A166) );
 a72315a <=( A167  and  a72314a );
 a72318a <=( (not A201)  and  A200 );
 a72321a <=( (not A265)  and  (not A202) );
 a72322a <=( a72321a  and  a72318a );
 a72323a <=( a72322a  and  a72315a );
 a72327a <=( (not A269)  and  (not A267) );
 a72328a <=( A266  and  a72327a );
 a72331a <=( (not A299)  and  A298 );
 a72334a <=( A302  and  (not A301) );
 a72335a <=( a72334a  and  a72331a );
 a72336a <=( a72335a  and  a72328a );
 a72340a <=( A199  and  (not A166) );
 a72341a <=( A167  and  a72340a );
 a72344a <=( (not A201)  and  A200 );
 a72347a <=( (not A265)  and  (not A202) );
 a72348a <=( a72347a  and  a72344a );
 a72349a <=( a72348a  and  a72341a );
 a72353a <=( (not A269)  and  (not A267) );
 a72354a <=( A266  and  a72353a );
 a72357a <=( A299  and  (not A298) );
 a72360a <=( A302  and  (not A301) );
 a72361a <=( a72360a  and  a72357a );
 a72362a <=( a72361a  and  a72354a );
 a72366a <=( A199  and  (not A166) );
 a72367a <=( A167  and  a72366a );
 a72370a <=( (not A201)  and  A200 );
 a72373a <=( (not A265)  and  (not A202) );
 a72374a <=( a72373a  and  a72370a );
 a72375a <=( a72374a  and  a72367a );
 a72379a <=( (not A269)  and  (not A267) );
 a72380a <=( A266  and  a72379a );
 a72383a <=( (not A299)  and  (not A298) );
 a72386a <=( (not A302)  and  A301 );
 a72387a <=( a72386a  and  a72383a );
 a72388a <=( a72387a  and  a72380a );
 a72392a <=( A199  and  (not A166) );
 a72393a <=( A167  and  a72392a );
 a72396a <=( (not A201)  and  A200 );
 a72399a <=( A265  and  (not A202) );
 a72400a <=( a72399a  and  a72396a );
 a72401a <=( a72400a  and  a72393a );
 a72405a <=( A268  and  (not A267) );
 a72406a <=( (not A266)  and  a72405a );
 a72409a <=( A299  and  A298 );
 a72412a <=( (not A302)  and  A301 );
 a72413a <=( a72412a  and  a72409a );
 a72414a <=( a72413a  and  a72406a );
 a72418a <=( A199  and  (not A166) );
 a72419a <=( A167  and  a72418a );
 a72422a <=( (not A201)  and  A200 );
 a72425a <=( A265  and  (not A202) );
 a72426a <=( a72425a  and  a72422a );
 a72427a <=( a72426a  and  a72419a );
 a72431a <=( A268  and  (not A267) );
 a72432a <=( (not A266)  and  a72431a );
 a72435a <=( (not A299)  and  A298 );
 a72438a <=( A302  and  (not A301) );
 a72439a <=( a72438a  and  a72435a );
 a72440a <=( a72439a  and  a72432a );
 a72444a <=( A199  and  (not A166) );
 a72445a <=( A167  and  a72444a );
 a72448a <=( (not A201)  and  A200 );
 a72451a <=( A265  and  (not A202) );
 a72452a <=( a72451a  and  a72448a );
 a72453a <=( a72452a  and  a72445a );
 a72457a <=( A268  and  (not A267) );
 a72458a <=( (not A266)  and  a72457a );
 a72461a <=( A299  and  (not A298) );
 a72464a <=( A302  and  (not A301) );
 a72465a <=( a72464a  and  a72461a );
 a72466a <=( a72465a  and  a72458a );
 a72470a <=( A199  and  (not A166) );
 a72471a <=( A167  and  a72470a );
 a72474a <=( (not A201)  and  A200 );
 a72477a <=( A265  and  (not A202) );
 a72478a <=( a72477a  and  a72474a );
 a72479a <=( a72478a  and  a72471a );
 a72483a <=( A268  and  (not A267) );
 a72484a <=( (not A266)  and  a72483a );
 a72487a <=( (not A299)  and  (not A298) );
 a72490a <=( (not A302)  and  A301 );
 a72491a <=( a72490a  and  a72487a );
 a72492a <=( a72491a  and  a72484a );
 a72496a <=( A199  and  (not A166) );
 a72497a <=( A167  and  a72496a );
 a72500a <=( (not A201)  and  A200 );
 a72503a <=( A265  and  (not A202) );
 a72504a <=( a72503a  and  a72500a );
 a72505a <=( a72504a  and  a72497a );
 a72509a <=( (not A269)  and  (not A267) );
 a72510a <=( (not A266)  and  a72509a );
 a72513a <=( A299  and  A298 );
 a72516a <=( (not A302)  and  A301 );
 a72517a <=( a72516a  and  a72513a );
 a72518a <=( a72517a  and  a72510a );
 a72522a <=( A199  and  (not A166) );
 a72523a <=( A167  and  a72522a );
 a72526a <=( (not A201)  and  A200 );
 a72529a <=( A265  and  (not A202) );
 a72530a <=( a72529a  and  a72526a );
 a72531a <=( a72530a  and  a72523a );
 a72535a <=( (not A269)  and  (not A267) );
 a72536a <=( (not A266)  and  a72535a );
 a72539a <=( (not A299)  and  A298 );
 a72542a <=( A302  and  (not A301) );
 a72543a <=( a72542a  and  a72539a );
 a72544a <=( a72543a  and  a72536a );
 a72548a <=( A199  and  (not A166) );
 a72549a <=( A167  and  a72548a );
 a72552a <=( (not A201)  and  A200 );
 a72555a <=( A265  and  (not A202) );
 a72556a <=( a72555a  and  a72552a );
 a72557a <=( a72556a  and  a72549a );
 a72561a <=( (not A269)  and  (not A267) );
 a72562a <=( (not A266)  and  a72561a );
 a72565a <=( A299  and  (not A298) );
 a72568a <=( A302  and  (not A301) );
 a72569a <=( a72568a  and  a72565a );
 a72570a <=( a72569a  and  a72562a );
 a72574a <=( A199  and  (not A166) );
 a72575a <=( A167  and  a72574a );
 a72578a <=( (not A201)  and  A200 );
 a72581a <=( A265  and  (not A202) );
 a72582a <=( a72581a  and  a72578a );
 a72583a <=( a72582a  and  a72575a );
 a72587a <=( (not A269)  and  (not A267) );
 a72588a <=( (not A266)  and  a72587a );
 a72591a <=( (not A299)  and  (not A298) );
 a72594a <=( (not A302)  and  A301 );
 a72595a <=( a72594a  and  a72591a );
 a72596a <=( a72595a  and  a72588a );
 a72600a <=( A199  and  (not A166) );
 a72601a <=( A167  and  a72600a );
 a72604a <=( (not A201)  and  A200 );
 a72607a <=( A265  and  A203 );
 a72608a <=( a72607a  and  a72604a );
 a72609a <=( a72608a  and  a72601a );
 a72613a <=( (not A268)  and  (not A267) );
 a72614a <=( A266  and  a72613a );
 a72617a <=( A299  and  A298 );
 a72620a <=( (not A302)  and  A301 );
 a72621a <=( a72620a  and  a72617a );
 a72622a <=( a72621a  and  a72614a );
 a72626a <=( A199  and  (not A166) );
 a72627a <=( A167  and  a72626a );
 a72630a <=( (not A201)  and  A200 );
 a72633a <=( A265  and  A203 );
 a72634a <=( a72633a  and  a72630a );
 a72635a <=( a72634a  and  a72627a );
 a72639a <=( (not A268)  and  (not A267) );
 a72640a <=( A266  and  a72639a );
 a72643a <=( (not A299)  and  A298 );
 a72646a <=( A302  and  (not A301) );
 a72647a <=( a72646a  and  a72643a );
 a72648a <=( a72647a  and  a72640a );
 a72652a <=( A199  and  (not A166) );
 a72653a <=( A167  and  a72652a );
 a72656a <=( (not A201)  and  A200 );
 a72659a <=( A265  and  A203 );
 a72660a <=( a72659a  and  a72656a );
 a72661a <=( a72660a  and  a72653a );
 a72665a <=( (not A268)  and  (not A267) );
 a72666a <=( A266  and  a72665a );
 a72669a <=( A299  and  (not A298) );
 a72672a <=( A302  and  (not A301) );
 a72673a <=( a72672a  and  a72669a );
 a72674a <=( a72673a  and  a72666a );
 a72678a <=( A199  and  (not A166) );
 a72679a <=( A167  and  a72678a );
 a72682a <=( (not A201)  and  A200 );
 a72685a <=( A265  and  A203 );
 a72686a <=( a72685a  and  a72682a );
 a72687a <=( a72686a  and  a72679a );
 a72691a <=( (not A268)  and  (not A267) );
 a72692a <=( A266  and  a72691a );
 a72695a <=( (not A299)  and  (not A298) );
 a72698a <=( (not A302)  and  A301 );
 a72699a <=( a72698a  and  a72695a );
 a72700a <=( a72699a  and  a72692a );
 a72704a <=( A199  and  (not A166) );
 a72705a <=( A167  and  a72704a );
 a72708a <=( (not A201)  and  A200 );
 a72711a <=( A265  and  A203 );
 a72712a <=( a72711a  and  a72708a );
 a72713a <=( a72712a  and  a72705a );
 a72717a <=( A269  and  (not A267) );
 a72718a <=( A266  and  a72717a );
 a72721a <=( A299  and  A298 );
 a72724a <=( (not A302)  and  A301 );
 a72725a <=( a72724a  and  a72721a );
 a72726a <=( a72725a  and  a72718a );
 a72730a <=( A199  and  (not A166) );
 a72731a <=( A167  and  a72730a );
 a72734a <=( (not A201)  and  A200 );
 a72737a <=( A265  and  A203 );
 a72738a <=( a72737a  and  a72734a );
 a72739a <=( a72738a  and  a72731a );
 a72743a <=( A269  and  (not A267) );
 a72744a <=( A266  and  a72743a );
 a72747a <=( (not A299)  and  A298 );
 a72750a <=( A302  and  (not A301) );
 a72751a <=( a72750a  and  a72747a );
 a72752a <=( a72751a  and  a72744a );
 a72756a <=( A199  and  (not A166) );
 a72757a <=( A167  and  a72756a );
 a72760a <=( (not A201)  and  A200 );
 a72763a <=( A265  and  A203 );
 a72764a <=( a72763a  and  a72760a );
 a72765a <=( a72764a  and  a72757a );
 a72769a <=( A269  and  (not A267) );
 a72770a <=( A266  and  a72769a );
 a72773a <=( A299  and  (not A298) );
 a72776a <=( A302  and  (not A301) );
 a72777a <=( a72776a  and  a72773a );
 a72778a <=( a72777a  and  a72770a );
 a72782a <=( A199  and  (not A166) );
 a72783a <=( A167  and  a72782a );
 a72786a <=( (not A201)  and  A200 );
 a72789a <=( A265  and  A203 );
 a72790a <=( a72789a  and  a72786a );
 a72791a <=( a72790a  and  a72783a );
 a72795a <=( A269  and  (not A267) );
 a72796a <=( A266  and  a72795a );
 a72799a <=( (not A299)  and  (not A298) );
 a72802a <=( (not A302)  and  A301 );
 a72803a <=( a72802a  and  a72799a );
 a72804a <=( a72803a  and  a72796a );
 a72808a <=( A199  and  (not A166) );
 a72809a <=( A167  and  a72808a );
 a72812a <=( (not A201)  and  A200 );
 a72815a <=( (not A265)  and  A203 );
 a72816a <=( a72815a  and  a72812a );
 a72817a <=( a72816a  and  a72809a );
 a72821a <=( A268  and  (not A267) );
 a72822a <=( A266  and  a72821a );
 a72825a <=( A299  and  A298 );
 a72828a <=( (not A302)  and  A301 );
 a72829a <=( a72828a  and  a72825a );
 a72830a <=( a72829a  and  a72822a );
 a72834a <=( A199  and  (not A166) );
 a72835a <=( A167  and  a72834a );
 a72838a <=( (not A201)  and  A200 );
 a72841a <=( (not A265)  and  A203 );
 a72842a <=( a72841a  and  a72838a );
 a72843a <=( a72842a  and  a72835a );
 a72847a <=( A268  and  (not A267) );
 a72848a <=( A266  and  a72847a );
 a72851a <=( (not A299)  and  A298 );
 a72854a <=( A302  and  (not A301) );
 a72855a <=( a72854a  and  a72851a );
 a72856a <=( a72855a  and  a72848a );
 a72860a <=( A199  and  (not A166) );
 a72861a <=( A167  and  a72860a );
 a72864a <=( (not A201)  and  A200 );
 a72867a <=( (not A265)  and  A203 );
 a72868a <=( a72867a  and  a72864a );
 a72869a <=( a72868a  and  a72861a );
 a72873a <=( A268  and  (not A267) );
 a72874a <=( A266  and  a72873a );
 a72877a <=( A299  and  (not A298) );
 a72880a <=( A302  and  (not A301) );
 a72881a <=( a72880a  and  a72877a );
 a72882a <=( a72881a  and  a72874a );
 a72886a <=( A199  and  (not A166) );
 a72887a <=( A167  and  a72886a );
 a72890a <=( (not A201)  and  A200 );
 a72893a <=( (not A265)  and  A203 );
 a72894a <=( a72893a  and  a72890a );
 a72895a <=( a72894a  and  a72887a );
 a72899a <=( A268  and  (not A267) );
 a72900a <=( A266  and  a72899a );
 a72903a <=( (not A299)  and  (not A298) );
 a72906a <=( (not A302)  and  A301 );
 a72907a <=( a72906a  and  a72903a );
 a72908a <=( a72907a  and  a72900a );
 a72912a <=( A199  and  (not A166) );
 a72913a <=( A167  and  a72912a );
 a72916a <=( (not A201)  and  A200 );
 a72919a <=( (not A265)  and  A203 );
 a72920a <=( a72919a  and  a72916a );
 a72921a <=( a72920a  and  a72913a );
 a72925a <=( (not A269)  and  (not A267) );
 a72926a <=( A266  and  a72925a );
 a72929a <=( A299  and  A298 );
 a72932a <=( (not A302)  and  A301 );
 a72933a <=( a72932a  and  a72929a );
 a72934a <=( a72933a  and  a72926a );
 a72938a <=( A199  and  (not A166) );
 a72939a <=( A167  and  a72938a );
 a72942a <=( (not A201)  and  A200 );
 a72945a <=( (not A265)  and  A203 );
 a72946a <=( a72945a  and  a72942a );
 a72947a <=( a72946a  and  a72939a );
 a72951a <=( (not A269)  and  (not A267) );
 a72952a <=( A266  and  a72951a );
 a72955a <=( (not A299)  and  A298 );
 a72958a <=( A302  and  (not A301) );
 a72959a <=( a72958a  and  a72955a );
 a72960a <=( a72959a  and  a72952a );
 a72964a <=( A199  and  (not A166) );
 a72965a <=( A167  and  a72964a );
 a72968a <=( (not A201)  and  A200 );
 a72971a <=( (not A265)  and  A203 );
 a72972a <=( a72971a  and  a72968a );
 a72973a <=( a72972a  and  a72965a );
 a72977a <=( (not A269)  and  (not A267) );
 a72978a <=( A266  and  a72977a );
 a72981a <=( A299  and  (not A298) );
 a72984a <=( A302  and  (not A301) );
 a72985a <=( a72984a  and  a72981a );
 a72986a <=( a72985a  and  a72978a );
 a72990a <=( A199  and  (not A166) );
 a72991a <=( A167  and  a72990a );
 a72994a <=( (not A201)  and  A200 );
 a72997a <=( (not A265)  and  A203 );
 a72998a <=( a72997a  and  a72994a );
 a72999a <=( a72998a  and  a72991a );
 a73003a <=( (not A269)  and  (not A267) );
 a73004a <=( A266  and  a73003a );
 a73007a <=( (not A299)  and  (not A298) );
 a73010a <=( (not A302)  and  A301 );
 a73011a <=( a73010a  and  a73007a );
 a73012a <=( a73011a  and  a73004a );
 a73016a <=( A199  and  (not A166) );
 a73017a <=( A167  and  a73016a );
 a73020a <=( (not A201)  and  A200 );
 a73023a <=( A265  and  A203 );
 a73024a <=( a73023a  and  a73020a );
 a73025a <=( a73024a  and  a73017a );
 a73029a <=( A268  and  (not A267) );
 a73030a <=( (not A266)  and  a73029a );
 a73033a <=( A299  and  A298 );
 a73036a <=( (not A302)  and  A301 );
 a73037a <=( a73036a  and  a73033a );
 a73038a <=( a73037a  and  a73030a );
 a73042a <=( A199  and  (not A166) );
 a73043a <=( A167  and  a73042a );
 a73046a <=( (not A201)  and  A200 );
 a73049a <=( A265  and  A203 );
 a73050a <=( a73049a  and  a73046a );
 a73051a <=( a73050a  and  a73043a );
 a73055a <=( A268  and  (not A267) );
 a73056a <=( (not A266)  and  a73055a );
 a73059a <=( (not A299)  and  A298 );
 a73062a <=( A302  and  (not A301) );
 a73063a <=( a73062a  and  a73059a );
 a73064a <=( a73063a  and  a73056a );
 a73068a <=( A199  and  (not A166) );
 a73069a <=( A167  and  a73068a );
 a73072a <=( (not A201)  and  A200 );
 a73075a <=( A265  and  A203 );
 a73076a <=( a73075a  and  a73072a );
 a73077a <=( a73076a  and  a73069a );
 a73081a <=( A268  and  (not A267) );
 a73082a <=( (not A266)  and  a73081a );
 a73085a <=( A299  and  (not A298) );
 a73088a <=( A302  and  (not A301) );
 a73089a <=( a73088a  and  a73085a );
 a73090a <=( a73089a  and  a73082a );
 a73094a <=( A199  and  (not A166) );
 a73095a <=( A167  and  a73094a );
 a73098a <=( (not A201)  and  A200 );
 a73101a <=( A265  and  A203 );
 a73102a <=( a73101a  and  a73098a );
 a73103a <=( a73102a  and  a73095a );
 a73107a <=( A268  and  (not A267) );
 a73108a <=( (not A266)  and  a73107a );
 a73111a <=( (not A299)  and  (not A298) );
 a73114a <=( (not A302)  and  A301 );
 a73115a <=( a73114a  and  a73111a );
 a73116a <=( a73115a  and  a73108a );
 a73120a <=( A199  and  (not A166) );
 a73121a <=( A167  and  a73120a );
 a73124a <=( (not A201)  and  A200 );
 a73127a <=( A265  and  A203 );
 a73128a <=( a73127a  and  a73124a );
 a73129a <=( a73128a  and  a73121a );
 a73133a <=( (not A269)  and  (not A267) );
 a73134a <=( (not A266)  and  a73133a );
 a73137a <=( A299  and  A298 );
 a73140a <=( (not A302)  and  A301 );
 a73141a <=( a73140a  and  a73137a );
 a73142a <=( a73141a  and  a73134a );
 a73146a <=( A199  and  (not A166) );
 a73147a <=( A167  and  a73146a );
 a73150a <=( (not A201)  and  A200 );
 a73153a <=( A265  and  A203 );
 a73154a <=( a73153a  and  a73150a );
 a73155a <=( a73154a  and  a73147a );
 a73159a <=( (not A269)  and  (not A267) );
 a73160a <=( (not A266)  and  a73159a );
 a73163a <=( (not A299)  and  A298 );
 a73166a <=( A302  and  (not A301) );
 a73167a <=( a73166a  and  a73163a );
 a73168a <=( a73167a  and  a73160a );
 a73172a <=( A199  and  (not A166) );
 a73173a <=( A167  and  a73172a );
 a73176a <=( (not A201)  and  A200 );
 a73179a <=( A265  and  A203 );
 a73180a <=( a73179a  and  a73176a );
 a73181a <=( a73180a  and  a73173a );
 a73185a <=( (not A269)  and  (not A267) );
 a73186a <=( (not A266)  and  a73185a );
 a73189a <=( A299  and  (not A298) );
 a73192a <=( A302  and  (not A301) );
 a73193a <=( a73192a  and  a73189a );
 a73194a <=( a73193a  and  a73186a );
 a73198a <=( A199  and  (not A166) );
 a73199a <=( A167  and  a73198a );
 a73202a <=( (not A201)  and  A200 );
 a73205a <=( A265  and  A203 );
 a73206a <=( a73205a  and  a73202a );
 a73207a <=( a73206a  and  a73199a );
 a73211a <=( (not A269)  and  (not A267) );
 a73212a <=( (not A266)  and  a73211a );
 a73215a <=( (not A299)  and  (not A298) );
 a73218a <=( (not A302)  and  A301 );
 a73219a <=( a73218a  and  a73215a );
 a73220a <=( a73219a  and  a73212a );
 a73224a <=( (not A199)  and  (not A166) );
 a73225a <=( A167  and  a73224a );
 a73228a <=( (not A202)  and  A200 );
 a73231a <=( A265  and  A203 );
 a73232a <=( a73231a  and  a73228a );
 a73233a <=( a73232a  and  a73225a );
 a73237a <=( (not A269)  and  A268 );
 a73238a <=( A266  and  a73237a );
 a73241a <=( A299  and  A298 );
 a73244a <=( (not A301)  and  (not A300) );
 a73245a <=( a73244a  and  a73241a );
 a73246a <=( a73245a  and  a73238a );
 a73250a <=( (not A199)  and  (not A166) );
 a73251a <=( A167  and  a73250a );
 a73254a <=( (not A202)  and  A200 );
 a73257a <=( A265  and  A203 );
 a73258a <=( a73257a  and  a73254a );
 a73259a <=( a73258a  and  a73251a );
 a73263a <=( (not A269)  and  A268 );
 a73264a <=( A266  and  a73263a );
 a73267a <=( A299  and  A298 );
 a73270a <=( A302  and  (not A300) );
 a73271a <=( a73270a  and  a73267a );
 a73272a <=( a73271a  and  a73264a );
 a73276a <=( (not A199)  and  (not A166) );
 a73277a <=( A167  and  a73276a );
 a73280a <=( (not A202)  and  A200 );
 a73283a <=( A265  and  A203 );
 a73284a <=( a73283a  and  a73280a );
 a73285a <=( a73284a  and  a73277a );
 a73289a <=( (not A269)  and  A268 );
 a73290a <=( A266  and  a73289a );
 a73293a <=( (not A299)  and  A298 );
 a73296a <=( A301  and  (not A300) );
 a73297a <=( a73296a  and  a73293a );
 a73298a <=( a73297a  and  a73290a );
 a73302a <=( (not A199)  and  (not A166) );
 a73303a <=( A167  and  a73302a );
 a73306a <=( (not A202)  and  A200 );
 a73309a <=( A265  and  A203 );
 a73310a <=( a73309a  and  a73306a );
 a73311a <=( a73310a  and  a73303a );
 a73315a <=( (not A269)  and  A268 );
 a73316a <=( A266  and  a73315a );
 a73319a <=( (not A299)  and  A298 );
 a73322a <=( (not A302)  and  (not A300) );
 a73323a <=( a73322a  and  a73319a );
 a73324a <=( a73323a  and  a73316a );
 a73328a <=( (not A199)  and  (not A166) );
 a73329a <=( A167  and  a73328a );
 a73332a <=( (not A202)  and  A200 );
 a73335a <=( A265  and  A203 );
 a73336a <=( a73335a  and  a73332a );
 a73337a <=( a73336a  and  a73329a );
 a73341a <=( (not A269)  and  A268 );
 a73342a <=( A266  and  a73341a );
 a73345a <=( A299  and  (not A298) );
 a73348a <=( A301  and  (not A300) );
 a73349a <=( a73348a  and  a73345a );
 a73350a <=( a73349a  and  a73342a );
 a73354a <=( (not A199)  and  (not A166) );
 a73355a <=( A167  and  a73354a );
 a73358a <=( (not A202)  and  A200 );
 a73361a <=( A265  and  A203 );
 a73362a <=( a73361a  and  a73358a );
 a73363a <=( a73362a  and  a73355a );
 a73367a <=( (not A269)  and  A268 );
 a73368a <=( A266  and  a73367a );
 a73371a <=( A299  and  (not A298) );
 a73374a <=( (not A302)  and  (not A300) );
 a73375a <=( a73374a  and  a73371a );
 a73376a <=( a73375a  and  a73368a );
 a73380a <=( (not A199)  and  (not A166) );
 a73381a <=( A167  and  a73380a );
 a73384a <=( (not A202)  and  A200 );
 a73387a <=( (not A265)  and  A203 );
 a73388a <=( a73387a  and  a73384a );
 a73389a <=( a73388a  and  a73381a );
 a73393a <=( A269  and  (not A268) );
 a73394a <=( A266  and  a73393a );
 a73397a <=( A299  and  A298 );
 a73400a <=( (not A301)  and  (not A300) );
 a73401a <=( a73400a  and  a73397a );
 a73402a <=( a73401a  and  a73394a );
 a73406a <=( (not A199)  and  (not A166) );
 a73407a <=( A167  and  a73406a );
 a73410a <=( (not A202)  and  A200 );
 a73413a <=( (not A265)  and  A203 );
 a73414a <=( a73413a  and  a73410a );
 a73415a <=( a73414a  and  a73407a );
 a73419a <=( A269  and  (not A268) );
 a73420a <=( A266  and  a73419a );
 a73423a <=( A299  and  A298 );
 a73426a <=( A302  and  (not A300) );
 a73427a <=( a73426a  and  a73423a );
 a73428a <=( a73427a  and  a73420a );
 a73432a <=( (not A199)  and  (not A166) );
 a73433a <=( A167  and  a73432a );
 a73436a <=( (not A202)  and  A200 );
 a73439a <=( (not A265)  and  A203 );
 a73440a <=( a73439a  and  a73436a );
 a73441a <=( a73440a  and  a73433a );
 a73445a <=( A269  and  (not A268) );
 a73446a <=( A266  and  a73445a );
 a73449a <=( (not A299)  and  A298 );
 a73452a <=( A301  and  (not A300) );
 a73453a <=( a73452a  and  a73449a );
 a73454a <=( a73453a  and  a73446a );
 a73458a <=( (not A199)  and  (not A166) );
 a73459a <=( A167  and  a73458a );
 a73462a <=( (not A202)  and  A200 );
 a73465a <=( (not A265)  and  A203 );
 a73466a <=( a73465a  and  a73462a );
 a73467a <=( a73466a  and  a73459a );
 a73471a <=( A269  and  (not A268) );
 a73472a <=( A266  and  a73471a );
 a73475a <=( (not A299)  and  A298 );
 a73478a <=( (not A302)  and  (not A300) );
 a73479a <=( a73478a  and  a73475a );
 a73480a <=( a73479a  and  a73472a );
 a73484a <=( (not A199)  and  (not A166) );
 a73485a <=( A167  and  a73484a );
 a73488a <=( (not A202)  and  A200 );
 a73491a <=( (not A265)  and  A203 );
 a73492a <=( a73491a  and  a73488a );
 a73493a <=( a73492a  and  a73485a );
 a73497a <=( A269  and  (not A268) );
 a73498a <=( A266  and  a73497a );
 a73501a <=( A299  and  (not A298) );
 a73504a <=( A301  and  (not A300) );
 a73505a <=( a73504a  and  a73501a );
 a73506a <=( a73505a  and  a73498a );
 a73510a <=( (not A199)  and  (not A166) );
 a73511a <=( A167  and  a73510a );
 a73514a <=( (not A202)  and  A200 );
 a73517a <=( (not A265)  and  A203 );
 a73518a <=( a73517a  and  a73514a );
 a73519a <=( a73518a  and  a73511a );
 a73523a <=( A269  and  (not A268) );
 a73524a <=( A266  and  a73523a );
 a73527a <=( A299  and  (not A298) );
 a73530a <=( (not A302)  and  (not A300) );
 a73531a <=( a73530a  and  a73527a );
 a73532a <=( a73531a  and  a73524a );
 a73536a <=( (not A199)  and  (not A166) );
 a73537a <=( A167  and  a73536a );
 a73540a <=( (not A202)  and  A200 );
 a73543a <=( A265  and  A203 );
 a73544a <=( a73543a  and  a73540a );
 a73545a <=( a73544a  and  a73537a );
 a73549a <=( A269  and  (not A268) );
 a73550a <=( (not A266)  and  a73549a );
 a73553a <=( A299  and  A298 );
 a73556a <=( (not A301)  and  (not A300) );
 a73557a <=( a73556a  and  a73553a );
 a73558a <=( a73557a  and  a73550a );
 a73562a <=( (not A199)  and  (not A166) );
 a73563a <=( A167  and  a73562a );
 a73566a <=( (not A202)  and  A200 );
 a73569a <=( A265  and  A203 );
 a73570a <=( a73569a  and  a73566a );
 a73571a <=( a73570a  and  a73563a );
 a73575a <=( A269  and  (not A268) );
 a73576a <=( (not A266)  and  a73575a );
 a73579a <=( A299  and  A298 );
 a73582a <=( A302  and  (not A300) );
 a73583a <=( a73582a  and  a73579a );
 a73584a <=( a73583a  and  a73576a );
 a73588a <=( (not A199)  and  (not A166) );
 a73589a <=( A167  and  a73588a );
 a73592a <=( (not A202)  and  A200 );
 a73595a <=( A265  and  A203 );
 a73596a <=( a73595a  and  a73592a );
 a73597a <=( a73596a  and  a73589a );
 a73601a <=( A269  and  (not A268) );
 a73602a <=( (not A266)  and  a73601a );
 a73605a <=( (not A299)  and  A298 );
 a73608a <=( A301  and  (not A300) );
 a73609a <=( a73608a  and  a73605a );
 a73610a <=( a73609a  and  a73602a );
 a73614a <=( (not A199)  and  (not A166) );
 a73615a <=( A167  and  a73614a );
 a73618a <=( (not A202)  and  A200 );
 a73621a <=( A265  and  A203 );
 a73622a <=( a73621a  and  a73618a );
 a73623a <=( a73622a  and  a73615a );
 a73627a <=( A269  and  (not A268) );
 a73628a <=( (not A266)  and  a73627a );
 a73631a <=( (not A299)  and  A298 );
 a73634a <=( (not A302)  and  (not A300) );
 a73635a <=( a73634a  and  a73631a );
 a73636a <=( a73635a  and  a73628a );
 a73640a <=( (not A199)  and  (not A166) );
 a73641a <=( A167  and  a73640a );
 a73644a <=( (not A202)  and  A200 );
 a73647a <=( A265  and  A203 );
 a73648a <=( a73647a  and  a73644a );
 a73649a <=( a73648a  and  a73641a );
 a73653a <=( A269  and  (not A268) );
 a73654a <=( (not A266)  and  a73653a );
 a73657a <=( A299  and  (not A298) );
 a73660a <=( A301  and  (not A300) );
 a73661a <=( a73660a  and  a73657a );
 a73662a <=( a73661a  and  a73654a );
 a73666a <=( (not A199)  and  (not A166) );
 a73667a <=( A167  and  a73666a );
 a73670a <=( (not A202)  and  A200 );
 a73673a <=( A265  and  A203 );
 a73674a <=( a73673a  and  a73670a );
 a73675a <=( a73674a  and  a73667a );
 a73679a <=( A269  and  (not A268) );
 a73680a <=( (not A266)  and  a73679a );
 a73683a <=( A299  and  (not A298) );
 a73686a <=( (not A302)  and  (not A300) );
 a73687a <=( a73686a  and  a73683a );
 a73688a <=( a73687a  and  a73680a );
 a73692a <=( (not A199)  and  (not A166) );
 a73693a <=( A167  and  a73692a );
 a73696a <=( (not A202)  and  A200 );
 a73699a <=( (not A265)  and  A203 );
 a73700a <=( a73699a  and  a73696a );
 a73701a <=( a73700a  and  a73693a );
 a73705a <=( (not A269)  and  A268 );
 a73706a <=( (not A266)  and  a73705a );
 a73709a <=( A299  and  A298 );
 a73712a <=( (not A301)  and  (not A300) );
 a73713a <=( a73712a  and  a73709a );
 a73714a <=( a73713a  and  a73706a );
 a73718a <=( (not A199)  and  (not A166) );
 a73719a <=( A167  and  a73718a );
 a73722a <=( (not A202)  and  A200 );
 a73725a <=( (not A265)  and  A203 );
 a73726a <=( a73725a  and  a73722a );
 a73727a <=( a73726a  and  a73719a );
 a73731a <=( (not A269)  and  A268 );
 a73732a <=( (not A266)  and  a73731a );
 a73735a <=( A299  and  A298 );
 a73738a <=( A302  and  (not A300) );
 a73739a <=( a73738a  and  a73735a );
 a73740a <=( a73739a  and  a73732a );
 a73744a <=( (not A199)  and  (not A166) );
 a73745a <=( A167  and  a73744a );
 a73748a <=( (not A202)  and  A200 );
 a73751a <=( (not A265)  and  A203 );
 a73752a <=( a73751a  and  a73748a );
 a73753a <=( a73752a  and  a73745a );
 a73757a <=( (not A269)  and  A268 );
 a73758a <=( (not A266)  and  a73757a );
 a73761a <=( (not A299)  and  A298 );
 a73764a <=( A301  and  (not A300) );
 a73765a <=( a73764a  and  a73761a );
 a73766a <=( a73765a  and  a73758a );
 a73770a <=( (not A199)  and  (not A166) );
 a73771a <=( A167  and  a73770a );
 a73774a <=( (not A202)  and  A200 );
 a73777a <=( (not A265)  and  A203 );
 a73778a <=( a73777a  and  a73774a );
 a73779a <=( a73778a  and  a73771a );
 a73783a <=( (not A269)  and  A268 );
 a73784a <=( (not A266)  and  a73783a );
 a73787a <=( (not A299)  and  A298 );
 a73790a <=( (not A302)  and  (not A300) );
 a73791a <=( a73790a  and  a73787a );
 a73792a <=( a73791a  and  a73784a );
 a73796a <=( (not A199)  and  (not A166) );
 a73797a <=( A167  and  a73796a );
 a73800a <=( (not A202)  and  A200 );
 a73803a <=( (not A265)  and  A203 );
 a73804a <=( a73803a  and  a73800a );
 a73805a <=( a73804a  and  a73797a );
 a73809a <=( (not A269)  and  A268 );
 a73810a <=( (not A266)  and  a73809a );
 a73813a <=( A299  and  (not A298) );
 a73816a <=( A301  and  (not A300) );
 a73817a <=( a73816a  and  a73813a );
 a73818a <=( a73817a  and  a73810a );
 a73822a <=( (not A199)  and  (not A166) );
 a73823a <=( A167  and  a73822a );
 a73826a <=( (not A202)  and  A200 );
 a73829a <=( (not A265)  and  A203 );
 a73830a <=( a73829a  and  a73826a );
 a73831a <=( a73830a  and  a73823a );
 a73835a <=( (not A269)  and  A268 );
 a73836a <=( (not A266)  and  a73835a );
 a73839a <=( A299  and  (not A298) );
 a73842a <=( (not A302)  and  (not A300) );
 a73843a <=( a73842a  and  a73839a );
 a73844a <=( a73843a  and  a73836a );
 a73848a <=( (not A199)  and  (not A166) );
 a73849a <=( A167  and  a73848a );
 a73852a <=( (not A201)  and  A200 );
 a73855a <=( A265  and  A202 );
 a73856a <=( a73855a  and  a73852a );
 a73857a <=( a73856a  and  a73849a );
 a73861a <=( (not A268)  and  (not A267) );
 a73862a <=( A266  and  a73861a );
 a73865a <=( A299  and  A298 );
 a73868a <=( (not A302)  and  A301 );
 a73869a <=( a73868a  and  a73865a );
 a73870a <=( a73869a  and  a73862a );
 a73874a <=( (not A199)  and  (not A166) );
 a73875a <=( A167  and  a73874a );
 a73878a <=( (not A201)  and  A200 );
 a73881a <=( A265  and  A202 );
 a73882a <=( a73881a  and  a73878a );
 a73883a <=( a73882a  and  a73875a );
 a73887a <=( (not A268)  and  (not A267) );
 a73888a <=( A266  and  a73887a );
 a73891a <=( (not A299)  and  A298 );
 a73894a <=( A302  and  (not A301) );
 a73895a <=( a73894a  and  a73891a );
 a73896a <=( a73895a  and  a73888a );
 a73900a <=( (not A199)  and  (not A166) );
 a73901a <=( A167  and  a73900a );
 a73904a <=( (not A201)  and  A200 );
 a73907a <=( A265  and  A202 );
 a73908a <=( a73907a  and  a73904a );
 a73909a <=( a73908a  and  a73901a );
 a73913a <=( (not A268)  and  (not A267) );
 a73914a <=( A266  and  a73913a );
 a73917a <=( A299  and  (not A298) );
 a73920a <=( A302  and  (not A301) );
 a73921a <=( a73920a  and  a73917a );
 a73922a <=( a73921a  and  a73914a );
 a73926a <=( (not A199)  and  (not A166) );
 a73927a <=( A167  and  a73926a );
 a73930a <=( (not A201)  and  A200 );
 a73933a <=( A265  and  A202 );
 a73934a <=( a73933a  and  a73930a );
 a73935a <=( a73934a  and  a73927a );
 a73939a <=( (not A268)  and  (not A267) );
 a73940a <=( A266  and  a73939a );
 a73943a <=( (not A299)  and  (not A298) );
 a73946a <=( (not A302)  and  A301 );
 a73947a <=( a73946a  and  a73943a );
 a73948a <=( a73947a  and  a73940a );
 a73952a <=( (not A199)  and  (not A166) );
 a73953a <=( A167  and  a73952a );
 a73956a <=( (not A201)  and  A200 );
 a73959a <=( A265  and  A202 );
 a73960a <=( a73959a  and  a73956a );
 a73961a <=( a73960a  and  a73953a );
 a73965a <=( A269  and  (not A267) );
 a73966a <=( A266  and  a73965a );
 a73969a <=( A299  and  A298 );
 a73972a <=( (not A302)  and  A301 );
 a73973a <=( a73972a  and  a73969a );
 a73974a <=( a73973a  and  a73966a );
 a73978a <=( (not A199)  and  (not A166) );
 a73979a <=( A167  and  a73978a );
 a73982a <=( (not A201)  and  A200 );
 a73985a <=( A265  and  A202 );
 a73986a <=( a73985a  and  a73982a );
 a73987a <=( a73986a  and  a73979a );
 a73991a <=( A269  and  (not A267) );
 a73992a <=( A266  and  a73991a );
 a73995a <=( (not A299)  and  A298 );
 a73998a <=( A302  and  (not A301) );
 a73999a <=( a73998a  and  a73995a );
 a74000a <=( a73999a  and  a73992a );
 a74004a <=( (not A199)  and  (not A166) );
 a74005a <=( A167  and  a74004a );
 a74008a <=( (not A201)  and  A200 );
 a74011a <=( A265  and  A202 );
 a74012a <=( a74011a  and  a74008a );
 a74013a <=( a74012a  and  a74005a );
 a74017a <=( A269  and  (not A267) );
 a74018a <=( A266  and  a74017a );
 a74021a <=( A299  and  (not A298) );
 a74024a <=( A302  and  (not A301) );
 a74025a <=( a74024a  and  a74021a );
 a74026a <=( a74025a  and  a74018a );
 a74030a <=( (not A199)  and  (not A166) );
 a74031a <=( A167  and  a74030a );
 a74034a <=( (not A201)  and  A200 );
 a74037a <=( A265  and  A202 );
 a74038a <=( a74037a  and  a74034a );
 a74039a <=( a74038a  and  a74031a );
 a74043a <=( A269  and  (not A267) );
 a74044a <=( A266  and  a74043a );
 a74047a <=( (not A299)  and  (not A298) );
 a74050a <=( (not A302)  and  A301 );
 a74051a <=( a74050a  and  a74047a );
 a74052a <=( a74051a  and  a74044a );
 a74056a <=( (not A199)  and  (not A166) );
 a74057a <=( A167  and  a74056a );
 a74060a <=( (not A201)  and  A200 );
 a74063a <=( (not A265)  and  A202 );
 a74064a <=( a74063a  and  a74060a );
 a74065a <=( a74064a  and  a74057a );
 a74069a <=( A268  and  (not A267) );
 a74070a <=( A266  and  a74069a );
 a74073a <=( A299  and  A298 );
 a74076a <=( (not A302)  and  A301 );
 a74077a <=( a74076a  and  a74073a );
 a74078a <=( a74077a  and  a74070a );
 a74082a <=( (not A199)  and  (not A166) );
 a74083a <=( A167  and  a74082a );
 a74086a <=( (not A201)  and  A200 );
 a74089a <=( (not A265)  and  A202 );
 a74090a <=( a74089a  and  a74086a );
 a74091a <=( a74090a  and  a74083a );
 a74095a <=( A268  and  (not A267) );
 a74096a <=( A266  and  a74095a );
 a74099a <=( (not A299)  and  A298 );
 a74102a <=( A302  and  (not A301) );
 a74103a <=( a74102a  and  a74099a );
 a74104a <=( a74103a  and  a74096a );
 a74108a <=( (not A199)  and  (not A166) );
 a74109a <=( A167  and  a74108a );
 a74112a <=( (not A201)  and  A200 );
 a74115a <=( (not A265)  and  A202 );
 a74116a <=( a74115a  and  a74112a );
 a74117a <=( a74116a  and  a74109a );
 a74121a <=( A268  and  (not A267) );
 a74122a <=( A266  and  a74121a );
 a74125a <=( A299  and  (not A298) );
 a74128a <=( A302  and  (not A301) );
 a74129a <=( a74128a  and  a74125a );
 a74130a <=( a74129a  and  a74122a );
 a74134a <=( (not A199)  and  (not A166) );
 a74135a <=( A167  and  a74134a );
 a74138a <=( (not A201)  and  A200 );
 a74141a <=( (not A265)  and  A202 );
 a74142a <=( a74141a  and  a74138a );
 a74143a <=( a74142a  and  a74135a );
 a74147a <=( A268  and  (not A267) );
 a74148a <=( A266  and  a74147a );
 a74151a <=( (not A299)  and  (not A298) );
 a74154a <=( (not A302)  and  A301 );
 a74155a <=( a74154a  and  a74151a );
 a74156a <=( a74155a  and  a74148a );
 a74160a <=( (not A199)  and  (not A166) );
 a74161a <=( A167  and  a74160a );
 a74164a <=( (not A201)  and  A200 );
 a74167a <=( (not A265)  and  A202 );
 a74168a <=( a74167a  and  a74164a );
 a74169a <=( a74168a  and  a74161a );
 a74173a <=( (not A269)  and  (not A267) );
 a74174a <=( A266  and  a74173a );
 a74177a <=( A299  and  A298 );
 a74180a <=( (not A302)  and  A301 );
 a74181a <=( a74180a  and  a74177a );
 a74182a <=( a74181a  and  a74174a );
 a74186a <=( (not A199)  and  (not A166) );
 a74187a <=( A167  and  a74186a );
 a74190a <=( (not A201)  and  A200 );
 a74193a <=( (not A265)  and  A202 );
 a74194a <=( a74193a  and  a74190a );
 a74195a <=( a74194a  and  a74187a );
 a74199a <=( (not A269)  and  (not A267) );
 a74200a <=( A266  and  a74199a );
 a74203a <=( (not A299)  and  A298 );
 a74206a <=( A302  and  (not A301) );
 a74207a <=( a74206a  and  a74203a );
 a74208a <=( a74207a  and  a74200a );
 a74212a <=( (not A199)  and  (not A166) );
 a74213a <=( A167  and  a74212a );
 a74216a <=( (not A201)  and  A200 );
 a74219a <=( (not A265)  and  A202 );
 a74220a <=( a74219a  and  a74216a );
 a74221a <=( a74220a  and  a74213a );
 a74225a <=( (not A269)  and  (not A267) );
 a74226a <=( A266  and  a74225a );
 a74229a <=( A299  and  (not A298) );
 a74232a <=( A302  and  (not A301) );
 a74233a <=( a74232a  and  a74229a );
 a74234a <=( a74233a  and  a74226a );
 a74238a <=( (not A199)  and  (not A166) );
 a74239a <=( A167  and  a74238a );
 a74242a <=( (not A201)  and  A200 );
 a74245a <=( (not A265)  and  A202 );
 a74246a <=( a74245a  and  a74242a );
 a74247a <=( a74246a  and  a74239a );
 a74251a <=( (not A269)  and  (not A267) );
 a74252a <=( A266  and  a74251a );
 a74255a <=( (not A299)  and  (not A298) );
 a74258a <=( (not A302)  and  A301 );
 a74259a <=( a74258a  and  a74255a );
 a74260a <=( a74259a  and  a74252a );
 a74264a <=( (not A199)  and  (not A166) );
 a74265a <=( A167  and  a74264a );
 a74268a <=( (not A201)  and  A200 );
 a74271a <=( A265  and  A202 );
 a74272a <=( a74271a  and  a74268a );
 a74273a <=( a74272a  and  a74265a );
 a74277a <=( A268  and  (not A267) );
 a74278a <=( (not A266)  and  a74277a );
 a74281a <=( A299  and  A298 );
 a74284a <=( (not A302)  and  A301 );
 a74285a <=( a74284a  and  a74281a );
 a74286a <=( a74285a  and  a74278a );
 a74290a <=( (not A199)  and  (not A166) );
 a74291a <=( A167  and  a74290a );
 a74294a <=( (not A201)  and  A200 );
 a74297a <=( A265  and  A202 );
 a74298a <=( a74297a  and  a74294a );
 a74299a <=( a74298a  and  a74291a );
 a74303a <=( A268  and  (not A267) );
 a74304a <=( (not A266)  and  a74303a );
 a74307a <=( (not A299)  and  A298 );
 a74310a <=( A302  and  (not A301) );
 a74311a <=( a74310a  and  a74307a );
 a74312a <=( a74311a  and  a74304a );
 a74316a <=( (not A199)  and  (not A166) );
 a74317a <=( A167  and  a74316a );
 a74320a <=( (not A201)  and  A200 );
 a74323a <=( A265  and  A202 );
 a74324a <=( a74323a  and  a74320a );
 a74325a <=( a74324a  and  a74317a );
 a74329a <=( A268  and  (not A267) );
 a74330a <=( (not A266)  and  a74329a );
 a74333a <=( A299  and  (not A298) );
 a74336a <=( A302  and  (not A301) );
 a74337a <=( a74336a  and  a74333a );
 a74338a <=( a74337a  and  a74330a );
 a74342a <=( (not A199)  and  (not A166) );
 a74343a <=( A167  and  a74342a );
 a74346a <=( (not A201)  and  A200 );
 a74349a <=( A265  and  A202 );
 a74350a <=( a74349a  and  a74346a );
 a74351a <=( a74350a  and  a74343a );
 a74355a <=( A268  and  (not A267) );
 a74356a <=( (not A266)  and  a74355a );
 a74359a <=( (not A299)  and  (not A298) );
 a74362a <=( (not A302)  and  A301 );
 a74363a <=( a74362a  and  a74359a );
 a74364a <=( a74363a  and  a74356a );
 a74368a <=( (not A199)  and  (not A166) );
 a74369a <=( A167  and  a74368a );
 a74372a <=( (not A201)  and  A200 );
 a74375a <=( A265  and  A202 );
 a74376a <=( a74375a  and  a74372a );
 a74377a <=( a74376a  and  a74369a );
 a74381a <=( (not A269)  and  (not A267) );
 a74382a <=( (not A266)  and  a74381a );
 a74385a <=( A299  and  A298 );
 a74388a <=( (not A302)  and  A301 );
 a74389a <=( a74388a  and  a74385a );
 a74390a <=( a74389a  and  a74382a );
 a74394a <=( (not A199)  and  (not A166) );
 a74395a <=( A167  and  a74394a );
 a74398a <=( (not A201)  and  A200 );
 a74401a <=( A265  and  A202 );
 a74402a <=( a74401a  and  a74398a );
 a74403a <=( a74402a  and  a74395a );
 a74407a <=( (not A269)  and  (not A267) );
 a74408a <=( (not A266)  and  a74407a );
 a74411a <=( (not A299)  and  A298 );
 a74414a <=( A302  and  (not A301) );
 a74415a <=( a74414a  and  a74411a );
 a74416a <=( a74415a  and  a74408a );
 a74420a <=( (not A199)  and  (not A166) );
 a74421a <=( A167  and  a74420a );
 a74424a <=( (not A201)  and  A200 );
 a74427a <=( A265  and  A202 );
 a74428a <=( a74427a  and  a74424a );
 a74429a <=( a74428a  and  a74421a );
 a74433a <=( (not A269)  and  (not A267) );
 a74434a <=( (not A266)  and  a74433a );
 a74437a <=( A299  and  (not A298) );
 a74440a <=( A302  and  (not A301) );
 a74441a <=( a74440a  and  a74437a );
 a74442a <=( a74441a  and  a74434a );
 a74446a <=( (not A199)  and  (not A166) );
 a74447a <=( A167  and  a74446a );
 a74450a <=( (not A201)  and  A200 );
 a74453a <=( A265  and  A202 );
 a74454a <=( a74453a  and  a74450a );
 a74455a <=( a74454a  and  a74447a );
 a74459a <=( (not A269)  and  (not A267) );
 a74460a <=( (not A266)  and  a74459a );
 a74463a <=( (not A299)  and  (not A298) );
 a74466a <=( (not A302)  and  A301 );
 a74467a <=( a74466a  and  a74463a );
 a74468a <=( a74467a  and  a74460a );
 a74472a <=( (not A199)  and  (not A166) );
 a74473a <=( A167  and  a74472a );
 a74476a <=( (not A201)  and  A200 );
 a74479a <=( A265  and  (not A203) );
 a74480a <=( a74479a  and  a74476a );
 a74481a <=( a74480a  and  a74473a );
 a74485a <=( (not A268)  and  (not A267) );
 a74486a <=( A266  and  a74485a );
 a74489a <=( A299  and  A298 );
 a74492a <=( (not A302)  and  A301 );
 a74493a <=( a74492a  and  a74489a );
 a74494a <=( a74493a  and  a74486a );
 a74498a <=( (not A199)  and  (not A166) );
 a74499a <=( A167  and  a74498a );
 a74502a <=( (not A201)  and  A200 );
 a74505a <=( A265  and  (not A203) );
 a74506a <=( a74505a  and  a74502a );
 a74507a <=( a74506a  and  a74499a );
 a74511a <=( (not A268)  and  (not A267) );
 a74512a <=( A266  and  a74511a );
 a74515a <=( (not A299)  and  A298 );
 a74518a <=( A302  and  (not A301) );
 a74519a <=( a74518a  and  a74515a );
 a74520a <=( a74519a  and  a74512a );
 a74524a <=( (not A199)  and  (not A166) );
 a74525a <=( A167  and  a74524a );
 a74528a <=( (not A201)  and  A200 );
 a74531a <=( A265  and  (not A203) );
 a74532a <=( a74531a  and  a74528a );
 a74533a <=( a74532a  and  a74525a );
 a74537a <=( (not A268)  and  (not A267) );
 a74538a <=( A266  and  a74537a );
 a74541a <=( A299  and  (not A298) );
 a74544a <=( A302  and  (not A301) );
 a74545a <=( a74544a  and  a74541a );
 a74546a <=( a74545a  and  a74538a );
 a74550a <=( (not A199)  and  (not A166) );
 a74551a <=( A167  and  a74550a );
 a74554a <=( (not A201)  and  A200 );
 a74557a <=( A265  and  (not A203) );
 a74558a <=( a74557a  and  a74554a );
 a74559a <=( a74558a  and  a74551a );
 a74563a <=( (not A268)  and  (not A267) );
 a74564a <=( A266  and  a74563a );
 a74567a <=( (not A299)  and  (not A298) );
 a74570a <=( (not A302)  and  A301 );
 a74571a <=( a74570a  and  a74567a );
 a74572a <=( a74571a  and  a74564a );
 a74576a <=( (not A199)  and  (not A166) );
 a74577a <=( A167  and  a74576a );
 a74580a <=( (not A201)  and  A200 );
 a74583a <=( A265  and  (not A203) );
 a74584a <=( a74583a  and  a74580a );
 a74585a <=( a74584a  and  a74577a );
 a74589a <=( A269  and  (not A267) );
 a74590a <=( A266  and  a74589a );
 a74593a <=( A299  and  A298 );
 a74596a <=( (not A302)  and  A301 );
 a74597a <=( a74596a  and  a74593a );
 a74598a <=( a74597a  and  a74590a );
 a74602a <=( (not A199)  and  (not A166) );
 a74603a <=( A167  and  a74602a );
 a74606a <=( (not A201)  and  A200 );
 a74609a <=( A265  and  (not A203) );
 a74610a <=( a74609a  and  a74606a );
 a74611a <=( a74610a  and  a74603a );
 a74615a <=( A269  and  (not A267) );
 a74616a <=( A266  and  a74615a );
 a74619a <=( (not A299)  and  A298 );
 a74622a <=( A302  and  (not A301) );
 a74623a <=( a74622a  and  a74619a );
 a74624a <=( a74623a  and  a74616a );
 a74628a <=( (not A199)  and  (not A166) );
 a74629a <=( A167  and  a74628a );
 a74632a <=( (not A201)  and  A200 );
 a74635a <=( A265  and  (not A203) );
 a74636a <=( a74635a  and  a74632a );
 a74637a <=( a74636a  and  a74629a );
 a74641a <=( A269  and  (not A267) );
 a74642a <=( A266  and  a74641a );
 a74645a <=( A299  and  (not A298) );
 a74648a <=( A302  and  (not A301) );
 a74649a <=( a74648a  and  a74645a );
 a74650a <=( a74649a  and  a74642a );
 a74654a <=( (not A199)  and  (not A166) );
 a74655a <=( A167  and  a74654a );
 a74658a <=( (not A201)  and  A200 );
 a74661a <=( A265  and  (not A203) );
 a74662a <=( a74661a  and  a74658a );
 a74663a <=( a74662a  and  a74655a );
 a74667a <=( A269  and  (not A267) );
 a74668a <=( A266  and  a74667a );
 a74671a <=( (not A299)  and  (not A298) );
 a74674a <=( (not A302)  and  A301 );
 a74675a <=( a74674a  and  a74671a );
 a74676a <=( a74675a  and  a74668a );
 a74680a <=( (not A199)  and  (not A166) );
 a74681a <=( A167  and  a74680a );
 a74684a <=( (not A201)  and  A200 );
 a74687a <=( (not A265)  and  (not A203) );
 a74688a <=( a74687a  and  a74684a );
 a74689a <=( a74688a  and  a74681a );
 a74693a <=( A268  and  (not A267) );
 a74694a <=( A266  and  a74693a );
 a74697a <=( A299  and  A298 );
 a74700a <=( (not A302)  and  A301 );
 a74701a <=( a74700a  and  a74697a );
 a74702a <=( a74701a  and  a74694a );
 a74706a <=( (not A199)  and  (not A166) );
 a74707a <=( A167  and  a74706a );
 a74710a <=( (not A201)  and  A200 );
 a74713a <=( (not A265)  and  (not A203) );
 a74714a <=( a74713a  and  a74710a );
 a74715a <=( a74714a  and  a74707a );
 a74719a <=( A268  and  (not A267) );
 a74720a <=( A266  and  a74719a );
 a74723a <=( (not A299)  and  A298 );
 a74726a <=( A302  and  (not A301) );
 a74727a <=( a74726a  and  a74723a );
 a74728a <=( a74727a  and  a74720a );
 a74732a <=( (not A199)  and  (not A166) );
 a74733a <=( A167  and  a74732a );
 a74736a <=( (not A201)  and  A200 );
 a74739a <=( (not A265)  and  (not A203) );
 a74740a <=( a74739a  and  a74736a );
 a74741a <=( a74740a  and  a74733a );
 a74745a <=( A268  and  (not A267) );
 a74746a <=( A266  and  a74745a );
 a74749a <=( A299  and  (not A298) );
 a74752a <=( A302  and  (not A301) );
 a74753a <=( a74752a  and  a74749a );
 a74754a <=( a74753a  and  a74746a );
 a74758a <=( (not A199)  and  (not A166) );
 a74759a <=( A167  and  a74758a );
 a74762a <=( (not A201)  and  A200 );
 a74765a <=( (not A265)  and  (not A203) );
 a74766a <=( a74765a  and  a74762a );
 a74767a <=( a74766a  and  a74759a );
 a74771a <=( A268  and  (not A267) );
 a74772a <=( A266  and  a74771a );
 a74775a <=( (not A299)  and  (not A298) );
 a74778a <=( (not A302)  and  A301 );
 a74779a <=( a74778a  and  a74775a );
 a74780a <=( a74779a  and  a74772a );
 a74784a <=( (not A199)  and  (not A166) );
 a74785a <=( A167  and  a74784a );
 a74788a <=( (not A201)  and  A200 );
 a74791a <=( (not A265)  and  (not A203) );
 a74792a <=( a74791a  and  a74788a );
 a74793a <=( a74792a  and  a74785a );
 a74797a <=( (not A269)  and  (not A267) );
 a74798a <=( A266  and  a74797a );
 a74801a <=( A299  and  A298 );
 a74804a <=( (not A302)  and  A301 );
 a74805a <=( a74804a  and  a74801a );
 a74806a <=( a74805a  and  a74798a );
 a74810a <=( (not A199)  and  (not A166) );
 a74811a <=( A167  and  a74810a );
 a74814a <=( (not A201)  and  A200 );
 a74817a <=( (not A265)  and  (not A203) );
 a74818a <=( a74817a  and  a74814a );
 a74819a <=( a74818a  and  a74811a );
 a74823a <=( (not A269)  and  (not A267) );
 a74824a <=( A266  and  a74823a );
 a74827a <=( (not A299)  and  A298 );
 a74830a <=( A302  and  (not A301) );
 a74831a <=( a74830a  and  a74827a );
 a74832a <=( a74831a  and  a74824a );
 a74836a <=( (not A199)  and  (not A166) );
 a74837a <=( A167  and  a74836a );
 a74840a <=( (not A201)  and  A200 );
 a74843a <=( (not A265)  and  (not A203) );
 a74844a <=( a74843a  and  a74840a );
 a74845a <=( a74844a  and  a74837a );
 a74849a <=( (not A269)  and  (not A267) );
 a74850a <=( A266  and  a74849a );
 a74853a <=( A299  and  (not A298) );
 a74856a <=( A302  and  (not A301) );
 a74857a <=( a74856a  and  a74853a );
 a74858a <=( a74857a  and  a74850a );
 a74862a <=( (not A199)  and  (not A166) );
 a74863a <=( A167  and  a74862a );
 a74866a <=( (not A201)  and  A200 );
 a74869a <=( (not A265)  and  (not A203) );
 a74870a <=( a74869a  and  a74866a );
 a74871a <=( a74870a  and  a74863a );
 a74875a <=( (not A269)  and  (not A267) );
 a74876a <=( A266  and  a74875a );
 a74879a <=( (not A299)  and  (not A298) );
 a74882a <=( (not A302)  and  A301 );
 a74883a <=( a74882a  and  a74879a );
 a74884a <=( a74883a  and  a74876a );
 a74888a <=( (not A199)  and  (not A166) );
 a74889a <=( A167  and  a74888a );
 a74892a <=( (not A201)  and  A200 );
 a74895a <=( A265  and  (not A203) );
 a74896a <=( a74895a  and  a74892a );
 a74897a <=( a74896a  and  a74889a );
 a74901a <=( A268  and  (not A267) );
 a74902a <=( (not A266)  and  a74901a );
 a74905a <=( A299  and  A298 );
 a74908a <=( (not A302)  and  A301 );
 a74909a <=( a74908a  and  a74905a );
 a74910a <=( a74909a  and  a74902a );
 a74914a <=( (not A199)  and  (not A166) );
 a74915a <=( A167  and  a74914a );
 a74918a <=( (not A201)  and  A200 );
 a74921a <=( A265  and  (not A203) );
 a74922a <=( a74921a  and  a74918a );
 a74923a <=( a74922a  and  a74915a );
 a74927a <=( A268  and  (not A267) );
 a74928a <=( (not A266)  and  a74927a );
 a74931a <=( (not A299)  and  A298 );
 a74934a <=( A302  and  (not A301) );
 a74935a <=( a74934a  and  a74931a );
 a74936a <=( a74935a  and  a74928a );
 a74940a <=( (not A199)  and  (not A166) );
 a74941a <=( A167  and  a74940a );
 a74944a <=( (not A201)  and  A200 );
 a74947a <=( A265  and  (not A203) );
 a74948a <=( a74947a  and  a74944a );
 a74949a <=( a74948a  and  a74941a );
 a74953a <=( A268  and  (not A267) );
 a74954a <=( (not A266)  and  a74953a );
 a74957a <=( A299  and  (not A298) );
 a74960a <=( A302  and  (not A301) );
 a74961a <=( a74960a  and  a74957a );
 a74962a <=( a74961a  and  a74954a );
 a74966a <=( (not A199)  and  (not A166) );
 a74967a <=( A167  and  a74966a );
 a74970a <=( (not A201)  and  A200 );
 a74973a <=( A265  and  (not A203) );
 a74974a <=( a74973a  and  a74970a );
 a74975a <=( a74974a  and  a74967a );
 a74979a <=( A268  and  (not A267) );
 a74980a <=( (not A266)  and  a74979a );
 a74983a <=( (not A299)  and  (not A298) );
 a74986a <=( (not A302)  and  A301 );
 a74987a <=( a74986a  and  a74983a );
 a74988a <=( a74987a  and  a74980a );
 a74992a <=( (not A199)  and  (not A166) );
 a74993a <=( A167  and  a74992a );
 a74996a <=( (not A201)  and  A200 );
 a74999a <=( A265  and  (not A203) );
 a75000a <=( a74999a  and  a74996a );
 a75001a <=( a75000a  and  a74993a );
 a75005a <=( (not A269)  and  (not A267) );
 a75006a <=( (not A266)  and  a75005a );
 a75009a <=( A299  and  A298 );
 a75012a <=( (not A302)  and  A301 );
 a75013a <=( a75012a  and  a75009a );
 a75014a <=( a75013a  and  a75006a );
 a75018a <=( (not A199)  and  (not A166) );
 a75019a <=( A167  and  a75018a );
 a75022a <=( (not A201)  and  A200 );
 a75025a <=( A265  and  (not A203) );
 a75026a <=( a75025a  and  a75022a );
 a75027a <=( a75026a  and  a75019a );
 a75031a <=( (not A269)  and  (not A267) );
 a75032a <=( (not A266)  and  a75031a );
 a75035a <=( (not A299)  and  A298 );
 a75038a <=( A302  and  (not A301) );
 a75039a <=( a75038a  and  a75035a );
 a75040a <=( a75039a  and  a75032a );
 a75044a <=( (not A199)  and  (not A166) );
 a75045a <=( A167  and  a75044a );
 a75048a <=( (not A201)  and  A200 );
 a75051a <=( A265  and  (not A203) );
 a75052a <=( a75051a  and  a75048a );
 a75053a <=( a75052a  and  a75045a );
 a75057a <=( (not A269)  and  (not A267) );
 a75058a <=( (not A266)  and  a75057a );
 a75061a <=( A299  and  (not A298) );
 a75064a <=( A302  and  (not A301) );
 a75065a <=( a75064a  and  a75061a );
 a75066a <=( a75065a  and  a75058a );
 a75070a <=( (not A199)  and  (not A166) );
 a75071a <=( A167  and  a75070a );
 a75074a <=( (not A201)  and  A200 );
 a75077a <=( A265  and  (not A203) );
 a75078a <=( a75077a  and  a75074a );
 a75079a <=( a75078a  and  a75071a );
 a75083a <=( (not A269)  and  (not A267) );
 a75084a <=( (not A266)  and  a75083a );
 a75087a <=( (not A299)  and  (not A298) );
 a75090a <=( (not A302)  and  A301 );
 a75091a <=( a75090a  and  a75087a );
 a75092a <=( a75091a  and  a75084a );
 a75096a <=( A199  and  (not A166) );
 a75097a <=( A167  and  a75096a );
 a75100a <=( (not A202)  and  (not A200) );
 a75103a <=( A265  and  A203 );
 a75104a <=( a75103a  and  a75100a );
 a75105a <=( a75104a  and  a75097a );
 a75109a <=( (not A269)  and  A268 );
 a75110a <=( A266  and  a75109a );
 a75113a <=( A299  and  A298 );
 a75116a <=( (not A301)  and  (not A300) );
 a75117a <=( a75116a  and  a75113a );
 a75118a <=( a75117a  and  a75110a );
 a75122a <=( A199  and  (not A166) );
 a75123a <=( A167  and  a75122a );
 a75126a <=( (not A202)  and  (not A200) );
 a75129a <=( A265  and  A203 );
 a75130a <=( a75129a  and  a75126a );
 a75131a <=( a75130a  and  a75123a );
 a75135a <=( (not A269)  and  A268 );
 a75136a <=( A266  and  a75135a );
 a75139a <=( A299  and  A298 );
 a75142a <=( A302  and  (not A300) );
 a75143a <=( a75142a  and  a75139a );
 a75144a <=( a75143a  and  a75136a );
 a75148a <=( A199  and  (not A166) );
 a75149a <=( A167  and  a75148a );
 a75152a <=( (not A202)  and  (not A200) );
 a75155a <=( A265  and  A203 );
 a75156a <=( a75155a  and  a75152a );
 a75157a <=( a75156a  and  a75149a );
 a75161a <=( (not A269)  and  A268 );
 a75162a <=( A266  and  a75161a );
 a75165a <=( (not A299)  and  A298 );
 a75168a <=( A301  and  (not A300) );
 a75169a <=( a75168a  and  a75165a );
 a75170a <=( a75169a  and  a75162a );
 a75174a <=( A199  and  (not A166) );
 a75175a <=( A167  and  a75174a );
 a75178a <=( (not A202)  and  (not A200) );
 a75181a <=( A265  and  A203 );
 a75182a <=( a75181a  and  a75178a );
 a75183a <=( a75182a  and  a75175a );
 a75187a <=( (not A269)  and  A268 );
 a75188a <=( A266  and  a75187a );
 a75191a <=( (not A299)  and  A298 );
 a75194a <=( (not A302)  and  (not A300) );
 a75195a <=( a75194a  and  a75191a );
 a75196a <=( a75195a  and  a75188a );
 a75200a <=( A199  and  (not A166) );
 a75201a <=( A167  and  a75200a );
 a75204a <=( (not A202)  and  (not A200) );
 a75207a <=( A265  and  A203 );
 a75208a <=( a75207a  and  a75204a );
 a75209a <=( a75208a  and  a75201a );
 a75213a <=( (not A269)  and  A268 );
 a75214a <=( A266  and  a75213a );
 a75217a <=( A299  and  (not A298) );
 a75220a <=( A301  and  (not A300) );
 a75221a <=( a75220a  and  a75217a );
 a75222a <=( a75221a  and  a75214a );
 a75226a <=( A199  and  (not A166) );
 a75227a <=( A167  and  a75226a );
 a75230a <=( (not A202)  and  (not A200) );
 a75233a <=( A265  and  A203 );
 a75234a <=( a75233a  and  a75230a );
 a75235a <=( a75234a  and  a75227a );
 a75239a <=( (not A269)  and  A268 );
 a75240a <=( A266  and  a75239a );
 a75243a <=( A299  and  (not A298) );
 a75246a <=( (not A302)  and  (not A300) );
 a75247a <=( a75246a  and  a75243a );
 a75248a <=( a75247a  and  a75240a );
 a75252a <=( A199  and  (not A166) );
 a75253a <=( A167  and  a75252a );
 a75256a <=( (not A202)  and  (not A200) );
 a75259a <=( (not A265)  and  A203 );
 a75260a <=( a75259a  and  a75256a );
 a75261a <=( a75260a  and  a75253a );
 a75265a <=( A269  and  (not A268) );
 a75266a <=( A266  and  a75265a );
 a75269a <=( A299  and  A298 );
 a75272a <=( (not A301)  and  (not A300) );
 a75273a <=( a75272a  and  a75269a );
 a75274a <=( a75273a  and  a75266a );
 a75278a <=( A199  and  (not A166) );
 a75279a <=( A167  and  a75278a );
 a75282a <=( (not A202)  and  (not A200) );
 a75285a <=( (not A265)  and  A203 );
 a75286a <=( a75285a  and  a75282a );
 a75287a <=( a75286a  and  a75279a );
 a75291a <=( A269  and  (not A268) );
 a75292a <=( A266  and  a75291a );
 a75295a <=( A299  and  A298 );
 a75298a <=( A302  and  (not A300) );
 a75299a <=( a75298a  and  a75295a );
 a75300a <=( a75299a  and  a75292a );
 a75304a <=( A199  and  (not A166) );
 a75305a <=( A167  and  a75304a );
 a75308a <=( (not A202)  and  (not A200) );
 a75311a <=( (not A265)  and  A203 );
 a75312a <=( a75311a  and  a75308a );
 a75313a <=( a75312a  and  a75305a );
 a75317a <=( A269  and  (not A268) );
 a75318a <=( A266  and  a75317a );
 a75321a <=( (not A299)  and  A298 );
 a75324a <=( A301  and  (not A300) );
 a75325a <=( a75324a  and  a75321a );
 a75326a <=( a75325a  and  a75318a );
 a75330a <=( A199  and  (not A166) );
 a75331a <=( A167  and  a75330a );
 a75334a <=( (not A202)  and  (not A200) );
 a75337a <=( (not A265)  and  A203 );
 a75338a <=( a75337a  and  a75334a );
 a75339a <=( a75338a  and  a75331a );
 a75343a <=( A269  and  (not A268) );
 a75344a <=( A266  and  a75343a );
 a75347a <=( (not A299)  and  A298 );
 a75350a <=( (not A302)  and  (not A300) );
 a75351a <=( a75350a  and  a75347a );
 a75352a <=( a75351a  and  a75344a );
 a75356a <=( A199  and  (not A166) );
 a75357a <=( A167  and  a75356a );
 a75360a <=( (not A202)  and  (not A200) );
 a75363a <=( (not A265)  and  A203 );
 a75364a <=( a75363a  and  a75360a );
 a75365a <=( a75364a  and  a75357a );
 a75369a <=( A269  and  (not A268) );
 a75370a <=( A266  and  a75369a );
 a75373a <=( A299  and  (not A298) );
 a75376a <=( A301  and  (not A300) );
 a75377a <=( a75376a  and  a75373a );
 a75378a <=( a75377a  and  a75370a );
 a75382a <=( A199  and  (not A166) );
 a75383a <=( A167  and  a75382a );
 a75386a <=( (not A202)  and  (not A200) );
 a75389a <=( (not A265)  and  A203 );
 a75390a <=( a75389a  and  a75386a );
 a75391a <=( a75390a  and  a75383a );
 a75395a <=( A269  and  (not A268) );
 a75396a <=( A266  and  a75395a );
 a75399a <=( A299  and  (not A298) );
 a75402a <=( (not A302)  and  (not A300) );
 a75403a <=( a75402a  and  a75399a );
 a75404a <=( a75403a  and  a75396a );
 a75408a <=( A199  and  (not A166) );
 a75409a <=( A167  and  a75408a );
 a75412a <=( (not A202)  and  (not A200) );
 a75415a <=( A265  and  A203 );
 a75416a <=( a75415a  and  a75412a );
 a75417a <=( a75416a  and  a75409a );
 a75421a <=( A269  and  (not A268) );
 a75422a <=( (not A266)  and  a75421a );
 a75425a <=( A299  and  A298 );
 a75428a <=( (not A301)  and  (not A300) );
 a75429a <=( a75428a  and  a75425a );
 a75430a <=( a75429a  and  a75422a );
 a75434a <=( A199  and  (not A166) );
 a75435a <=( A167  and  a75434a );
 a75438a <=( (not A202)  and  (not A200) );
 a75441a <=( A265  and  A203 );
 a75442a <=( a75441a  and  a75438a );
 a75443a <=( a75442a  and  a75435a );
 a75447a <=( A269  and  (not A268) );
 a75448a <=( (not A266)  and  a75447a );
 a75451a <=( A299  and  A298 );
 a75454a <=( A302  and  (not A300) );
 a75455a <=( a75454a  and  a75451a );
 a75456a <=( a75455a  and  a75448a );
 a75460a <=( A199  and  (not A166) );
 a75461a <=( A167  and  a75460a );
 a75464a <=( (not A202)  and  (not A200) );
 a75467a <=( A265  and  A203 );
 a75468a <=( a75467a  and  a75464a );
 a75469a <=( a75468a  and  a75461a );
 a75473a <=( A269  and  (not A268) );
 a75474a <=( (not A266)  and  a75473a );
 a75477a <=( (not A299)  and  A298 );
 a75480a <=( A301  and  (not A300) );
 a75481a <=( a75480a  and  a75477a );
 a75482a <=( a75481a  and  a75474a );
 a75486a <=( A199  and  (not A166) );
 a75487a <=( A167  and  a75486a );
 a75490a <=( (not A202)  and  (not A200) );
 a75493a <=( A265  and  A203 );
 a75494a <=( a75493a  and  a75490a );
 a75495a <=( a75494a  and  a75487a );
 a75499a <=( A269  and  (not A268) );
 a75500a <=( (not A266)  and  a75499a );
 a75503a <=( (not A299)  and  A298 );
 a75506a <=( (not A302)  and  (not A300) );
 a75507a <=( a75506a  and  a75503a );
 a75508a <=( a75507a  and  a75500a );
 a75512a <=( A199  and  (not A166) );
 a75513a <=( A167  and  a75512a );
 a75516a <=( (not A202)  and  (not A200) );
 a75519a <=( A265  and  A203 );
 a75520a <=( a75519a  and  a75516a );
 a75521a <=( a75520a  and  a75513a );
 a75525a <=( A269  and  (not A268) );
 a75526a <=( (not A266)  and  a75525a );
 a75529a <=( A299  and  (not A298) );
 a75532a <=( A301  and  (not A300) );
 a75533a <=( a75532a  and  a75529a );
 a75534a <=( a75533a  and  a75526a );
 a75538a <=( A199  and  (not A166) );
 a75539a <=( A167  and  a75538a );
 a75542a <=( (not A202)  and  (not A200) );
 a75545a <=( A265  and  A203 );
 a75546a <=( a75545a  and  a75542a );
 a75547a <=( a75546a  and  a75539a );
 a75551a <=( A269  and  (not A268) );
 a75552a <=( (not A266)  and  a75551a );
 a75555a <=( A299  and  (not A298) );
 a75558a <=( (not A302)  and  (not A300) );
 a75559a <=( a75558a  and  a75555a );
 a75560a <=( a75559a  and  a75552a );
 a75564a <=( A199  and  (not A166) );
 a75565a <=( A167  and  a75564a );
 a75568a <=( (not A202)  and  (not A200) );
 a75571a <=( (not A265)  and  A203 );
 a75572a <=( a75571a  and  a75568a );
 a75573a <=( a75572a  and  a75565a );
 a75577a <=( (not A269)  and  A268 );
 a75578a <=( (not A266)  and  a75577a );
 a75581a <=( A299  and  A298 );
 a75584a <=( (not A301)  and  (not A300) );
 a75585a <=( a75584a  and  a75581a );
 a75586a <=( a75585a  and  a75578a );
 a75590a <=( A199  and  (not A166) );
 a75591a <=( A167  and  a75590a );
 a75594a <=( (not A202)  and  (not A200) );
 a75597a <=( (not A265)  and  A203 );
 a75598a <=( a75597a  and  a75594a );
 a75599a <=( a75598a  and  a75591a );
 a75603a <=( (not A269)  and  A268 );
 a75604a <=( (not A266)  and  a75603a );
 a75607a <=( A299  and  A298 );
 a75610a <=( A302  and  (not A300) );
 a75611a <=( a75610a  and  a75607a );
 a75612a <=( a75611a  and  a75604a );
 a75616a <=( A199  and  (not A166) );
 a75617a <=( A167  and  a75616a );
 a75620a <=( (not A202)  and  (not A200) );
 a75623a <=( (not A265)  and  A203 );
 a75624a <=( a75623a  and  a75620a );
 a75625a <=( a75624a  and  a75617a );
 a75629a <=( (not A269)  and  A268 );
 a75630a <=( (not A266)  and  a75629a );
 a75633a <=( (not A299)  and  A298 );
 a75636a <=( A301  and  (not A300) );
 a75637a <=( a75636a  and  a75633a );
 a75638a <=( a75637a  and  a75630a );
 a75642a <=( A199  and  (not A166) );
 a75643a <=( A167  and  a75642a );
 a75646a <=( (not A202)  and  (not A200) );
 a75649a <=( (not A265)  and  A203 );
 a75650a <=( a75649a  and  a75646a );
 a75651a <=( a75650a  and  a75643a );
 a75655a <=( (not A269)  and  A268 );
 a75656a <=( (not A266)  and  a75655a );
 a75659a <=( (not A299)  and  A298 );
 a75662a <=( (not A302)  and  (not A300) );
 a75663a <=( a75662a  and  a75659a );
 a75664a <=( a75663a  and  a75656a );
 a75668a <=( A199  and  (not A166) );
 a75669a <=( A167  and  a75668a );
 a75672a <=( (not A202)  and  (not A200) );
 a75675a <=( (not A265)  and  A203 );
 a75676a <=( a75675a  and  a75672a );
 a75677a <=( a75676a  and  a75669a );
 a75681a <=( (not A269)  and  A268 );
 a75682a <=( (not A266)  and  a75681a );
 a75685a <=( A299  and  (not A298) );
 a75688a <=( A301  and  (not A300) );
 a75689a <=( a75688a  and  a75685a );
 a75690a <=( a75689a  and  a75682a );
 a75694a <=( A199  and  (not A166) );
 a75695a <=( A167  and  a75694a );
 a75698a <=( (not A202)  and  (not A200) );
 a75701a <=( (not A265)  and  A203 );
 a75702a <=( a75701a  and  a75698a );
 a75703a <=( a75702a  and  a75695a );
 a75707a <=( (not A269)  and  A268 );
 a75708a <=( (not A266)  and  a75707a );
 a75711a <=( A299  and  (not A298) );
 a75714a <=( (not A302)  and  (not A300) );
 a75715a <=( a75714a  and  a75711a );
 a75716a <=( a75715a  and  a75708a );
 a75720a <=( A199  and  (not A166) );
 a75721a <=( A167  and  a75720a );
 a75724a <=( (not A201)  and  (not A200) );
 a75727a <=( A265  and  A202 );
 a75728a <=( a75727a  and  a75724a );
 a75729a <=( a75728a  and  a75721a );
 a75733a <=( (not A268)  and  (not A267) );
 a75734a <=( A266  and  a75733a );
 a75737a <=( A299  and  A298 );
 a75740a <=( (not A302)  and  A301 );
 a75741a <=( a75740a  and  a75737a );
 a75742a <=( a75741a  and  a75734a );
 a75746a <=( A199  and  (not A166) );
 a75747a <=( A167  and  a75746a );
 a75750a <=( (not A201)  and  (not A200) );
 a75753a <=( A265  and  A202 );
 a75754a <=( a75753a  and  a75750a );
 a75755a <=( a75754a  and  a75747a );
 a75759a <=( (not A268)  and  (not A267) );
 a75760a <=( A266  and  a75759a );
 a75763a <=( (not A299)  and  A298 );
 a75766a <=( A302  and  (not A301) );
 a75767a <=( a75766a  and  a75763a );
 a75768a <=( a75767a  and  a75760a );
 a75772a <=( A199  and  (not A166) );
 a75773a <=( A167  and  a75772a );
 a75776a <=( (not A201)  and  (not A200) );
 a75779a <=( A265  and  A202 );
 a75780a <=( a75779a  and  a75776a );
 a75781a <=( a75780a  and  a75773a );
 a75785a <=( (not A268)  and  (not A267) );
 a75786a <=( A266  and  a75785a );
 a75789a <=( A299  and  (not A298) );
 a75792a <=( A302  and  (not A301) );
 a75793a <=( a75792a  and  a75789a );
 a75794a <=( a75793a  and  a75786a );
 a75798a <=( A199  and  (not A166) );
 a75799a <=( A167  and  a75798a );
 a75802a <=( (not A201)  and  (not A200) );
 a75805a <=( A265  and  A202 );
 a75806a <=( a75805a  and  a75802a );
 a75807a <=( a75806a  and  a75799a );
 a75811a <=( (not A268)  and  (not A267) );
 a75812a <=( A266  and  a75811a );
 a75815a <=( (not A299)  and  (not A298) );
 a75818a <=( (not A302)  and  A301 );
 a75819a <=( a75818a  and  a75815a );
 a75820a <=( a75819a  and  a75812a );
 a75824a <=( A199  and  (not A166) );
 a75825a <=( A167  and  a75824a );
 a75828a <=( (not A201)  and  (not A200) );
 a75831a <=( A265  and  A202 );
 a75832a <=( a75831a  and  a75828a );
 a75833a <=( a75832a  and  a75825a );
 a75837a <=( A269  and  (not A267) );
 a75838a <=( A266  and  a75837a );
 a75841a <=( A299  and  A298 );
 a75844a <=( (not A302)  and  A301 );
 a75845a <=( a75844a  and  a75841a );
 a75846a <=( a75845a  and  a75838a );
 a75850a <=( A199  and  (not A166) );
 a75851a <=( A167  and  a75850a );
 a75854a <=( (not A201)  and  (not A200) );
 a75857a <=( A265  and  A202 );
 a75858a <=( a75857a  and  a75854a );
 a75859a <=( a75858a  and  a75851a );
 a75863a <=( A269  and  (not A267) );
 a75864a <=( A266  and  a75863a );
 a75867a <=( (not A299)  and  A298 );
 a75870a <=( A302  and  (not A301) );
 a75871a <=( a75870a  and  a75867a );
 a75872a <=( a75871a  and  a75864a );
 a75876a <=( A199  and  (not A166) );
 a75877a <=( A167  and  a75876a );
 a75880a <=( (not A201)  and  (not A200) );
 a75883a <=( A265  and  A202 );
 a75884a <=( a75883a  and  a75880a );
 a75885a <=( a75884a  and  a75877a );
 a75889a <=( A269  and  (not A267) );
 a75890a <=( A266  and  a75889a );
 a75893a <=( A299  and  (not A298) );
 a75896a <=( A302  and  (not A301) );
 a75897a <=( a75896a  and  a75893a );
 a75898a <=( a75897a  and  a75890a );
 a75902a <=( A199  and  (not A166) );
 a75903a <=( A167  and  a75902a );
 a75906a <=( (not A201)  and  (not A200) );
 a75909a <=( A265  and  A202 );
 a75910a <=( a75909a  and  a75906a );
 a75911a <=( a75910a  and  a75903a );
 a75915a <=( A269  and  (not A267) );
 a75916a <=( A266  and  a75915a );
 a75919a <=( (not A299)  and  (not A298) );
 a75922a <=( (not A302)  and  A301 );
 a75923a <=( a75922a  and  a75919a );
 a75924a <=( a75923a  and  a75916a );
 a75928a <=( A199  and  (not A166) );
 a75929a <=( A167  and  a75928a );
 a75932a <=( (not A201)  and  (not A200) );
 a75935a <=( (not A265)  and  A202 );
 a75936a <=( a75935a  and  a75932a );
 a75937a <=( a75936a  and  a75929a );
 a75941a <=( A268  and  (not A267) );
 a75942a <=( A266  and  a75941a );
 a75945a <=( A299  and  A298 );
 a75948a <=( (not A302)  and  A301 );
 a75949a <=( a75948a  and  a75945a );
 a75950a <=( a75949a  and  a75942a );
 a75954a <=( A199  and  (not A166) );
 a75955a <=( A167  and  a75954a );
 a75958a <=( (not A201)  and  (not A200) );
 a75961a <=( (not A265)  and  A202 );
 a75962a <=( a75961a  and  a75958a );
 a75963a <=( a75962a  and  a75955a );
 a75967a <=( A268  and  (not A267) );
 a75968a <=( A266  and  a75967a );
 a75971a <=( (not A299)  and  A298 );
 a75974a <=( A302  and  (not A301) );
 a75975a <=( a75974a  and  a75971a );
 a75976a <=( a75975a  and  a75968a );
 a75980a <=( A199  and  (not A166) );
 a75981a <=( A167  and  a75980a );
 a75984a <=( (not A201)  and  (not A200) );
 a75987a <=( (not A265)  and  A202 );
 a75988a <=( a75987a  and  a75984a );
 a75989a <=( a75988a  and  a75981a );
 a75993a <=( A268  and  (not A267) );
 a75994a <=( A266  and  a75993a );
 a75997a <=( A299  and  (not A298) );
 a76000a <=( A302  and  (not A301) );
 a76001a <=( a76000a  and  a75997a );
 a76002a <=( a76001a  and  a75994a );
 a76006a <=( A199  and  (not A166) );
 a76007a <=( A167  and  a76006a );
 a76010a <=( (not A201)  and  (not A200) );
 a76013a <=( (not A265)  and  A202 );
 a76014a <=( a76013a  and  a76010a );
 a76015a <=( a76014a  and  a76007a );
 a76019a <=( A268  and  (not A267) );
 a76020a <=( A266  and  a76019a );
 a76023a <=( (not A299)  and  (not A298) );
 a76026a <=( (not A302)  and  A301 );
 a76027a <=( a76026a  and  a76023a );
 a76028a <=( a76027a  and  a76020a );
 a76032a <=( A199  and  (not A166) );
 a76033a <=( A167  and  a76032a );
 a76036a <=( (not A201)  and  (not A200) );
 a76039a <=( (not A265)  and  A202 );
 a76040a <=( a76039a  and  a76036a );
 a76041a <=( a76040a  and  a76033a );
 a76045a <=( (not A269)  and  (not A267) );
 a76046a <=( A266  and  a76045a );
 a76049a <=( A299  and  A298 );
 a76052a <=( (not A302)  and  A301 );
 a76053a <=( a76052a  and  a76049a );
 a76054a <=( a76053a  and  a76046a );
 a76058a <=( A199  and  (not A166) );
 a76059a <=( A167  and  a76058a );
 a76062a <=( (not A201)  and  (not A200) );
 a76065a <=( (not A265)  and  A202 );
 a76066a <=( a76065a  and  a76062a );
 a76067a <=( a76066a  and  a76059a );
 a76071a <=( (not A269)  and  (not A267) );
 a76072a <=( A266  and  a76071a );
 a76075a <=( (not A299)  and  A298 );
 a76078a <=( A302  and  (not A301) );
 a76079a <=( a76078a  and  a76075a );
 a76080a <=( a76079a  and  a76072a );
 a76084a <=( A199  and  (not A166) );
 a76085a <=( A167  and  a76084a );
 a76088a <=( (not A201)  and  (not A200) );
 a76091a <=( (not A265)  and  A202 );
 a76092a <=( a76091a  and  a76088a );
 a76093a <=( a76092a  and  a76085a );
 a76097a <=( (not A269)  and  (not A267) );
 a76098a <=( A266  and  a76097a );
 a76101a <=( A299  and  (not A298) );
 a76104a <=( A302  and  (not A301) );
 a76105a <=( a76104a  and  a76101a );
 a76106a <=( a76105a  and  a76098a );
 a76110a <=( A199  and  (not A166) );
 a76111a <=( A167  and  a76110a );
 a76114a <=( (not A201)  and  (not A200) );
 a76117a <=( (not A265)  and  A202 );
 a76118a <=( a76117a  and  a76114a );
 a76119a <=( a76118a  and  a76111a );
 a76123a <=( (not A269)  and  (not A267) );
 a76124a <=( A266  and  a76123a );
 a76127a <=( (not A299)  and  (not A298) );
 a76130a <=( (not A302)  and  A301 );
 a76131a <=( a76130a  and  a76127a );
 a76132a <=( a76131a  and  a76124a );
 a76136a <=( A199  and  (not A166) );
 a76137a <=( A167  and  a76136a );
 a76140a <=( (not A201)  and  (not A200) );
 a76143a <=( A265  and  A202 );
 a76144a <=( a76143a  and  a76140a );
 a76145a <=( a76144a  and  a76137a );
 a76149a <=( A268  and  (not A267) );
 a76150a <=( (not A266)  and  a76149a );
 a76153a <=( A299  and  A298 );
 a76156a <=( (not A302)  and  A301 );
 a76157a <=( a76156a  and  a76153a );
 a76158a <=( a76157a  and  a76150a );
 a76162a <=( A199  and  (not A166) );
 a76163a <=( A167  and  a76162a );
 a76166a <=( (not A201)  and  (not A200) );
 a76169a <=( A265  and  A202 );
 a76170a <=( a76169a  and  a76166a );
 a76171a <=( a76170a  and  a76163a );
 a76175a <=( A268  and  (not A267) );
 a76176a <=( (not A266)  and  a76175a );
 a76179a <=( (not A299)  and  A298 );
 a76182a <=( A302  and  (not A301) );
 a76183a <=( a76182a  and  a76179a );
 a76184a <=( a76183a  and  a76176a );
 a76188a <=( A199  and  (not A166) );
 a76189a <=( A167  and  a76188a );
 a76192a <=( (not A201)  and  (not A200) );
 a76195a <=( A265  and  A202 );
 a76196a <=( a76195a  and  a76192a );
 a76197a <=( a76196a  and  a76189a );
 a76201a <=( A268  and  (not A267) );
 a76202a <=( (not A266)  and  a76201a );
 a76205a <=( A299  and  (not A298) );
 a76208a <=( A302  and  (not A301) );
 a76209a <=( a76208a  and  a76205a );
 a76210a <=( a76209a  and  a76202a );
 a76214a <=( A199  and  (not A166) );
 a76215a <=( A167  and  a76214a );
 a76218a <=( (not A201)  and  (not A200) );
 a76221a <=( A265  and  A202 );
 a76222a <=( a76221a  and  a76218a );
 a76223a <=( a76222a  and  a76215a );
 a76227a <=( A268  and  (not A267) );
 a76228a <=( (not A266)  and  a76227a );
 a76231a <=( (not A299)  and  (not A298) );
 a76234a <=( (not A302)  and  A301 );
 a76235a <=( a76234a  and  a76231a );
 a76236a <=( a76235a  and  a76228a );
 a76240a <=( A199  and  (not A166) );
 a76241a <=( A167  and  a76240a );
 a76244a <=( (not A201)  and  (not A200) );
 a76247a <=( A265  and  A202 );
 a76248a <=( a76247a  and  a76244a );
 a76249a <=( a76248a  and  a76241a );
 a76253a <=( (not A269)  and  (not A267) );
 a76254a <=( (not A266)  and  a76253a );
 a76257a <=( A299  and  A298 );
 a76260a <=( (not A302)  and  A301 );
 a76261a <=( a76260a  and  a76257a );
 a76262a <=( a76261a  and  a76254a );
 a76266a <=( A199  and  (not A166) );
 a76267a <=( A167  and  a76266a );
 a76270a <=( (not A201)  and  (not A200) );
 a76273a <=( A265  and  A202 );
 a76274a <=( a76273a  and  a76270a );
 a76275a <=( a76274a  and  a76267a );
 a76279a <=( (not A269)  and  (not A267) );
 a76280a <=( (not A266)  and  a76279a );
 a76283a <=( (not A299)  and  A298 );
 a76286a <=( A302  and  (not A301) );
 a76287a <=( a76286a  and  a76283a );
 a76288a <=( a76287a  and  a76280a );
 a76292a <=( A199  and  (not A166) );
 a76293a <=( A167  and  a76292a );
 a76296a <=( (not A201)  and  (not A200) );
 a76299a <=( A265  and  A202 );
 a76300a <=( a76299a  and  a76296a );
 a76301a <=( a76300a  and  a76293a );
 a76305a <=( (not A269)  and  (not A267) );
 a76306a <=( (not A266)  and  a76305a );
 a76309a <=( A299  and  (not A298) );
 a76312a <=( A302  and  (not A301) );
 a76313a <=( a76312a  and  a76309a );
 a76314a <=( a76313a  and  a76306a );
 a76318a <=( A199  and  (not A166) );
 a76319a <=( A167  and  a76318a );
 a76322a <=( (not A201)  and  (not A200) );
 a76325a <=( A265  and  A202 );
 a76326a <=( a76325a  and  a76322a );
 a76327a <=( a76326a  and  a76319a );
 a76331a <=( (not A269)  and  (not A267) );
 a76332a <=( (not A266)  and  a76331a );
 a76335a <=( (not A299)  and  (not A298) );
 a76338a <=( (not A302)  and  A301 );
 a76339a <=( a76338a  and  a76335a );
 a76340a <=( a76339a  and  a76332a );
 a76344a <=( A199  and  (not A166) );
 a76345a <=( A167  and  a76344a );
 a76348a <=( (not A201)  and  (not A200) );
 a76351a <=( A265  and  (not A203) );
 a76352a <=( a76351a  and  a76348a );
 a76353a <=( a76352a  and  a76345a );
 a76357a <=( (not A268)  and  (not A267) );
 a76358a <=( A266  and  a76357a );
 a76361a <=( A299  and  A298 );
 a76364a <=( (not A302)  and  A301 );
 a76365a <=( a76364a  and  a76361a );
 a76366a <=( a76365a  and  a76358a );
 a76370a <=( A199  and  (not A166) );
 a76371a <=( A167  and  a76370a );
 a76374a <=( (not A201)  and  (not A200) );
 a76377a <=( A265  and  (not A203) );
 a76378a <=( a76377a  and  a76374a );
 a76379a <=( a76378a  and  a76371a );
 a76383a <=( (not A268)  and  (not A267) );
 a76384a <=( A266  and  a76383a );
 a76387a <=( (not A299)  and  A298 );
 a76390a <=( A302  and  (not A301) );
 a76391a <=( a76390a  and  a76387a );
 a76392a <=( a76391a  and  a76384a );
 a76396a <=( A199  and  (not A166) );
 a76397a <=( A167  and  a76396a );
 a76400a <=( (not A201)  and  (not A200) );
 a76403a <=( A265  and  (not A203) );
 a76404a <=( a76403a  and  a76400a );
 a76405a <=( a76404a  and  a76397a );
 a76409a <=( (not A268)  and  (not A267) );
 a76410a <=( A266  and  a76409a );
 a76413a <=( A299  and  (not A298) );
 a76416a <=( A302  and  (not A301) );
 a76417a <=( a76416a  and  a76413a );
 a76418a <=( a76417a  and  a76410a );
 a76422a <=( A199  and  (not A166) );
 a76423a <=( A167  and  a76422a );
 a76426a <=( (not A201)  and  (not A200) );
 a76429a <=( A265  and  (not A203) );
 a76430a <=( a76429a  and  a76426a );
 a76431a <=( a76430a  and  a76423a );
 a76435a <=( (not A268)  and  (not A267) );
 a76436a <=( A266  and  a76435a );
 a76439a <=( (not A299)  and  (not A298) );
 a76442a <=( (not A302)  and  A301 );
 a76443a <=( a76442a  and  a76439a );
 a76444a <=( a76443a  and  a76436a );
 a76448a <=( A199  and  (not A166) );
 a76449a <=( A167  and  a76448a );
 a76452a <=( (not A201)  and  (not A200) );
 a76455a <=( A265  and  (not A203) );
 a76456a <=( a76455a  and  a76452a );
 a76457a <=( a76456a  and  a76449a );
 a76461a <=( A269  and  (not A267) );
 a76462a <=( A266  and  a76461a );
 a76465a <=( A299  and  A298 );
 a76468a <=( (not A302)  and  A301 );
 a76469a <=( a76468a  and  a76465a );
 a76470a <=( a76469a  and  a76462a );
 a76474a <=( A199  and  (not A166) );
 a76475a <=( A167  and  a76474a );
 a76478a <=( (not A201)  and  (not A200) );
 a76481a <=( A265  and  (not A203) );
 a76482a <=( a76481a  and  a76478a );
 a76483a <=( a76482a  and  a76475a );
 a76487a <=( A269  and  (not A267) );
 a76488a <=( A266  and  a76487a );
 a76491a <=( (not A299)  and  A298 );
 a76494a <=( A302  and  (not A301) );
 a76495a <=( a76494a  and  a76491a );
 a76496a <=( a76495a  and  a76488a );
 a76500a <=( A199  and  (not A166) );
 a76501a <=( A167  and  a76500a );
 a76504a <=( (not A201)  and  (not A200) );
 a76507a <=( A265  and  (not A203) );
 a76508a <=( a76507a  and  a76504a );
 a76509a <=( a76508a  and  a76501a );
 a76513a <=( A269  and  (not A267) );
 a76514a <=( A266  and  a76513a );
 a76517a <=( A299  and  (not A298) );
 a76520a <=( A302  and  (not A301) );
 a76521a <=( a76520a  and  a76517a );
 a76522a <=( a76521a  and  a76514a );
 a76526a <=( A199  and  (not A166) );
 a76527a <=( A167  and  a76526a );
 a76530a <=( (not A201)  and  (not A200) );
 a76533a <=( A265  and  (not A203) );
 a76534a <=( a76533a  and  a76530a );
 a76535a <=( a76534a  and  a76527a );
 a76539a <=( A269  and  (not A267) );
 a76540a <=( A266  and  a76539a );
 a76543a <=( (not A299)  and  (not A298) );
 a76546a <=( (not A302)  and  A301 );
 a76547a <=( a76546a  and  a76543a );
 a76548a <=( a76547a  and  a76540a );
 a76552a <=( A199  and  (not A166) );
 a76553a <=( A167  and  a76552a );
 a76556a <=( (not A201)  and  (not A200) );
 a76559a <=( (not A265)  and  (not A203) );
 a76560a <=( a76559a  and  a76556a );
 a76561a <=( a76560a  and  a76553a );
 a76565a <=( A268  and  (not A267) );
 a76566a <=( A266  and  a76565a );
 a76569a <=( A299  and  A298 );
 a76572a <=( (not A302)  and  A301 );
 a76573a <=( a76572a  and  a76569a );
 a76574a <=( a76573a  and  a76566a );
 a76578a <=( A199  and  (not A166) );
 a76579a <=( A167  and  a76578a );
 a76582a <=( (not A201)  and  (not A200) );
 a76585a <=( (not A265)  and  (not A203) );
 a76586a <=( a76585a  and  a76582a );
 a76587a <=( a76586a  and  a76579a );
 a76591a <=( A268  and  (not A267) );
 a76592a <=( A266  and  a76591a );
 a76595a <=( (not A299)  and  A298 );
 a76598a <=( A302  and  (not A301) );
 a76599a <=( a76598a  and  a76595a );
 a76600a <=( a76599a  and  a76592a );
 a76604a <=( A199  and  (not A166) );
 a76605a <=( A167  and  a76604a );
 a76608a <=( (not A201)  and  (not A200) );
 a76611a <=( (not A265)  and  (not A203) );
 a76612a <=( a76611a  and  a76608a );
 a76613a <=( a76612a  and  a76605a );
 a76617a <=( A268  and  (not A267) );
 a76618a <=( A266  and  a76617a );
 a76621a <=( A299  and  (not A298) );
 a76624a <=( A302  and  (not A301) );
 a76625a <=( a76624a  and  a76621a );
 a76626a <=( a76625a  and  a76618a );
 a76630a <=( A199  and  (not A166) );
 a76631a <=( A167  and  a76630a );
 a76634a <=( (not A201)  and  (not A200) );
 a76637a <=( (not A265)  and  (not A203) );
 a76638a <=( a76637a  and  a76634a );
 a76639a <=( a76638a  and  a76631a );
 a76643a <=( A268  and  (not A267) );
 a76644a <=( A266  and  a76643a );
 a76647a <=( (not A299)  and  (not A298) );
 a76650a <=( (not A302)  and  A301 );
 a76651a <=( a76650a  and  a76647a );
 a76652a <=( a76651a  and  a76644a );
 a76656a <=( A199  and  (not A166) );
 a76657a <=( A167  and  a76656a );
 a76660a <=( (not A201)  and  (not A200) );
 a76663a <=( (not A265)  and  (not A203) );
 a76664a <=( a76663a  and  a76660a );
 a76665a <=( a76664a  and  a76657a );
 a76669a <=( (not A269)  and  (not A267) );
 a76670a <=( A266  and  a76669a );
 a76673a <=( A299  and  A298 );
 a76676a <=( (not A302)  and  A301 );
 a76677a <=( a76676a  and  a76673a );
 a76678a <=( a76677a  and  a76670a );
 a76682a <=( A199  and  (not A166) );
 a76683a <=( A167  and  a76682a );
 a76686a <=( (not A201)  and  (not A200) );
 a76689a <=( (not A265)  and  (not A203) );
 a76690a <=( a76689a  and  a76686a );
 a76691a <=( a76690a  and  a76683a );
 a76695a <=( (not A269)  and  (not A267) );
 a76696a <=( A266  and  a76695a );
 a76699a <=( (not A299)  and  A298 );
 a76702a <=( A302  and  (not A301) );
 a76703a <=( a76702a  and  a76699a );
 a76704a <=( a76703a  and  a76696a );
 a76708a <=( A199  and  (not A166) );
 a76709a <=( A167  and  a76708a );
 a76712a <=( (not A201)  and  (not A200) );
 a76715a <=( (not A265)  and  (not A203) );
 a76716a <=( a76715a  and  a76712a );
 a76717a <=( a76716a  and  a76709a );
 a76721a <=( (not A269)  and  (not A267) );
 a76722a <=( A266  and  a76721a );
 a76725a <=( A299  and  (not A298) );
 a76728a <=( A302  and  (not A301) );
 a76729a <=( a76728a  and  a76725a );
 a76730a <=( a76729a  and  a76722a );
 a76734a <=( A199  and  (not A166) );
 a76735a <=( A167  and  a76734a );
 a76738a <=( (not A201)  and  (not A200) );
 a76741a <=( (not A265)  and  (not A203) );
 a76742a <=( a76741a  and  a76738a );
 a76743a <=( a76742a  and  a76735a );
 a76747a <=( (not A269)  and  (not A267) );
 a76748a <=( A266  and  a76747a );
 a76751a <=( (not A299)  and  (not A298) );
 a76754a <=( (not A302)  and  A301 );
 a76755a <=( a76754a  and  a76751a );
 a76756a <=( a76755a  and  a76748a );
 a76760a <=( A199  and  (not A166) );
 a76761a <=( A167  and  a76760a );
 a76764a <=( (not A201)  and  (not A200) );
 a76767a <=( A265  and  (not A203) );
 a76768a <=( a76767a  and  a76764a );
 a76769a <=( a76768a  and  a76761a );
 a76773a <=( A268  and  (not A267) );
 a76774a <=( (not A266)  and  a76773a );
 a76777a <=( A299  and  A298 );
 a76780a <=( (not A302)  and  A301 );
 a76781a <=( a76780a  and  a76777a );
 a76782a <=( a76781a  and  a76774a );
 a76786a <=( A199  and  (not A166) );
 a76787a <=( A167  and  a76786a );
 a76790a <=( (not A201)  and  (not A200) );
 a76793a <=( A265  and  (not A203) );
 a76794a <=( a76793a  and  a76790a );
 a76795a <=( a76794a  and  a76787a );
 a76799a <=( A268  and  (not A267) );
 a76800a <=( (not A266)  and  a76799a );
 a76803a <=( (not A299)  and  A298 );
 a76806a <=( A302  and  (not A301) );
 a76807a <=( a76806a  and  a76803a );
 a76808a <=( a76807a  and  a76800a );
 a76812a <=( A199  and  (not A166) );
 a76813a <=( A167  and  a76812a );
 a76816a <=( (not A201)  and  (not A200) );
 a76819a <=( A265  and  (not A203) );
 a76820a <=( a76819a  and  a76816a );
 a76821a <=( a76820a  and  a76813a );
 a76825a <=( A268  and  (not A267) );
 a76826a <=( (not A266)  and  a76825a );
 a76829a <=( A299  and  (not A298) );
 a76832a <=( A302  and  (not A301) );
 a76833a <=( a76832a  and  a76829a );
 a76834a <=( a76833a  and  a76826a );
 a76838a <=( A199  and  (not A166) );
 a76839a <=( A167  and  a76838a );
 a76842a <=( (not A201)  and  (not A200) );
 a76845a <=( A265  and  (not A203) );
 a76846a <=( a76845a  and  a76842a );
 a76847a <=( a76846a  and  a76839a );
 a76851a <=( A268  and  (not A267) );
 a76852a <=( (not A266)  and  a76851a );
 a76855a <=( (not A299)  and  (not A298) );
 a76858a <=( (not A302)  and  A301 );
 a76859a <=( a76858a  and  a76855a );
 a76860a <=( a76859a  and  a76852a );
 a76864a <=( A199  and  (not A166) );
 a76865a <=( A167  and  a76864a );
 a76868a <=( (not A201)  and  (not A200) );
 a76871a <=( A265  and  (not A203) );
 a76872a <=( a76871a  and  a76868a );
 a76873a <=( a76872a  and  a76865a );
 a76877a <=( (not A269)  and  (not A267) );
 a76878a <=( (not A266)  and  a76877a );
 a76881a <=( A299  and  A298 );
 a76884a <=( (not A302)  and  A301 );
 a76885a <=( a76884a  and  a76881a );
 a76886a <=( a76885a  and  a76878a );
 a76890a <=( A199  and  (not A166) );
 a76891a <=( A167  and  a76890a );
 a76894a <=( (not A201)  and  (not A200) );
 a76897a <=( A265  and  (not A203) );
 a76898a <=( a76897a  and  a76894a );
 a76899a <=( a76898a  and  a76891a );
 a76903a <=( (not A269)  and  (not A267) );
 a76904a <=( (not A266)  and  a76903a );
 a76907a <=( (not A299)  and  A298 );
 a76910a <=( A302  and  (not A301) );
 a76911a <=( a76910a  and  a76907a );
 a76912a <=( a76911a  and  a76904a );
 a76916a <=( A199  and  (not A166) );
 a76917a <=( A167  and  a76916a );
 a76920a <=( (not A201)  and  (not A200) );
 a76923a <=( A265  and  (not A203) );
 a76924a <=( a76923a  and  a76920a );
 a76925a <=( a76924a  and  a76917a );
 a76929a <=( (not A269)  and  (not A267) );
 a76930a <=( (not A266)  and  a76929a );
 a76933a <=( A299  and  (not A298) );
 a76936a <=( A302  and  (not A301) );
 a76937a <=( a76936a  and  a76933a );
 a76938a <=( a76937a  and  a76930a );
 a76942a <=( A199  and  (not A166) );
 a76943a <=( A167  and  a76942a );
 a76946a <=( (not A201)  and  (not A200) );
 a76949a <=( A265  and  (not A203) );
 a76950a <=( a76949a  and  a76946a );
 a76951a <=( a76950a  and  a76943a );
 a76955a <=( (not A269)  and  (not A267) );
 a76956a <=( (not A266)  and  a76955a );
 a76959a <=( (not A299)  and  (not A298) );
 a76962a <=( (not A302)  and  A301 );
 a76963a <=( a76962a  and  a76959a );
 a76964a <=( a76963a  and  a76956a );
 a76968a <=( (not A199)  and  (not A166) );
 a76969a <=( A167  and  a76968a );
 a76972a <=( A202  and  (not A200) );
 a76975a <=( A265  and  (not A203) );
 a76976a <=( a76975a  and  a76972a );
 a76977a <=( a76976a  and  a76969a );
 a76981a <=( (not A269)  and  A268 );
 a76982a <=( A266  and  a76981a );
 a76985a <=( A299  and  A298 );
 a76988a <=( (not A301)  and  (not A300) );
 a76989a <=( a76988a  and  a76985a );
 a76990a <=( a76989a  and  a76982a );
 a76994a <=( (not A199)  and  (not A166) );
 a76995a <=( A167  and  a76994a );
 a76998a <=( A202  and  (not A200) );
 a77001a <=( A265  and  (not A203) );
 a77002a <=( a77001a  and  a76998a );
 a77003a <=( a77002a  and  a76995a );
 a77007a <=( (not A269)  and  A268 );
 a77008a <=( A266  and  a77007a );
 a77011a <=( A299  and  A298 );
 a77014a <=( A302  and  (not A300) );
 a77015a <=( a77014a  and  a77011a );
 a77016a <=( a77015a  and  a77008a );
 a77020a <=( (not A199)  and  (not A166) );
 a77021a <=( A167  and  a77020a );
 a77024a <=( A202  and  (not A200) );
 a77027a <=( A265  and  (not A203) );
 a77028a <=( a77027a  and  a77024a );
 a77029a <=( a77028a  and  a77021a );
 a77033a <=( (not A269)  and  A268 );
 a77034a <=( A266  and  a77033a );
 a77037a <=( (not A299)  and  A298 );
 a77040a <=( A301  and  (not A300) );
 a77041a <=( a77040a  and  a77037a );
 a77042a <=( a77041a  and  a77034a );
 a77046a <=( (not A199)  and  (not A166) );
 a77047a <=( A167  and  a77046a );
 a77050a <=( A202  and  (not A200) );
 a77053a <=( A265  and  (not A203) );
 a77054a <=( a77053a  and  a77050a );
 a77055a <=( a77054a  and  a77047a );
 a77059a <=( (not A269)  and  A268 );
 a77060a <=( A266  and  a77059a );
 a77063a <=( (not A299)  and  A298 );
 a77066a <=( (not A302)  and  (not A300) );
 a77067a <=( a77066a  and  a77063a );
 a77068a <=( a77067a  and  a77060a );
 a77072a <=( (not A199)  and  (not A166) );
 a77073a <=( A167  and  a77072a );
 a77076a <=( A202  and  (not A200) );
 a77079a <=( A265  and  (not A203) );
 a77080a <=( a77079a  and  a77076a );
 a77081a <=( a77080a  and  a77073a );
 a77085a <=( (not A269)  and  A268 );
 a77086a <=( A266  and  a77085a );
 a77089a <=( A299  and  (not A298) );
 a77092a <=( A301  and  (not A300) );
 a77093a <=( a77092a  and  a77089a );
 a77094a <=( a77093a  and  a77086a );
 a77098a <=( (not A199)  and  (not A166) );
 a77099a <=( A167  and  a77098a );
 a77102a <=( A202  and  (not A200) );
 a77105a <=( A265  and  (not A203) );
 a77106a <=( a77105a  and  a77102a );
 a77107a <=( a77106a  and  a77099a );
 a77111a <=( (not A269)  and  A268 );
 a77112a <=( A266  and  a77111a );
 a77115a <=( A299  and  (not A298) );
 a77118a <=( (not A302)  and  (not A300) );
 a77119a <=( a77118a  and  a77115a );
 a77120a <=( a77119a  and  a77112a );
 a77124a <=( (not A199)  and  (not A166) );
 a77125a <=( A167  and  a77124a );
 a77128a <=( A202  and  (not A200) );
 a77131a <=( (not A265)  and  (not A203) );
 a77132a <=( a77131a  and  a77128a );
 a77133a <=( a77132a  and  a77125a );
 a77137a <=( A269  and  (not A268) );
 a77138a <=( A266  and  a77137a );
 a77141a <=( A299  and  A298 );
 a77144a <=( (not A301)  and  (not A300) );
 a77145a <=( a77144a  and  a77141a );
 a77146a <=( a77145a  and  a77138a );
 a77150a <=( (not A199)  and  (not A166) );
 a77151a <=( A167  and  a77150a );
 a77154a <=( A202  and  (not A200) );
 a77157a <=( (not A265)  and  (not A203) );
 a77158a <=( a77157a  and  a77154a );
 a77159a <=( a77158a  and  a77151a );
 a77163a <=( A269  and  (not A268) );
 a77164a <=( A266  and  a77163a );
 a77167a <=( A299  and  A298 );
 a77170a <=( A302  and  (not A300) );
 a77171a <=( a77170a  and  a77167a );
 a77172a <=( a77171a  and  a77164a );
 a77176a <=( (not A199)  and  (not A166) );
 a77177a <=( A167  and  a77176a );
 a77180a <=( A202  and  (not A200) );
 a77183a <=( (not A265)  and  (not A203) );
 a77184a <=( a77183a  and  a77180a );
 a77185a <=( a77184a  and  a77177a );
 a77189a <=( A269  and  (not A268) );
 a77190a <=( A266  and  a77189a );
 a77193a <=( (not A299)  and  A298 );
 a77196a <=( A301  and  (not A300) );
 a77197a <=( a77196a  and  a77193a );
 a77198a <=( a77197a  and  a77190a );
 a77202a <=( (not A199)  and  (not A166) );
 a77203a <=( A167  and  a77202a );
 a77206a <=( A202  and  (not A200) );
 a77209a <=( (not A265)  and  (not A203) );
 a77210a <=( a77209a  and  a77206a );
 a77211a <=( a77210a  and  a77203a );
 a77215a <=( A269  and  (not A268) );
 a77216a <=( A266  and  a77215a );
 a77219a <=( (not A299)  and  A298 );
 a77222a <=( (not A302)  and  (not A300) );
 a77223a <=( a77222a  and  a77219a );
 a77224a <=( a77223a  and  a77216a );
 a77228a <=( (not A199)  and  (not A166) );
 a77229a <=( A167  and  a77228a );
 a77232a <=( A202  and  (not A200) );
 a77235a <=( (not A265)  and  (not A203) );
 a77236a <=( a77235a  and  a77232a );
 a77237a <=( a77236a  and  a77229a );
 a77241a <=( A269  and  (not A268) );
 a77242a <=( A266  and  a77241a );
 a77245a <=( A299  and  (not A298) );
 a77248a <=( A301  and  (not A300) );
 a77249a <=( a77248a  and  a77245a );
 a77250a <=( a77249a  and  a77242a );
 a77254a <=( (not A199)  and  (not A166) );
 a77255a <=( A167  and  a77254a );
 a77258a <=( A202  and  (not A200) );
 a77261a <=( (not A265)  and  (not A203) );
 a77262a <=( a77261a  and  a77258a );
 a77263a <=( a77262a  and  a77255a );
 a77267a <=( A269  and  (not A268) );
 a77268a <=( A266  and  a77267a );
 a77271a <=( A299  and  (not A298) );
 a77274a <=( (not A302)  and  (not A300) );
 a77275a <=( a77274a  and  a77271a );
 a77276a <=( a77275a  and  a77268a );
 a77280a <=( (not A199)  and  (not A166) );
 a77281a <=( A167  and  a77280a );
 a77284a <=( A202  and  (not A200) );
 a77287a <=( A265  and  (not A203) );
 a77288a <=( a77287a  and  a77284a );
 a77289a <=( a77288a  and  a77281a );
 a77293a <=( A269  and  (not A268) );
 a77294a <=( (not A266)  and  a77293a );
 a77297a <=( A299  and  A298 );
 a77300a <=( (not A301)  and  (not A300) );
 a77301a <=( a77300a  and  a77297a );
 a77302a <=( a77301a  and  a77294a );
 a77306a <=( (not A199)  and  (not A166) );
 a77307a <=( A167  and  a77306a );
 a77310a <=( A202  and  (not A200) );
 a77313a <=( A265  and  (not A203) );
 a77314a <=( a77313a  and  a77310a );
 a77315a <=( a77314a  and  a77307a );
 a77319a <=( A269  and  (not A268) );
 a77320a <=( (not A266)  and  a77319a );
 a77323a <=( A299  and  A298 );
 a77326a <=( A302  and  (not A300) );
 a77327a <=( a77326a  and  a77323a );
 a77328a <=( a77327a  and  a77320a );
 a77332a <=( (not A199)  and  (not A166) );
 a77333a <=( A167  and  a77332a );
 a77336a <=( A202  and  (not A200) );
 a77339a <=( A265  and  (not A203) );
 a77340a <=( a77339a  and  a77336a );
 a77341a <=( a77340a  and  a77333a );
 a77345a <=( A269  and  (not A268) );
 a77346a <=( (not A266)  and  a77345a );
 a77349a <=( (not A299)  and  A298 );
 a77352a <=( A301  and  (not A300) );
 a77353a <=( a77352a  and  a77349a );
 a77354a <=( a77353a  and  a77346a );
 a77358a <=( (not A199)  and  (not A166) );
 a77359a <=( A167  and  a77358a );
 a77362a <=( A202  and  (not A200) );
 a77365a <=( A265  and  (not A203) );
 a77366a <=( a77365a  and  a77362a );
 a77367a <=( a77366a  and  a77359a );
 a77371a <=( A269  and  (not A268) );
 a77372a <=( (not A266)  and  a77371a );
 a77375a <=( (not A299)  and  A298 );
 a77378a <=( (not A302)  and  (not A300) );
 a77379a <=( a77378a  and  a77375a );
 a77380a <=( a77379a  and  a77372a );
 a77384a <=( (not A199)  and  (not A166) );
 a77385a <=( A167  and  a77384a );
 a77388a <=( A202  and  (not A200) );
 a77391a <=( A265  and  (not A203) );
 a77392a <=( a77391a  and  a77388a );
 a77393a <=( a77392a  and  a77385a );
 a77397a <=( A269  and  (not A268) );
 a77398a <=( (not A266)  and  a77397a );
 a77401a <=( A299  and  (not A298) );
 a77404a <=( A301  and  (not A300) );
 a77405a <=( a77404a  and  a77401a );
 a77406a <=( a77405a  and  a77398a );
 a77410a <=( (not A199)  and  (not A166) );
 a77411a <=( A167  and  a77410a );
 a77414a <=( A202  and  (not A200) );
 a77417a <=( A265  and  (not A203) );
 a77418a <=( a77417a  and  a77414a );
 a77419a <=( a77418a  and  a77411a );
 a77423a <=( A269  and  (not A268) );
 a77424a <=( (not A266)  and  a77423a );
 a77427a <=( A299  and  (not A298) );
 a77430a <=( (not A302)  and  (not A300) );
 a77431a <=( a77430a  and  a77427a );
 a77432a <=( a77431a  and  a77424a );
 a77436a <=( (not A199)  and  (not A166) );
 a77437a <=( A167  and  a77436a );
 a77440a <=( A202  and  (not A200) );
 a77443a <=( (not A265)  and  (not A203) );
 a77444a <=( a77443a  and  a77440a );
 a77445a <=( a77444a  and  a77437a );
 a77449a <=( (not A269)  and  A268 );
 a77450a <=( (not A266)  and  a77449a );
 a77453a <=( A299  and  A298 );
 a77456a <=( (not A301)  and  (not A300) );
 a77457a <=( a77456a  and  a77453a );
 a77458a <=( a77457a  and  a77450a );
 a77462a <=( (not A199)  and  (not A166) );
 a77463a <=( A167  and  a77462a );
 a77466a <=( A202  and  (not A200) );
 a77469a <=( (not A265)  and  (not A203) );
 a77470a <=( a77469a  and  a77466a );
 a77471a <=( a77470a  and  a77463a );
 a77475a <=( (not A269)  and  A268 );
 a77476a <=( (not A266)  and  a77475a );
 a77479a <=( A299  and  A298 );
 a77482a <=( A302  and  (not A300) );
 a77483a <=( a77482a  and  a77479a );
 a77484a <=( a77483a  and  a77476a );
 a77488a <=( (not A199)  and  (not A166) );
 a77489a <=( A167  and  a77488a );
 a77492a <=( A202  and  (not A200) );
 a77495a <=( (not A265)  and  (not A203) );
 a77496a <=( a77495a  and  a77492a );
 a77497a <=( a77496a  and  a77489a );
 a77501a <=( (not A269)  and  A268 );
 a77502a <=( (not A266)  and  a77501a );
 a77505a <=( (not A299)  and  A298 );
 a77508a <=( A301  and  (not A300) );
 a77509a <=( a77508a  and  a77505a );
 a77510a <=( a77509a  and  a77502a );
 a77514a <=( (not A199)  and  (not A166) );
 a77515a <=( A167  and  a77514a );
 a77518a <=( A202  and  (not A200) );
 a77521a <=( (not A265)  and  (not A203) );
 a77522a <=( a77521a  and  a77518a );
 a77523a <=( a77522a  and  a77515a );
 a77527a <=( (not A269)  and  A268 );
 a77528a <=( (not A266)  and  a77527a );
 a77531a <=( (not A299)  and  A298 );
 a77534a <=( (not A302)  and  (not A300) );
 a77535a <=( a77534a  and  a77531a );
 a77536a <=( a77535a  and  a77528a );
 a77540a <=( (not A199)  and  (not A166) );
 a77541a <=( A167  and  a77540a );
 a77544a <=( A202  and  (not A200) );
 a77547a <=( (not A265)  and  (not A203) );
 a77548a <=( a77547a  and  a77544a );
 a77549a <=( a77548a  and  a77541a );
 a77553a <=( (not A269)  and  A268 );
 a77554a <=( (not A266)  and  a77553a );
 a77557a <=( A299  and  (not A298) );
 a77560a <=( A301  and  (not A300) );
 a77561a <=( a77560a  and  a77557a );
 a77562a <=( a77561a  and  a77554a );
 a77566a <=( (not A199)  and  (not A166) );
 a77567a <=( A167  and  a77566a );
 a77570a <=( A202  and  (not A200) );
 a77573a <=( (not A265)  and  (not A203) );
 a77574a <=( a77573a  and  a77570a );
 a77575a <=( a77574a  and  a77567a );
 a77579a <=( (not A269)  and  A268 );
 a77580a <=( (not A266)  and  a77579a );
 a77583a <=( A299  and  (not A298) );
 a77586a <=( (not A302)  and  (not A300) );
 a77587a <=( a77586a  and  a77583a );
 a77588a <=( a77587a  and  a77580a );
 a77592a <=( A199  and  (not A166) );
 a77593a <=( (not A167)  and  a77592a );
 a77596a <=( A202  and  A200 );
 a77599a <=( A265  and  (not A203) );
 a77600a <=( a77599a  and  a77596a );
 a77601a <=( a77600a  and  a77593a );
 a77605a <=( (not A268)  and  (not A267) );
 a77606a <=( A266  and  a77605a );
 a77609a <=( A299  and  A298 );
 a77612a <=( (not A302)  and  A301 );
 a77613a <=( a77612a  and  a77609a );
 a77614a <=( a77613a  and  a77606a );
 a77618a <=( A199  and  (not A166) );
 a77619a <=( (not A167)  and  a77618a );
 a77622a <=( A202  and  A200 );
 a77625a <=( A265  and  (not A203) );
 a77626a <=( a77625a  and  a77622a );
 a77627a <=( a77626a  and  a77619a );
 a77631a <=( (not A268)  and  (not A267) );
 a77632a <=( A266  and  a77631a );
 a77635a <=( (not A299)  and  A298 );
 a77638a <=( A302  and  (not A301) );
 a77639a <=( a77638a  and  a77635a );
 a77640a <=( a77639a  and  a77632a );
 a77644a <=( A199  and  (not A166) );
 a77645a <=( (not A167)  and  a77644a );
 a77648a <=( A202  and  A200 );
 a77651a <=( A265  and  (not A203) );
 a77652a <=( a77651a  and  a77648a );
 a77653a <=( a77652a  and  a77645a );
 a77657a <=( (not A268)  and  (not A267) );
 a77658a <=( A266  and  a77657a );
 a77661a <=( A299  and  (not A298) );
 a77664a <=( A302  and  (not A301) );
 a77665a <=( a77664a  and  a77661a );
 a77666a <=( a77665a  and  a77658a );
 a77670a <=( A199  and  (not A166) );
 a77671a <=( (not A167)  and  a77670a );
 a77674a <=( A202  and  A200 );
 a77677a <=( A265  and  (not A203) );
 a77678a <=( a77677a  and  a77674a );
 a77679a <=( a77678a  and  a77671a );
 a77683a <=( (not A268)  and  (not A267) );
 a77684a <=( A266  and  a77683a );
 a77687a <=( (not A299)  and  (not A298) );
 a77690a <=( (not A302)  and  A301 );
 a77691a <=( a77690a  and  a77687a );
 a77692a <=( a77691a  and  a77684a );
 a77696a <=( A199  and  (not A166) );
 a77697a <=( (not A167)  and  a77696a );
 a77700a <=( A202  and  A200 );
 a77703a <=( A265  and  (not A203) );
 a77704a <=( a77703a  and  a77700a );
 a77705a <=( a77704a  and  a77697a );
 a77709a <=( A269  and  (not A267) );
 a77710a <=( A266  and  a77709a );
 a77713a <=( A299  and  A298 );
 a77716a <=( (not A302)  and  A301 );
 a77717a <=( a77716a  and  a77713a );
 a77718a <=( a77717a  and  a77710a );
 a77722a <=( A199  and  (not A166) );
 a77723a <=( (not A167)  and  a77722a );
 a77726a <=( A202  and  A200 );
 a77729a <=( A265  and  (not A203) );
 a77730a <=( a77729a  and  a77726a );
 a77731a <=( a77730a  and  a77723a );
 a77735a <=( A269  and  (not A267) );
 a77736a <=( A266  and  a77735a );
 a77739a <=( (not A299)  and  A298 );
 a77742a <=( A302  and  (not A301) );
 a77743a <=( a77742a  and  a77739a );
 a77744a <=( a77743a  and  a77736a );
 a77748a <=( A199  and  (not A166) );
 a77749a <=( (not A167)  and  a77748a );
 a77752a <=( A202  and  A200 );
 a77755a <=( A265  and  (not A203) );
 a77756a <=( a77755a  and  a77752a );
 a77757a <=( a77756a  and  a77749a );
 a77761a <=( A269  and  (not A267) );
 a77762a <=( A266  and  a77761a );
 a77765a <=( A299  and  (not A298) );
 a77768a <=( A302  and  (not A301) );
 a77769a <=( a77768a  and  a77765a );
 a77770a <=( a77769a  and  a77762a );
 a77774a <=( A199  and  (not A166) );
 a77775a <=( (not A167)  and  a77774a );
 a77778a <=( A202  and  A200 );
 a77781a <=( A265  and  (not A203) );
 a77782a <=( a77781a  and  a77778a );
 a77783a <=( a77782a  and  a77775a );
 a77787a <=( A269  and  (not A267) );
 a77788a <=( A266  and  a77787a );
 a77791a <=( (not A299)  and  (not A298) );
 a77794a <=( (not A302)  and  A301 );
 a77795a <=( a77794a  and  a77791a );
 a77796a <=( a77795a  and  a77788a );
 a77800a <=( A199  and  (not A166) );
 a77801a <=( (not A167)  and  a77800a );
 a77804a <=( A202  and  A200 );
 a77807a <=( (not A265)  and  (not A203) );
 a77808a <=( a77807a  and  a77804a );
 a77809a <=( a77808a  and  a77801a );
 a77813a <=( A268  and  (not A267) );
 a77814a <=( A266  and  a77813a );
 a77817a <=( A299  and  A298 );
 a77820a <=( (not A302)  and  A301 );
 a77821a <=( a77820a  and  a77817a );
 a77822a <=( a77821a  and  a77814a );
 a77826a <=( A199  and  (not A166) );
 a77827a <=( (not A167)  and  a77826a );
 a77830a <=( A202  and  A200 );
 a77833a <=( (not A265)  and  (not A203) );
 a77834a <=( a77833a  and  a77830a );
 a77835a <=( a77834a  and  a77827a );
 a77839a <=( A268  and  (not A267) );
 a77840a <=( A266  and  a77839a );
 a77843a <=( (not A299)  and  A298 );
 a77846a <=( A302  and  (not A301) );
 a77847a <=( a77846a  and  a77843a );
 a77848a <=( a77847a  and  a77840a );
 a77852a <=( A199  and  (not A166) );
 a77853a <=( (not A167)  and  a77852a );
 a77856a <=( A202  and  A200 );
 a77859a <=( (not A265)  and  (not A203) );
 a77860a <=( a77859a  and  a77856a );
 a77861a <=( a77860a  and  a77853a );
 a77865a <=( A268  and  (not A267) );
 a77866a <=( A266  and  a77865a );
 a77869a <=( A299  and  (not A298) );
 a77872a <=( A302  and  (not A301) );
 a77873a <=( a77872a  and  a77869a );
 a77874a <=( a77873a  and  a77866a );
 a77878a <=( A199  and  (not A166) );
 a77879a <=( (not A167)  and  a77878a );
 a77882a <=( A202  and  A200 );
 a77885a <=( (not A265)  and  (not A203) );
 a77886a <=( a77885a  and  a77882a );
 a77887a <=( a77886a  and  a77879a );
 a77891a <=( A268  and  (not A267) );
 a77892a <=( A266  and  a77891a );
 a77895a <=( (not A299)  and  (not A298) );
 a77898a <=( (not A302)  and  A301 );
 a77899a <=( a77898a  and  a77895a );
 a77900a <=( a77899a  and  a77892a );
 a77904a <=( A199  and  (not A166) );
 a77905a <=( (not A167)  and  a77904a );
 a77908a <=( A202  and  A200 );
 a77911a <=( (not A265)  and  (not A203) );
 a77912a <=( a77911a  and  a77908a );
 a77913a <=( a77912a  and  a77905a );
 a77917a <=( (not A269)  and  (not A267) );
 a77918a <=( A266  and  a77917a );
 a77921a <=( A299  and  A298 );
 a77924a <=( (not A302)  and  A301 );
 a77925a <=( a77924a  and  a77921a );
 a77926a <=( a77925a  and  a77918a );
 a77930a <=( A199  and  (not A166) );
 a77931a <=( (not A167)  and  a77930a );
 a77934a <=( A202  and  A200 );
 a77937a <=( (not A265)  and  (not A203) );
 a77938a <=( a77937a  and  a77934a );
 a77939a <=( a77938a  and  a77931a );
 a77943a <=( (not A269)  and  (not A267) );
 a77944a <=( A266  and  a77943a );
 a77947a <=( (not A299)  and  A298 );
 a77950a <=( A302  and  (not A301) );
 a77951a <=( a77950a  and  a77947a );
 a77952a <=( a77951a  and  a77944a );
 a77956a <=( A199  and  (not A166) );
 a77957a <=( (not A167)  and  a77956a );
 a77960a <=( A202  and  A200 );
 a77963a <=( (not A265)  and  (not A203) );
 a77964a <=( a77963a  and  a77960a );
 a77965a <=( a77964a  and  a77957a );
 a77969a <=( (not A269)  and  (not A267) );
 a77970a <=( A266  and  a77969a );
 a77973a <=( A299  and  (not A298) );
 a77976a <=( A302  and  (not A301) );
 a77977a <=( a77976a  and  a77973a );
 a77978a <=( a77977a  and  a77970a );
 a77982a <=( A199  and  (not A166) );
 a77983a <=( (not A167)  and  a77982a );
 a77986a <=( A202  and  A200 );
 a77989a <=( (not A265)  and  (not A203) );
 a77990a <=( a77989a  and  a77986a );
 a77991a <=( a77990a  and  a77983a );
 a77995a <=( (not A269)  and  (not A267) );
 a77996a <=( A266  and  a77995a );
 a77999a <=( (not A299)  and  (not A298) );
 a78002a <=( (not A302)  and  A301 );
 a78003a <=( a78002a  and  a77999a );
 a78004a <=( a78003a  and  a77996a );
 a78008a <=( A199  and  (not A166) );
 a78009a <=( (not A167)  and  a78008a );
 a78012a <=( A202  and  A200 );
 a78015a <=( A265  and  (not A203) );
 a78016a <=( a78015a  and  a78012a );
 a78017a <=( a78016a  and  a78009a );
 a78021a <=( A268  and  (not A267) );
 a78022a <=( (not A266)  and  a78021a );
 a78025a <=( A299  and  A298 );
 a78028a <=( (not A302)  and  A301 );
 a78029a <=( a78028a  and  a78025a );
 a78030a <=( a78029a  and  a78022a );
 a78034a <=( A199  and  (not A166) );
 a78035a <=( (not A167)  and  a78034a );
 a78038a <=( A202  and  A200 );
 a78041a <=( A265  and  (not A203) );
 a78042a <=( a78041a  and  a78038a );
 a78043a <=( a78042a  and  a78035a );
 a78047a <=( A268  and  (not A267) );
 a78048a <=( (not A266)  and  a78047a );
 a78051a <=( (not A299)  and  A298 );
 a78054a <=( A302  and  (not A301) );
 a78055a <=( a78054a  and  a78051a );
 a78056a <=( a78055a  and  a78048a );
 a78060a <=( A199  and  (not A166) );
 a78061a <=( (not A167)  and  a78060a );
 a78064a <=( A202  and  A200 );
 a78067a <=( A265  and  (not A203) );
 a78068a <=( a78067a  and  a78064a );
 a78069a <=( a78068a  and  a78061a );
 a78073a <=( A268  and  (not A267) );
 a78074a <=( (not A266)  and  a78073a );
 a78077a <=( A299  and  (not A298) );
 a78080a <=( A302  and  (not A301) );
 a78081a <=( a78080a  and  a78077a );
 a78082a <=( a78081a  and  a78074a );
 a78086a <=( A199  and  (not A166) );
 a78087a <=( (not A167)  and  a78086a );
 a78090a <=( A202  and  A200 );
 a78093a <=( A265  and  (not A203) );
 a78094a <=( a78093a  and  a78090a );
 a78095a <=( a78094a  and  a78087a );
 a78099a <=( A268  and  (not A267) );
 a78100a <=( (not A266)  and  a78099a );
 a78103a <=( (not A299)  and  (not A298) );
 a78106a <=( (not A302)  and  A301 );
 a78107a <=( a78106a  and  a78103a );
 a78108a <=( a78107a  and  a78100a );
 a78112a <=( A199  and  (not A166) );
 a78113a <=( (not A167)  and  a78112a );
 a78116a <=( A202  and  A200 );
 a78119a <=( A265  and  (not A203) );
 a78120a <=( a78119a  and  a78116a );
 a78121a <=( a78120a  and  a78113a );
 a78125a <=( (not A269)  and  (not A267) );
 a78126a <=( (not A266)  and  a78125a );
 a78129a <=( A299  and  A298 );
 a78132a <=( (not A302)  and  A301 );
 a78133a <=( a78132a  and  a78129a );
 a78134a <=( a78133a  and  a78126a );
 a78138a <=( A199  and  (not A166) );
 a78139a <=( (not A167)  and  a78138a );
 a78142a <=( A202  and  A200 );
 a78145a <=( A265  and  (not A203) );
 a78146a <=( a78145a  and  a78142a );
 a78147a <=( a78146a  and  a78139a );
 a78151a <=( (not A269)  and  (not A267) );
 a78152a <=( (not A266)  and  a78151a );
 a78155a <=( (not A299)  and  A298 );
 a78158a <=( A302  and  (not A301) );
 a78159a <=( a78158a  and  a78155a );
 a78160a <=( a78159a  and  a78152a );
 a78164a <=( A199  and  (not A166) );
 a78165a <=( (not A167)  and  a78164a );
 a78168a <=( A202  and  A200 );
 a78171a <=( A265  and  (not A203) );
 a78172a <=( a78171a  and  a78168a );
 a78173a <=( a78172a  and  a78165a );
 a78177a <=( (not A269)  and  (not A267) );
 a78178a <=( (not A266)  and  a78177a );
 a78181a <=( A299  and  (not A298) );
 a78184a <=( A302  and  (not A301) );
 a78185a <=( a78184a  and  a78181a );
 a78186a <=( a78185a  and  a78178a );
 a78190a <=( A199  and  (not A166) );
 a78191a <=( (not A167)  and  a78190a );
 a78194a <=( A202  and  A200 );
 a78197a <=( A265  and  (not A203) );
 a78198a <=( a78197a  and  a78194a );
 a78199a <=( a78198a  and  a78191a );
 a78203a <=( (not A269)  and  (not A267) );
 a78204a <=( (not A266)  and  a78203a );
 a78207a <=( (not A299)  and  (not A298) );
 a78210a <=( (not A302)  and  A301 );
 a78211a <=( a78210a  and  a78207a );
 a78212a <=( a78211a  and  a78204a );
 a78216a <=( A199  and  (not A166) );
 a78217a <=( (not A167)  and  a78216a );
 a78220a <=( (not A201)  and  A200 );
 a78223a <=( A265  and  (not A202) );
 a78224a <=( a78223a  and  a78220a );
 a78225a <=( a78224a  and  a78217a );
 a78229a <=( (not A269)  and  A268 );
 a78230a <=( A266  and  a78229a );
 a78233a <=( A299  and  A298 );
 a78236a <=( (not A301)  and  (not A300) );
 a78237a <=( a78236a  and  a78233a );
 a78238a <=( a78237a  and  a78230a );
 a78242a <=( A199  and  (not A166) );
 a78243a <=( (not A167)  and  a78242a );
 a78246a <=( (not A201)  and  A200 );
 a78249a <=( A265  and  (not A202) );
 a78250a <=( a78249a  and  a78246a );
 a78251a <=( a78250a  and  a78243a );
 a78255a <=( (not A269)  and  A268 );
 a78256a <=( A266  and  a78255a );
 a78259a <=( A299  and  A298 );
 a78262a <=( A302  and  (not A300) );
 a78263a <=( a78262a  and  a78259a );
 a78264a <=( a78263a  and  a78256a );
 a78268a <=( A199  and  (not A166) );
 a78269a <=( (not A167)  and  a78268a );
 a78272a <=( (not A201)  and  A200 );
 a78275a <=( A265  and  (not A202) );
 a78276a <=( a78275a  and  a78272a );
 a78277a <=( a78276a  and  a78269a );
 a78281a <=( (not A269)  and  A268 );
 a78282a <=( A266  and  a78281a );
 a78285a <=( (not A299)  and  A298 );
 a78288a <=( A301  and  (not A300) );
 a78289a <=( a78288a  and  a78285a );
 a78290a <=( a78289a  and  a78282a );
 a78294a <=( A199  and  (not A166) );
 a78295a <=( (not A167)  and  a78294a );
 a78298a <=( (not A201)  and  A200 );
 a78301a <=( A265  and  (not A202) );
 a78302a <=( a78301a  and  a78298a );
 a78303a <=( a78302a  and  a78295a );
 a78307a <=( (not A269)  and  A268 );
 a78308a <=( A266  and  a78307a );
 a78311a <=( (not A299)  and  A298 );
 a78314a <=( (not A302)  and  (not A300) );
 a78315a <=( a78314a  and  a78311a );
 a78316a <=( a78315a  and  a78308a );
 a78320a <=( A199  and  (not A166) );
 a78321a <=( (not A167)  and  a78320a );
 a78324a <=( (not A201)  and  A200 );
 a78327a <=( A265  and  (not A202) );
 a78328a <=( a78327a  and  a78324a );
 a78329a <=( a78328a  and  a78321a );
 a78333a <=( (not A269)  and  A268 );
 a78334a <=( A266  and  a78333a );
 a78337a <=( A299  and  (not A298) );
 a78340a <=( A301  and  (not A300) );
 a78341a <=( a78340a  and  a78337a );
 a78342a <=( a78341a  and  a78334a );
 a78346a <=( A199  and  (not A166) );
 a78347a <=( (not A167)  and  a78346a );
 a78350a <=( (not A201)  and  A200 );
 a78353a <=( A265  and  (not A202) );
 a78354a <=( a78353a  and  a78350a );
 a78355a <=( a78354a  and  a78347a );
 a78359a <=( (not A269)  and  A268 );
 a78360a <=( A266  and  a78359a );
 a78363a <=( A299  and  (not A298) );
 a78366a <=( (not A302)  and  (not A300) );
 a78367a <=( a78366a  and  a78363a );
 a78368a <=( a78367a  and  a78360a );
 a78372a <=( A199  and  (not A166) );
 a78373a <=( (not A167)  and  a78372a );
 a78376a <=( (not A201)  and  A200 );
 a78379a <=( (not A265)  and  (not A202) );
 a78380a <=( a78379a  and  a78376a );
 a78381a <=( a78380a  and  a78373a );
 a78385a <=( A269  and  (not A268) );
 a78386a <=( A266  and  a78385a );
 a78389a <=( A299  and  A298 );
 a78392a <=( (not A301)  and  (not A300) );
 a78393a <=( a78392a  and  a78389a );
 a78394a <=( a78393a  and  a78386a );
 a78398a <=( A199  and  (not A166) );
 a78399a <=( (not A167)  and  a78398a );
 a78402a <=( (not A201)  and  A200 );
 a78405a <=( (not A265)  and  (not A202) );
 a78406a <=( a78405a  and  a78402a );
 a78407a <=( a78406a  and  a78399a );
 a78411a <=( A269  and  (not A268) );
 a78412a <=( A266  and  a78411a );
 a78415a <=( A299  and  A298 );
 a78418a <=( A302  and  (not A300) );
 a78419a <=( a78418a  and  a78415a );
 a78420a <=( a78419a  and  a78412a );
 a78424a <=( A199  and  (not A166) );
 a78425a <=( (not A167)  and  a78424a );
 a78428a <=( (not A201)  and  A200 );
 a78431a <=( (not A265)  and  (not A202) );
 a78432a <=( a78431a  and  a78428a );
 a78433a <=( a78432a  and  a78425a );
 a78437a <=( A269  and  (not A268) );
 a78438a <=( A266  and  a78437a );
 a78441a <=( (not A299)  and  A298 );
 a78444a <=( A301  and  (not A300) );
 a78445a <=( a78444a  and  a78441a );
 a78446a <=( a78445a  and  a78438a );
 a78450a <=( A199  and  (not A166) );
 a78451a <=( (not A167)  and  a78450a );
 a78454a <=( (not A201)  and  A200 );
 a78457a <=( (not A265)  and  (not A202) );
 a78458a <=( a78457a  and  a78454a );
 a78459a <=( a78458a  and  a78451a );
 a78463a <=( A269  and  (not A268) );
 a78464a <=( A266  and  a78463a );
 a78467a <=( (not A299)  and  A298 );
 a78470a <=( (not A302)  and  (not A300) );
 a78471a <=( a78470a  and  a78467a );
 a78472a <=( a78471a  and  a78464a );
 a78476a <=( A199  and  (not A166) );
 a78477a <=( (not A167)  and  a78476a );
 a78480a <=( (not A201)  and  A200 );
 a78483a <=( (not A265)  and  (not A202) );
 a78484a <=( a78483a  and  a78480a );
 a78485a <=( a78484a  and  a78477a );
 a78489a <=( A269  and  (not A268) );
 a78490a <=( A266  and  a78489a );
 a78493a <=( A299  and  (not A298) );
 a78496a <=( A301  and  (not A300) );
 a78497a <=( a78496a  and  a78493a );
 a78498a <=( a78497a  and  a78490a );
 a78502a <=( A199  and  (not A166) );
 a78503a <=( (not A167)  and  a78502a );
 a78506a <=( (not A201)  and  A200 );
 a78509a <=( (not A265)  and  (not A202) );
 a78510a <=( a78509a  and  a78506a );
 a78511a <=( a78510a  and  a78503a );
 a78515a <=( A269  and  (not A268) );
 a78516a <=( A266  and  a78515a );
 a78519a <=( A299  and  (not A298) );
 a78522a <=( (not A302)  and  (not A300) );
 a78523a <=( a78522a  and  a78519a );
 a78524a <=( a78523a  and  a78516a );
 a78528a <=( A199  and  (not A166) );
 a78529a <=( (not A167)  and  a78528a );
 a78532a <=( (not A201)  and  A200 );
 a78535a <=( A265  and  (not A202) );
 a78536a <=( a78535a  and  a78532a );
 a78537a <=( a78536a  and  a78529a );
 a78541a <=( A269  and  (not A268) );
 a78542a <=( (not A266)  and  a78541a );
 a78545a <=( A299  and  A298 );
 a78548a <=( (not A301)  and  (not A300) );
 a78549a <=( a78548a  and  a78545a );
 a78550a <=( a78549a  and  a78542a );
 a78554a <=( A199  and  (not A166) );
 a78555a <=( (not A167)  and  a78554a );
 a78558a <=( (not A201)  and  A200 );
 a78561a <=( A265  and  (not A202) );
 a78562a <=( a78561a  and  a78558a );
 a78563a <=( a78562a  and  a78555a );
 a78567a <=( A269  and  (not A268) );
 a78568a <=( (not A266)  and  a78567a );
 a78571a <=( A299  and  A298 );
 a78574a <=( A302  and  (not A300) );
 a78575a <=( a78574a  and  a78571a );
 a78576a <=( a78575a  and  a78568a );
 a78580a <=( A199  and  (not A166) );
 a78581a <=( (not A167)  and  a78580a );
 a78584a <=( (not A201)  and  A200 );
 a78587a <=( A265  and  (not A202) );
 a78588a <=( a78587a  and  a78584a );
 a78589a <=( a78588a  and  a78581a );
 a78593a <=( A269  and  (not A268) );
 a78594a <=( (not A266)  and  a78593a );
 a78597a <=( (not A299)  and  A298 );
 a78600a <=( A301  and  (not A300) );
 a78601a <=( a78600a  and  a78597a );
 a78602a <=( a78601a  and  a78594a );
 a78606a <=( A199  and  (not A166) );
 a78607a <=( (not A167)  and  a78606a );
 a78610a <=( (not A201)  and  A200 );
 a78613a <=( A265  and  (not A202) );
 a78614a <=( a78613a  and  a78610a );
 a78615a <=( a78614a  and  a78607a );
 a78619a <=( A269  and  (not A268) );
 a78620a <=( (not A266)  and  a78619a );
 a78623a <=( (not A299)  and  A298 );
 a78626a <=( (not A302)  and  (not A300) );
 a78627a <=( a78626a  and  a78623a );
 a78628a <=( a78627a  and  a78620a );
 a78632a <=( A199  and  (not A166) );
 a78633a <=( (not A167)  and  a78632a );
 a78636a <=( (not A201)  and  A200 );
 a78639a <=( A265  and  (not A202) );
 a78640a <=( a78639a  and  a78636a );
 a78641a <=( a78640a  and  a78633a );
 a78645a <=( A269  and  (not A268) );
 a78646a <=( (not A266)  and  a78645a );
 a78649a <=( A299  and  (not A298) );
 a78652a <=( A301  and  (not A300) );
 a78653a <=( a78652a  and  a78649a );
 a78654a <=( a78653a  and  a78646a );
 a78658a <=( A199  and  (not A166) );
 a78659a <=( (not A167)  and  a78658a );
 a78662a <=( (not A201)  and  A200 );
 a78665a <=( A265  and  (not A202) );
 a78666a <=( a78665a  and  a78662a );
 a78667a <=( a78666a  and  a78659a );
 a78671a <=( A269  and  (not A268) );
 a78672a <=( (not A266)  and  a78671a );
 a78675a <=( A299  and  (not A298) );
 a78678a <=( (not A302)  and  (not A300) );
 a78679a <=( a78678a  and  a78675a );
 a78680a <=( a78679a  and  a78672a );
 a78684a <=( A199  and  (not A166) );
 a78685a <=( (not A167)  and  a78684a );
 a78688a <=( (not A201)  and  A200 );
 a78691a <=( (not A265)  and  (not A202) );
 a78692a <=( a78691a  and  a78688a );
 a78693a <=( a78692a  and  a78685a );
 a78697a <=( (not A269)  and  A268 );
 a78698a <=( (not A266)  and  a78697a );
 a78701a <=( A299  and  A298 );
 a78704a <=( (not A301)  and  (not A300) );
 a78705a <=( a78704a  and  a78701a );
 a78706a <=( a78705a  and  a78698a );
 a78710a <=( A199  and  (not A166) );
 a78711a <=( (not A167)  and  a78710a );
 a78714a <=( (not A201)  and  A200 );
 a78717a <=( (not A265)  and  (not A202) );
 a78718a <=( a78717a  and  a78714a );
 a78719a <=( a78718a  and  a78711a );
 a78723a <=( (not A269)  and  A268 );
 a78724a <=( (not A266)  and  a78723a );
 a78727a <=( A299  and  A298 );
 a78730a <=( A302  and  (not A300) );
 a78731a <=( a78730a  and  a78727a );
 a78732a <=( a78731a  and  a78724a );
 a78736a <=( A199  and  (not A166) );
 a78737a <=( (not A167)  and  a78736a );
 a78740a <=( (not A201)  and  A200 );
 a78743a <=( (not A265)  and  (not A202) );
 a78744a <=( a78743a  and  a78740a );
 a78745a <=( a78744a  and  a78737a );
 a78749a <=( (not A269)  and  A268 );
 a78750a <=( (not A266)  and  a78749a );
 a78753a <=( (not A299)  and  A298 );
 a78756a <=( A301  and  (not A300) );
 a78757a <=( a78756a  and  a78753a );
 a78758a <=( a78757a  and  a78750a );
 a78762a <=( A199  and  (not A166) );
 a78763a <=( (not A167)  and  a78762a );
 a78766a <=( (not A201)  and  A200 );
 a78769a <=( (not A265)  and  (not A202) );
 a78770a <=( a78769a  and  a78766a );
 a78771a <=( a78770a  and  a78763a );
 a78775a <=( (not A269)  and  A268 );
 a78776a <=( (not A266)  and  a78775a );
 a78779a <=( (not A299)  and  A298 );
 a78782a <=( (not A302)  and  (not A300) );
 a78783a <=( a78782a  and  a78779a );
 a78784a <=( a78783a  and  a78776a );
 a78788a <=( A199  and  (not A166) );
 a78789a <=( (not A167)  and  a78788a );
 a78792a <=( (not A201)  and  A200 );
 a78795a <=( (not A265)  and  (not A202) );
 a78796a <=( a78795a  and  a78792a );
 a78797a <=( a78796a  and  a78789a );
 a78801a <=( (not A269)  and  A268 );
 a78802a <=( (not A266)  and  a78801a );
 a78805a <=( A299  and  (not A298) );
 a78808a <=( A301  and  (not A300) );
 a78809a <=( a78808a  and  a78805a );
 a78810a <=( a78809a  and  a78802a );
 a78814a <=( A199  and  (not A166) );
 a78815a <=( (not A167)  and  a78814a );
 a78818a <=( (not A201)  and  A200 );
 a78821a <=( (not A265)  and  (not A202) );
 a78822a <=( a78821a  and  a78818a );
 a78823a <=( a78822a  and  a78815a );
 a78827a <=( (not A269)  and  A268 );
 a78828a <=( (not A266)  and  a78827a );
 a78831a <=( A299  and  (not A298) );
 a78834a <=( (not A302)  and  (not A300) );
 a78835a <=( a78834a  and  a78831a );
 a78836a <=( a78835a  and  a78828a );
 a78840a <=( A199  and  (not A166) );
 a78841a <=( (not A167)  and  a78840a );
 a78844a <=( (not A201)  and  A200 );
 a78847a <=( A265  and  A203 );
 a78848a <=( a78847a  and  a78844a );
 a78849a <=( a78848a  and  a78841a );
 a78853a <=( (not A269)  and  A268 );
 a78854a <=( A266  and  a78853a );
 a78857a <=( A299  and  A298 );
 a78860a <=( (not A301)  and  (not A300) );
 a78861a <=( a78860a  and  a78857a );
 a78862a <=( a78861a  and  a78854a );
 a78866a <=( A199  and  (not A166) );
 a78867a <=( (not A167)  and  a78866a );
 a78870a <=( (not A201)  and  A200 );
 a78873a <=( A265  and  A203 );
 a78874a <=( a78873a  and  a78870a );
 a78875a <=( a78874a  and  a78867a );
 a78879a <=( (not A269)  and  A268 );
 a78880a <=( A266  and  a78879a );
 a78883a <=( A299  and  A298 );
 a78886a <=( A302  and  (not A300) );
 a78887a <=( a78886a  and  a78883a );
 a78888a <=( a78887a  and  a78880a );
 a78892a <=( A199  and  (not A166) );
 a78893a <=( (not A167)  and  a78892a );
 a78896a <=( (not A201)  and  A200 );
 a78899a <=( A265  and  A203 );
 a78900a <=( a78899a  and  a78896a );
 a78901a <=( a78900a  and  a78893a );
 a78905a <=( (not A269)  and  A268 );
 a78906a <=( A266  and  a78905a );
 a78909a <=( (not A299)  and  A298 );
 a78912a <=( A301  and  (not A300) );
 a78913a <=( a78912a  and  a78909a );
 a78914a <=( a78913a  and  a78906a );
 a78918a <=( A199  and  (not A166) );
 a78919a <=( (not A167)  and  a78918a );
 a78922a <=( (not A201)  and  A200 );
 a78925a <=( A265  and  A203 );
 a78926a <=( a78925a  and  a78922a );
 a78927a <=( a78926a  and  a78919a );
 a78931a <=( (not A269)  and  A268 );
 a78932a <=( A266  and  a78931a );
 a78935a <=( (not A299)  and  A298 );
 a78938a <=( (not A302)  and  (not A300) );
 a78939a <=( a78938a  and  a78935a );
 a78940a <=( a78939a  and  a78932a );
 a78944a <=( A199  and  (not A166) );
 a78945a <=( (not A167)  and  a78944a );
 a78948a <=( (not A201)  and  A200 );
 a78951a <=( A265  and  A203 );
 a78952a <=( a78951a  and  a78948a );
 a78953a <=( a78952a  and  a78945a );
 a78957a <=( (not A269)  and  A268 );
 a78958a <=( A266  and  a78957a );
 a78961a <=( A299  and  (not A298) );
 a78964a <=( A301  and  (not A300) );
 a78965a <=( a78964a  and  a78961a );
 a78966a <=( a78965a  and  a78958a );
 a78970a <=( A199  and  (not A166) );
 a78971a <=( (not A167)  and  a78970a );
 a78974a <=( (not A201)  and  A200 );
 a78977a <=( A265  and  A203 );
 a78978a <=( a78977a  and  a78974a );
 a78979a <=( a78978a  and  a78971a );
 a78983a <=( (not A269)  and  A268 );
 a78984a <=( A266  and  a78983a );
 a78987a <=( A299  and  (not A298) );
 a78990a <=( (not A302)  and  (not A300) );
 a78991a <=( a78990a  and  a78987a );
 a78992a <=( a78991a  and  a78984a );
 a78996a <=( A199  and  (not A166) );
 a78997a <=( (not A167)  and  a78996a );
 a79000a <=( (not A201)  and  A200 );
 a79003a <=( (not A265)  and  A203 );
 a79004a <=( a79003a  and  a79000a );
 a79005a <=( a79004a  and  a78997a );
 a79009a <=( A269  and  (not A268) );
 a79010a <=( A266  and  a79009a );
 a79013a <=( A299  and  A298 );
 a79016a <=( (not A301)  and  (not A300) );
 a79017a <=( a79016a  and  a79013a );
 a79018a <=( a79017a  and  a79010a );
 a79022a <=( A199  and  (not A166) );
 a79023a <=( (not A167)  and  a79022a );
 a79026a <=( (not A201)  and  A200 );
 a79029a <=( (not A265)  and  A203 );
 a79030a <=( a79029a  and  a79026a );
 a79031a <=( a79030a  and  a79023a );
 a79035a <=( A269  and  (not A268) );
 a79036a <=( A266  and  a79035a );
 a79039a <=( A299  and  A298 );
 a79042a <=( A302  and  (not A300) );
 a79043a <=( a79042a  and  a79039a );
 a79044a <=( a79043a  and  a79036a );
 a79048a <=( A199  and  (not A166) );
 a79049a <=( (not A167)  and  a79048a );
 a79052a <=( (not A201)  and  A200 );
 a79055a <=( (not A265)  and  A203 );
 a79056a <=( a79055a  and  a79052a );
 a79057a <=( a79056a  and  a79049a );
 a79061a <=( A269  and  (not A268) );
 a79062a <=( A266  and  a79061a );
 a79065a <=( (not A299)  and  A298 );
 a79068a <=( A301  and  (not A300) );
 a79069a <=( a79068a  and  a79065a );
 a79070a <=( a79069a  and  a79062a );
 a79074a <=( A199  and  (not A166) );
 a79075a <=( (not A167)  and  a79074a );
 a79078a <=( (not A201)  and  A200 );
 a79081a <=( (not A265)  and  A203 );
 a79082a <=( a79081a  and  a79078a );
 a79083a <=( a79082a  and  a79075a );
 a79087a <=( A269  and  (not A268) );
 a79088a <=( A266  and  a79087a );
 a79091a <=( (not A299)  and  A298 );
 a79094a <=( (not A302)  and  (not A300) );
 a79095a <=( a79094a  and  a79091a );
 a79096a <=( a79095a  and  a79088a );
 a79100a <=( A199  and  (not A166) );
 a79101a <=( (not A167)  and  a79100a );
 a79104a <=( (not A201)  and  A200 );
 a79107a <=( (not A265)  and  A203 );
 a79108a <=( a79107a  and  a79104a );
 a79109a <=( a79108a  and  a79101a );
 a79113a <=( A269  and  (not A268) );
 a79114a <=( A266  and  a79113a );
 a79117a <=( A299  and  (not A298) );
 a79120a <=( A301  and  (not A300) );
 a79121a <=( a79120a  and  a79117a );
 a79122a <=( a79121a  and  a79114a );
 a79126a <=( A199  and  (not A166) );
 a79127a <=( (not A167)  and  a79126a );
 a79130a <=( (not A201)  and  A200 );
 a79133a <=( (not A265)  and  A203 );
 a79134a <=( a79133a  and  a79130a );
 a79135a <=( a79134a  and  a79127a );
 a79139a <=( A269  and  (not A268) );
 a79140a <=( A266  and  a79139a );
 a79143a <=( A299  and  (not A298) );
 a79146a <=( (not A302)  and  (not A300) );
 a79147a <=( a79146a  and  a79143a );
 a79148a <=( a79147a  and  a79140a );
 a79152a <=( A199  and  (not A166) );
 a79153a <=( (not A167)  and  a79152a );
 a79156a <=( (not A201)  and  A200 );
 a79159a <=( A265  and  A203 );
 a79160a <=( a79159a  and  a79156a );
 a79161a <=( a79160a  and  a79153a );
 a79165a <=( A269  and  (not A268) );
 a79166a <=( (not A266)  and  a79165a );
 a79169a <=( A299  and  A298 );
 a79172a <=( (not A301)  and  (not A300) );
 a79173a <=( a79172a  and  a79169a );
 a79174a <=( a79173a  and  a79166a );
 a79178a <=( A199  and  (not A166) );
 a79179a <=( (not A167)  and  a79178a );
 a79182a <=( (not A201)  and  A200 );
 a79185a <=( A265  and  A203 );
 a79186a <=( a79185a  and  a79182a );
 a79187a <=( a79186a  and  a79179a );
 a79191a <=( A269  and  (not A268) );
 a79192a <=( (not A266)  and  a79191a );
 a79195a <=( A299  and  A298 );
 a79198a <=( A302  and  (not A300) );
 a79199a <=( a79198a  and  a79195a );
 a79200a <=( a79199a  and  a79192a );
 a79204a <=( A199  and  (not A166) );
 a79205a <=( (not A167)  and  a79204a );
 a79208a <=( (not A201)  and  A200 );
 a79211a <=( A265  and  A203 );
 a79212a <=( a79211a  and  a79208a );
 a79213a <=( a79212a  and  a79205a );
 a79217a <=( A269  and  (not A268) );
 a79218a <=( (not A266)  and  a79217a );
 a79221a <=( (not A299)  and  A298 );
 a79224a <=( A301  and  (not A300) );
 a79225a <=( a79224a  and  a79221a );
 a79226a <=( a79225a  and  a79218a );
 a79230a <=( A199  and  (not A166) );
 a79231a <=( (not A167)  and  a79230a );
 a79234a <=( (not A201)  and  A200 );
 a79237a <=( A265  and  A203 );
 a79238a <=( a79237a  and  a79234a );
 a79239a <=( a79238a  and  a79231a );
 a79243a <=( A269  and  (not A268) );
 a79244a <=( (not A266)  and  a79243a );
 a79247a <=( (not A299)  and  A298 );
 a79250a <=( (not A302)  and  (not A300) );
 a79251a <=( a79250a  and  a79247a );
 a79252a <=( a79251a  and  a79244a );
 a79256a <=( A199  and  (not A166) );
 a79257a <=( (not A167)  and  a79256a );
 a79260a <=( (not A201)  and  A200 );
 a79263a <=( A265  and  A203 );
 a79264a <=( a79263a  and  a79260a );
 a79265a <=( a79264a  and  a79257a );
 a79269a <=( A269  and  (not A268) );
 a79270a <=( (not A266)  and  a79269a );
 a79273a <=( A299  and  (not A298) );
 a79276a <=( A301  and  (not A300) );
 a79277a <=( a79276a  and  a79273a );
 a79278a <=( a79277a  and  a79270a );
 a79282a <=( A199  and  (not A166) );
 a79283a <=( (not A167)  and  a79282a );
 a79286a <=( (not A201)  and  A200 );
 a79289a <=( A265  and  A203 );
 a79290a <=( a79289a  and  a79286a );
 a79291a <=( a79290a  and  a79283a );
 a79295a <=( A269  and  (not A268) );
 a79296a <=( (not A266)  and  a79295a );
 a79299a <=( A299  and  (not A298) );
 a79302a <=( (not A302)  and  (not A300) );
 a79303a <=( a79302a  and  a79299a );
 a79304a <=( a79303a  and  a79296a );
 a79308a <=( A199  and  (not A166) );
 a79309a <=( (not A167)  and  a79308a );
 a79312a <=( (not A201)  and  A200 );
 a79315a <=( (not A265)  and  A203 );
 a79316a <=( a79315a  and  a79312a );
 a79317a <=( a79316a  and  a79309a );
 a79321a <=( (not A269)  and  A268 );
 a79322a <=( (not A266)  and  a79321a );
 a79325a <=( A299  and  A298 );
 a79328a <=( (not A301)  and  (not A300) );
 a79329a <=( a79328a  and  a79325a );
 a79330a <=( a79329a  and  a79322a );
 a79334a <=( A199  and  (not A166) );
 a79335a <=( (not A167)  and  a79334a );
 a79338a <=( (not A201)  and  A200 );
 a79341a <=( (not A265)  and  A203 );
 a79342a <=( a79341a  and  a79338a );
 a79343a <=( a79342a  and  a79335a );
 a79347a <=( (not A269)  and  A268 );
 a79348a <=( (not A266)  and  a79347a );
 a79351a <=( A299  and  A298 );
 a79354a <=( A302  and  (not A300) );
 a79355a <=( a79354a  and  a79351a );
 a79356a <=( a79355a  and  a79348a );
 a79360a <=( A199  and  (not A166) );
 a79361a <=( (not A167)  and  a79360a );
 a79364a <=( (not A201)  and  A200 );
 a79367a <=( (not A265)  and  A203 );
 a79368a <=( a79367a  and  a79364a );
 a79369a <=( a79368a  and  a79361a );
 a79373a <=( (not A269)  and  A268 );
 a79374a <=( (not A266)  and  a79373a );
 a79377a <=( (not A299)  and  A298 );
 a79380a <=( A301  and  (not A300) );
 a79381a <=( a79380a  and  a79377a );
 a79382a <=( a79381a  and  a79374a );
 a79386a <=( A199  and  (not A166) );
 a79387a <=( (not A167)  and  a79386a );
 a79390a <=( (not A201)  and  A200 );
 a79393a <=( (not A265)  and  A203 );
 a79394a <=( a79393a  and  a79390a );
 a79395a <=( a79394a  and  a79387a );
 a79399a <=( (not A269)  and  A268 );
 a79400a <=( (not A266)  and  a79399a );
 a79403a <=( (not A299)  and  A298 );
 a79406a <=( (not A302)  and  (not A300) );
 a79407a <=( a79406a  and  a79403a );
 a79408a <=( a79407a  and  a79400a );
 a79412a <=( A199  and  (not A166) );
 a79413a <=( (not A167)  and  a79412a );
 a79416a <=( (not A201)  and  A200 );
 a79419a <=( (not A265)  and  A203 );
 a79420a <=( a79419a  and  a79416a );
 a79421a <=( a79420a  and  a79413a );
 a79425a <=( (not A269)  and  A268 );
 a79426a <=( (not A266)  and  a79425a );
 a79429a <=( A299  and  (not A298) );
 a79432a <=( A301  and  (not A300) );
 a79433a <=( a79432a  and  a79429a );
 a79434a <=( a79433a  and  a79426a );
 a79438a <=( A199  and  (not A166) );
 a79439a <=( (not A167)  and  a79438a );
 a79442a <=( (not A201)  and  A200 );
 a79445a <=( (not A265)  and  A203 );
 a79446a <=( a79445a  and  a79442a );
 a79447a <=( a79446a  and  a79439a );
 a79451a <=( (not A269)  and  A268 );
 a79452a <=( (not A266)  and  a79451a );
 a79455a <=( A299  and  (not A298) );
 a79458a <=( (not A302)  and  (not A300) );
 a79459a <=( a79458a  and  a79455a );
 a79460a <=( a79459a  and  a79452a );
 a79464a <=( (not A199)  and  (not A166) );
 a79465a <=( (not A167)  and  a79464a );
 a79468a <=( (not A202)  and  A200 );
 a79471a <=( A265  and  A203 );
 a79472a <=( a79471a  and  a79468a );
 a79473a <=( a79472a  and  a79465a );
 a79477a <=( (not A268)  and  (not A267) );
 a79478a <=( A266  and  a79477a );
 a79481a <=( A299  and  A298 );
 a79484a <=( (not A302)  and  A301 );
 a79485a <=( a79484a  and  a79481a );
 a79486a <=( a79485a  and  a79478a );
 a79490a <=( (not A199)  and  (not A166) );
 a79491a <=( (not A167)  and  a79490a );
 a79494a <=( (not A202)  and  A200 );
 a79497a <=( A265  and  A203 );
 a79498a <=( a79497a  and  a79494a );
 a79499a <=( a79498a  and  a79491a );
 a79503a <=( (not A268)  and  (not A267) );
 a79504a <=( A266  and  a79503a );
 a79507a <=( (not A299)  and  A298 );
 a79510a <=( A302  and  (not A301) );
 a79511a <=( a79510a  and  a79507a );
 a79512a <=( a79511a  and  a79504a );
 a79516a <=( (not A199)  and  (not A166) );
 a79517a <=( (not A167)  and  a79516a );
 a79520a <=( (not A202)  and  A200 );
 a79523a <=( A265  and  A203 );
 a79524a <=( a79523a  and  a79520a );
 a79525a <=( a79524a  and  a79517a );
 a79529a <=( (not A268)  and  (not A267) );
 a79530a <=( A266  and  a79529a );
 a79533a <=( A299  and  (not A298) );
 a79536a <=( A302  and  (not A301) );
 a79537a <=( a79536a  and  a79533a );
 a79538a <=( a79537a  and  a79530a );
 a79542a <=( (not A199)  and  (not A166) );
 a79543a <=( (not A167)  and  a79542a );
 a79546a <=( (not A202)  and  A200 );
 a79549a <=( A265  and  A203 );
 a79550a <=( a79549a  and  a79546a );
 a79551a <=( a79550a  and  a79543a );
 a79555a <=( (not A268)  and  (not A267) );
 a79556a <=( A266  and  a79555a );
 a79559a <=( (not A299)  and  (not A298) );
 a79562a <=( (not A302)  and  A301 );
 a79563a <=( a79562a  and  a79559a );
 a79564a <=( a79563a  and  a79556a );
 a79568a <=( (not A199)  and  (not A166) );
 a79569a <=( (not A167)  and  a79568a );
 a79572a <=( (not A202)  and  A200 );
 a79575a <=( A265  and  A203 );
 a79576a <=( a79575a  and  a79572a );
 a79577a <=( a79576a  and  a79569a );
 a79581a <=( A269  and  (not A267) );
 a79582a <=( A266  and  a79581a );
 a79585a <=( A299  and  A298 );
 a79588a <=( (not A302)  and  A301 );
 a79589a <=( a79588a  and  a79585a );
 a79590a <=( a79589a  and  a79582a );
 a79594a <=( (not A199)  and  (not A166) );
 a79595a <=( (not A167)  and  a79594a );
 a79598a <=( (not A202)  and  A200 );
 a79601a <=( A265  and  A203 );
 a79602a <=( a79601a  and  a79598a );
 a79603a <=( a79602a  and  a79595a );
 a79607a <=( A269  and  (not A267) );
 a79608a <=( A266  and  a79607a );
 a79611a <=( (not A299)  and  A298 );
 a79614a <=( A302  and  (not A301) );
 a79615a <=( a79614a  and  a79611a );
 a79616a <=( a79615a  and  a79608a );
 a79620a <=( (not A199)  and  (not A166) );
 a79621a <=( (not A167)  and  a79620a );
 a79624a <=( (not A202)  and  A200 );
 a79627a <=( A265  and  A203 );
 a79628a <=( a79627a  and  a79624a );
 a79629a <=( a79628a  and  a79621a );
 a79633a <=( A269  and  (not A267) );
 a79634a <=( A266  and  a79633a );
 a79637a <=( A299  and  (not A298) );
 a79640a <=( A302  and  (not A301) );
 a79641a <=( a79640a  and  a79637a );
 a79642a <=( a79641a  and  a79634a );
 a79646a <=( (not A199)  and  (not A166) );
 a79647a <=( (not A167)  and  a79646a );
 a79650a <=( (not A202)  and  A200 );
 a79653a <=( A265  and  A203 );
 a79654a <=( a79653a  and  a79650a );
 a79655a <=( a79654a  and  a79647a );
 a79659a <=( A269  and  (not A267) );
 a79660a <=( A266  and  a79659a );
 a79663a <=( (not A299)  and  (not A298) );
 a79666a <=( (not A302)  and  A301 );
 a79667a <=( a79666a  and  a79663a );
 a79668a <=( a79667a  and  a79660a );
 a79672a <=( (not A199)  and  (not A166) );
 a79673a <=( (not A167)  and  a79672a );
 a79676a <=( (not A202)  and  A200 );
 a79679a <=( (not A265)  and  A203 );
 a79680a <=( a79679a  and  a79676a );
 a79681a <=( a79680a  and  a79673a );
 a79685a <=( A268  and  (not A267) );
 a79686a <=( A266  and  a79685a );
 a79689a <=( A299  and  A298 );
 a79692a <=( (not A302)  and  A301 );
 a79693a <=( a79692a  and  a79689a );
 a79694a <=( a79693a  and  a79686a );
 a79698a <=( (not A199)  and  (not A166) );
 a79699a <=( (not A167)  and  a79698a );
 a79702a <=( (not A202)  and  A200 );
 a79705a <=( (not A265)  and  A203 );
 a79706a <=( a79705a  and  a79702a );
 a79707a <=( a79706a  and  a79699a );
 a79711a <=( A268  and  (not A267) );
 a79712a <=( A266  and  a79711a );
 a79715a <=( (not A299)  and  A298 );
 a79718a <=( A302  and  (not A301) );
 a79719a <=( a79718a  and  a79715a );
 a79720a <=( a79719a  and  a79712a );
 a79724a <=( (not A199)  and  (not A166) );
 a79725a <=( (not A167)  and  a79724a );
 a79728a <=( (not A202)  and  A200 );
 a79731a <=( (not A265)  and  A203 );
 a79732a <=( a79731a  and  a79728a );
 a79733a <=( a79732a  and  a79725a );
 a79737a <=( A268  and  (not A267) );
 a79738a <=( A266  and  a79737a );
 a79741a <=( A299  and  (not A298) );
 a79744a <=( A302  and  (not A301) );
 a79745a <=( a79744a  and  a79741a );
 a79746a <=( a79745a  and  a79738a );
 a79750a <=( (not A199)  and  (not A166) );
 a79751a <=( (not A167)  and  a79750a );
 a79754a <=( (not A202)  and  A200 );
 a79757a <=( (not A265)  and  A203 );
 a79758a <=( a79757a  and  a79754a );
 a79759a <=( a79758a  and  a79751a );
 a79763a <=( A268  and  (not A267) );
 a79764a <=( A266  and  a79763a );
 a79767a <=( (not A299)  and  (not A298) );
 a79770a <=( (not A302)  and  A301 );
 a79771a <=( a79770a  and  a79767a );
 a79772a <=( a79771a  and  a79764a );
 a79776a <=( (not A199)  and  (not A166) );
 a79777a <=( (not A167)  and  a79776a );
 a79780a <=( (not A202)  and  A200 );
 a79783a <=( (not A265)  and  A203 );
 a79784a <=( a79783a  and  a79780a );
 a79785a <=( a79784a  and  a79777a );
 a79789a <=( (not A269)  and  (not A267) );
 a79790a <=( A266  and  a79789a );
 a79793a <=( A299  and  A298 );
 a79796a <=( (not A302)  and  A301 );
 a79797a <=( a79796a  and  a79793a );
 a79798a <=( a79797a  and  a79790a );
 a79802a <=( (not A199)  and  (not A166) );
 a79803a <=( (not A167)  and  a79802a );
 a79806a <=( (not A202)  and  A200 );
 a79809a <=( (not A265)  and  A203 );
 a79810a <=( a79809a  and  a79806a );
 a79811a <=( a79810a  and  a79803a );
 a79815a <=( (not A269)  and  (not A267) );
 a79816a <=( A266  and  a79815a );
 a79819a <=( (not A299)  and  A298 );
 a79822a <=( A302  and  (not A301) );
 a79823a <=( a79822a  and  a79819a );
 a79824a <=( a79823a  and  a79816a );
 a79828a <=( (not A199)  and  (not A166) );
 a79829a <=( (not A167)  and  a79828a );
 a79832a <=( (not A202)  and  A200 );
 a79835a <=( (not A265)  and  A203 );
 a79836a <=( a79835a  and  a79832a );
 a79837a <=( a79836a  and  a79829a );
 a79841a <=( (not A269)  and  (not A267) );
 a79842a <=( A266  and  a79841a );
 a79845a <=( A299  and  (not A298) );
 a79848a <=( A302  and  (not A301) );
 a79849a <=( a79848a  and  a79845a );
 a79850a <=( a79849a  and  a79842a );
 a79854a <=( (not A199)  and  (not A166) );
 a79855a <=( (not A167)  and  a79854a );
 a79858a <=( (not A202)  and  A200 );
 a79861a <=( (not A265)  and  A203 );
 a79862a <=( a79861a  and  a79858a );
 a79863a <=( a79862a  and  a79855a );
 a79867a <=( (not A269)  and  (not A267) );
 a79868a <=( A266  and  a79867a );
 a79871a <=( (not A299)  and  (not A298) );
 a79874a <=( (not A302)  and  A301 );
 a79875a <=( a79874a  and  a79871a );
 a79876a <=( a79875a  and  a79868a );
 a79880a <=( (not A199)  and  (not A166) );
 a79881a <=( (not A167)  and  a79880a );
 a79884a <=( (not A202)  and  A200 );
 a79887a <=( A265  and  A203 );
 a79888a <=( a79887a  and  a79884a );
 a79889a <=( a79888a  and  a79881a );
 a79893a <=( A268  and  (not A267) );
 a79894a <=( (not A266)  and  a79893a );
 a79897a <=( A299  and  A298 );
 a79900a <=( (not A302)  and  A301 );
 a79901a <=( a79900a  and  a79897a );
 a79902a <=( a79901a  and  a79894a );
 a79906a <=( (not A199)  and  (not A166) );
 a79907a <=( (not A167)  and  a79906a );
 a79910a <=( (not A202)  and  A200 );
 a79913a <=( A265  and  A203 );
 a79914a <=( a79913a  and  a79910a );
 a79915a <=( a79914a  and  a79907a );
 a79919a <=( A268  and  (not A267) );
 a79920a <=( (not A266)  and  a79919a );
 a79923a <=( (not A299)  and  A298 );
 a79926a <=( A302  and  (not A301) );
 a79927a <=( a79926a  and  a79923a );
 a79928a <=( a79927a  and  a79920a );
 a79932a <=( (not A199)  and  (not A166) );
 a79933a <=( (not A167)  and  a79932a );
 a79936a <=( (not A202)  and  A200 );
 a79939a <=( A265  and  A203 );
 a79940a <=( a79939a  and  a79936a );
 a79941a <=( a79940a  and  a79933a );
 a79945a <=( A268  and  (not A267) );
 a79946a <=( (not A266)  and  a79945a );
 a79949a <=( A299  and  (not A298) );
 a79952a <=( A302  and  (not A301) );
 a79953a <=( a79952a  and  a79949a );
 a79954a <=( a79953a  and  a79946a );
 a79958a <=( (not A199)  and  (not A166) );
 a79959a <=( (not A167)  and  a79958a );
 a79962a <=( (not A202)  and  A200 );
 a79965a <=( A265  and  A203 );
 a79966a <=( a79965a  and  a79962a );
 a79967a <=( a79966a  and  a79959a );
 a79971a <=( A268  and  (not A267) );
 a79972a <=( (not A266)  and  a79971a );
 a79975a <=( (not A299)  and  (not A298) );
 a79978a <=( (not A302)  and  A301 );
 a79979a <=( a79978a  and  a79975a );
 a79980a <=( a79979a  and  a79972a );
 a79984a <=( (not A199)  and  (not A166) );
 a79985a <=( (not A167)  and  a79984a );
 a79988a <=( (not A202)  and  A200 );
 a79991a <=( A265  and  A203 );
 a79992a <=( a79991a  and  a79988a );
 a79993a <=( a79992a  and  a79985a );
 a79997a <=( (not A269)  and  (not A267) );
 a79998a <=( (not A266)  and  a79997a );
 a80001a <=( A299  and  A298 );
 a80004a <=( (not A302)  and  A301 );
 a80005a <=( a80004a  and  a80001a );
 a80006a <=( a80005a  and  a79998a );
 a80010a <=( (not A199)  and  (not A166) );
 a80011a <=( (not A167)  and  a80010a );
 a80014a <=( (not A202)  and  A200 );
 a80017a <=( A265  and  A203 );
 a80018a <=( a80017a  and  a80014a );
 a80019a <=( a80018a  and  a80011a );
 a80023a <=( (not A269)  and  (not A267) );
 a80024a <=( (not A266)  and  a80023a );
 a80027a <=( (not A299)  and  A298 );
 a80030a <=( A302  and  (not A301) );
 a80031a <=( a80030a  and  a80027a );
 a80032a <=( a80031a  and  a80024a );
 a80036a <=( (not A199)  and  (not A166) );
 a80037a <=( (not A167)  and  a80036a );
 a80040a <=( (not A202)  and  A200 );
 a80043a <=( A265  and  A203 );
 a80044a <=( a80043a  and  a80040a );
 a80045a <=( a80044a  and  a80037a );
 a80049a <=( (not A269)  and  (not A267) );
 a80050a <=( (not A266)  and  a80049a );
 a80053a <=( A299  and  (not A298) );
 a80056a <=( A302  and  (not A301) );
 a80057a <=( a80056a  and  a80053a );
 a80058a <=( a80057a  and  a80050a );
 a80062a <=( (not A199)  and  (not A166) );
 a80063a <=( (not A167)  and  a80062a );
 a80066a <=( (not A202)  and  A200 );
 a80069a <=( A265  and  A203 );
 a80070a <=( a80069a  and  a80066a );
 a80071a <=( a80070a  and  a80063a );
 a80075a <=( (not A269)  and  (not A267) );
 a80076a <=( (not A266)  and  a80075a );
 a80079a <=( (not A299)  and  (not A298) );
 a80082a <=( (not A302)  and  A301 );
 a80083a <=( a80082a  and  a80079a );
 a80084a <=( a80083a  and  a80076a );
 a80088a <=( (not A199)  and  (not A166) );
 a80089a <=( (not A167)  and  a80088a );
 a80092a <=( (not A201)  and  A200 );
 a80095a <=( A265  and  A202 );
 a80096a <=( a80095a  and  a80092a );
 a80097a <=( a80096a  and  a80089a );
 a80101a <=( (not A269)  and  A268 );
 a80102a <=( A266  and  a80101a );
 a80105a <=( A299  and  A298 );
 a80108a <=( (not A301)  and  (not A300) );
 a80109a <=( a80108a  and  a80105a );
 a80110a <=( a80109a  and  a80102a );
 a80114a <=( (not A199)  and  (not A166) );
 a80115a <=( (not A167)  and  a80114a );
 a80118a <=( (not A201)  and  A200 );
 a80121a <=( A265  and  A202 );
 a80122a <=( a80121a  and  a80118a );
 a80123a <=( a80122a  and  a80115a );
 a80127a <=( (not A269)  and  A268 );
 a80128a <=( A266  and  a80127a );
 a80131a <=( A299  and  A298 );
 a80134a <=( A302  and  (not A300) );
 a80135a <=( a80134a  and  a80131a );
 a80136a <=( a80135a  and  a80128a );
 a80140a <=( (not A199)  and  (not A166) );
 a80141a <=( (not A167)  and  a80140a );
 a80144a <=( (not A201)  and  A200 );
 a80147a <=( A265  and  A202 );
 a80148a <=( a80147a  and  a80144a );
 a80149a <=( a80148a  and  a80141a );
 a80153a <=( (not A269)  and  A268 );
 a80154a <=( A266  and  a80153a );
 a80157a <=( (not A299)  and  A298 );
 a80160a <=( A301  and  (not A300) );
 a80161a <=( a80160a  and  a80157a );
 a80162a <=( a80161a  and  a80154a );
 a80166a <=( (not A199)  and  (not A166) );
 a80167a <=( (not A167)  and  a80166a );
 a80170a <=( (not A201)  and  A200 );
 a80173a <=( A265  and  A202 );
 a80174a <=( a80173a  and  a80170a );
 a80175a <=( a80174a  and  a80167a );
 a80179a <=( (not A269)  and  A268 );
 a80180a <=( A266  and  a80179a );
 a80183a <=( (not A299)  and  A298 );
 a80186a <=( (not A302)  and  (not A300) );
 a80187a <=( a80186a  and  a80183a );
 a80188a <=( a80187a  and  a80180a );
 a80192a <=( (not A199)  and  (not A166) );
 a80193a <=( (not A167)  and  a80192a );
 a80196a <=( (not A201)  and  A200 );
 a80199a <=( A265  and  A202 );
 a80200a <=( a80199a  and  a80196a );
 a80201a <=( a80200a  and  a80193a );
 a80205a <=( (not A269)  and  A268 );
 a80206a <=( A266  and  a80205a );
 a80209a <=( A299  and  (not A298) );
 a80212a <=( A301  and  (not A300) );
 a80213a <=( a80212a  and  a80209a );
 a80214a <=( a80213a  and  a80206a );
 a80218a <=( (not A199)  and  (not A166) );
 a80219a <=( (not A167)  and  a80218a );
 a80222a <=( (not A201)  and  A200 );
 a80225a <=( A265  and  A202 );
 a80226a <=( a80225a  and  a80222a );
 a80227a <=( a80226a  and  a80219a );
 a80231a <=( (not A269)  and  A268 );
 a80232a <=( A266  and  a80231a );
 a80235a <=( A299  and  (not A298) );
 a80238a <=( (not A302)  and  (not A300) );
 a80239a <=( a80238a  and  a80235a );
 a80240a <=( a80239a  and  a80232a );
 a80244a <=( (not A199)  and  (not A166) );
 a80245a <=( (not A167)  and  a80244a );
 a80248a <=( (not A201)  and  A200 );
 a80251a <=( (not A265)  and  A202 );
 a80252a <=( a80251a  and  a80248a );
 a80253a <=( a80252a  and  a80245a );
 a80257a <=( A269  and  (not A268) );
 a80258a <=( A266  and  a80257a );
 a80261a <=( A299  and  A298 );
 a80264a <=( (not A301)  and  (not A300) );
 a80265a <=( a80264a  and  a80261a );
 a80266a <=( a80265a  and  a80258a );
 a80270a <=( (not A199)  and  (not A166) );
 a80271a <=( (not A167)  and  a80270a );
 a80274a <=( (not A201)  and  A200 );
 a80277a <=( (not A265)  and  A202 );
 a80278a <=( a80277a  and  a80274a );
 a80279a <=( a80278a  and  a80271a );
 a80283a <=( A269  and  (not A268) );
 a80284a <=( A266  and  a80283a );
 a80287a <=( A299  and  A298 );
 a80290a <=( A302  and  (not A300) );
 a80291a <=( a80290a  and  a80287a );
 a80292a <=( a80291a  and  a80284a );
 a80296a <=( (not A199)  and  (not A166) );
 a80297a <=( (not A167)  and  a80296a );
 a80300a <=( (not A201)  and  A200 );
 a80303a <=( (not A265)  and  A202 );
 a80304a <=( a80303a  and  a80300a );
 a80305a <=( a80304a  and  a80297a );
 a80309a <=( A269  and  (not A268) );
 a80310a <=( A266  and  a80309a );
 a80313a <=( (not A299)  and  A298 );
 a80316a <=( A301  and  (not A300) );
 a80317a <=( a80316a  and  a80313a );
 a80318a <=( a80317a  and  a80310a );
 a80322a <=( (not A199)  and  (not A166) );
 a80323a <=( (not A167)  and  a80322a );
 a80326a <=( (not A201)  and  A200 );
 a80329a <=( (not A265)  and  A202 );
 a80330a <=( a80329a  and  a80326a );
 a80331a <=( a80330a  and  a80323a );
 a80335a <=( A269  and  (not A268) );
 a80336a <=( A266  and  a80335a );
 a80339a <=( (not A299)  and  A298 );
 a80342a <=( (not A302)  and  (not A300) );
 a80343a <=( a80342a  and  a80339a );
 a80344a <=( a80343a  and  a80336a );
 a80348a <=( (not A199)  and  (not A166) );
 a80349a <=( (not A167)  and  a80348a );
 a80352a <=( (not A201)  and  A200 );
 a80355a <=( (not A265)  and  A202 );
 a80356a <=( a80355a  and  a80352a );
 a80357a <=( a80356a  and  a80349a );
 a80361a <=( A269  and  (not A268) );
 a80362a <=( A266  and  a80361a );
 a80365a <=( A299  and  (not A298) );
 a80368a <=( A301  and  (not A300) );
 a80369a <=( a80368a  and  a80365a );
 a80370a <=( a80369a  and  a80362a );
 a80374a <=( (not A199)  and  (not A166) );
 a80375a <=( (not A167)  and  a80374a );
 a80378a <=( (not A201)  and  A200 );
 a80381a <=( (not A265)  and  A202 );
 a80382a <=( a80381a  and  a80378a );
 a80383a <=( a80382a  and  a80375a );
 a80387a <=( A269  and  (not A268) );
 a80388a <=( A266  and  a80387a );
 a80391a <=( A299  and  (not A298) );
 a80394a <=( (not A302)  and  (not A300) );
 a80395a <=( a80394a  and  a80391a );
 a80396a <=( a80395a  and  a80388a );
 a80400a <=( (not A199)  and  (not A166) );
 a80401a <=( (not A167)  and  a80400a );
 a80404a <=( (not A201)  and  A200 );
 a80407a <=( A265  and  A202 );
 a80408a <=( a80407a  and  a80404a );
 a80409a <=( a80408a  and  a80401a );
 a80413a <=( A269  and  (not A268) );
 a80414a <=( (not A266)  and  a80413a );
 a80417a <=( A299  and  A298 );
 a80420a <=( (not A301)  and  (not A300) );
 a80421a <=( a80420a  and  a80417a );
 a80422a <=( a80421a  and  a80414a );
 a80426a <=( (not A199)  and  (not A166) );
 a80427a <=( (not A167)  and  a80426a );
 a80430a <=( (not A201)  and  A200 );
 a80433a <=( A265  and  A202 );
 a80434a <=( a80433a  and  a80430a );
 a80435a <=( a80434a  and  a80427a );
 a80439a <=( A269  and  (not A268) );
 a80440a <=( (not A266)  and  a80439a );
 a80443a <=( A299  and  A298 );
 a80446a <=( A302  and  (not A300) );
 a80447a <=( a80446a  and  a80443a );
 a80448a <=( a80447a  and  a80440a );
 a80452a <=( (not A199)  and  (not A166) );
 a80453a <=( (not A167)  and  a80452a );
 a80456a <=( (not A201)  and  A200 );
 a80459a <=( A265  and  A202 );
 a80460a <=( a80459a  and  a80456a );
 a80461a <=( a80460a  and  a80453a );
 a80465a <=( A269  and  (not A268) );
 a80466a <=( (not A266)  and  a80465a );
 a80469a <=( (not A299)  and  A298 );
 a80472a <=( A301  and  (not A300) );
 a80473a <=( a80472a  and  a80469a );
 a80474a <=( a80473a  and  a80466a );
 a80478a <=( (not A199)  and  (not A166) );
 a80479a <=( (not A167)  and  a80478a );
 a80482a <=( (not A201)  and  A200 );
 a80485a <=( A265  and  A202 );
 a80486a <=( a80485a  and  a80482a );
 a80487a <=( a80486a  and  a80479a );
 a80491a <=( A269  and  (not A268) );
 a80492a <=( (not A266)  and  a80491a );
 a80495a <=( (not A299)  and  A298 );
 a80498a <=( (not A302)  and  (not A300) );
 a80499a <=( a80498a  and  a80495a );
 a80500a <=( a80499a  and  a80492a );
 a80504a <=( (not A199)  and  (not A166) );
 a80505a <=( (not A167)  and  a80504a );
 a80508a <=( (not A201)  and  A200 );
 a80511a <=( A265  and  A202 );
 a80512a <=( a80511a  and  a80508a );
 a80513a <=( a80512a  and  a80505a );
 a80517a <=( A269  and  (not A268) );
 a80518a <=( (not A266)  and  a80517a );
 a80521a <=( A299  and  (not A298) );
 a80524a <=( A301  and  (not A300) );
 a80525a <=( a80524a  and  a80521a );
 a80526a <=( a80525a  and  a80518a );
 a80530a <=( (not A199)  and  (not A166) );
 a80531a <=( (not A167)  and  a80530a );
 a80534a <=( (not A201)  and  A200 );
 a80537a <=( A265  and  A202 );
 a80538a <=( a80537a  and  a80534a );
 a80539a <=( a80538a  and  a80531a );
 a80543a <=( A269  and  (not A268) );
 a80544a <=( (not A266)  and  a80543a );
 a80547a <=( A299  and  (not A298) );
 a80550a <=( (not A302)  and  (not A300) );
 a80551a <=( a80550a  and  a80547a );
 a80552a <=( a80551a  and  a80544a );
 a80556a <=( (not A199)  and  (not A166) );
 a80557a <=( (not A167)  and  a80556a );
 a80560a <=( (not A201)  and  A200 );
 a80563a <=( (not A265)  and  A202 );
 a80564a <=( a80563a  and  a80560a );
 a80565a <=( a80564a  and  a80557a );
 a80569a <=( (not A269)  and  A268 );
 a80570a <=( (not A266)  and  a80569a );
 a80573a <=( A299  and  A298 );
 a80576a <=( (not A301)  and  (not A300) );
 a80577a <=( a80576a  and  a80573a );
 a80578a <=( a80577a  and  a80570a );
 a80582a <=( (not A199)  and  (not A166) );
 a80583a <=( (not A167)  and  a80582a );
 a80586a <=( (not A201)  and  A200 );
 a80589a <=( (not A265)  and  A202 );
 a80590a <=( a80589a  and  a80586a );
 a80591a <=( a80590a  and  a80583a );
 a80595a <=( (not A269)  and  A268 );
 a80596a <=( (not A266)  and  a80595a );
 a80599a <=( A299  and  A298 );
 a80602a <=( A302  and  (not A300) );
 a80603a <=( a80602a  and  a80599a );
 a80604a <=( a80603a  and  a80596a );
 a80608a <=( (not A199)  and  (not A166) );
 a80609a <=( (not A167)  and  a80608a );
 a80612a <=( (not A201)  and  A200 );
 a80615a <=( (not A265)  and  A202 );
 a80616a <=( a80615a  and  a80612a );
 a80617a <=( a80616a  and  a80609a );
 a80621a <=( (not A269)  and  A268 );
 a80622a <=( (not A266)  and  a80621a );
 a80625a <=( (not A299)  and  A298 );
 a80628a <=( A301  and  (not A300) );
 a80629a <=( a80628a  and  a80625a );
 a80630a <=( a80629a  and  a80622a );
 a80634a <=( (not A199)  and  (not A166) );
 a80635a <=( (not A167)  and  a80634a );
 a80638a <=( (not A201)  and  A200 );
 a80641a <=( (not A265)  and  A202 );
 a80642a <=( a80641a  and  a80638a );
 a80643a <=( a80642a  and  a80635a );
 a80647a <=( (not A269)  and  A268 );
 a80648a <=( (not A266)  and  a80647a );
 a80651a <=( (not A299)  and  A298 );
 a80654a <=( (not A302)  and  (not A300) );
 a80655a <=( a80654a  and  a80651a );
 a80656a <=( a80655a  and  a80648a );
 a80660a <=( (not A199)  and  (not A166) );
 a80661a <=( (not A167)  and  a80660a );
 a80664a <=( (not A201)  and  A200 );
 a80667a <=( (not A265)  and  A202 );
 a80668a <=( a80667a  and  a80664a );
 a80669a <=( a80668a  and  a80661a );
 a80673a <=( (not A269)  and  A268 );
 a80674a <=( (not A266)  and  a80673a );
 a80677a <=( A299  and  (not A298) );
 a80680a <=( A301  and  (not A300) );
 a80681a <=( a80680a  and  a80677a );
 a80682a <=( a80681a  and  a80674a );
 a80686a <=( (not A199)  and  (not A166) );
 a80687a <=( (not A167)  and  a80686a );
 a80690a <=( (not A201)  and  A200 );
 a80693a <=( (not A265)  and  A202 );
 a80694a <=( a80693a  and  a80690a );
 a80695a <=( a80694a  and  a80687a );
 a80699a <=( (not A269)  and  A268 );
 a80700a <=( (not A266)  and  a80699a );
 a80703a <=( A299  and  (not A298) );
 a80706a <=( (not A302)  and  (not A300) );
 a80707a <=( a80706a  and  a80703a );
 a80708a <=( a80707a  and  a80700a );
 a80712a <=( (not A199)  and  (not A166) );
 a80713a <=( (not A167)  and  a80712a );
 a80716a <=( (not A201)  and  A200 );
 a80719a <=( A265  and  (not A203) );
 a80720a <=( a80719a  and  a80716a );
 a80721a <=( a80720a  and  a80713a );
 a80725a <=( (not A269)  and  A268 );
 a80726a <=( A266  and  a80725a );
 a80729a <=( A299  and  A298 );
 a80732a <=( (not A301)  and  (not A300) );
 a80733a <=( a80732a  and  a80729a );
 a80734a <=( a80733a  and  a80726a );
 a80738a <=( (not A199)  and  (not A166) );
 a80739a <=( (not A167)  and  a80738a );
 a80742a <=( (not A201)  and  A200 );
 a80745a <=( A265  and  (not A203) );
 a80746a <=( a80745a  and  a80742a );
 a80747a <=( a80746a  and  a80739a );
 a80751a <=( (not A269)  and  A268 );
 a80752a <=( A266  and  a80751a );
 a80755a <=( A299  and  A298 );
 a80758a <=( A302  and  (not A300) );
 a80759a <=( a80758a  and  a80755a );
 a80760a <=( a80759a  and  a80752a );
 a80764a <=( (not A199)  and  (not A166) );
 a80765a <=( (not A167)  and  a80764a );
 a80768a <=( (not A201)  and  A200 );
 a80771a <=( A265  and  (not A203) );
 a80772a <=( a80771a  and  a80768a );
 a80773a <=( a80772a  and  a80765a );
 a80777a <=( (not A269)  and  A268 );
 a80778a <=( A266  and  a80777a );
 a80781a <=( (not A299)  and  A298 );
 a80784a <=( A301  and  (not A300) );
 a80785a <=( a80784a  and  a80781a );
 a80786a <=( a80785a  and  a80778a );
 a80790a <=( (not A199)  and  (not A166) );
 a80791a <=( (not A167)  and  a80790a );
 a80794a <=( (not A201)  and  A200 );
 a80797a <=( A265  and  (not A203) );
 a80798a <=( a80797a  and  a80794a );
 a80799a <=( a80798a  and  a80791a );
 a80803a <=( (not A269)  and  A268 );
 a80804a <=( A266  and  a80803a );
 a80807a <=( (not A299)  and  A298 );
 a80810a <=( (not A302)  and  (not A300) );
 a80811a <=( a80810a  and  a80807a );
 a80812a <=( a80811a  and  a80804a );
 a80816a <=( (not A199)  and  (not A166) );
 a80817a <=( (not A167)  and  a80816a );
 a80820a <=( (not A201)  and  A200 );
 a80823a <=( A265  and  (not A203) );
 a80824a <=( a80823a  and  a80820a );
 a80825a <=( a80824a  and  a80817a );
 a80829a <=( (not A269)  and  A268 );
 a80830a <=( A266  and  a80829a );
 a80833a <=( A299  and  (not A298) );
 a80836a <=( A301  and  (not A300) );
 a80837a <=( a80836a  and  a80833a );
 a80838a <=( a80837a  and  a80830a );
 a80842a <=( (not A199)  and  (not A166) );
 a80843a <=( (not A167)  and  a80842a );
 a80846a <=( (not A201)  and  A200 );
 a80849a <=( A265  and  (not A203) );
 a80850a <=( a80849a  and  a80846a );
 a80851a <=( a80850a  and  a80843a );
 a80855a <=( (not A269)  and  A268 );
 a80856a <=( A266  and  a80855a );
 a80859a <=( A299  and  (not A298) );
 a80862a <=( (not A302)  and  (not A300) );
 a80863a <=( a80862a  and  a80859a );
 a80864a <=( a80863a  and  a80856a );
 a80868a <=( (not A199)  and  (not A166) );
 a80869a <=( (not A167)  and  a80868a );
 a80872a <=( (not A201)  and  A200 );
 a80875a <=( (not A265)  and  (not A203) );
 a80876a <=( a80875a  and  a80872a );
 a80877a <=( a80876a  and  a80869a );
 a80881a <=( A269  and  (not A268) );
 a80882a <=( A266  and  a80881a );
 a80885a <=( A299  and  A298 );
 a80888a <=( (not A301)  and  (not A300) );
 a80889a <=( a80888a  and  a80885a );
 a80890a <=( a80889a  and  a80882a );
 a80894a <=( (not A199)  and  (not A166) );
 a80895a <=( (not A167)  and  a80894a );
 a80898a <=( (not A201)  and  A200 );
 a80901a <=( (not A265)  and  (not A203) );
 a80902a <=( a80901a  and  a80898a );
 a80903a <=( a80902a  and  a80895a );
 a80907a <=( A269  and  (not A268) );
 a80908a <=( A266  and  a80907a );
 a80911a <=( A299  and  A298 );
 a80914a <=( A302  and  (not A300) );
 a80915a <=( a80914a  and  a80911a );
 a80916a <=( a80915a  and  a80908a );
 a80920a <=( (not A199)  and  (not A166) );
 a80921a <=( (not A167)  and  a80920a );
 a80924a <=( (not A201)  and  A200 );
 a80927a <=( (not A265)  and  (not A203) );
 a80928a <=( a80927a  and  a80924a );
 a80929a <=( a80928a  and  a80921a );
 a80933a <=( A269  and  (not A268) );
 a80934a <=( A266  and  a80933a );
 a80937a <=( (not A299)  and  A298 );
 a80940a <=( A301  and  (not A300) );
 a80941a <=( a80940a  and  a80937a );
 a80942a <=( a80941a  and  a80934a );
 a80946a <=( (not A199)  and  (not A166) );
 a80947a <=( (not A167)  and  a80946a );
 a80950a <=( (not A201)  and  A200 );
 a80953a <=( (not A265)  and  (not A203) );
 a80954a <=( a80953a  and  a80950a );
 a80955a <=( a80954a  and  a80947a );
 a80959a <=( A269  and  (not A268) );
 a80960a <=( A266  and  a80959a );
 a80963a <=( (not A299)  and  A298 );
 a80966a <=( (not A302)  and  (not A300) );
 a80967a <=( a80966a  and  a80963a );
 a80968a <=( a80967a  and  a80960a );
 a80972a <=( (not A199)  and  (not A166) );
 a80973a <=( (not A167)  and  a80972a );
 a80976a <=( (not A201)  and  A200 );
 a80979a <=( (not A265)  and  (not A203) );
 a80980a <=( a80979a  and  a80976a );
 a80981a <=( a80980a  and  a80973a );
 a80985a <=( A269  and  (not A268) );
 a80986a <=( A266  and  a80985a );
 a80989a <=( A299  and  (not A298) );
 a80992a <=( A301  and  (not A300) );
 a80993a <=( a80992a  and  a80989a );
 a80994a <=( a80993a  and  a80986a );
 a80998a <=( (not A199)  and  (not A166) );
 a80999a <=( (not A167)  and  a80998a );
 a81002a <=( (not A201)  and  A200 );
 a81005a <=( (not A265)  and  (not A203) );
 a81006a <=( a81005a  and  a81002a );
 a81007a <=( a81006a  and  a80999a );
 a81011a <=( A269  and  (not A268) );
 a81012a <=( A266  and  a81011a );
 a81015a <=( A299  and  (not A298) );
 a81018a <=( (not A302)  and  (not A300) );
 a81019a <=( a81018a  and  a81015a );
 a81020a <=( a81019a  and  a81012a );
 a81024a <=( (not A199)  and  (not A166) );
 a81025a <=( (not A167)  and  a81024a );
 a81028a <=( (not A201)  and  A200 );
 a81031a <=( A265  and  (not A203) );
 a81032a <=( a81031a  and  a81028a );
 a81033a <=( a81032a  and  a81025a );
 a81037a <=( A269  and  (not A268) );
 a81038a <=( (not A266)  and  a81037a );
 a81041a <=( A299  and  A298 );
 a81044a <=( (not A301)  and  (not A300) );
 a81045a <=( a81044a  and  a81041a );
 a81046a <=( a81045a  and  a81038a );
 a81050a <=( (not A199)  and  (not A166) );
 a81051a <=( (not A167)  and  a81050a );
 a81054a <=( (not A201)  and  A200 );
 a81057a <=( A265  and  (not A203) );
 a81058a <=( a81057a  and  a81054a );
 a81059a <=( a81058a  and  a81051a );
 a81063a <=( A269  and  (not A268) );
 a81064a <=( (not A266)  and  a81063a );
 a81067a <=( A299  and  A298 );
 a81070a <=( A302  and  (not A300) );
 a81071a <=( a81070a  and  a81067a );
 a81072a <=( a81071a  and  a81064a );
 a81076a <=( (not A199)  and  (not A166) );
 a81077a <=( (not A167)  and  a81076a );
 a81080a <=( (not A201)  and  A200 );
 a81083a <=( A265  and  (not A203) );
 a81084a <=( a81083a  and  a81080a );
 a81085a <=( a81084a  and  a81077a );
 a81089a <=( A269  and  (not A268) );
 a81090a <=( (not A266)  and  a81089a );
 a81093a <=( (not A299)  and  A298 );
 a81096a <=( A301  and  (not A300) );
 a81097a <=( a81096a  and  a81093a );
 a81098a <=( a81097a  and  a81090a );
 a81102a <=( (not A199)  and  (not A166) );
 a81103a <=( (not A167)  and  a81102a );
 a81106a <=( (not A201)  and  A200 );
 a81109a <=( A265  and  (not A203) );
 a81110a <=( a81109a  and  a81106a );
 a81111a <=( a81110a  and  a81103a );
 a81115a <=( A269  and  (not A268) );
 a81116a <=( (not A266)  and  a81115a );
 a81119a <=( (not A299)  and  A298 );
 a81122a <=( (not A302)  and  (not A300) );
 a81123a <=( a81122a  and  a81119a );
 a81124a <=( a81123a  and  a81116a );
 a81128a <=( (not A199)  and  (not A166) );
 a81129a <=( (not A167)  and  a81128a );
 a81132a <=( (not A201)  and  A200 );
 a81135a <=( A265  and  (not A203) );
 a81136a <=( a81135a  and  a81132a );
 a81137a <=( a81136a  and  a81129a );
 a81141a <=( A269  and  (not A268) );
 a81142a <=( (not A266)  and  a81141a );
 a81145a <=( A299  and  (not A298) );
 a81148a <=( A301  and  (not A300) );
 a81149a <=( a81148a  and  a81145a );
 a81150a <=( a81149a  and  a81142a );
 a81154a <=( (not A199)  and  (not A166) );
 a81155a <=( (not A167)  and  a81154a );
 a81158a <=( (not A201)  and  A200 );
 a81161a <=( A265  and  (not A203) );
 a81162a <=( a81161a  and  a81158a );
 a81163a <=( a81162a  and  a81155a );
 a81167a <=( A269  and  (not A268) );
 a81168a <=( (not A266)  and  a81167a );
 a81171a <=( A299  and  (not A298) );
 a81174a <=( (not A302)  and  (not A300) );
 a81175a <=( a81174a  and  a81171a );
 a81176a <=( a81175a  and  a81168a );
 a81180a <=( (not A199)  and  (not A166) );
 a81181a <=( (not A167)  and  a81180a );
 a81184a <=( (not A201)  and  A200 );
 a81187a <=( (not A265)  and  (not A203) );
 a81188a <=( a81187a  and  a81184a );
 a81189a <=( a81188a  and  a81181a );
 a81193a <=( (not A269)  and  A268 );
 a81194a <=( (not A266)  and  a81193a );
 a81197a <=( A299  and  A298 );
 a81200a <=( (not A301)  and  (not A300) );
 a81201a <=( a81200a  and  a81197a );
 a81202a <=( a81201a  and  a81194a );
 a81206a <=( (not A199)  and  (not A166) );
 a81207a <=( (not A167)  and  a81206a );
 a81210a <=( (not A201)  and  A200 );
 a81213a <=( (not A265)  and  (not A203) );
 a81214a <=( a81213a  and  a81210a );
 a81215a <=( a81214a  and  a81207a );
 a81219a <=( (not A269)  and  A268 );
 a81220a <=( (not A266)  and  a81219a );
 a81223a <=( A299  and  A298 );
 a81226a <=( A302  and  (not A300) );
 a81227a <=( a81226a  and  a81223a );
 a81228a <=( a81227a  and  a81220a );
 a81232a <=( (not A199)  and  (not A166) );
 a81233a <=( (not A167)  and  a81232a );
 a81236a <=( (not A201)  and  A200 );
 a81239a <=( (not A265)  and  (not A203) );
 a81240a <=( a81239a  and  a81236a );
 a81241a <=( a81240a  and  a81233a );
 a81245a <=( (not A269)  and  A268 );
 a81246a <=( (not A266)  and  a81245a );
 a81249a <=( (not A299)  and  A298 );
 a81252a <=( A301  and  (not A300) );
 a81253a <=( a81252a  and  a81249a );
 a81254a <=( a81253a  and  a81246a );
 a81258a <=( (not A199)  and  (not A166) );
 a81259a <=( (not A167)  and  a81258a );
 a81262a <=( (not A201)  and  A200 );
 a81265a <=( (not A265)  and  (not A203) );
 a81266a <=( a81265a  and  a81262a );
 a81267a <=( a81266a  and  a81259a );
 a81271a <=( (not A269)  and  A268 );
 a81272a <=( (not A266)  and  a81271a );
 a81275a <=( (not A299)  and  A298 );
 a81278a <=( (not A302)  and  (not A300) );
 a81279a <=( a81278a  and  a81275a );
 a81280a <=( a81279a  and  a81272a );
 a81284a <=( (not A199)  and  (not A166) );
 a81285a <=( (not A167)  and  a81284a );
 a81288a <=( (not A201)  and  A200 );
 a81291a <=( (not A265)  and  (not A203) );
 a81292a <=( a81291a  and  a81288a );
 a81293a <=( a81292a  and  a81285a );
 a81297a <=( (not A269)  and  A268 );
 a81298a <=( (not A266)  and  a81297a );
 a81301a <=( A299  and  (not A298) );
 a81304a <=( A301  and  (not A300) );
 a81305a <=( a81304a  and  a81301a );
 a81306a <=( a81305a  and  a81298a );
 a81310a <=( (not A199)  and  (not A166) );
 a81311a <=( (not A167)  and  a81310a );
 a81314a <=( (not A201)  and  A200 );
 a81317a <=( (not A265)  and  (not A203) );
 a81318a <=( a81317a  and  a81314a );
 a81319a <=( a81318a  and  a81311a );
 a81323a <=( (not A269)  and  A268 );
 a81324a <=( (not A266)  and  a81323a );
 a81327a <=( A299  and  (not A298) );
 a81330a <=( (not A302)  and  (not A300) );
 a81331a <=( a81330a  and  a81327a );
 a81332a <=( a81331a  and  a81324a );
 a81336a <=( A199  and  (not A166) );
 a81337a <=( (not A167)  and  a81336a );
 a81340a <=( (not A202)  and  (not A200) );
 a81343a <=( A265  and  A203 );
 a81344a <=( a81343a  and  a81340a );
 a81345a <=( a81344a  and  a81337a );
 a81349a <=( (not A268)  and  (not A267) );
 a81350a <=( A266  and  a81349a );
 a81353a <=( A299  and  A298 );
 a81356a <=( (not A302)  and  A301 );
 a81357a <=( a81356a  and  a81353a );
 a81358a <=( a81357a  and  a81350a );
 a81362a <=( A199  and  (not A166) );
 a81363a <=( (not A167)  and  a81362a );
 a81366a <=( (not A202)  and  (not A200) );
 a81369a <=( A265  and  A203 );
 a81370a <=( a81369a  and  a81366a );
 a81371a <=( a81370a  and  a81363a );
 a81375a <=( (not A268)  and  (not A267) );
 a81376a <=( A266  and  a81375a );
 a81379a <=( (not A299)  and  A298 );
 a81382a <=( A302  and  (not A301) );
 a81383a <=( a81382a  and  a81379a );
 a81384a <=( a81383a  and  a81376a );
 a81388a <=( A199  and  (not A166) );
 a81389a <=( (not A167)  and  a81388a );
 a81392a <=( (not A202)  and  (not A200) );
 a81395a <=( A265  and  A203 );
 a81396a <=( a81395a  and  a81392a );
 a81397a <=( a81396a  and  a81389a );
 a81401a <=( (not A268)  and  (not A267) );
 a81402a <=( A266  and  a81401a );
 a81405a <=( A299  and  (not A298) );
 a81408a <=( A302  and  (not A301) );
 a81409a <=( a81408a  and  a81405a );
 a81410a <=( a81409a  and  a81402a );
 a81414a <=( A199  and  (not A166) );
 a81415a <=( (not A167)  and  a81414a );
 a81418a <=( (not A202)  and  (not A200) );
 a81421a <=( A265  and  A203 );
 a81422a <=( a81421a  and  a81418a );
 a81423a <=( a81422a  and  a81415a );
 a81427a <=( (not A268)  and  (not A267) );
 a81428a <=( A266  and  a81427a );
 a81431a <=( (not A299)  and  (not A298) );
 a81434a <=( (not A302)  and  A301 );
 a81435a <=( a81434a  and  a81431a );
 a81436a <=( a81435a  and  a81428a );
 a81440a <=( A199  and  (not A166) );
 a81441a <=( (not A167)  and  a81440a );
 a81444a <=( (not A202)  and  (not A200) );
 a81447a <=( A265  and  A203 );
 a81448a <=( a81447a  and  a81444a );
 a81449a <=( a81448a  and  a81441a );
 a81453a <=( A269  and  (not A267) );
 a81454a <=( A266  and  a81453a );
 a81457a <=( A299  and  A298 );
 a81460a <=( (not A302)  and  A301 );
 a81461a <=( a81460a  and  a81457a );
 a81462a <=( a81461a  and  a81454a );
 a81466a <=( A199  and  (not A166) );
 a81467a <=( (not A167)  and  a81466a );
 a81470a <=( (not A202)  and  (not A200) );
 a81473a <=( A265  and  A203 );
 a81474a <=( a81473a  and  a81470a );
 a81475a <=( a81474a  and  a81467a );
 a81479a <=( A269  and  (not A267) );
 a81480a <=( A266  and  a81479a );
 a81483a <=( (not A299)  and  A298 );
 a81486a <=( A302  and  (not A301) );
 a81487a <=( a81486a  and  a81483a );
 a81488a <=( a81487a  and  a81480a );
 a81492a <=( A199  and  (not A166) );
 a81493a <=( (not A167)  and  a81492a );
 a81496a <=( (not A202)  and  (not A200) );
 a81499a <=( A265  and  A203 );
 a81500a <=( a81499a  and  a81496a );
 a81501a <=( a81500a  and  a81493a );
 a81505a <=( A269  and  (not A267) );
 a81506a <=( A266  and  a81505a );
 a81509a <=( A299  and  (not A298) );
 a81512a <=( A302  and  (not A301) );
 a81513a <=( a81512a  and  a81509a );
 a81514a <=( a81513a  and  a81506a );
 a81518a <=( A199  and  (not A166) );
 a81519a <=( (not A167)  and  a81518a );
 a81522a <=( (not A202)  and  (not A200) );
 a81525a <=( A265  and  A203 );
 a81526a <=( a81525a  and  a81522a );
 a81527a <=( a81526a  and  a81519a );
 a81531a <=( A269  and  (not A267) );
 a81532a <=( A266  and  a81531a );
 a81535a <=( (not A299)  and  (not A298) );
 a81538a <=( (not A302)  and  A301 );
 a81539a <=( a81538a  and  a81535a );
 a81540a <=( a81539a  and  a81532a );
 a81544a <=( A199  and  (not A166) );
 a81545a <=( (not A167)  and  a81544a );
 a81548a <=( (not A202)  and  (not A200) );
 a81551a <=( (not A265)  and  A203 );
 a81552a <=( a81551a  and  a81548a );
 a81553a <=( a81552a  and  a81545a );
 a81557a <=( A268  and  (not A267) );
 a81558a <=( A266  and  a81557a );
 a81561a <=( A299  and  A298 );
 a81564a <=( (not A302)  and  A301 );
 a81565a <=( a81564a  and  a81561a );
 a81566a <=( a81565a  and  a81558a );
 a81570a <=( A199  and  (not A166) );
 a81571a <=( (not A167)  and  a81570a );
 a81574a <=( (not A202)  and  (not A200) );
 a81577a <=( (not A265)  and  A203 );
 a81578a <=( a81577a  and  a81574a );
 a81579a <=( a81578a  and  a81571a );
 a81583a <=( A268  and  (not A267) );
 a81584a <=( A266  and  a81583a );
 a81587a <=( (not A299)  and  A298 );
 a81590a <=( A302  and  (not A301) );
 a81591a <=( a81590a  and  a81587a );
 a81592a <=( a81591a  and  a81584a );
 a81596a <=( A199  and  (not A166) );
 a81597a <=( (not A167)  and  a81596a );
 a81600a <=( (not A202)  and  (not A200) );
 a81603a <=( (not A265)  and  A203 );
 a81604a <=( a81603a  and  a81600a );
 a81605a <=( a81604a  and  a81597a );
 a81609a <=( A268  and  (not A267) );
 a81610a <=( A266  and  a81609a );
 a81613a <=( A299  and  (not A298) );
 a81616a <=( A302  and  (not A301) );
 a81617a <=( a81616a  and  a81613a );
 a81618a <=( a81617a  and  a81610a );
 a81622a <=( A199  and  (not A166) );
 a81623a <=( (not A167)  and  a81622a );
 a81626a <=( (not A202)  and  (not A200) );
 a81629a <=( (not A265)  and  A203 );
 a81630a <=( a81629a  and  a81626a );
 a81631a <=( a81630a  and  a81623a );
 a81635a <=( A268  and  (not A267) );
 a81636a <=( A266  and  a81635a );
 a81639a <=( (not A299)  and  (not A298) );
 a81642a <=( (not A302)  and  A301 );
 a81643a <=( a81642a  and  a81639a );
 a81644a <=( a81643a  and  a81636a );
 a81648a <=( A199  and  (not A166) );
 a81649a <=( (not A167)  and  a81648a );
 a81652a <=( (not A202)  and  (not A200) );
 a81655a <=( (not A265)  and  A203 );
 a81656a <=( a81655a  and  a81652a );
 a81657a <=( a81656a  and  a81649a );
 a81661a <=( (not A269)  and  (not A267) );
 a81662a <=( A266  and  a81661a );
 a81665a <=( A299  and  A298 );
 a81668a <=( (not A302)  and  A301 );
 a81669a <=( a81668a  and  a81665a );
 a81670a <=( a81669a  and  a81662a );
 a81674a <=( A199  and  (not A166) );
 a81675a <=( (not A167)  and  a81674a );
 a81678a <=( (not A202)  and  (not A200) );
 a81681a <=( (not A265)  and  A203 );
 a81682a <=( a81681a  and  a81678a );
 a81683a <=( a81682a  and  a81675a );
 a81687a <=( (not A269)  and  (not A267) );
 a81688a <=( A266  and  a81687a );
 a81691a <=( (not A299)  and  A298 );
 a81694a <=( A302  and  (not A301) );
 a81695a <=( a81694a  and  a81691a );
 a81696a <=( a81695a  and  a81688a );
 a81700a <=( A199  and  (not A166) );
 a81701a <=( (not A167)  and  a81700a );
 a81704a <=( (not A202)  and  (not A200) );
 a81707a <=( (not A265)  and  A203 );
 a81708a <=( a81707a  and  a81704a );
 a81709a <=( a81708a  and  a81701a );
 a81713a <=( (not A269)  and  (not A267) );
 a81714a <=( A266  and  a81713a );
 a81717a <=( A299  and  (not A298) );
 a81720a <=( A302  and  (not A301) );
 a81721a <=( a81720a  and  a81717a );
 a81722a <=( a81721a  and  a81714a );
 a81726a <=( A199  and  (not A166) );
 a81727a <=( (not A167)  and  a81726a );
 a81730a <=( (not A202)  and  (not A200) );
 a81733a <=( (not A265)  and  A203 );
 a81734a <=( a81733a  and  a81730a );
 a81735a <=( a81734a  and  a81727a );
 a81739a <=( (not A269)  and  (not A267) );
 a81740a <=( A266  and  a81739a );
 a81743a <=( (not A299)  and  (not A298) );
 a81746a <=( (not A302)  and  A301 );
 a81747a <=( a81746a  and  a81743a );
 a81748a <=( a81747a  and  a81740a );
 a81752a <=( A199  and  (not A166) );
 a81753a <=( (not A167)  and  a81752a );
 a81756a <=( (not A202)  and  (not A200) );
 a81759a <=( A265  and  A203 );
 a81760a <=( a81759a  and  a81756a );
 a81761a <=( a81760a  and  a81753a );
 a81765a <=( A268  and  (not A267) );
 a81766a <=( (not A266)  and  a81765a );
 a81769a <=( A299  and  A298 );
 a81772a <=( (not A302)  and  A301 );
 a81773a <=( a81772a  and  a81769a );
 a81774a <=( a81773a  and  a81766a );
 a81778a <=( A199  and  (not A166) );
 a81779a <=( (not A167)  and  a81778a );
 a81782a <=( (not A202)  and  (not A200) );
 a81785a <=( A265  and  A203 );
 a81786a <=( a81785a  and  a81782a );
 a81787a <=( a81786a  and  a81779a );
 a81791a <=( A268  and  (not A267) );
 a81792a <=( (not A266)  and  a81791a );
 a81795a <=( (not A299)  and  A298 );
 a81798a <=( A302  and  (not A301) );
 a81799a <=( a81798a  and  a81795a );
 a81800a <=( a81799a  and  a81792a );
 a81804a <=( A199  and  (not A166) );
 a81805a <=( (not A167)  and  a81804a );
 a81808a <=( (not A202)  and  (not A200) );
 a81811a <=( A265  and  A203 );
 a81812a <=( a81811a  and  a81808a );
 a81813a <=( a81812a  and  a81805a );
 a81817a <=( A268  and  (not A267) );
 a81818a <=( (not A266)  and  a81817a );
 a81821a <=( A299  and  (not A298) );
 a81824a <=( A302  and  (not A301) );
 a81825a <=( a81824a  and  a81821a );
 a81826a <=( a81825a  and  a81818a );
 a81830a <=( A199  and  (not A166) );
 a81831a <=( (not A167)  and  a81830a );
 a81834a <=( (not A202)  and  (not A200) );
 a81837a <=( A265  and  A203 );
 a81838a <=( a81837a  and  a81834a );
 a81839a <=( a81838a  and  a81831a );
 a81843a <=( A268  and  (not A267) );
 a81844a <=( (not A266)  and  a81843a );
 a81847a <=( (not A299)  and  (not A298) );
 a81850a <=( (not A302)  and  A301 );
 a81851a <=( a81850a  and  a81847a );
 a81852a <=( a81851a  and  a81844a );
 a81856a <=( A199  and  (not A166) );
 a81857a <=( (not A167)  and  a81856a );
 a81860a <=( (not A202)  and  (not A200) );
 a81863a <=( A265  and  A203 );
 a81864a <=( a81863a  and  a81860a );
 a81865a <=( a81864a  and  a81857a );
 a81869a <=( (not A269)  and  (not A267) );
 a81870a <=( (not A266)  and  a81869a );
 a81873a <=( A299  and  A298 );
 a81876a <=( (not A302)  and  A301 );
 a81877a <=( a81876a  and  a81873a );
 a81878a <=( a81877a  and  a81870a );
 a81882a <=( A199  and  (not A166) );
 a81883a <=( (not A167)  and  a81882a );
 a81886a <=( (not A202)  and  (not A200) );
 a81889a <=( A265  and  A203 );
 a81890a <=( a81889a  and  a81886a );
 a81891a <=( a81890a  and  a81883a );
 a81895a <=( (not A269)  and  (not A267) );
 a81896a <=( (not A266)  and  a81895a );
 a81899a <=( (not A299)  and  A298 );
 a81902a <=( A302  and  (not A301) );
 a81903a <=( a81902a  and  a81899a );
 a81904a <=( a81903a  and  a81896a );
 a81908a <=( A199  and  (not A166) );
 a81909a <=( (not A167)  and  a81908a );
 a81912a <=( (not A202)  and  (not A200) );
 a81915a <=( A265  and  A203 );
 a81916a <=( a81915a  and  a81912a );
 a81917a <=( a81916a  and  a81909a );
 a81921a <=( (not A269)  and  (not A267) );
 a81922a <=( (not A266)  and  a81921a );
 a81925a <=( A299  and  (not A298) );
 a81928a <=( A302  and  (not A301) );
 a81929a <=( a81928a  and  a81925a );
 a81930a <=( a81929a  and  a81922a );
 a81934a <=( A199  and  (not A166) );
 a81935a <=( (not A167)  and  a81934a );
 a81938a <=( (not A202)  and  (not A200) );
 a81941a <=( A265  and  A203 );
 a81942a <=( a81941a  and  a81938a );
 a81943a <=( a81942a  and  a81935a );
 a81947a <=( (not A269)  and  (not A267) );
 a81948a <=( (not A266)  and  a81947a );
 a81951a <=( (not A299)  and  (not A298) );
 a81954a <=( (not A302)  and  A301 );
 a81955a <=( a81954a  and  a81951a );
 a81956a <=( a81955a  and  a81948a );
 a81960a <=( A199  and  (not A166) );
 a81961a <=( (not A167)  and  a81960a );
 a81964a <=( (not A201)  and  (not A200) );
 a81967a <=( A265  and  A202 );
 a81968a <=( a81967a  and  a81964a );
 a81969a <=( a81968a  and  a81961a );
 a81973a <=( (not A269)  and  A268 );
 a81974a <=( A266  and  a81973a );
 a81977a <=( A299  and  A298 );
 a81980a <=( (not A301)  and  (not A300) );
 a81981a <=( a81980a  and  a81977a );
 a81982a <=( a81981a  and  a81974a );
 a81986a <=( A199  and  (not A166) );
 a81987a <=( (not A167)  and  a81986a );
 a81990a <=( (not A201)  and  (not A200) );
 a81993a <=( A265  and  A202 );
 a81994a <=( a81993a  and  a81990a );
 a81995a <=( a81994a  and  a81987a );
 a81999a <=( (not A269)  and  A268 );
 a82000a <=( A266  and  a81999a );
 a82003a <=( A299  and  A298 );
 a82006a <=( A302  and  (not A300) );
 a82007a <=( a82006a  and  a82003a );
 a82008a <=( a82007a  and  a82000a );
 a82012a <=( A199  and  (not A166) );
 a82013a <=( (not A167)  and  a82012a );
 a82016a <=( (not A201)  and  (not A200) );
 a82019a <=( A265  and  A202 );
 a82020a <=( a82019a  and  a82016a );
 a82021a <=( a82020a  and  a82013a );
 a82025a <=( (not A269)  and  A268 );
 a82026a <=( A266  and  a82025a );
 a82029a <=( (not A299)  and  A298 );
 a82032a <=( A301  and  (not A300) );
 a82033a <=( a82032a  and  a82029a );
 a82034a <=( a82033a  and  a82026a );
 a82038a <=( A199  and  (not A166) );
 a82039a <=( (not A167)  and  a82038a );
 a82042a <=( (not A201)  and  (not A200) );
 a82045a <=( A265  and  A202 );
 a82046a <=( a82045a  and  a82042a );
 a82047a <=( a82046a  and  a82039a );
 a82051a <=( (not A269)  and  A268 );
 a82052a <=( A266  and  a82051a );
 a82055a <=( (not A299)  and  A298 );
 a82058a <=( (not A302)  and  (not A300) );
 a82059a <=( a82058a  and  a82055a );
 a82060a <=( a82059a  and  a82052a );
 a82064a <=( A199  and  (not A166) );
 a82065a <=( (not A167)  and  a82064a );
 a82068a <=( (not A201)  and  (not A200) );
 a82071a <=( A265  and  A202 );
 a82072a <=( a82071a  and  a82068a );
 a82073a <=( a82072a  and  a82065a );
 a82077a <=( (not A269)  and  A268 );
 a82078a <=( A266  and  a82077a );
 a82081a <=( A299  and  (not A298) );
 a82084a <=( A301  and  (not A300) );
 a82085a <=( a82084a  and  a82081a );
 a82086a <=( a82085a  and  a82078a );
 a82090a <=( A199  and  (not A166) );
 a82091a <=( (not A167)  and  a82090a );
 a82094a <=( (not A201)  and  (not A200) );
 a82097a <=( A265  and  A202 );
 a82098a <=( a82097a  and  a82094a );
 a82099a <=( a82098a  and  a82091a );
 a82103a <=( (not A269)  and  A268 );
 a82104a <=( A266  and  a82103a );
 a82107a <=( A299  and  (not A298) );
 a82110a <=( (not A302)  and  (not A300) );
 a82111a <=( a82110a  and  a82107a );
 a82112a <=( a82111a  and  a82104a );
 a82116a <=( A199  and  (not A166) );
 a82117a <=( (not A167)  and  a82116a );
 a82120a <=( (not A201)  and  (not A200) );
 a82123a <=( (not A265)  and  A202 );
 a82124a <=( a82123a  and  a82120a );
 a82125a <=( a82124a  and  a82117a );
 a82129a <=( A269  and  (not A268) );
 a82130a <=( A266  and  a82129a );
 a82133a <=( A299  and  A298 );
 a82136a <=( (not A301)  and  (not A300) );
 a82137a <=( a82136a  and  a82133a );
 a82138a <=( a82137a  and  a82130a );
 a82142a <=( A199  and  (not A166) );
 a82143a <=( (not A167)  and  a82142a );
 a82146a <=( (not A201)  and  (not A200) );
 a82149a <=( (not A265)  and  A202 );
 a82150a <=( a82149a  and  a82146a );
 a82151a <=( a82150a  and  a82143a );
 a82155a <=( A269  and  (not A268) );
 a82156a <=( A266  and  a82155a );
 a82159a <=( A299  and  A298 );
 a82162a <=( A302  and  (not A300) );
 a82163a <=( a82162a  and  a82159a );
 a82164a <=( a82163a  and  a82156a );
 a82168a <=( A199  and  (not A166) );
 a82169a <=( (not A167)  and  a82168a );
 a82172a <=( (not A201)  and  (not A200) );
 a82175a <=( (not A265)  and  A202 );
 a82176a <=( a82175a  and  a82172a );
 a82177a <=( a82176a  and  a82169a );
 a82181a <=( A269  and  (not A268) );
 a82182a <=( A266  and  a82181a );
 a82185a <=( (not A299)  and  A298 );
 a82188a <=( A301  and  (not A300) );
 a82189a <=( a82188a  and  a82185a );
 a82190a <=( a82189a  and  a82182a );
 a82194a <=( A199  and  (not A166) );
 a82195a <=( (not A167)  and  a82194a );
 a82198a <=( (not A201)  and  (not A200) );
 a82201a <=( (not A265)  and  A202 );
 a82202a <=( a82201a  and  a82198a );
 a82203a <=( a82202a  and  a82195a );
 a82207a <=( A269  and  (not A268) );
 a82208a <=( A266  and  a82207a );
 a82211a <=( (not A299)  and  A298 );
 a82214a <=( (not A302)  and  (not A300) );
 a82215a <=( a82214a  and  a82211a );
 a82216a <=( a82215a  and  a82208a );
 a82220a <=( A199  and  (not A166) );
 a82221a <=( (not A167)  and  a82220a );
 a82224a <=( (not A201)  and  (not A200) );
 a82227a <=( (not A265)  and  A202 );
 a82228a <=( a82227a  and  a82224a );
 a82229a <=( a82228a  and  a82221a );
 a82233a <=( A269  and  (not A268) );
 a82234a <=( A266  and  a82233a );
 a82237a <=( A299  and  (not A298) );
 a82240a <=( A301  and  (not A300) );
 a82241a <=( a82240a  and  a82237a );
 a82242a <=( a82241a  and  a82234a );
 a82246a <=( A199  and  (not A166) );
 a82247a <=( (not A167)  and  a82246a );
 a82250a <=( (not A201)  and  (not A200) );
 a82253a <=( (not A265)  and  A202 );
 a82254a <=( a82253a  and  a82250a );
 a82255a <=( a82254a  and  a82247a );
 a82259a <=( A269  and  (not A268) );
 a82260a <=( A266  and  a82259a );
 a82263a <=( A299  and  (not A298) );
 a82266a <=( (not A302)  and  (not A300) );
 a82267a <=( a82266a  and  a82263a );
 a82268a <=( a82267a  and  a82260a );
 a82272a <=( A199  and  (not A166) );
 a82273a <=( (not A167)  and  a82272a );
 a82276a <=( (not A201)  and  (not A200) );
 a82279a <=( A265  and  A202 );
 a82280a <=( a82279a  and  a82276a );
 a82281a <=( a82280a  and  a82273a );
 a82285a <=( A269  and  (not A268) );
 a82286a <=( (not A266)  and  a82285a );
 a82289a <=( A299  and  A298 );
 a82292a <=( (not A301)  and  (not A300) );
 a82293a <=( a82292a  and  a82289a );
 a82294a <=( a82293a  and  a82286a );
 a82298a <=( A199  and  (not A166) );
 a82299a <=( (not A167)  and  a82298a );
 a82302a <=( (not A201)  and  (not A200) );
 a82305a <=( A265  and  A202 );
 a82306a <=( a82305a  and  a82302a );
 a82307a <=( a82306a  and  a82299a );
 a82311a <=( A269  and  (not A268) );
 a82312a <=( (not A266)  and  a82311a );
 a82315a <=( A299  and  A298 );
 a82318a <=( A302  and  (not A300) );
 a82319a <=( a82318a  and  a82315a );
 a82320a <=( a82319a  and  a82312a );
 a82324a <=( A199  and  (not A166) );
 a82325a <=( (not A167)  and  a82324a );
 a82328a <=( (not A201)  and  (not A200) );
 a82331a <=( A265  and  A202 );
 a82332a <=( a82331a  and  a82328a );
 a82333a <=( a82332a  and  a82325a );
 a82337a <=( A269  and  (not A268) );
 a82338a <=( (not A266)  and  a82337a );
 a82341a <=( (not A299)  and  A298 );
 a82344a <=( A301  and  (not A300) );
 a82345a <=( a82344a  and  a82341a );
 a82346a <=( a82345a  and  a82338a );
 a82350a <=( A199  and  (not A166) );
 a82351a <=( (not A167)  and  a82350a );
 a82354a <=( (not A201)  and  (not A200) );
 a82357a <=( A265  and  A202 );
 a82358a <=( a82357a  and  a82354a );
 a82359a <=( a82358a  and  a82351a );
 a82363a <=( A269  and  (not A268) );
 a82364a <=( (not A266)  and  a82363a );
 a82367a <=( (not A299)  and  A298 );
 a82370a <=( (not A302)  and  (not A300) );
 a82371a <=( a82370a  and  a82367a );
 a82372a <=( a82371a  and  a82364a );
 a82376a <=( A199  and  (not A166) );
 a82377a <=( (not A167)  and  a82376a );
 a82380a <=( (not A201)  and  (not A200) );
 a82383a <=( A265  and  A202 );
 a82384a <=( a82383a  and  a82380a );
 a82385a <=( a82384a  and  a82377a );
 a82389a <=( A269  and  (not A268) );
 a82390a <=( (not A266)  and  a82389a );
 a82393a <=( A299  and  (not A298) );
 a82396a <=( A301  and  (not A300) );
 a82397a <=( a82396a  and  a82393a );
 a82398a <=( a82397a  and  a82390a );
 a82402a <=( A199  and  (not A166) );
 a82403a <=( (not A167)  and  a82402a );
 a82406a <=( (not A201)  and  (not A200) );
 a82409a <=( A265  and  A202 );
 a82410a <=( a82409a  and  a82406a );
 a82411a <=( a82410a  and  a82403a );
 a82415a <=( A269  and  (not A268) );
 a82416a <=( (not A266)  and  a82415a );
 a82419a <=( A299  and  (not A298) );
 a82422a <=( (not A302)  and  (not A300) );
 a82423a <=( a82422a  and  a82419a );
 a82424a <=( a82423a  and  a82416a );
 a82428a <=( A199  and  (not A166) );
 a82429a <=( (not A167)  and  a82428a );
 a82432a <=( (not A201)  and  (not A200) );
 a82435a <=( (not A265)  and  A202 );
 a82436a <=( a82435a  and  a82432a );
 a82437a <=( a82436a  and  a82429a );
 a82441a <=( (not A269)  and  A268 );
 a82442a <=( (not A266)  and  a82441a );
 a82445a <=( A299  and  A298 );
 a82448a <=( (not A301)  and  (not A300) );
 a82449a <=( a82448a  and  a82445a );
 a82450a <=( a82449a  and  a82442a );
 a82454a <=( A199  and  (not A166) );
 a82455a <=( (not A167)  and  a82454a );
 a82458a <=( (not A201)  and  (not A200) );
 a82461a <=( (not A265)  and  A202 );
 a82462a <=( a82461a  and  a82458a );
 a82463a <=( a82462a  and  a82455a );
 a82467a <=( (not A269)  and  A268 );
 a82468a <=( (not A266)  and  a82467a );
 a82471a <=( A299  and  A298 );
 a82474a <=( A302  and  (not A300) );
 a82475a <=( a82474a  and  a82471a );
 a82476a <=( a82475a  and  a82468a );
 a82480a <=( A199  and  (not A166) );
 a82481a <=( (not A167)  and  a82480a );
 a82484a <=( (not A201)  and  (not A200) );
 a82487a <=( (not A265)  and  A202 );
 a82488a <=( a82487a  and  a82484a );
 a82489a <=( a82488a  and  a82481a );
 a82493a <=( (not A269)  and  A268 );
 a82494a <=( (not A266)  and  a82493a );
 a82497a <=( (not A299)  and  A298 );
 a82500a <=( A301  and  (not A300) );
 a82501a <=( a82500a  and  a82497a );
 a82502a <=( a82501a  and  a82494a );
 a82506a <=( A199  and  (not A166) );
 a82507a <=( (not A167)  and  a82506a );
 a82510a <=( (not A201)  and  (not A200) );
 a82513a <=( (not A265)  and  A202 );
 a82514a <=( a82513a  and  a82510a );
 a82515a <=( a82514a  and  a82507a );
 a82519a <=( (not A269)  and  A268 );
 a82520a <=( (not A266)  and  a82519a );
 a82523a <=( (not A299)  and  A298 );
 a82526a <=( (not A302)  and  (not A300) );
 a82527a <=( a82526a  and  a82523a );
 a82528a <=( a82527a  and  a82520a );
 a82532a <=( A199  and  (not A166) );
 a82533a <=( (not A167)  and  a82532a );
 a82536a <=( (not A201)  and  (not A200) );
 a82539a <=( (not A265)  and  A202 );
 a82540a <=( a82539a  and  a82536a );
 a82541a <=( a82540a  and  a82533a );
 a82545a <=( (not A269)  and  A268 );
 a82546a <=( (not A266)  and  a82545a );
 a82549a <=( A299  and  (not A298) );
 a82552a <=( A301  and  (not A300) );
 a82553a <=( a82552a  and  a82549a );
 a82554a <=( a82553a  and  a82546a );
 a82558a <=( A199  and  (not A166) );
 a82559a <=( (not A167)  and  a82558a );
 a82562a <=( (not A201)  and  (not A200) );
 a82565a <=( (not A265)  and  A202 );
 a82566a <=( a82565a  and  a82562a );
 a82567a <=( a82566a  and  a82559a );
 a82571a <=( (not A269)  and  A268 );
 a82572a <=( (not A266)  and  a82571a );
 a82575a <=( A299  and  (not A298) );
 a82578a <=( (not A302)  and  (not A300) );
 a82579a <=( a82578a  and  a82575a );
 a82580a <=( a82579a  and  a82572a );
 a82584a <=( A199  and  (not A166) );
 a82585a <=( (not A167)  and  a82584a );
 a82588a <=( (not A201)  and  (not A200) );
 a82591a <=( A265  and  (not A203) );
 a82592a <=( a82591a  and  a82588a );
 a82593a <=( a82592a  and  a82585a );
 a82597a <=( (not A269)  and  A268 );
 a82598a <=( A266  and  a82597a );
 a82601a <=( A299  and  A298 );
 a82604a <=( (not A301)  and  (not A300) );
 a82605a <=( a82604a  and  a82601a );
 a82606a <=( a82605a  and  a82598a );
 a82610a <=( A199  and  (not A166) );
 a82611a <=( (not A167)  and  a82610a );
 a82614a <=( (not A201)  and  (not A200) );
 a82617a <=( A265  and  (not A203) );
 a82618a <=( a82617a  and  a82614a );
 a82619a <=( a82618a  and  a82611a );
 a82623a <=( (not A269)  and  A268 );
 a82624a <=( A266  and  a82623a );
 a82627a <=( A299  and  A298 );
 a82630a <=( A302  and  (not A300) );
 a82631a <=( a82630a  and  a82627a );
 a82632a <=( a82631a  and  a82624a );
 a82636a <=( A199  and  (not A166) );
 a82637a <=( (not A167)  and  a82636a );
 a82640a <=( (not A201)  and  (not A200) );
 a82643a <=( A265  and  (not A203) );
 a82644a <=( a82643a  and  a82640a );
 a82645a <=( a82644a  and  a82637a );
 a82649a <=( (not A269)  and  A268 );
 a82650a <=( A266  and  a82649a );
 a82653a <=( (not A299)  and  A298 );
 a82656a <=( A301  and  (not A300) );
 a82657a <=( a82656a  and  a82653a );
 a82658a <=( a82657a  and  a82650a );
 a82662a <=( A199  and  (not A166) );
 a82663a <=( (not A167)  and  a82662a );
 a82666a <=( (not A201)  and  (not A200) );
 a82669a <=( A265  and  (not A203) );
 a82670a <=( a82669a  and  a82666a );
 a82671a <=( a82670a  and  a82663a );
 a82675a <=( (not A269)  and  A268 );
 a82676a <=( A266  and  a82675a );
 a82679a <=( (not A299)  and  A298 );
 a82682a <=( (not A302)  and  (not A300) );
 a82683a <=( a82682a  and  a82679a );
 a82684a <=( a82683a  and  a82676a );
 a82688a <=( A199  and  (not A166) );
 a82689a <=( (not A167)  and  a82688a );
 a82692a <=( (not A201)  and  (not A200) );
 a82695a <=( A265  and  (not A203) );
 a82696a <=( a82695a  and  a82692a );
 a82697a <=( a82696a  and  a82689a );
 a82701a <=( (not A269)  and  A268 );
 a82702a <=( A266  and  a82701a );
 a82705a <=( A299  and  (not A298) );
 a82708a <=( A301  and  (not A300) );
 a82709a <=( a82708a  and  a82705a );
 a82710a <=( a82709a  and  a82702a );
 a82714a <=( A199  and  (not A166) );
 a82715a <=( (not A167)  and  a82714a );
 a82718a <=( (not A201)  and  (not A200) );
 a82721a <=( A265  and  (not A203) );
 a82722a <=( a82721a  and  a82718a );
 a82723a <=( a82722a  and  a82715a );
 a82727a <=( (not A269)  and  A268 );
 a82728a <=( A266  and  a82727a );
 a82731a <=( A299  and  (not A298) );
 a82734a <=( (not A302)  and  (not A300) );
 a82735a <=( a82734a  and  a82731a );
 a82736a <=( a82735a  and  a82728a );
 a82740a <=( A199  and  (not A166) );
 a82741a <=( (not A167)  and  a82740a );
 a82744a <=( (not A201)  and  (not A200) );
 a82747a <=( (not A265)  and  (not A203) );
 a82748a <=( a82747a  and  a82744a );
 a82749a <=( a82748a  and  a82741a );
 a82753a <=( A269  and  (not A268) );
 a82754a <=( A266  and  a82753a );
 a82757a <=( A299  and  A298 );
 a82760a <=( (not A301)  and  (not A300) );
 a82761a <=( a82760a  and  a82757a );
 a82762a <=( a82761a  and  a82754a );
 a82766a <=( A199  and  (not A166) );
 a82767a <=( (not A167)  and  a82766a );
 a82770a <=( (not A201)  and  (not A200) );
 a82773a <=( (not A265)  and  (not A203) );
 a82774a <=( a82773a  and  a82770a );
 a82775a <=( a82774a  and  a82767a );
 a82779a <=( A269  and  (not A268) );
 a82780a <=( A266  and  a82779a );
 a82783a <=( A299  and  A298 );
 a82786a <=( A302  and  (not A300) );
 a82787a <=( a82786a  and  a82783a );
 a82788a <=( a82787a  and  a82780a );
 a82792a <=( A199  and  (not A166) );
 a82793a <=( (not A167)  and  a82792a );
 a82796a <=( (not A201)  and  (not A200) );
 a82799a <=( (not A265)  and  (not A203) );
 a82800a <=( a82799a  and  a82796a );
 a82801a <=( a82800a  and  a82793a );
 a82805a <=( A269  and  (not A268) );
 a82806a <=( A266  and  a82805a );
 a82809a <=( (not A299)  and  A298 );
 a82812a <=( A301  and  (not A300) );
 a82813a <=( a82812a  and  a82809a );
 a82814a <=( a82813a  and  a82806a );
 a82818a <=( A199  and  (not A166) );
 a82819a <=( (not A167)  and  a82818a );
 a82822a <=( (not A201)  and  (not A200) );
 a82825a <=( (not A265)  and  (not A203) );
 a82826a <=( a82825a  and  a82822a );
 a82827a <=( a82826a  and  a82819a );
 a82831a <=( A269  and  (not A268) );
 a82832a <=( A266  and  a82831a );
 a82835a <=( (not A299)  and  A298 );
 a82838a <=( (not A302)  and  (not A300) );
 a82839a <=( a82838a  and  a82835a );
 a82840a <=( a82839a  and  a82832a );
 a82844a <=( A199  and  (not A166) );
 a82845a <=( (not A167)  and  a82844a );
 a82848a <=( (not A201)  and  (not A200) );
 a82851a <=( (not A265)  and  (not A203) );
 a82852a <=( a82851a  and  a82848a );
 a82853a <=( a82852a  and  a82845a );
 a82857a <=( A269  and  (not A268) );
 a82858a <=( A266  and  a82857a );
 a82861a <=( A299  and  (not A298) );
 a82864a <=( A301  and  (not A300) );
 a82865a <=( a82864a  and  a82861a );
 a82866a <=( a82865a  and  a82858a );
 a82870a <=( A199  and  (not A166) );
 a82871a <=( (not A167)  and  a82870a );
 a82874a <=( (not A201)  and  (not A200) );
 a82877a <=( (not A265)  and  (not A203) );
 a82878a <=( a82877a  and  a82874a );
 a82879a <=( a82878a  and  a82871a );
 a82883a <=( A269  and  (not A268) );
 a82884a <=( A266  and  a82883a );
 a82887a <=( A299  and  (not A298) );
 a82890a <=( (not A302)  and  (not A300) );
 a82891a <=( a82890a  and  a82887a );
 a82892a <=( a82891a  and  a82884a );
 a82896a <=( A199  and  (not A166) );
 a82897a <=( (not A167)  and  a82896a );
 a82900a <=( (not A201)  and  (not A200) );
 a82903a <=( A265  and  (not A203) );
 a82904a <=( a82903a  and  a82900a );
 a82905a <=( a82904a  and  a82897a );
 a82909a <=( A269  and  (not A268) );
 a82910a <=( (not A266)  and  a82909a );
 a82913a <=( A299  and  A298 );
 a82916a <=( (not A301)  and  (not A300) );
 a82917a <=( a82916a  and  a82913a );
 a82918a <=( a82917a  and  a82910a );
 a82922a <=( A199  and  (not A166) );
 a82923a <=( (not A167)  and  a82922a );
 a82926a <=( (not A201)  and  (not A200) );
 a82929a <=( A265  and  (not A203) );
 a82930a <=( a82929a  and  a82926a );
 a82931a <=( a82930a  and  a82923a );
 a82935a <=( A269  and  (not A268) );
 a82936a <=( (not A266)  and  a82935a );
 a82939a <=( A299  and  A298 );
 a82942a <=( A302  and  (not A300) );
 a82943a <=( a82942a  and  a82939a );
 a82944a <=( a82943a  and  a82936a );
 a82948a <=( A199  and  (not A166) );
 a82949a <=( (not A167)  and  a82948a );
 a82952a <=( (not A201)  and  (not A200) );
 a82955a <=( A265  and  (not A203) );
 a82956a <=( a82955a  and  a82952a );
 a82957a <=( a82956a  and  a82949a );
 a82961a <=( A269  and  (not A268) );
 a82962a <=( (not A266)  and  a82961a );
 a82965a <=( (not A299)  and  A298 );
 a82968a <=( A301  and  (not A300) );
 a82969a <=( a82968a  and  a82965a );
 a82970a <=( a82969a  and  a82962a );
 a82974a <=( A199  and  (not A166) );
 a82975a <=( (not A167)  and  a82974a );
 a82978a <=( (not A201)  and  (not A200) );
 a82981a <=( A265  and  (not A203) );
 a82982a <=( a82981a  and  a82978a );
 a82983a <=( a82982a  and  a82975a );
 a82987a <=( A269  and  (not A268) );
 a82988a <=( (not A266)  and  a82987a );
 a82991a <=( (not A299)  and  A298 );
 a82994a <=( (not A302)  and  (not A300) );
 a82995a <=( a82994a  and  a82991a );
 a82996a <=( a82995a  and  a82988a );
 a83000a <=( A199  and  (not A166) );
 a83001a <=( (not A167)  and  a83000a );
 a83004a <=( (not A201)  and  (not A200) );
 a83007a <=( A265  and  (not A203) );
 a83008a <=( a83007a  and  a83004a );
 a83009a <=( a83008a  and  a83001a );
 a83013a <=( A269  and  (not A268) );
 a83014a <=( (not A266)  and  a83013a );
 a83017a <=( A299  and  (not A298) );
 a83020a <=( A301  and  (not A300) );
 a83021a <=( a83020a  and  a83017a );
 a83022a <=( a83021a  and  a83014a );
 a83026a <=( A199  and  (not A166) );
 a83027a <=( (not A167)  and  a83026a );
 a83030a <=( (not A201)  and  (not A200) );
 a83033a <=( A265  and  (not A203) );
 a83034a <=( a83033a  and  a83030a );
 a83035a <=( a83034a  and  a83027a );
 a83039a <=( A269  and  (not A268) );
 a83040a <=( (not A266)  and  a83039a );
 a83043a <=( A299  and  (not A298) );
 a83046a <=( (not A302)  and  (not A300) );
 a83047a <=( a83046a  and  a83043a );
 a83048a <=( a83047a  and  a83040a );
 a83052a <=( A199  and  (not A166) );
 a83053a <=( (not A167)  and  a83052a );
 a83056a <=( (not A201)  and  (not A200) );
 a83059a <=( (not A265)  and  (not A203) );
 a83060a <=( a83059a  and  a83056a );
 a83061a <=( a83060a  and  a83053a );
 a83065a <=( (not A269)  and  A268 );
 a83066a <=( (not A266)  and  a83065a );
 a83069a <=( A299  and  A298 );
 a83072a <=( (not A301)  and  (not A300) );
 a83073a <=( a83072a  and  a83069a );
 a83074a <=( a83073a  and  a83066a );
 a83078a <=( A199  and  (not A166) );
 a83079a <=( (not A167)  and  a83078a );
 a83082a <=( (not A201)  and  (not A200) );
 a83085a <=( (not A265)  and  (not A203) );
 a83086a <=( a83085a  and  a83082a );
 a83087a <=( a83086a  and  a83079a );
 a83091a <=( (not A269)  and  A268 );
 a83092a <=( (not A266)  and  a83091a );
 a83095a <=( A299  and  A298 );
 a83098a <=( A302  and  (not A300) );
 a83099a <=( a83098a  and  a83095a );
 a83100a <=( a83099a  and  a83092a );
 a83104a <=( A199  and  (not A166) );
 a83105a <=( (not A167)  and  a83104a );
 a83108a <=( (not A201)  and  (not A200) );
 a83111a <=( (not A265)  and  (not A203) );
 a83112a <=( a83111a  and  a83108a );
 a83113a <=( a83112a  and  a83105a );
 a83117a <=( (not A269)  and  A268 );
 a83118a <=( (not A266)  and  a83117a );
 a83121a <=( (not A299)  and  A298 );
 a83124a <=( A301  and  (not A300) );
 a83125a <=( a83124a  and  a83121a );
 a83126a <=( a83125a  and  a83118a );
 a83130a <=( A199  and  (not A166) );
 a83131a <=( (not A167)  and  a83130a );
 a83134a <=( (not A201)  and  (not A200) );
 a83137a <=( (not A265)  and  (not A203) );
 a83138a <=( a83137a  and  a83134a );
 a83139a <=( a83138a  and  a83131a );
 a83143a <=( (not A269)  and  A268 );
 a83144a <=( (not A266)  and  a83143a );
 a83147a <=( (not A299)  and  A298 );
 a83150a <=( (not A302)  and  (not A300) );
 a83151a <=( a83150a  and  a83147a );
 a83152a <=( a83151a  and  a83144a );
 a83156a <=( A199  and  (not A166) );
 a83157a <=( (not A167)  and  a83156a );
 a83160a <=( (not A201)  and  (not A200) );
 a83163a <=( (not A265)  and  (not A203) );
 a83164a <=( a83163a  and  a83160a );
 a83165a <=( a83164a  and  a83157a );
 a83169a <=( (not A269)  and  A268 );
 a83170a <=( (not A266)  and  a83169a );
 a83173a <=( A299  and  (not A298) );
 a83176a <=( A301  and  (not A300) );
 a83177a <=( a83176a  and  a83173a );
 a83178a <=( a83177a  and  a83170a );
 a83182a <=( A199  and  (not A166) );
 a83183a <=( (not A167)  and  a83182a );
 a83186a <=( (not A201)  and  (not A200) );
 a83189a <=( (not A265)  and  (not A203) );
 a83190a <=( a83189a  and  a83186a );
 a83191a <=( a83190a  and  a83183a );
 a83195a <=( (not A269)  and  A268 );
 a83196a <=( (not A266)  and  a83195a );
 a83199a <=( A299  and  (not A298) );
 a83202a <=( (not A302)  and  (not A300) );
 a83203a <=( a83202a  and  a83199a );
 a83204a <=( a83203a  and  a83196a );
 a83208a <=( (not A199)  and  (not A166) );
 a83209a <=( (not A167)  and  a83208a );
 a83212a <=( A202  and  (not A200) );
 a83215a <=( A265  and  (not A203) );
 a83216a <=( a83215a  and  a83212a );
 a83217a <=( a83216a  and  a83209a );
 a83221a <=( (not A268)  and  (not A267) );
 a83222a <=( A266  and  a83221a );
 a83225a <=( A299  and  A298 );
 a83228a <=( (not A302)  and  A301 );
 a83229a <=( a83228a  and  a83225a );
 a83230a <=( a83229a  and  a83222a );
 a83234a <=( (not A199)  and  (not A166) );
 a83235a <=( (not A167)  and  a83234a );
 a83238a <=( A202  and  (not A200) );
 a83241a <=( A265  and  (not A203) );
 a83242a <=( a83241a  and  a83238a );
 a83243a <=( a83242a  and  a83235a );
 a83247a <=( (not A268)  and  (not A267) );
 a83248a <=( A266  and  a83247a );
 a83251a <=( (not A299)  and  A298 );
 a83254a <=( A302  and  (not A301) );
 a83255a <=( a83254a  and  a83251a );
 a83256a <=( a83255a  and  a83248a );
 a83260a <=( (not A199)  and  (not A166) );
 a83261a <=( (not A167)  and  a83260a );
 a83264a <=( A202  and  (not A200) );
 a83267a <=( A265  and  (not A203) );
 a83268a <=( a83267a  and  a83264a );
 a83269a <=( a83268a  and  a83261a );
 a83273a <=( (not A268)  and  (not A267) );
 a83274a <=( A266  and  a83273a );
 a83277a <=( A299  and  (not A298) );
 a83280a <=( A302  and  (not A301) );
 a83281a <=( a83280a  and  a83277a );
 a83282a <=( a83281a  and  a83274a );
 a83286a <=( (not A199)  and  (not A166) );
 a83287a <=( (not A167)  and  a83286a );
 a83290a <=( A202  and  (not A200) );
 a83293a <=( A265  and  (not A203) );
 a83294a <=( a83293a  and  a83290a );
 a83295a <=( a83294a  and  a83287a );
 a83299a <=( (not A268)  and  (not A267) );
 a83300a <=( A266  and  a83299a );
 a83303a <=( (not A299)  and  (not A298) );
 a83306a <=( (not A302)  and  A301 );
 a83307a <=( a83306a  and  a83303a );
 a83308a <=( a83307a  and  a83300a );
 a83312a <=( (not A199)  and  (not A166) );
 a83313a <=( (not A167)  and  a83312a );
 a83316a <=( A202  and  (not A200) );
 a83319a <=( A265  and  (not A203) );
 a83320a <=( a83319a  and  a83316a );
 a83321a <=( a83320a  and  a83313a );
 a83325a <=( A269  and  (not A267) );
 a83326a <=( A266  and  a83325a );
 a83329a <=( A299  and  A298 );
 a83332a <=( (not A302)  and  A301 );
 a83333a <=( a83332a  and  a83329a );
 a83334a <=( a83333a  and  a83326a );
 a83338a <=( (not A199)  and  (not A166) );
 a83339a <=( (not A167)  and  a83338a );
 a83342a <=( A202  and  (not A200) );
 a83345a <=( A265  and  (not A203) );
 a83346a <=( a83345a  and  a83342a );
 a83347a <=( a83346a  and  a83339a );
 a83351a <=( A269  and  (not A267) );
 a83352a <=( A266  and  a83351a );
 a83355a <=( (not A299)  and  A298 );
 a83358a <=( A302  and  (not A301) );
 a83359a <=( a83358a  and  a83355a );
 a83360a <=( a83359a  and  a83352a );
 a83364a <=( (not A199)  and  (not A166) );
 a83365a <=( (not A167)  and  a83364a );
 a83368a <=( A202  and  (not A200) );
 a83371a <=( A265  and  (not A203) );
 a83372a <=( a83371a  and  a83368a );
 a83373a <=( a83372a  and  a83365a );
 a83377a <=( A269  and  (not A267) );
 a83378a <=( A266  and  a83377a );
 a83381a <=( A299  and  (not A298) );
 a83384a <=( A302  and  (not A301) );
 a83385a <=( a83384a  and  a83381a );
 a83386a <=( a83385a  and  a83378a );
 a83390a <=( (not A199)  and  (not A166) );
 a83391a <=( (not A167)  and  a83390a );
 a83394a <=( A202  and  (not A200) );
 a83397a <=( A265  and  (not A203) );
 a83398a <=( a83397a  and  a83394a );
 a83399a <=( a83398a  and  a83391a );
 a83403a <=( A269  and  (not A267) );
 a83404a <=( A266  and  a83403a );
 a83407a <=( (not A299)  and  (not A298) );
 a83410a <=( (not A302)  and  A301 );
 a83411a <=( a83410a  and  a83407a );
 a83412a <=( a83411a  and  a83404a );
 a83416a <=( (not A199)  and  (not A166) );
 a83417a <=( (not A167)  and  a83416a );
 a83420a <=( A202  and  (not A200) );
 a83423a <=( (not A265)  and  (not A203) );
 a83424a <=( a83423a  and  a83420a );
 a83425a <=( a83424a  and  a83417a );
 a83429a <=( A268  and  (not A267) );
 a83430a <=( A266  and  a83429a );
 a83433a <=( A299  and  A298 );
 a83436a <=( (not A302)  and  A301 );
 a83437a <=( a83436a  and  a83433a );
 a83438a <=( a83437a  and  a83430a );
 a83442a <=( (not A199)  and  (not A166) );
 a83443a <=( (not A167)  and  a83442a );
 a83446a <=( A202  and  (not A200) );
 a83449a <=( (not A265)  and  (not A203) );
 a83450a <=( a83449a  and  a83446a );
 a83451a <=( a83450a  and  a83443a );
 a83455a <=( A268  and  (not A267) );
 a83456a <=( A266  and  a83455a );
 a83459a <=( (not A299)  and  A298 );
 a83462a <=( A302  and  (not A301) );
 a83463a <=( a83462a  and  a83459a );
 a83464a <=( a83463a  and  a83456a );
 a83468a <=( (not A199)  and  (not A166) );
 a83469a <=( (not A167)  and  a83468a );
 a83472a <=( A202  and  (not A200) );
 a83475a <=( (not A265)  and  (not A203) );
 a83476a <=( a83475a  and  a83472a );
 a83477a <=( a83476a  and  a83469a );
 a83481a <=( A268  and  (not A267) );
 a83482a <=( A266  and  a83481a );
 a83485a <=( A299  and  (not A298) );
 a83488a <=( A302  and  (not A301) );
 a83489a <=( a83488a  and  a83485a );
 a83490a <=( a83489a  and  a83482a );
 a83494a <=( (not A199)  and  (not A166) );
 a83495a <=( (not A167)  and  a83494a );
 a83498a <=( A202  and  (not A200) );
 a83501a <=( (not A265)  and  (not A203) );
 a83502a <=( a83501a  and  a83498a );
 a83503a <=( a83502a  and  a83495a );
 a83507a <=( A268  and  (not A267) );
 a83508a <=( A266  and  a83507a );
 a83511a <=( (not A299)  and  (not A298) );
 a83514a <=( (not A302)  and  A301 );
 a83515a <=( a83514a  and  a83511a );
 a83516a <=( a83515a  and  a83508a );
 a83520a <=( (not A199)  and  (not A166) );
 a83521a <=( (not A167)  and  a83520a );
 a83524a <=( A202  and  (not A200) );
 a83527a <=( (not A265)  and  (not A203) );
 a83528a <=( a83527a  and  a83524a );
 a83529a <=( a83528a  and  a83521a );
 a83533a <=( (not A269)  and  (not A267) );
 a83534a <=( A266  and  a83533a );
 a83537a <=( A299  and  A298 );
 a83540a <=( (not A302)  and  A301 );
 a83541a <=( a83540a  and  a83537a );
 a83542a <=( a83541a  and  a83534a );
 a83546a <=( (not A199)  and  (not A166) );
 a83547a <=( (not A167)  and  a83546a );
 a83550a <=( A202  and  (not A200) );
 a83553a <=( (not A265)  and  (not A203) );
 a83554a <=( a83553a  and  a83550a );
 a83555a <=( a83554a  and  a83547a );
 a83559a <=( (not A269)  and  (not A267) );
 a83560a <=( A266  and  a83559a );
 a83563a <=( (not A299)  and  A298 );
 a83566a <=( A302  and  (not A301) );
 a83567a <=( a83566a  and  a83563a );
 a83568a <=( a83567a  and  a83560a );
 a83572a <=( (not A199)  and  (not A166) );
 a83573a <=( (not A167)  and  a83572a );
 a83576a <=( A202  and  (not A200) );
 a83579a <=( (not A265)  and  (not A203) );
 a83580a <=( a83579a  and  a83576a );
 a83581a <=( a83580a  and  a83573a );
 a83585a <=( (not A269)  and  (not A267) );
 a83586a <=( A266  and  a83585a );
 a83589a <=( A299  and  (not A298) );
 a83592a <=( A302  and  (not A301) );
 a83593a <=( a83592a  and  a83589a );
 a83594a <=( a83593a  and  a83586a );
 a83598a <=( (not A199)  and  (not A166) );
 a83599a <=( (not A167)  and  a83598a );
 a83602a <=( A202  and  (not A200) );
 a83605a <=( (not A265)  and  (not A203) );
 a83606a <=( a83605a  and  a83602a );
 a83607a <=( a83606a  and  a83599a );
 a83611a <=( (not A269)  and  (not A267) );
 a83612a <=( A266  and  a83611a );
 a83615a <=( (not A299)  and  (not A298) );
 a83618a <=( (not A302)  and  A301 );
 a83619a <=( a83618a  and  a83615a );
 a83620a <=( a83619a  and  a83612a );
 a83624a <=( (not A199)  and  (not A166) );
 a83625a <=( (not A167)  and  a83624a );
 a83628a <=( A202  and  (not A200) );
 a83631a <=( A265  and  (not A203) );
 a83632a <=( a83631a  and  a83628a );
 a83633a <=( a83632a  and  a83625a );
 a83637a <=( A268  and  (not A267) );
 a83638a <=( (not A266)  and  a83637a );
 a83641a <=( A299  and  A298 );
 a83644a <=( (not A302)  and  A301 );
 a83645a <=( a83644a  and  a83641a );
 a83646a <=( a83645a  and  a83638a );
 a83650a <=( (not A199)  and  (not A166) );
 a83651a <=( (not A167)  and  a83650a );
 a83654a <=( A202  and  (not A200) );
 a83657a <=( A265  and  (not A203) );
 a83658a <=( a83657a  and  a83654a );
 a83659a <=( a83658a  and  a83651a );
 a83663a <=( A268  and  (not A267) );
 a83664a <=( (not A266)  and  a83663a );
 a83667a <=( (not A299)  and  A298 );
 a83670a <=( A302  and  (not A301) );
 a83671a <=( a83670a  and  a83667a );
 a83672a <=( a83671a  and  a83664a );
 a83676a <=( (not A199)  and  (not A166) );
 a83677a <=( (not A167)  and  a83676a );
 a83680a <=( A202  and  (not A200) );
 a83683a <=( A265  and  (not A203) );
 a83684a <=( a83683a  and  a83680a );
 a83685a <=( a83684a  and  a83677a );
 a83689a <=( A268  and  (not A267) );
 a83690a <=( (not A266)  and  a83689a );
 a83693a <=( A299  and  (not A298) );
 a83696a <=( A302  and  (not A301) );
 a83697a <=( a83696a  and  a83693a );
 a83698a <=( a83697a  and  a83690a );
 a83702a <=( (not A199)  and  (not A166) );
 a83703a <=( (not A167)  and  a83702a );
 a83706a <=( A202  and  (not A200) );
 a83709a <=( A265  and  (not A203) );
 a83710a <=( a83709a  and  a83706a );
 a83711a <=( a83710a  and  a83703a );
 a83715a <=( A268  and  (not A267) );
 a83716a <=( (not A266)  and  a83715a );
 a83719a <=( (not A299)  and  (not A298) );
 a83722a <=( (not A302)  and  A301 );
 a83723a <=( a83722a  and  a83719a );
 a83724a <=( a83723a  and  a83716a );
 a83728a <=( (not A199)  and  (not A166) );
 a83729a <=( (not A167)  and  a83728a );
 a83732a <=( A202  and  (not A200) );
 a83735a <=( A265  and  (not A203) );
 a83736a <=( a83735a  and  a83732a );
 a83737a <=( a83736a  and  a83729a );
 a83741a <=( (not A269)  and  (not A267) );
 a83742a <=( (not A266)  and  a83741a );
 a83745a <=( A299  and  A298 );
 a83748a <=( (not A302)  and  A301 );
 a83749a <=( a83748a  and  a83745a );
 a83750a <=( a83749a  and  a83742a );
 a83754a <=( (not A199)  and  (not A166) );
 a83755a <=( (not A167)  and  a83754a );
 a83758a <=( A202  and  (not A200) );
 a83761a <=( A265  and  (not A203) );
 a83762a <=( a83761a  and  a83758a );
 a83763a <=( a83762a  and  a83755a );
 a83767a <=( (not A269)  and  (not A267) );
 a83768a <=( (not A266)  and  a83767a );
 a83771a <=( (not A299)  and  A298 );
 a83774a <=( A302  and  (not A301) );
 a83775a <=( a83774a  and  a83771a );
 a83776a <=( a83775a  and  a83768a );
 a83780a <=( (not A199)  and  (not A166) );
 a83781a <=( (not A167)  and  a83780a );
 a83784a <=( A202  and  (not A200) );
 a83787a <=( A265  and  (not A203) );
 a83788a <=( a83787a  and  a83784a );
 a83789a <=( a83788a  and  a83781a );
 a83793a <=( (not A269)  and  (not A267) );
 a83794a <=( (not A266)  and  a83793a );
 a83797a <=( A299  and  (not A298) );
 a83800a <=( A302  and  (not A301) );
 a83801a <=( a83800a  and  a83797a );
 a83802a <=( a83801a  and  a83794a );
 a83806a <=( (not A199)  and  (not A166) );
 a83807a <=( (not A167)  and  a83806a );
 a83810a <=( A202  and  (not A200) );
 a83813a <=( A265  and  (not A203) );
 a83814a <=( a83813a  and  a83810a );
 a83815a <=( a83814a  and  a83807a );
 a83819a <=( (not A269)  and  (not A267) );
 a83820a <=( (not A266)  and  a83819a );
 a83823a <=( (not A299)  and  (not A298) );
 a83826a <=( (not A302)  and  A301 );
 a83827a <=( a83826a  and  a83823a );
 a83828a <=( a83827a  and  a83820a );
 a83832a <=( A199  and  (not A167) );
 a83833a <=( (not A168)  and  a83832a );
 a83836a <=( A202  and  A200 );
 a83839a <=( A265  and  (not A203) );
 a83840a <=( a83839a  and  a83836a );
 a83841a <=( a83840a  and  a83833a );
 a83845a <=( (not A268)  and  (not A267) );
 a83846a <=( A266  and  a83845a );
 a83849a <=( A299  and  A298 );
 a83852a <=( (not A302)  and  A301 );
 a83853a <=( a83852a  and  a83849a );
 a83854a <=( a83853a  and  a83846a );
 a83858a <=( A199  and  (not A167) );
 a83859a <=( (not A168)  and  a83858a );
 a83862a <=( A202  and  A200 );
 a83865a <=( A265  and  (not A203) );
 a83866a <=( a83865a  and  a83862a );
 a83867a <=( a83866a  and  a83859a );
 a83871a <=( (not A268)  and  (not A267) );
 a83872a <=( A266  and  a83871a );
 a83875a <=( (not A299)  and  A298 );
 a83878a <=( A302  and  (not A301) );
 a83879a <=( a83878a  and  a83875a );
 a83880a <=( a83879a  and  a83872a );
 a83884a <=( A199  and  (not A167) );
 a83885a <=( (not A168)  and  a83884a );
 a83888a <=( A202  and  A200 );
 a83891a <=( A265  and  (not A203) );
 a83892a <=( a83891a  and  a83888a );
 a83893a <=( a83892a  and  a83885a );
 a83897a <=( (not A268)  and  (not A267) );
 a83898a <=( A266  and  a83897a );
 a83901a <=( A299  and  (not A298) );
 a83904a <=( A302  and  (not A301) );
 a83905a <=( a83904a  and  a83901a );
 a83906a <=( a83905a  and  a83898a );
 a83910a <=( A199  and  (not A167) );
 a83911a <=( (not A168)  and  a83910a );
 a83914a <=( A202  and  A200 );
 a83917a <=( A265  and  (not A203) );
 a83918a <=( a83917a  and  a83914a );
 a83919a <=( a83918a  and  a83911a );
 a83923a <=( (not A268)  and  (not A267) );
 a83924a <=( A266  and  a83923a );
 a83927a <=( (not A299)  and  (not A298) );
 a83930a <=( (not A302)  and  A301 );
 a83931a <=( a83930a  and  a83927a );
 a83932a <=( a83931a  and  a83924a );
 a83936a <=( A199  and  (not A167) );
 a83937a <=( (not A168)  and  a83936a );
 a83940a <=( A202  and  A200 );
 a83943a <=( A265  and  (not A203) );
 a83944a <=( a83943a  and  a83940a );
 a83945a <=( a83944a  and  a83937a );
 a83949a <=( A269  and  (not A267) );
 a83950a <=( A266  and  a83949a );
 a83953a <=( A299  and  A298 );
 a83956a <=( (not A302)  and  A301 );
 a83957a <=( a83956a  and  a83953a );
 a83958a <=( a83957a  and  a83950a );
 a83962a <=( A199  and  (not A167) );
 a83963a <=( (not A168)  and  a83962a );
 a83966a <=( A202  and  A200 );
 a83969a <=( A265  and  (not A203) );
 a83970a <=( a83969a  and  a83966a );
 a83971a <=( a83970a  and  a83963a );
 a83975a <=( A269  and  (not A267) );
 a83976a <=( A266  and  a83975a );
 a83979a <=( (not A299)  and  A298 );
 a83982a <=( A302  and  (not A301) );
 a83983a <=( a83982a  and  a83979a );
 a83984a <=( a83983a  and  a83976a );
 a83988a <=( A199  and  (not A167) );
 a83989a <=( (not A168)  and  a83988a );
 a83992a <=( A202  and  A200 );
 a83995a <=( A265  and  (not A203) );
 a83996a <=( a83995a  and  a83992a );
 a83997a <=( a83996a  and  a83989a );
 a84001a <=( A269  and  (not A267) );
 a84002a <=( A266  and  a84001a );
 a84005a <=( A299  and  (not A298) );
 a84008a <=( A302  and  (not A301) );
 a84009a <=( a84008a  and  a84005a );
 a84010a <=( a84009a  and  a84002a );
 a84014a <=( A199  and  (not A167) );
 a84015a <=( (not A168)  and  a84014a );
 a84018a <=( A202  and  A200 );
 a84021a <=( A265  and  (not A203) );
 a84022a <=( a84021a  and  a84018a );
 a84023a <=( a84022a  and  a84015a );
 a84027a <=( A269  and  (not A267) );
 a84028a <=( A266  and  a84027a );
 a84031a <=( (not A299)  and  (not A298) );
 a84034a <=( (not A302)  and  A301 );
 a84035a <=( a84034a  and  a84031a );
 a84036a <=( a84035a  and  a84028a );
 a84040a <=( A199  and  (not A167) );
 a84041a <=( (not A168)  and  a84040a );
 a84044a <=( A202  and  A200 );
 a84047a <=( (not A265)  and  (not A203) );
 a84048a <=( a84047a  and  a84044a );
 a84049a <=( a84048a  and  a84041a );
 a84053a <=( A268  and  (not A267) );
 a84054a <=( A266  and  a84053a );
 a84057a <=( A299  and  A298 );
 a84060a <=( (not A302)  and  A301 );
 a84061a <=( a84060a  and  a84057a );
 a84062a <=( a84061a  and  a84054a );
 a84066a <=( A199  and  (not A167) );
 a84067a <=( (not A168)  and  a84066a );
 a84070a <=( A202  and  A200 );
 a84073a <=( (not A265)  and  (not A203) );
 a84074a <=( a84073a  and  a84070a );
 a84075a <=( a84074a  and  a84067a );
 a84079a <=( A268  and  (not A267) );
 a84080a <=( A266  and  a84079a );
 a84083a <=( (not A299)  and  A298 );
 a84086a <=( A302  and  (not A301) );
 a84087a <=( a84086a  and  a84083a );
 a84088a <=( a84087a  and  a84080a );
 a84092a <=( A199  and  (not A167) );
 a84093a <=( (not A168)  and  a84092a );
 a84096a <=( A202  and  A200 );
 a84099a <=( (not A265)  and  (not A203) );
 a84100a <=( a84099a  and  a84096a );
 a84101a <=( a84100a  and  a84093a );
 a84105a <=( A268  and  (not A267) );
 a84106a <=( A266  and  a84105a );
 a84109a <=( A299  and  (not A298) );
 a84112a <=( A302  and  (not A301) );
 a84113a <=( a84112a  and  a84109a );
 a84114a <=( a84113a  and  a84106a );
 a84118a <=( A199  and  (not A167) );
 a84119a <=( (not A168)  and  a84118a );
 a84122a <=( A202  and  A200 );
 a84125a <=( (not A265)  and  (not A203) );
 a84126a <=( a84125a  and  a84122a );
 a84127a <=( a84126a  and  a84119a );
 a84131a <=( A268  and  (not A267) );
 a84132a <=( A266  and  a84131a );
 a84135a <=( (not A299)  and  (not A298) );
 a84138a <=( (not A302)  and  A301 );
 a84139a <=( a84138a  and  a84135a );
 a84140a <=( a84139a  and  a84132a );
 a84144a <=( A199  and  (not A167) );
 a84145a <=( (not A168)  and  a84144a );
 a84148a <=( A202  and  A200 );
 a84151a <=( (not A265)  and  (not A203) );
 a84152a <=( a84151a  and  a84148a );
 a84153a <=( a84152a  and  a84145a );
 a84157a <=( (not A269)  and  (not A267) );
 a84158a <=( A266  and  a84157a );
 a84161a <=( A299  and  A298 );
 a84164a <=( (not A302)  and  A301 );
 a84165a <=( a84164a  and  a84161a );
 a84166a <=( a84165a  and  a84158a );
 a84170a <=( A199  and  (not A167) );
 a84171a <=( (not A168)  and  a84170a );
 a84174a <=( A202  and  A200 );
 a84177a <=( (not A265)  and  (not A203) );
 a84178a <=( a84177a  and  a84174a );
 a84179a <=( a84178a  and  a84171a );
 a84183a <=( (not A269)  and  (not A267) );
 a84184a <=( A266  and  a84183a );
 a84187a <=( (not A299)  and  A298 );
 a84190a <=( A302  and  (not A301) );
 a84191a <=( a84190a  and  a84187a );
 a84192a <=( a84191a  and  a84184a );
 a84196a <=( A199  and  (not A167) );
 a84197a <=( (not A168)  and  a84196a );
 a84200a <=( A202  and  A200 );
 a84203a <=( (not A265)  and  (not A203) );
 a84204a <=( a84203a  and  a84200a );
 a84205a <=( a84204a  and  a84197a );
 a84209a <=( (not A269)  and  (not A267) );
 a84210a <=( A266  and  a84209a );
 a84213a <=( A299  and  (not A298) );
 a84216a <=( A302  and  (not A301) );
 a84217a <=( a84216a  and  a84213a );
 a84218a <=( a84217a  and  a84210a );
 a84222a <=( A199  and  (not A167) );
 a84223a <=( (not A168)  and  a84222a );
 a84226a <=( A202  and  A200 );
 a84229a <=( (not A265)  and  (not A203) );
 a84230a <=( a84229a  and  a84226a );
 a84231a <=( a84230a  and  a84223a );
 a84235a <=( (not A269)  and  (not A267) );
 a84236a <=( A266  and  a84235a );
 a84239a <=( (not A299)  and  (not A298) );
 a84242a <=( (not A302)  and  A301 );
 a84243a <=( a84242a  and  a84239a );
 a84244a <=( a84243a  and  a84236a );
 a84248a <=( A199  and  (not A167) );
 a84249a <=( (not A168)  and  a84248a );
 a84252a <=( A202  and  A200 );
 a84255a <=( A265  and  (not A203) );
 a84256a <=( a84255a  and  a84252a );
 a84257a <=( a84256a  and  a84249a );
 a84261a <=( A268  and  (not A267) );
 a84262a <=( (not A266)  and  a84261a );
 a84265a <=( A299  and  A298 );
 a84268a <=( (not A302)  and  A301 );
 a84269a <=( a84268a  and  a84265a );
 a84270a <=( a84269a  and  a84262a );
 a84274a <=( A199  and  (not A167) );
 a84275a <=( (not A168)  and  a84274a );
 a84278a <=( A202  and  A200 );
 a84281a <=( A265  and  (not A203) );
 a84282a <=( a84281a  and  a84278a );
 a84283a <=( a84282a  and  a84275a );
 a84287a <=( A268  and  (not A267) );
 a84288a <=( (not A266)  and  a84287a );
 a84291a <=( (not A299)  and  A298 );
 a84294a <=( A302  and  (not A301) );
 a84295a <=( a84294a  and  a84291a );
 a84296a <=( a84295a  and  a84288a );
 a84300a <=( A199  and  (not A167) );
 a84301a <=( (not A168)  and  a84300a );
 a84304a <=( A202  and  A200 );
 a84307a <=( A265  and  (not A203) );
 a84308a <=( a84307a  and  a84304a );
 a84309a <=( a84308a  and  a84301a );
 a84313a <=( A268  and  (not A267) );
 a84314a <=( (not A266)  and  a84313a );
 a84317a <=( A299  and  (not A298) );
 a84320a <=( A302  and  (not A301) );
 a84321a <=( a84320a  and  a84317a );
 a84322a <=( a84321a  and  a84314a );
 a84326a <=( A199  and  (not A167) );
 a84327a <=( (not A168)  and  a84326a );
 a84330a <=( A202  and  A200 );
 a84333a <=( A265  and  (not A203) );
 a84334a <=( a84333a  and  a84330a );
 a84335a <=( a84334a  and  a84327a );
 a84339a <=( A268  and  (not A267) );
 a84340a <=( (not A266)  and  a84339a );
 a84343a <=( (not A299)  and  (not A298) );
 a84346a <=( (not A302)  and  A301 );
 a84347a <=( a84346a  and  a84343a );
 a84348a <=( a84347a  and  a84340a );
 a84352a <=( A199  and  (not A167) );
 a84353a <=( (not A168)  and  a84352a );
 a84356a <=( A202  and  A200 );
 a84359a <=( A265  and  (not A203) );
 a84360a <=( a84359a  and  a84356a );
 a84361a <=( a84360a  and  a84353a );
 a84365a <=( (not A269)  and  (not A267) );
 a84366a <=( (not A266)  and  a84365a );
 a84369a <=( A299  and  A298 );
 a84372a <=( (not A302)  and  A301 );
 a84373a <=( a84372a  and  a84369a );
 a84374a <=( a84373a  and  a84366a );
 a84378a <=( A199  and  (not A167) );
 a84379a <=( (not A168)  and  a84378a );
 a84382a <=( A202  and  A200 );
 a84385a <=( A265  and  (not A203) );
 a84386a <=( a84385a  and  a84382a );
 a84387a <=( a84386a  and  a84379a );
 a84391a <=( (not A269)  and  (not A267) );
 a84392a <=( (not A266)  and  a84391a );
 a84395a <=( (not A299)  and  A298 );
 a84398a <=( A302  and  (not A301) );
 a84399a <=( a84398a  and  a84395a );
 a84400a <=( a84399a  and  a84392a );
 a84404a <=( A199  and  (not A167) );
 a84405a <=( (not A168)  and  a84404a );
 a84408a <=( A202  and  A200 );
 a84411a <=( A265  and  (not A203) );
 a84412a <=( a84411a  and  a84408a );
 a84413a <=( a84412a  and  a84405a );
 a84417a <=( (not A269)  and  (not A267) );
 a84418a <=( (not A266)  and  a84417a );
 a84421a <=( A299  and  (not A298) );
 a84424a <=( A302  and  (not A301) );
 a84425a <=( a84424a  and  a84421a );
 a84426a <=( a84425a  and  a84418a );
 a84430a <=( A199  and  (not A167) );
 a84431a <=( (not A168)  and  a84430a );
 a84434a <=( A202  and  A200 );
 a84437a <=( A265  and  (not A203) );
 a84438a <=( a84437a  and  a84434a );
 a84439a <=( a84438a  and  a84431a );
 a84443a <=( (not A269)  and  (not A267) );
 a84444a <=( (not A266)  and  a84443a );
 a84447a <=( (not A299)  and  (not A298) );
 a84450a <=( (not A302)  and  A301 );
 a84451a <=( a84450a  and  a84447a );
 a84452a <=( a84451a  and  a84444a );
 a84456a <=( A199  and  (not A167) );
 a84457a <=( (not A168)  and  a84456a );
 a84460a <=( (not A201)  and  A200 );
 a84463a <=( A265  and  (not A202) );
 a84464a <=( a84463a  and  a84460a );
 a84465a <=( a84464a  and  a84457a );
 a84469a <=( (not A269)  and  A268 );
 a84470a <=( A266  and  a84469a );
 a84473a <=( A299  and  A298 );
 a84476a <=( (not A301)  and  (not A300) );
 a84477a <=( a84476a  and  a84473a );
 a84478a <=( a84477a  and  a84470a );
 a84482a <=( A199  and  (not A167) );
 a84483a <=( (not A168)  and  a84482a );
 a84486a <=( (not A201)  and  A200 );
 a84489a <=( A265  and  (not A202) );
 a84490a <=( a84489a  and  a84486a );
 a84491a <=( a84490a  and  a84483a );
 a84495a <=( (not A269)  and  A268 );
 a84496a <=( A266  and  a84495a );
 a84499a <=( A299  and  A298 );
 a84502a <=( A302  and  (not A300) );
 a84503a <=( a84502a  and  a84499a );
 a84504a <=( a84503a  and  a84496a );
 a84508a <=( A199  and  (not A167) );
 a84509a <=( (not A168)  and  a84508a );
 a84512a <=( (not A201)  and  A200 );
 a84515a <=( A265  and  (not A202) );
 a84516a <=( a84515a  and  a84512a );
 a84517a <=( a84516a  and  a84509a );
 a84521a <=( (not A269)  and  A268 );
 a84522a <=( A266  and  a84521a );
 a84525a <=( (not A299)  and  A298 );
 a84528a <=( A301  and  (not A300) );
 a84529a <=( a84528a  and  a84525a );
 a84530a <=( a84529a  and  a84522a );
 a84534a <=( A199  and  (not A167) );
 a84535a <=( (not A168)  and  a84534a );
 a84538a <=( (not A201)  and  A200 );
 a84541a <=( A265  and  (not A202) );
 a84542a <=( a84541a  and  a84538a );
 a84543a <=( a84542a  and  a84535a );
 a84547a <=( (not A269)  and  A268 );
 a84548a <=( A266  and  a84547a );
 a84551a <=( (not A299)  and  A298 );
 a84554a <=( (not A302)  and  (not A300) );
 a84555a <=( a84554a  and  a84551a );
 a84556a <=( a84555a  and  a84548a );
 a84560a <=( A199  and  (not A167) );
 a84561a <=( (not A168)  and  a84560a );
 a84564a <=( (not A201)  and  A200 );
 a84567a <=( A265  and  (not A202) );
 a84568a <=( a84567a  and  a84564a );
 a84569a <=( a84568a  and  a84561a );
 a84573a <=( (not A269)  and  A268 );
 a84574a <=( A266  and  a84573a );
 a84577a <=( A299  and  (not A298) );
 a84580a <=( A301  and  (not A300) );
 a84581a <=( a84580a  and  a84577a );
 a84582a <=( a84581a  and  a84574a );
 a84586a <=( A199  and  (not A167) );
 a84587a <=( (not A168)  and  a84586a );
 a84590a <=( (not A201)  and  A200 );
 a84593a <=( A265  and  (not A202) );
 a84594a <=( a84593a  and  a84590a );
 a84595a <=( a84594a  and  a84587a );
 a84599a <=( (not A269)  and  A268 );
 a84600a <=( A266  and  a84599a );
 a84603a <=( A299  and  (not A298) );
 a84606a <=( (not A302)  and  (not A300) );
 a84607a <=( a84606a  and  a84603a );
 a84608a <=( a84607a  and  a84600a );
 a84612a <=( A199  and  (not A167) );
 a84613a <=( (not A168)  and  a84612a );
 a84616a <=( (not A201)  and  A200 );
 a84619a <=( (not A265)  and  (not A202) );
 a84620a <=( a84619a  and  a84616a );
 a84621a <=( a84620a  and  a84613a );
 a84625a <=( A269  and  (not A268) );
 a84626a <=( A266  and  a84625a );
 a84629a <=( A299  and  A298 );
 a84632a <=( (not A301)  and  (not A300) );
 a84633a <=( a84632a  and  a84629a );
 a84634a <=( a84633a  and  a84626a );
 a84638a <=( A199  and  (not A167) );
 a84639a <=( (not A168)  and  a84638a );
 a84642a <=( (not A201)  and  A200 );
 a84645a <=( (not A265)  and  (not A202) );
 a84646a <=( a84645a  and  a84642a );
 a84647a <=( a84646a  and  a84639a );
 a84651a <=( A269  and  (not A268) );
 a84652a <=( A266  and  a84651a );
 a84655a <=( A299  and  A298 );
 a84658a <=( A302  and  (not A300) );
 a84659a <=( a84658a  and  a84655a );
 a84660a <=( a84659a  and  a84652a );
 a84664a <=( A199  and  (not A167) );
 a84665a <=( (not A168)  and  a84664a );
 a84668a <=( (not A201)  and  A200 );
 a84671a <=( (not A265)  and  (not A202) );
 a84672a <=( a84671a  and  a84668a );
 a84673a <=( a84672a  and  a84665a );
 a84677a <=( A269  and  (not A268) );
 a84678a <=( A266  and  a84677a );
 a84681a <=( (not A299)  and  A298 );
 a84684a <=( A301  and  (not A300) );
 a84685a <=( a84684a  and  a84681a );
 a84686a <=( a84685a  and  a84678a );
 a84690a <=( A199  and  (not A167) );
 a84691a <=( (not A168)  and  a84690a );
 a84694a <=( (not A201)  and  A200 );
 a84697a <=( (not A265)  and  (not A202) );
 a84698a <=( a84697a  and  a84694a );
 a84699a <=( a84698a  and  a84691a );
 a84703a <=( A269  and  (not A268) );
 a84704a <=( A266  and  a84703a );
 a84707a <=( (not A299)  and  A298 );
 a84710a <=( (not A302)  and  (not A300) );
 a84711a <=( a84710a  and  a84707a );
 a84712a <=( a84711a  and  a84704a );
 a84716a <=( A199  and  (not A167) );
 a84717a <=( (not A168)  and  a84716a );
 a84720a <=( (not A201)  and  A200 );
 a84723a <=( (not A265)  and  (not A202) );
 a84724a <=( a84723a  and  a84720a );
 a84725a <=( a84724a  and  a84717a );
 a84729a <=( A269  and  (not A268) );
 a84730a <=( A266  and  a84729a );
 a84733a <=( A299  and  (not A298) );
 a84736a <=( A301  and  (not A300) );
 a84737a <=( a84736a  and  a84733a );
 a84738a <=( a84737a  and  a84730a );
 a84742a <=( A199  and  (not A167) );
 a84743a <=( (not A168)  and  a84742a );
 a84746a <=( (not A201)  and  A200 );
 a84749a <=( (not A265)  and  (not A202) );
 a84750a <=( a84749a  and  a84746a );
 a84751a <=( a84750a  and  a84743a );
 a84755a <=( A269  and  (not A268) );
 a84756a <=( A266  and  a84755a );
 a84759a <=( A299  and  (not A298) );
 a84762a <=( (not A302)  and  (not A300) );
 a84763a <=( a84762a  and  a84759a );
 a84764a <=( a84763a  and  a84756a );
 a84768a <=( A199  and  (not A167) );
 a84769a <=( (not A168)  and  a84768a );
 a84772a <=( (not A201)  and  A200 );
 a84775a <=( A265  and  (not A202) );
 a84776a <=( a84775a  and  a84772a );
 a84777a <=( a84776a  and  a84769a );
 a84781a <=( A269  and  (not A268) );
 a84782a <=( (not A266)  and  a84781a );
 a84785a <=( A299  and  A298 );
 a84788a <=( (not A301)  and  (not A300) );
 a84789a <=( a84788a  and  a84785a );
 a84790a <=( a84789a  and  a84782a );
 a84794a <=( A199  and  (not A167) );
 a84795a <=( (not A168)  and  a84794a );
 a84798a <=( (not A201)  and  A200 );
 a84801a <=( A265  and  (not A202) );
 a84802a <=( a84801a  and  a84798a );
 a84803a <=( a84802a  and  a84795a );
 a84807a <=( A269  and  (not A268) );
 a84808a <=( (not A266)  and  a84807a );
 a84811a <=( A299  and  A298 );
 a84814a <=( A302  and  (not A300) );
 a84815a <=( a84814a  and  a84811a );
 a84816a <=( a84815a  and  a84808a );
 a84820a <=( A199  and  (not A167) );
 a84821a <=( (not A168)  and  a84820a );
 a84824a <=( (not A201)  and  A200 );
 a84827a <=( A265  and  (not A202) );
 a84828a <=( a84827a  and  a84824a );
 a84829a <=( a84828a  and  a84821a );
 a84833a <=( A269  and  (not A268) );
 a84834a <=( (not A266)  and  a84833a );
 a84837a <=( (not A299)  and  A298 );
 a84840a <=( A301  and  (not A300) );
 a84841a <=( a84840a  and  a84837a );
 a84842a <=( a84841a  and  a84834a );
 a84846a <=( A199  and  (not A167) );
 a84847a <=( (not A168)  and  a84846a );
 a84850a <=( (not A201)  and  A200 );
 a84853a <=( A265  and  (not A202) );
 a84854a <=( a84853a  and  a84850a );
 a84855a <=( a84854a  and  a84847a );
 a84859a <=( A269  and  (not A268) );
 a84860a <=( (not A266)  and  a84859a );
 a84863a <=( (not A299)  and  A298 );
 a84866a <=( (not A302)  and  (not A300) );
 a84867a <=( a84866a  and  a84863a );
 a84868a <=( a84867a  and  a84860a );
 a84872a <=( A199  and  (not A167) );
 a84873a <=( (not A168)  and  a84872a );
 a84876a <=( (not A201)  and  A200 );
 a84879a <=( A265  and  (not A202) );
 a84880a <=( a84879a  and  a84876a );
 a84881a <=( a84880a  and  a84873a );
 a84885a <=( A269  and  (not A268) );
 a84886a <=( (not A266)  and  a84885a );
 a84889a <=( A299  and  (not A298) );
 a84892a <=( A301  and  (not A300) );
 a84893a <=( a84892a  and  a84889a );
 a84894a <=( a84893a  and  a84886a );
 a84898a <=( A199  and  (not A167) );
 a84899a <=( (not A168)  and  a84898a );
 a84902a <=( (not A201)  and  A200 );
 a84905a <=( A265  and  (not A202) );
 a84906a <=( a84905a  and  a84902a );
 a84907a <=( a84906a  and  a84899a );
 a84911a <=( A269  and  (not A268) );
 a84912a <=( (not A266)  and  a84911a );
 a84915a <=( A299  and  (not A298) );
 a84918a <=( (not A302)  and  (not A300) );
 a84919a <=( a84918a  and  a84915a );
 a84920a <=( a84919a  and  a84912a );
 a84924a <=( A199  and  (not A167) );
 a84925a <=( (not A168)  and  a84924a );
 a84928a <=( (not A201)  and  A200 );
 a84931a <=( (not A265)  and  (not A202) );
 a84932a <=( a84931a  and  a84928a );
 a84933a <=( a84932a  and  a84925a );
 a84937a <=( (not A269)  and  A268 );
 a84938a <=( (not A266)  and  a84937a );
 a84941a <=( A299  and  A298 );
 a84944a <=( (not A301)  and  (not A300) );
 a84945a <=( a84944a  and  a84941a );
 a84946a <=( a84945a  and  a84938a );
 a84950a <=( A199  and  (not A167) );
 a84951a <=( (not A168)  and  a84950a );
 a84954a <=( (not A201)  and  A200 );
 a84957a <=( (not A265)  and  (not A202) );
 a84958a <=( a84957a  and  a84954a );
 a84959a <=( a84958a  and  a84951a );
 a84963a <=( (not A269)  and  A268 );
 a84964a <=( (not A266)  and  a84963a );
 a84967a <=( A299  and  A298 );
 a84970a <=( A302  and  (not A300) );
 a84971a <=( a84970a  and  a84967a );
 a84972a <=( a84971a  and  a84964a );
 a84976a <=( A199  and  (not A167) );
 a84977a <=( (not A168)  and  a84976a );
 a84980a <=( (not A201)  and  A200 );
 a84983a <=( (not A265)  and  (not A202) );
 a84984a <=( a84983a  and  a84980a );
 a84985a <=( a84984a  and  a84977a );
 a84989a <=( (not A269)  and  A268 );
 a84990a <=( (not A266)  and  a84989a );
 a84993a <=( (not A299)  and  A298 );
 a84996a <=( A301  and  (not A300) );
 a84997a <=( a84996a  and  a84993a );
 a84998a <=( a84997a  and  a84990a );
 a85002a <=( A199  and  (not A167) );
 a85003a <=( (not A168)  and  a85002a );
 a85006a <=( (not A201)  and  A200 );
 a85009a <=( (not A265)  and  (not A202) );
 a85010a <=( a85009a  and  a85006a );
 a85011a <=( a85010a  and  a85003a );
 a85015a <=( (not A269)  and  A268 );
 a85016a <=( (not A266)  and  a85015a );
 a85019a <=( (not A299)  and  A298 );
 a85022a <=( (not A302)  and  (not A300) );
 a85023a <=( a85022a  and  a85019a );
 a85024a <=( a85023a  and  a85016a );
 a85028a <=( A199  and  (not A167) );
 a85029a <=( (not A168)  and  a85028a );
 a85032a <=( (not A201)  and  A200 );
 a85035a <=( (not A265)  and  (not A202) );
 a85036a <=( a85035a  and  a85032a );
 a85037a <=( a85036a  and  a85029a );
 a85041a <=( (not A269)  and  A268 );
 a85042a <=( (not A266)  and  a85041a );
 a85045a <=( A299  and  (not A298) );
 a85048a <=( A301  and  (not A300) );
 a85049a <=( a85048a  and  a85045a );
 a85050a <=( a85049a  and  a85042a );
 a85054a <=( A199  and  (not A167) );
 a85055a <=( (not A168)  and  a85054a );
 a85058a <=( (not A201)  and  A200 );
 a85061a <=( (not A265)  and  (not A202) );
 a85062a <=( a85061a  and  a85058a );
 a85063a <=( a85062a  and  a85055a );
 a85067a <=( (not A269)  and  A268 );
 a85068a <=( (not A266)  and  a85067a );
 a85071a <=( A299  and  (not A298) );
 a85074a <=( (not A302)  and  (not A300) );
 a85075a <=( a85074a  and  a85071a );
 a85076a <=( a85075a  and  a85068a );
 a85080a <=( A199  and  (not A167) );
 a85081a <=( (not A168)  and  a85080a );
 a85084a <=( (not A201)  and  A200 );
 a85087a <=( A265  and  A203 );
 a85088a <=( a85087a  and  a85084a );
 a85089a <=( a85088a  and  a85081a );
 a85093a <=( (not A269)  and  A268 );
 a85094a <=( A266  and  a85093a );
 a85097a <=( A299  and  A298 );
 a85100a <=( (not A301)  and  (not A300) );
 a85101a <=( a85100a  and  a85097a );
 a85102a <=( a85101a  and  a85094a );
 a85106a <=( A199  and  (not A167) );
 a85107a <=( (not A168)  and  a85106a );
 a85110a <=( (not A201)  and  A200 );
 a85113a <=( A265  and  A203 );
 a85114a <=( a85113a  and  a85110a );
 a85115a <=( a85114a  and  a85107a );
 a85119a <=( (not A269)  and  A268 );
 a85120a <=( A266  and  a85119a );
 a85123a <=( A299  and  A298 );
 a85126a <=( A302  and  (not A300) );
 a85127a <=( a85126a  and  a85123a );
 a85128a <=( a85127a  and  a85120a );
 a85132a <=( A199  and  (not A167) );
 a85133a <=( (not A168)  and  a85132a );
 a85136a <=( (not A201)  and  A200 );
 a85139a <=( A265  and  A203 );
 a85140a <=( a85139a  and  a85136a );
 a85141a <=( a85140a  and  a85133a );
 a85145a <=( (not A269)  and  A268 );
 a85146a <=( A266  and  a85145a );
 a85149a <=( (not A299)  and  A298 );
 a85152a <=( A301  and  (not A300) );
 a85153a <=( a85152a  and  a85149a );
 a85154a <=( a85153a  and  a85146a );
 a85158a <=( A199  and  (not A167) );
 a85159a <=( (not A168)  and  a85158a );
 a85162a <=( (not A201)  and  A200 );
 a85165a <=( A265  and  A203 );
 a85166a <=( a85165a  and  a85162a );
 a85167a <=( a85166a  and  a85159a );
 a85171a <=( (not A269)  and  A268 );
 a85172a <=( A266  and  a85171a );
 a85175a <=( (not A299)  and  A298 );
 a85178a <=( (not A302)  and  (not A300) );
 a85179a <=( a85178a  and  a85175a );
 a85180a <=( a85179a  and  a85172a );
 a85184a <=( A199  and  (not A167) );
 a85185a <=( (not A168)  and  a85184a );
 a85188a <=( (not A201)  and  A200 );
 a85191a <=( A265  and  A203 );
 a85192a <=( a85191a  and  a85188a );
 a85193a <=( a85192a  and  a85185a );
 a85197a <=( (not A269)  and  A268 );
 a85198a <=( A266  and  a85197a );
 a85201a <=( A299  and  (not A298) );
 a85204a <=( A301  and  (not A300) );
 a85205a <=( a85204a  and  a85201a );
 a85206a <=( a85205a  and  a85198a );
 a85210a <=( A199  and  (not A167) );
 a85211a <=( (not A168)  and  a85210a );
 a85214a <=( (not A201)  and  A200 );
 a85217a <=( A265  and  A203 );
 a85218a <=( a85217a  and  a85214a );
 a85219a <=( a85218a  and  a85211a );
 a85223a <=( (not A269)  and  A268 );
 a85224a <=( A266  and  a85223a );
 a85227a <=( A299  and  (not A298) );
 a85230a <=( (not A302)  and  (not A300) );
 a85231a <=( a85230a  and  a85227a );
 a85232a <=( a85231a  and  a85224a );
 a85236a <=( A199  and  (not A167) );
 a85237a <=( (not A168)  and  a85236a );
 a85240a <=( (not A201)  and  A200 );
 a85243a <=( (not A265)  and  A203 );
 a85244a <=( a85243a  and  a85240a );
 a85245a <=( a85244a  and  a85237a );
 a85249a <=( A269  and  (not A268) );
 a85250a <=( A266  and  a85249a );
 a85253a <=( A299  and  A298 );
 a85256a <=( (not A301)  and  (not A300) );
 a85257a <=( a85256a  and  a85253a );
 a85258a <=( a85257a  and  a85250a );
 a85262a <=( A199  and  (not A167) );
 a85263a <=( (not A168)  and  a85262a );
 a85266a <=( (not A201)  and  A200 );
 a85269a <=( (not A265)  and  A203 );
 a85270a <=( a85269a  and  a85266a );
 a85271a <=( a85270a  and  a85263a );
 a85275a <=( A269  and  (not A268) );
 a85276a <=( A266  and  a85275a );
 a85279a <=( A299  and  A298 );
 a85282a <=( A302  and  (not A300) );
 a85283a <=( a85282a  and  a85279a );
 a85284a <=( a85283a  and  a85276a );
 a85288a <=( A199  and  (not A167) );
 a85289a <=( (not A168)  and  a85288a );
 a85292a <=( (not A201)  and  A200 );
 a85295a <=( (not A265)  and  A203 );
 a85296a <=( a85295a  and  a85292a );
 a85297a <=( a85296a  and  a85289a );
 a85301a <=( A269  and  (not A268) );
 a85302a <=( A266  and  a85301a );
 a85305a <=( (not A299)  and  A298 );
 a85308a <=( A301  and  (not A300) );
 a85309a <=( a85308a  and  a85305a );
 a85310a <=( a85309a  and  a85302a );
 a85314a <=( A199  and  (not A167) );
 a85315a <=( (not A168)  and  a85314a );
 a85318a <=( (not A201)  and  A200 );
 a85321a <=( (not A265)  and  A203 );
 a85322a <=( a85321a  and  a85318a );
 a85323a <=( a85322a  and  a85315a );
 a85327a <=( A269  and  (not A268) );
 a85328a <=( A266  and  a85327a );
 a85331a <=( (not A299)  and  A298 );
 a85334a <=( (not A302)  and  (not A300) );
 a85335a <=( a85334a  and  a85331a );
 a85336a <=( a85335a  and  a85328a );
 a85340a <=( A199  and  (not A167) );
 a85341a <=( (not A168)  and  a85340a );
 a85344a <=( (not A201)  and  A200 );
 a85347a <=( (not A265)  and  A203 );
 a85348a <=( a85347a  and  a85344a );
 a85349a <=( a85348a  and  a85341a );
 a85353a <=( A269  and  (not A268) );
 a85354a <=( A266  and  a85353a );
 a85357a <=( A299  and  (not A298) );
 a85360a <=( A301  and  (not A300) );
 a85361a <=( a85360a  and  a85357a );
 a85362a <=( a85361a  and  a85354a );
 a85366a <=( A199  and  (not A167) );
 a85367a <=( (not A168)  and  a85366a );
 a85370a <=( (not A201)  and  A200 );
 a85373a <=( (not A265)  and  A203 );
 a85374a <=( a85373a  and  a85370a );
 a85375a <=( a85374a  and  a85367a );
 a85379a <=( A269  and  (not A268) );
 a85380a <=( A266  and  a85379a );
 a85383a <=( A299  and  (not A298) );
 a85386a <=( (not A302)  and  (not A300) );
 a85387a <=( a85386a  and  a85383a );
 a85388a <=( a85387a  and  a85380a );
 a85392a <=( A199  and  (not A167) );
 a85393a <=( (not A168)  and  a85392a );
 a85396a <=( (not A201)  and  A200 );
 a85399a <=( A265  and  A203 );
 a85400a <=( a85399a  and  a85396a );
 a85401a <=( a85400a  and  a85393a );
 a85405a <=( A269  and  (not A268) );
 a85406a <=( (not A266)  and  a85405a );
 a85409a <=( A299  and  A298 );
 a85412a <=( (not A301)  and  (not A300) );
 a85413a <=( a85412a  and  a85409a );
 a85414a <=( a85413a  and  a85406a );
 a85418a <=( A199  and  (not A167) );
 a85419a <=( (not A168)  and  a85418a );
 a85422a <=( (not A201)  and  A200 );
 a85425a <=( A265  and  A203 );
 a85426a <=( a85425a  and  a85422a );
 a85427a <=( a85426a  and  a85419a );
 a85431a <=( A269  and  (not A268) );
 a85432a <=( (not A266)  and  a85431a );
 a85435a <=( A299  and  A298 );
 a85438a <=( A302  and  (not A300) );
 a85439a <=( a85438a  and  a85435a );
 a85440a <=( a85439a  and  a85432a );
 a85444a <=( A199  and  (not A167) );
 a85445a <=( (not A168)  and  a85444a );
 a85448a <=( (not A201)  and  A200 );
 a85451a <=( A265  and  A203 );
 a85452a <=( a85451a  and  a85448a );
 a85453a <=( a85452a  and  a85445a );
 a85457a <=( A269  and  (not A268) );
 a85458a <=( (not A266)  and  a85457a );
 a85461a <=( (not A299)  and  A298 );
 a85464a <=( A301  and  (not A300) );
 a85465a <=( a85464a  and  a85461a );
 a85466a <=( a85465a  and  a85458a );
 a85470a <=( A199  and  (not A167) );
 a85471a <=( (not A168)  and  a85470a );
 a85474a <=( (not A201)  and  A200 );
 a85477a <=( A265  and  A203 );
 a85478a <=( a85477a  and  a85474a );
 a85479a <=( a85478a  and  a85471a );
 a85483a <=( A269  and  (not A268) );
 a85484a <=( (not A266)  and  a85483a );
 a85487a <=( (not A299)  and  A298 );
 a85490a <=( (not A302)  and  (not A300) );
 a85491a <=( a85490a  and  a85487a );
 a85492a <=( a85491a  and  a85484a );
 a85496a <=( A199  and  (not A167) );
 a85497a <=( (not A168)  and  a85496a );
 a85500a <=( (not A201)  and  A200 );
 a85503a <=( A265  and  A203 );
 a85504a <=( a85503a  and  a85500a );
 a85505a <=( a85504a  and  a85497a );
 a85509a <=( A269  and  (not A268) );
 a85510a <=( (not A266)  and  a85509a );
 a85513a <=( A299  and  (not A298) );
 a85516a <=( A301  and  (not A300) );
 a85517a <=( a85516a  and  a85513a );
 a85518a <=( a85517a  and  a85510a );
 a85522a <=( A199  and  (not A167) );
 a85523a <=( (not A168)  and  a85522a );
 a85526a <=( (not A201)  and  A200 );
 a85529a <=( A265  and  A203 );
 a85530a <=( a85529a  and  a85526a );
 a85531a <=( a85530a  and  a85523a );
 a85535a <=( A269  and  (not A268) );
 a85536a <=( (not A266)  and  a85535a );
 a85539a <=( A299  and  (not A298) );
 a85542a <=( (not A302)  and  (not A300) );
 a85543a <=( a85542a  and  a85539a );
 a85544a <=( a85543a  and  a85536a );
 a85548a <=( A199  and  (not A167) );
 a85549a <=( (not A168)  and  a85548a );
 a85552a <=( (not A201)  and  A200 );
 a85555a <=( (not A265)  and  A203 );
 a85556a <=( a85555a  and  a85552a );
 a85557a <=( a85556a  and  a85549a );
 a85561a <=( (not A269)  and  A268 );
 a85562a <=( (not A266)  and  a85561a );
 a85565a <=( A299  and  A298 );
 a85568a <=( (not A301)  and  (not A300) );
 a85569a <=( a85568a  and  a85565a );
 a85570a <=( a85569a  and  a85562a );
 a85574a <=( A199  and  (not A167) );
 a85575a <=( (not A168)  and  a85574a );
 a85578a <=( (not A201)  and  A200 );
 a85581a <=( (not A265)  and  A203 );
 a85582a <=( a85581a  and  a85578a );
 a85583a <=( a85582a  and  a85575a );
 a85587a <=( (not A269)  and  A268 );
 a85588a <=( (not A266)  and  a85587a );
 a85591a <=( A299  and  A298 );
 a85594a <=( A302  and  (not A300) );
 a85595a <=( a85594a  and  a85591a );
 a85596a <=( a85595a  and  a85588a );
 a85600a <=( A199  and  (not A167) );
 a85601a <=( (not A168)  and  a85600a );
 a85604a <=( (not A201)  and  A200 );
 a85607a <=( (not A265)  and  A203 );
 a85608a <=( a85607a  and  a85604a );
 a85609a <=( a85608a  and  a85601a );
 a85613a <=( (not A269)  and  A268 );
 a85614a <=( (not A266)  and  a85613a );
 a85617a <=( (not A299)  and  A298 );
 a85620a <=( A301  and  (not A300) );
 a85621a <=( a85620a  and  a85617a );
 a85622a <=( a85621a  and  a85614a );
 a85626a <=( A199  and  (not A167) );
 a85627a <=( (not A168)  and  a85626a );
 a85630a <=( (not A201)  and  A200 );
 a85633a <=( (not A265)  and  A203 );
 a85634a <=( a85633a  and  a85630a );
 a85635a <=( a85634a  and  a85627a );
 a85639a <=( (not A269)  and  A268 );
 a85640a <=( (not A266)  and  a85639a );
 a85643a <=( (not A299)  and  A298 );
 a85646a <=( (not A302)  and  (not A300) );
 a85647a <=( a85646a  and  a85643a );
 a85648a <=( a85647a  and  a85640a );
 a85652a <=( A199  and  (not A167) );
 a85653a <=( (not A168)  and  a85652a );
 a85656a <=( (not A201)  and  A200 );
 a85659a <=( (not A265)  and  A203 );
 a85660a <=( a85659a  and  a85656a );
 a85661a <=( a85660a  and  a85653a );
 a85665a <=( (not A269)  and  A268 );
 a85666a <=( (not A266)  and  a85665a );
 a85669a <=( A299  and  (not A298) );
 a85672a <=( A301  and  (not A300) );
 a85673a <=( a85672a  and  a85669a );
 a85674a <=( a85673a  and  a85666a );
 a85678a <=( A199  and  (not A167) );
 a85679a <=( (not A168)  and  a85678a );
 a85682a <=( (not A201)  and  A200 );
 a85685a <=( (not A265)  and  A203 );
 a85686a <=( a85685a  and  a85682a );
 a85687a <=( a85686a  and  a85679a );
 a85691a <=( (not A269)  and  A268 );
 a85692a <=( (not A266)  and  a85691a );
 a85695a <=( A299  and  (not A298) );
 a85698a <=( (not A302)  and  (not A300) );
 a85699a <=( a85698a  and  a85695a );
 a85700a <=( a85699a  and  a85692a );
 a85704a <=( (not A199)  and  (not A167) );
 a85705a <=( (not A168)  and  a85704a );
 a85708a <=( (not A202)  and  A200 );
 a85711a <=( A265  and  A203 );
 a85712a <=( a85711a  and  a85708a );
 a85713a <=( a85712a  and  a85705a );
 a85717a <=( (not A268)  and  (not A267) );
 a85718a <=( A266  and  a85717a );
 a85721a <=( A299  and  A298 );
 a85724a <=( (not A302)  and  A301 );
 a85725a <=( a85724a  and  a85721a );
 a85726a <=( a85725a  and  a85718a );
 a85730a <=( (not A199)  and  (not A167) );
 a85731a <=( (not A168)  and  a85730a );
 a85734a <=( (not A202)  and  A200 );
 a85737a <=( A265  and  A203 );
 a85738a <=( a85737a  and  a85734a );
 a85739a <=( a85738a  and  a85731a );
 a85743a <=( (not A268)  and  (not A267) );
 a85744a <=( A266  and  a85743a );
 a85747a <=( (not A299)  and  A298 );
 a85750a <=( A302  and  (not A301) );
 a85751a <=( a85750a  and  a85747a );
 a85752a <=( a85751a  and  a85744a );
 a85756a <=( (not A199)  and  (not A167) );
 a85757a <=( (not A168)  and  a85756a );
 a85760a <=( (not A202)  and  A200 );
 a85763a <=( A265  and  A203 );
 a85764a <=( a85763a  and  a85760a );
 a85765a <=( a85764a  and  a85757a );
 a85769a <=( (not A268)  and  (not A267) );
 a85770a <=( A266  and  a85769a );
 a85773a <=( A299  and  (not A298) );
 a85776a <=( A302  and  (not A301) );
 a85777a <=( a85776a  and  a85773a );
 a85778a <=( a85777a  and  a85770a );
 a85782a <=( (not A199)  and  (not A167) );
 a85783a <=( (not A168)  and  a85782a );
 a85786a <=( (not A202)  and  A200 );
 a85789a <=( A265  and  A203 );
 a85790a <=( a85789a  and  a85786a );
 a85791a <=( a85790a  and  a85783a );
 a85795a <=( (not A268)  and  (not A267) );
 a85796a <=( A266  and  a85795a );
 a85799a <=( (not A299)  and  (not A298) );
 a85802a <=( (not A302)  and  A301 );
 a85803a <=( a85802a  and  a85799a );
 a85804a <=( a85803a  and  a85796a );
 a85808a <=( (not A199)  and  (not A167) );
 a85809a <=( (not A168)  and  a85808a );
 a85812a <=( (not A202)  and  A200 );
 a85815a <=( A265  and  A203 );
 a85816a <=( a85815a  and  a85812a );
 a85817a <=( a85816a  and  a85809a );
 a85821a <=( A269  and  (not A267) );
 a85822a <=( A266  and  a85821a );
 a85825a <=( A299  and  A298 );
 a85828a <=( (not A302)  and  A301 );
 a85829a <=( a85828a  and  a85825a );
 a85830a <=( a85829a  and  a85822a );
 a85834a <=( (not A199)  and  (not A167) );
 a85835a <=( (not A168)  and  a85834a );
 a85838a <=( (not A202)  and  A200 );
 a85841a <=( A265  and  A203 );
 a85842a <=( a85841a  and  a85838a );
 a85843a <=( a85842a  and  a85835a );
 a85847a <=( A269  and  (not A267) );
 a85848a <=( A266  and  a85847a );
 a85851a <=( (not A299)  and  A298 );
 a85854a <=( A302  and  (not A301) );
 a85855a <=( a85854a  and  a85851a );
 a85856a <=( a85855a  and  a85848a );
 a85860a <=( (not A199)  and  (not A167) );
 a85861a <=( (not A168)  and  a85860a );
 a85864a <=( (not A202)  and  A200 );
 a85867a <=( A265  and  A203 );
 a85868a <=( a85867a  and  a85864a );
 a85869a <=( a85868a  and  a85861a );
 a85873a <=( A269  and  (not A267) );
 a85874a <=( A266  and  a85873a );
 a85877a <=( A299  and  (not A298) );
 a85880a <=( A302  and  (not A301) );
 a85881a <=( a85880a  and  a85877a );
 a85882a <=( a85881a  and  a85874a );
 a85886a <=( (not A199)  and  (not A167) );
 a85887a <=( (not A168)  and  a85886a );
 a85890a <=( (not A202)  and  A200 );
 a85893a <=( A265  and  A203 );
 a85894a <=( a85893a  and  a85890a );
 a85895a <=( a85894a  and  a85887a );
 a85899a <=( A269  and  (not A267) );
 a85900a <=( A266  and  a85899a );
 a85903a <=( (not A299)  and  (not A298) );
 a85906a <=( (not A302)  and  A301 );
 a85907a <=( a85906a  and  a85903a );
 a85908a <=( a85907a  and  a85900a );
 a85912a <=( (not A199)  and  (not A167) );
 a85913a <=( (not A168)  and  a85912a );
 a85916a <=( (not A202)  and  A200 );
 a85919a <=( (not A265)  and  A203 );
 a85920a <=( a85919a  and  a85916a );
 a85921a <=( a85920a  and  a85913a );
 a85925a <=( A268  and  (not A267) );
 a85926a <=( A266  and  a85925a );
 a85929a <=( A299  and  A298 );
 a85932a <=( (not A302)  and  A301 );
 a85933a <=( a85932a  and  a85929a );
 a85934a <=( a85933a  and  a85926a );
 a85938a <=( (not A199)  and  (not A167) );
 a85939a <=( (not A168)  and  a85938a );
 a85942a <=( (not A202)  and  A200 );
 a85945a <=( (not A265)  and  A203 );
 a85946a <=( a85945a  and  a85942a );
 a85947a <=( a85946a  and  a85939a );
 a85951a <=( A268  and  (not A267) );
 a85952a <=( A266  and  a85951a );
 a85955a <=( (not A299)  and  A298 );
 a85958a <=( A302  and  (not A301) );
 a85959a <=( a85958a  and  a85955a );
 a85960a <=( a85959a  and  a85952a );
 a85964a <=( (not A199)  and  (not A167) );
 a85965a <=( (not A168)  and  a85964a );
 a85968a <=( (not A202)  and  A200 );
 a85971a <=( (not A265)  and  A203 );
 a85972a <=( a85971a  and  a85968a );
 a85973a <=( a85972a  and  a85965a );
 a85977a <=( A268  and  (not A267) );
 a85978a <=( A266  and  a85977a );
 a85981a <=( A299  and  (not A298) );
 a85984a <=( A302  and  (not A301) );
 a85985a <=( a85984a  and  a85981a );
 a85986a <=( a85985a  and  a85978a );
 a85990a <=( (not A199)  and  (not A167) );
 a85991a <=( (not A168)  and  a85990a );
 a85994a <=( (not A202)  and  A200 );
 a85997a <=( (not A265)  and  A203 );
 a85998a <=( a85997a  and  a85994a );
 a85999a <=( a85998a  and  a85991a );
 a86003a <=( A268  and  (not A267) );
 a86004a <=( A266  and  a86003a );
 a86007a <=( (not A299)  and  (not A298) );
 a86010a <=( (not A302)  and  A301 );
 a86011a <=( a86010a  and  a86007a );
 a86012a <=( a86011a  and  a86004a );
 a86016a <=( (not A199)  and  (not A167) );
 a86017a <=( (not A168)  and  a86016a );
 a86020a <=( (not A202)  and  A200 );
 a86023a <=( (not A265)  and  A203 );
 a86024a <=( a86023a  and  a86020a );
 a86025a <=( a86024a  and  a86017a );
 a86029a <=( (not A269)  and  (not A267) );
 a86030a <=( A266  and  a86029a );
 a86033a <=( A299  and  A298 );
 a86036a <=( (not A302)  and  A301 );
 a86037a <=( a86036a  and  a86033a );
 a86038a <=( a86037a  and  a86030a );
 a86042a <=( (not A199)  and  (not A167) );
 a86043a <=( (not A168)  and  a86042a );
 a86046a <=( (not A202)  and  A200 );
 a86049a <=( (not A265)  and  A203 );
 a86050a <=( a86049a  and  a86046a );
 a86051a <=( a86050a  and  a86043a );
 a86055a <=( (not A269)  and  (not A267) );
 a86056a <=( A266  and  a86055a );
 a86059a <=( (not A299)  and  A298 );
 a86062a <=( A302  and  (not A301) );
 a86063a <=( a86062a  and  a86059a );
 a86064a <=( a86063a  and  a86056a );
 a86068a <=( (not A199)  and  (not A167) );
 a86069a <=( (not A168)  and  a86068a );
 a86072a <=( (not A202)  and  A200 );
 a86075a <=( (not A265)  and  A203 );
 a86076a <=( a86075a  and  a86072a );
 a86077a <=( a86076a  and  a86069a );
 a86081a <=( (not A269)  and  (not A267) );
 a86082a <=( A266  and  a86081a );
 a86085a <=( A299  and  (not A298) );
 a86088a <=( A302  and  (not A301) );
 a86089a <=( a86088a  and  a86085a );
 a86090a <=( a86089a  and  a86082a );
 a86094a <=( (not A199)  and  (not A167) );
 a86095a <=( (not A168)  and  a86094a );
 a86098a <=( (not A202)  and  A200 );
 a86101a <=( (not A265)  and  A203 );
 a86102a <=( a86101a  and  a86098a );
 a86103a <=( a86102a  and  a86095a );
 a86107a <=( (not A269)  and  (not A267) );
 a86108a <=( A266  and  a86107a );
 a86111a <=( (not A299)  and  (not A298) );
 a86114a <=( (not A302)  and  A301 );
 a86115a <=( a86114a  and  a86111a );
 a86116a <=( a86115a  and  a86108a );
 a86120a <=( (not A199)  and  (not A167) );
 a86121a <=( (not A168)  and  a86120a );
 a86124a <=( (not A202)  and  A200 );
 a86127a <=( A265  and  A203 );
 a86128a <=( a86127a  and  a86124a );
 a86129a <=( a86128a  and  a86121a );
 a86133a <=( A268  and  (not A267) );
 a86134a <=( (not A266)  and  a86133a );
 a86137a <=( A299  and  A298 );
 a86140a <=( (not A302)  and  A301 );
 a86141a <=( a86140a  and  a86137a );
 a86142a <=( a86141a  and  a86134a );
 a86146a <=( (not A199)  and  (not A167) );
 a86147a <=( (not A168)  and  a86146a );
 a86150a <=( (not A202)  and  A200 );
 a86153a <=( A265  and  A203 );
 a86154a <=( a86153a  and  a86150a );
 a86155a <=( a86154a  and  a86147a );
 a86159a <=( A268  and  (not A267) );
 a86160a <=( (not A266)  and  a86159a );
 a86163a <=( (not A299)  and  A298 );
 a86166a <=( A302  and  (not A301) );
 a86167a <=( a86166a  and  a86163a );
 a86168a <=( a86167a  and  a86160a );
 a86172a <=( (not A199)  and  (not A167) );
 a86173a <=( (not A168)  and  a86172a );
 a86176a <=( (not A202)  and  A200 );
 a86179a <=( A265  and  A203 );
 a86180a <=( a86179a  and  a86176a );
 a86181a <=( a86180a  and  a86173a );
 a86185a <=( A268  and  (not A267) );
 a86186a <=( (not A266)  and  a86185a );
 a86189a <=( A299  and  (not A298) );
 a86192a <=( A302  and  (not A301) );
 a86193a <=( a86192a  and  a86189a );
 a86194a <=( a86193a  and  a86186a );
 a86198a <=( (not A199)  and  (not A167) );
 a86199a <=( (not A168)  and  a86198a );
 a86202a <=( (not A202)  and  A200 );
 a86205a <=( A265  and  A203 );
 a86206a <=( a86205a  and  a86202a );
 a86207a <=( a86206a  and  a86199a );
 a86211a <=( A268  and  (not A267) );
 a86212a <=( (not A266)  and  a86211a );
 a86215a <=( (not A299)  and  (not A298) );
 a86218a <=( (not A302)  and  A301 );
 a86219a <=( a86218a  and  a86215a );
 a86220a <=( a86219a  and  a86212a );
 a86224a <=( (not A199)  and  (not A167) );
 a86225a <=( (not A168)  and  a86224a );
 a86228a <=( (not A202)  and  A200 );
 a86231a <=( A265  and  A203 );
 a86232a <=( a86231a  and  a86228a );
 a86233a <=( a86232a  and  a86225a );
 a86237a <=( (not A269)  and  (not A267) );
 a86238a <=( (not A266)  and  a86237a );
 a86241a <=( A299  and  A298 );
 a86244a <=( (not A302)  and  A301 );
 a86245a <=( a86244a  and  a86241a );
 a86246a <=( a86245a  and  a86238a );
 a86250a <=( (not A199)  and  (not A167) );
 a86251a <=( (not A168)  and  a86250a );
 a86254a <=( (not A202)  and  A200 );
 a86257a <=( A265  and  A203 );
 a86258a <=( a86257a  and  a86254a );
 a86259a <=( a86258a  and  a86251a );
 a86263a <=( (not A269)  and  (not A267) );
 a86264a <=( (not A266)  and  a86263a );
 a86267a <=( (not A299)  and  A298 );
 a86270a <=( A302  and  (not A301) );
 a86271a <=( a86270a  and  a86267a );
 a86272a <=( a86271a  and  a86264a );
 a86276a <=( (not A199)  and  (not A167) );
 a86277a <=( (not A168)  and  a86276a );
 a86280a <=( (not A202)  and  A200 );
 a86283a <=( A265  and  A203 );
 a86284a <=( a86283a  and  a86280a );
 a86285a <=( a86284a  and  a86277a );
 a86289a <=( (not A269)  and  (not A267) );
 a86290a <=( (not A266)  and  a86289a );
 a86293a <=( A299  and  (not A298) );
 a86296a <=( A302  and  (not A301) );
 a86297a <=( a86296a  and  a86293a );
 a86298a <=( a86297a  and  a86290a );
 a86302a <=( (not A199)  and  (not A167) );
 a86303a <=( (not A168)  and  a86302a );
 a86306a <=( (not A202)  and  A200 );
 a86309a <=( A265  and  A203 );
 a86310a <=( a86309a  and  a86306a );
 a86311a <=( a86310a  and  a86303a );
 a86315a <=( (not A269)  and  (not A267) );
 a86316a <=( (not A266)  and  a86315a );
 a86319a <=( (not A299)  and  (not A298) );
 a86322a <=( (not A302)  and  A301 );
 a86323a <=( a86322a  and  a86319a );
 a86324a <=( a86323a  and  a86316a );
 a86328a <=( (not A199)  and  (not A167) );
 a86329a <=( (not A168)  and  a86328a );
 a86332a <=( (not A201)  and  A200 );
 a86335a <=( A265  and  A202 );
 a86336a <=( a86335a  and  a86332a );
 a86337a <=( a86336a  and  a86329a );
 a86341a <=( (not A269)  and  A268 );
 a86342a <=( A266  and  a86341a );
 a86345a <=( A299  and  A298 );
 a86348a <=( (not A301)  and  (not A300) );
 a86349a <=( a86348a  and  a86345a );
 a86350a <=( a86349a  and  a86342a );
 a86354a <=( (not A199)  and  (not A167) );
 a86355a <=( (not A168)  and  a86354a );
 a86358a <=( (not A201)  and  A200 );
 a86361a <=( A265  and  A202 );
 a86362a <=( a86361a  and  a86358a );
 a86363a <=( a86362a  and  a86355a );
 a86367a <=( (not A269)  and  A268 );
 a86368a <=( A266  and  a86367a );
 a86371a <=( A299  and  A298 );
 a86374a <=( A302  and  (not A300) );
 a86375a <=( a86374a  and  a86371a );
 a86376a <=( a86375a  and  a86368a );
 a86380a <=( (not A199)  and  (not A167) );
 a86381a <=( (not A168)  and  a86380a );
 a86384a <=( (not A201)  and  A200 );
 a86387a <=( A265  and  A202 );
 a86388a <=( a86387a  and  a86384a );
 a86389a <=( a86388a  and  a86381a );
 a86393a <=( (not A269)  and  A268 );
 a86394a <=( A266  and  a86393a );
 a86397a <=( (not A299)  and  A298 );
 a86400a <=( A301  and  (not A300) );
 a86401a <=( a86400a  and  a86397a );
 a86402a <=( a86401a  and  a86394a );
 a86406a <=( (not A199)  and  (not A167) );
 a86407a <=( (not A168)  and  a86406a );
 a86410a <=( (not A201)  and  A200 );
 a86413a <=( A265  and  A202 );
 a86414a <=( a86413a  and  a86410a );
 a86415a <=( a86414a  and  a86407a );
 a86419a <=( (not A269)  and  A268 );
 a86420a <=( A266  and  a86419a );
 a86423a <=( (not A299)  and  A298 );
 a86426a <=( (not A302)  and  (not A300) );
 a86427a <=( a86426a  and  a86423a );
 a86428a <=( a86427a  and  a86420a );
 a86432a <=( (not A199)  and  (not A167) );
 a86433a <=( (not A168)  and  a86432a );
 a86436a <=( (not A201)  and  A200 );
 a86439a <=( A265  and  A202 );
 a86440a <=( a86439a  and  a86436a );
 a86441a <=( a86440a  and  a86433a );
 a86445a <=( (not A269)  and  A268 );
 a86446a <=( A266  and  a86445a );
 a86449a <=( A299  and  (not A298) );
 a86452a <=( A301  and  (not A300) );
 a86453a <=( a86452a  and  a86449a );
 a86454a <=( a86453a  and  a86446a );
 a86458a <=( (not A199)  and  (not A167) );
 a86459a <=( (not A168)  and  a86458a );
 a86462a <=( (not A201)  and  A200 );
 a86465a <=( A265  and  A202 );
 a86466a <=( a86465a  and  a86462a );
 a86467a <=( a86466a  and  a86459a );
 a86471a <=( (not A269)  and  A268 );
 a86472a <=( A266  and  a86471a );
 a86475a <=( A299  and  (not A298) );
 a86478a <=( (not A302)  and  (not A300) );
 a86479a <=( a86478a  and  a86475a );
 a86480a <=( a86479a  and  a86472a );
 a86484a <=( (not A199)  and  (not A167) );
 a86485a <=( (not A168)  and  a86484a );
 a86488a <=( (not A201)  and  A200 );
 a86491a <=( (not A265)  and  A202 );
 a86492a <=( a86491a  and  a86488a );
 a86493a <=( a86492a  and  a86485a );
 a86497a <=( A269  and  (not A268) );
 a86498a <=( A266  and  a86497a );
 a86501a <=( A299  and  A298 );
 a86504a <=( (not A301)  and  (not A300) );
 a86505a <=( a86504a  and  a86501a );
 a86506a <=( a86505a  and  a86498a );
 a86510a <=( (not A199)  and  (not A167) );
 a86511a <=( (not A168)  and  a86510a );
 a86514a <=( (not A201)  and  A200 );
 a86517a <=( (not A265)  and  A202 );
 a86518a <=( a86517a  and  a86514a );
 a86519a <=( a86518a  and  a86511a );
 a86523a <=( A269  and  (not A268) );
 a86524a <=( A266  and  a86523a );
 a86527a <=( A299  and  A298 );
 a86530a <=( A302  and  (not A300) );
 a86531a <=( a86530a  and  a86527a );
 a86532a <=( a86531a  and  a86524a );
 a86536a <=( (not A199)  and  (not A167) );
 a86537a <=( (not A168)  and  a86536a );
 a86540a <=( (not A201)  and  A200 );
 a86543a <=( (not A265)  and  A202 );
 a86544a <=( a86543a  and  a86540a );
 a86545a <=( a86544a  and  a86537a );
 a86549a <=( A269  and  (not A268) );
 a86550a <=( A266  and  a86549a );
 a86553a <=( (not A299)  and  A298 );
 a86556a <=( A301  and  (not A300) );
 a86557a <=( a86556a  and  a86553a );
 a86558a <=( a86557a  and  a86550a );
 a86562a <=( (not A199)  and  (not A167) );
 a86563a <=( (not A168)  and  a86562a );
 a86566a <=( (not A201)  and  A200 );
 a86569a <=( (not A265)  and  A202 );
 a86570a <=( a86569a  and  a86566a );
 a86571a <=( a86570a  and  a86563a );
 a86575a <=( A269  and  (not A268) );
 a86576a <=( A266  and  a86575a );
 a86579a <=( (not A299)  and  A298 );
 a86582a <=( (not A302)  and  (not A300) );
 a86583a <=( a86582a  and  a86579a );
 a86584a <=( a86583a  and  a86576a );
 a86588a <=( (not A199)  and  (not A167) );
 a86589a <=( (not A168)  and  a86588a );
 a86592a <=( (not A201)  and  A200 );
 a86595a <=( (not A265)  and  A202 );
 a86596a <=( a86595a  and  a86592a );
 a86597a <=( a86596a  and  a86589a );
 a86601a <=( A269  and  (not A268) );
 a86602a <=( A266  and  a86601a );
 a86605a <=( A299  and  (not A298) );
 a86608a <=( A301  and  (not A300) );
 a86609a <=( a86608a  and  a86605a );
 a86610a <=( a86609a  and  a86602a );
 a86614a <=( (not A199)  and  (not A167) );
 a86615a <=( (not A168)  and  a86614a );
 a86618a <=( (not A201)  and  A200 );
 a86621a <=( (not A265)  and  A202 );
 a86622a <=( a86621a  and  a86618a );
 a86623a <=( a86622a  and  a86615a );
 a86627a <=( A269  and  (not A268) );
 a86628a <=( A266  and  a86627a );
 a86631a <=( A299  and  (not A298) );
 a86634a <=( (not A302)  and  (not A300) );
 a86635a <=( a86634a  and  a86631a );
 a86636a <=( a86635a  and  a86628a );
 a86640a <=( (not A199)  and  (not A167) );
 a86641a <=( (not A168)  and  a86640a );
 a86644a <=( (not A201)  and  A200 );
 a86647a <=( A265  and  A202 );
 a86648a <=( a86647a  and  a86644a );
 a86649a <=( a86648a  and  a86641a );
 a86653a <=( A269  and  (not A268) );
 a86654a <=( (not A266)  and  a86653a );
 a86657a <=( A299  and  A298 );
 a86660a <=( (not A301)  and  (not A300) );
 a86661a <=( a86660a  and  a86657a );
 a86662a <=( a86661a  and  a86654a );
 a86666a <=( (not A199)  and  (not A167) );
 a86667a <=( (not A168)  and  a86666a );
 a86670a <=( (not A201)  and  A200 );
 a86673a <=( A265  and  A202 );
 a86674a <=( a86673a  and  a86670a );
 a86675a <=( a86674a  and  a86667a );
 a86679a <=( A269  and  (not A268) );
 a86680a <=( (not A266)  and  a86679a );
 a86683a <=( A299  and  A298 );
 a86686a <=( A302  and  (not A300) );
 a86687a <=( a86686a  and  a86683a );
 a86688a <=( a86687a  and  a86680a );
 a86692a <=( (not A199)  and  (not A167) );
 a86693a <=( (not A168)  and  a86692a );
 a86696a <=( (not A201)  and  A200 );
 a86699a <=( A265  and  A202 );
 a86700a <=( a86699a  and  a86696a );
 a86701a <=( a86700a  and  a86693a );
 a86705a <=( A269  and  (not A268) );
 a86706a <=( (not A266)  and  a86705a );
 a86709a <=( (not A299)  and  A298 );
 a86712a <=( A301  and  (not A300) );
 a86713a <=( a86712a  and  a86709a );
 a86714a <=( a86713a  and  a86706a );
 a86718a <=( (not A199)  and  (not A167) );
 a86719a <=( (not A168)  and  a86718a );
 a86722a <=( (not A201)  and  A200 );
 a86725a <=( A265  and  A202 );
 a86726a <=( a86725a  and  a86722a );
 a86727a <=( a86726a  and  a86719a );
 a86731a <=( A269  and  (not A268) );
 a86732a <=( (not A266)  and  a86731a );
 a86735a <=( (not A299)  and  A298 );
 a86738a <=( (not A302)  and  (not A300) );
 a86739a <=( a86738a  and  a86735a );
 a86740a <=( a86739a  and  a86732a );
 a86744a <=( (not A199)  and  (not A167) );
 a86745a <=( (not A168)  and  a86744a );
 a86748a <=( (not A201)  and  A200 );
 a86751a <=( A265  and  A202 );
 a86752a <=( a86751a  and  a86748a );
 a86753a <=( a86752a  and  a86745a );
 a86757a <=( A269  and  (not A268) );
 a86758a <=( (not A266)  and  a86757a );
 a86761a <=( A299  and  (not A298) );
 a86764a <=( A301  and  (not A300) );
 a86765a <=( a86764a  and  a86761a );
 a86766a <=( a86765a  and  a86758a );
 a86770a <=( (not A199)  and  (not A167) );
 a86771a <=( (not A168)  and  a86770a );
 a86774a <=( (not A201)  and  A200 );
 a86777a <=( A265  and  A202 );
 a86778a <=( a86777a  and  a86774a );
 a86779a <=( a86778a  and  a86771a );
 a86783a <=( A269  and  (not A268) );
 a86784a <=( (not A266)  and  a86783a );
 a86787a <=( A299  and  (not A298) );
 a86790a <=( (not A302)  and  (not A300) );
 a86791a <=( a86790a  and  a86787a );
 a86792a <=( a86791a  and  a86784a );
 a86796a <=( (not A199)  and  (not A167) );
 a86797a <=( (not A168)  and  a86796a );
 a86800a <=( (not A201)  and  A200 );
 a86803a <=( (not A265)  and  A202 );
 a86804a <=( a86803a  and  a86800a );
 a86805a <=( a86804a  and  a86797a );
 a86809a <=( (not A269)  and  A268 );
 a86810a <=( (not A266)  and  a86809a );
 a86813a <=( A299  and  A298 );
 a86816a <=( (not A301)  and  (not A300) );
 a86817a <=( a86816a  and  a86813a );
 a86818a <=( a86817a  and  a86810a );
 a86822a <=( (not A199)  and  (not A167) );
 a86823a <=( (not A168)  and  a86822a );
 a86826a <=( (not A201)  and  A200 );
 a86829a <=( (not A265)  and  A202 );
 a86830a <=( a86829a  and  a86826a );
 a86831a <=( a86830a  and  a86823a );
 a86835a <=( (not A269)  and  A268 );
 a86836a <=( (not A266)  and  a86835a );
 a86839a <=( A299  and  A298 );
 a86842a <=( A302  and  (not A300) );
 a86843a <=( a86842a  and  a86839a );
 a86844a <=( a86843a  and  a86836a );
 a86848a <=( (not A199)  and  (not A167) );
 a86849a <=( (not A168)  and  a86848a );
 a86852a <=( (not A201)  and  A200 );
 a86855a <=( (not A265)  and  A202 );
 a86856a <=( a86855a  and  a86852a );
 a86857a <=( a86856a  and  a86849a );
 a86861a <=( (not A269)  and  A268 );
 a86862a <=( (not A266)  and  a86861a );
 a86865a <=( (not A299)  and  A298 );
 a86868a <=( A301  and  (not A300) );
 a86869a <=( a86868a  and  a86865a );
 a86870a <=( a86869a  and  a86862a );
 a86874a <=( (not A199)  and  (not A167) );
 a86875a <=( (not A168)  and  a86874a );
 a86878a <=( (not A201)  and  A200 );
 a86881a <=( (not A265)  and  A202 );
 a86882a <=( a86881a  and  a86878a );
 a86883a <=( a86882a  and  a86875a );
 a86887a <=( (not A269)  and  A268 );
 a86888a <=( (not A266)  and  a86887a );
 a86891a <=( (not A299)  and  A298 );
 a86894a <=( (not A302)  and  (not A300) );
 a86895a <=( a86894a  and  a86891a );
 a86896a <=( a86895a  and  a86888a );
 a86900a <=( (not A199)  and  (not A167) );
 a86901a <=( (not A168)  and  a86900a );
 a86904a <=( (not A201)  and  A200 );
 a86907a <=( (not A265)  and  A202 );
 a86908a <=( a86907a  and  a86904a );
 a86909a <=( a86908a  and  a86901a );
 a86913a <=( (not A269)  and  A268 );
 a86914a <=( (not A266)  and  a86913a );
 a86917a <=( A299  and  (not A298) );
 a86920a <=( A301  and  (not A300) );
 a86921a <=( a86920a  and  a86917a );
 a86922a <=( a86921a  and  a86914a );
 a86926a <=( (not A199)  and  (not A167) );
 a86927a <=( (not A168)  and  a86926a );
 a86930a <=( (not A201)  and  A200 );
 a86933a <=( (not A265)  and  A202 );
 a86934a <=( a86933a  and  a86930a );
 a86935a <=( a86934a  and  a86927a );
 a86939a <=( (not A269)  and  A268 );
 a86940a <=( (not A266)  and  a86939a );
 a86943a <=( A299  and  (not A298) );
 a86946a <=( (not A302)  and  (not A300) );
 a86947a <=( a86946a  and  a86943a );
 a86948a <=( a86947a  and  a86940a );
 a86952a <=( (not A199)  and  (not A167) );
 a86953a <=( (not A168)  and  a86952a );
 a86956a <=( (not A201)  and  A200 );
 a86959a <=( A265  and  (not A203) );
 a86960a <=( a86959a  and  a86956a );
 a86961a <=( a86960a  and  a86953a );
 a86965a <=( (not A269)  and  A268 );
 a86966a <=( A266  and  a86965a );
 a86969a <=( A299  and  A298 );
 a86972a <=( (not A301)  and  (not A300) );
 a86973a <=( a86972a  and  a86969a );
 a86974a <=( a86973a  and  a86966a );
 a86978a <=( (not A199)  and  (not A167) );
 a86979a <=( (not A168)  and  a86978a );
 a86982a <=( (not A201)  and  A200 );
 a86985a <=( A265  and  (not A203) );
 a86986a <=( a86985a  and  a86982a );
 a86987a <=( a86986a  and  a86979a );
 a86991a <=( (not A269)  and  A268 );
 a86992a <=( A266  and  a86991a );
 a86995a <=( A299  and  A298 );
 a86998a <=( A302  and  (not A300) );
 a86999a <=( a86998a  and  a86995a );
 a87000a <=( a86999a  and  a86992a );
 a87004a <=( (not A199)  and  (not A167) );
 a87005a <=( (not A168)  and  a87004a );
 a87008a <=( (not A201)  and  A200 );
 a87011a <=( A265  and  (not A203) );
 a87012a <=( a87011a  and  a87008a );
 a87013a <=( a87012a  and  a87005a );
 a87017a <=( (not A269)  and  A268 );
 a87018a <=( A266  and  a87017a );
 a87021a <=( (not A299)  and  A298 );
 a87024a <=( A301  and  (not A300) );
 a87025a <=( a87024a  and  a87021a );
 a87026a <=( a87025a  and  a87018a );
 a87030a <=( (not A199)  and  (not A167) );
 a87031a <=( (not A168)  and  a87030a );
 a87034a <=( (not A201)  and  A200 );
 a87037a <=( A265  and  (not A203) );
 a87038a <=( a87037a  and  a87034a );
 a87039a <=( a87038a  and  a87031a );
 a87043a <=( (not A269)  and  A268 );
 a87044a <=( A266  and  a87043a );
 a87047a <=( (not A299)  and  A298 );
 a87050a <=( (not A302)  and  (not A300) );
 a87051a <=( a87050a  and  a87047a );
 a87052a <=( a87051a  and  a87044a );
 a87056a <=( (not A199)  and  (not A167) );
 a87057a <=( (not A168)  and  a87056a );
 a87060a <=( (not A201)  and  A200 );
 a87063a <=( A265  and  (not A203) );
 a87064a <=( a87063a  and  a87060a );
 a87065a <=( a87064a  and  a87057a );
 a87069a <=( (not A269)  and  A268 );
 a87070a <=( A266  and  a87069a );
 a87073a <=( A299  and  (not A298) );
 a87076a <=( A301  and  (not A300) );
 a87077a <=( a87076a  and  a87073a );
 a87078a <=( a87077a  and  a87070a );
 a87082a <=( (not A199)  and  (not A167) );
 a87083a <=( (not A168)  and  a87082a );
 a87086a <=( (not A201)  and  A200 );
 a87089a <=( A265  and  (not A203) );
 a87090a <=( a87089a  and  a87086a );
 a87091a <=( a87090a  and  a87083a );
 a87095a <=( (not A269)  and  A268 );
 a87096a <=( A266  and  a87095a );
 a87099a <=( A299  and  (not A298) );
 a87102a <=( (not A302)  and  (not A300) );
 a87103a <=( a87102a  and  a87099a );
 a87104a <=( a87103a  and  a87096a );
 a87108a <=( (not A199)  and  (not A167) );
 a87109a <=( (not A168)  and  a87108a );
 a87112a <=( (not A201)  and  A200 );
 a87115a <=( (not A265)  and  (not A203) );
 a87116a <=( a87115a  and  a87112a );
 a87117a <=( a87116a  and  a87109a );
 a87121a <=( A269  and  (not A268) );
 a87122a <=( A266  and  a87121a );
 a87125a <=( A299  and  A298 );
 a87128a <=( (not A301)  and  (not A300) );
 a87129a <=( a87128a  and  a87125a );
 a87130a <=( a87129a  and  a87122a );
 a87134a <=( (not A199)  and  (not A167) );
 a87135a <=( (not A168)  and  a87134a );
 a87138a <=( (not A201)  and  A200 );
 a87141a <=( (not A265)  and  (not A203) );
 a87142a <=( a87141a  and  a87138a );
 a87143a <=( a87142a  and  a87135a );
 a87147a <=( A269  and  (not A268) );
 a87148a <=( A266  and  a87147a );
 a87151a <=( A299  and  A298 );
 a87154a <=( A302  and  (not A300) );
 a87155a <=( a87154a  and  a87151a );
 a87156a <=( a87155a  and  a87148a );
 a87160a <=( (not A199)  and  (not A167) );
 a87161a <=( (not A168)  and  a87160a );
 a87164a <=( (not A201)  and  A200 );
 a87167a <=( (not A265)  and  (not A203) );
 a87168a <=( a87167a  and  a87164a );
 a87169a <=( a87168a  and  a87161a );
 a87173a <=( A269  and  (not A268) );
 a87174a <=( A266  and  a87173a );
 a87177a <=( (not A299)  and  A298 );
 a87180a <=( A301  and  (not A300) );
 a87181a <=( a87180a  and  a87177a );
 a87182a <=( a87181a  and  a87174a );
 a87186a <=( (not A199)  and  (not A167) );
 a87187a <=( (not A168)  and  a87186a );
 a87190a <=( (not A201)  and  A200 );
 a87193a <=( (not A265)  and  (not A203) );
 a87194a <=( a87193a  and  a87190a );
 a87195a <=( a87194a  and  a87187a );
 a87199a <=( A269  and  (not A268) );
 a87200a <=( A266  and  a87199a );
 a87203a <=( (not A299)  and  A298 );
 a87206a <=( (not A302)  and  (not A300) );
 a87207a <=( a87206a  and  a87203a );
 a87208a <=( a87207a  and  a87200a );
 a87212a <=( (not A199)  and  (not A167) );
 a87213a <=( (not A168)  and  a87212a );
 a87216a <=( (not A201)  and  A200 );
 a87219a <=( (not A265)  and  (not A203) );
 a87220a <=( a87219a  and  a87216a );
 a87221a <=( a87220a  and  a87213a );
 a87225a <=( A269  and  (not A268) );
 a87226a <=( A266  and  a87225a );
 a87229a <=( A299  and  (not A298) );
 a87232a <=( A301  and  (not A300) );
 a87233a <=( a87232a  and  a87229a );
 a87234a <=( a87233a  and  a87226a );
 a87238a <=( (not A199)  and  (not A167) );
 a87239a <=( (not A168)  and  a87238a );
 a87242a <=( (not A201)  and  A200 );
 a87245a <=( (not A265)  and  (not A203) );
 a87246a <=( a87245a  and  a87242a );
 a87247a <=( a87246a  and  a87239a );
 a87251a <=( A269  and  (not A268) );
 a87252a <=( A266  and  a87251a );
 a87255a <=( A299  and  (not A298) );
 a87258a <=( (not A302)  and  (not A300) );
 a87259a <=( a87258a  and  a87255a );
 a87260a <=( a87259a  and  a87252a );
 a87264a <=( (not A199)  and  (not A167) );
 a87265a <=( (not A168)  and  a87264a );
 a87268a <=( (not A201)  and  A200 );
 a87271a <=( A265  and  (not A203) );
 a87272a <=( a87271a  and  a87268a );
 a87273a <=( a87272a  and  a87265a );
 a87277a <=( A269  and  (not A268) );
 a87278a <=( (not A266)  and  a87277a );
 a87281a <=( A299  and  A298 );
 a87284a <=( (not A301)  and  (not A300) );
 a87285a <=( a87284a  and  a87281a );
 a87286a <=( a87285a  and  a87278a );
 a87290a <=( (not A199)  and  (not A167) );
 a87291a <=( (not A168)  and  a87290a );
 a87294a <=( (not A201)  and  A200 );
 a87297a <=( A265  and  (not A203) );
 a87298a <=( a87297a  and  a87294a );
 a87299a <=( a87298a  and  a87291a );
 a87303a <=( A269  and  (not A268) );
 a87304a <=( (not A266)  and  a87303a );
 a87307a <=( A299  and  A298 );
 a87310a <=( A302  and  (not A300) );
 a87311a <=( a87310a  and  a87307a );
 a87312a <=( a87311a  and  a87304a );
 a87316a <=( (not A199)  and  (not A167) );
 a87317a <=( (not A168)  and  a87316a );
 a87320a <=( (not A201)  and  A200 );
 a87323a <=( A265  and  (not A203) );
 a87324a <=( a87323a  and  a87320a );
 a87325a <=( a87324a  and  a87317a );
 a87329a <=( A269  and  (not A268) );
 a87330a <=( (not A266)  and  a87329a );
 a87333a <=( (not A299)  and  A298 );
 a87336a <=( A301  and  (not A300) );
 a87337a <=( a87336a  and  a87333a );
 a87338a <=( a87337a  and  a87330a );
 a87342a <=( (not A199)  and  (not A167) );
 a87343a <=( (not A168)  and  a87342a );
 a87346a <=( (not A201)  and  A200 );
 a87349a <=( A265  and  (not A203) );
 a87350a <=( a87349a  and  a87346a );
 a87351a <=( a87350a  and  a87343a );
 a87355a <=( A269  and  (not A268) );
 a87356a <=( (not A266)  and  a87355a );
 a87359a <=( (not A299)  and  A298 );
 a87362a <=( (not A302)  and  (not A300) );
 a87363a <=( a87362a  and  a87359a );
 a87364a <=( a87363a  and  a87356a );
 a87368a <=( (not A199)  and  (not A167) );
 a87369a <=( (not A168)  and  a87368a );
 a87372a <=( (not A201)  and  A200 );
 a87375a <=( A265  and  (not A203) );
 a87376a <=( a87375a  and  a87372a );
 a87377a <=( a87376a  and  a87369a );
 a87381a <=( A269  and  (not A268) );
 a87382a <=( (not A266)  and  a87381a );
 a87385a <=( A299  and  (not A298) );
 a87388a <=( A301  and  (not A300) );
 a87389a <=( a87388a  and  a87385a );
 a87390a <=( a87389a  and  a87382a );
 a87394a <=( (not A199)  and  (not A167) );
 a87395a <=( (not A168)  and  a87394a );
 a87398a <=( (not A201)  and  A200 );
 a87401a <=( A265  and  (not A203) );
 a87402a <=( a87401a  and  a87398a );
 a87403a <=( a87402a  and  a87395a );
 a87407a <=( A269  and  (not A268) );
 a87408a <=( (not A266)  and  a87407a );
 a87411a <=( A299  and  (not A298) );
 a87414a <=( (not A302)  and  (not A300) );
 a87415a <=( a87414a  and  a87411a );
 a87416a <=( a87415a  and  a87408a );
 a87420a <=( (not A199)  and  (not A167) );
 a87421a <=( (not A168)  and  a87420a );
 a87424a <=( (not A201)  and  A200 );
 a87427a <=( (not A265)  and  (not A203) );
 a87428a <=( a87427a  and  a87424a );
 a87429a <=( a87428a  and  a87421a );
 a87433a <=( (not A269)  and  A268 );
 a87434a <=( (not A266)  and  a87433a );
 a87437a <=( A299  and  A298 );
 a87440a <=( (not A301)  and  (not A300) );
 a87441a <=( a87440a  and  a87437a );
 a87442a <=( a87441a  and  a87434a );
 a87446a <=( (not A199)  and  (not A167) );
 a87447a <=( (not A168)  and  a87446a );
 a87450a <=( (not A201)  and  A200 );
 a87453a <=( (not A265)  and  (not A203) );
 a87454a <=( a87453a  and  a87450a );
 a87455a <=( a87454a  and  a87447a );
 a87459a <=( (not A269)  and  A268 );
 a87460a <=( (not A266)  and  a87459a );
 a87463a <=( A299  and  A298 );
 a87466a <=( A302  and  (not A300) );
 a87467a <=( a87466a  and  a87463a );
 a87468a <=( a87467a  and  a87460a );
 a87472a <=( (not A199)  and  (not A167) );
 a87473a <=( (not A168)  and  a87472a );
 a87476a <=( (not A201)  and  A200 );
 a87479a <=( (not A265)  and  (not A203) );
 a87480a <=( a87479a  and  a87476a );
 a87481a <=( a87480a  and  a87473a );
 a87485a <=( (not A269)  and  A268 );
 a87486a <=( (not A266)  and  a87485a );
 a87489a <=( (not A299)  and  A298 );
 a87492a <=( A301  and  (not A300) );
 a87493a <=( a87492a  and  a87489a );
 a87494a <=( a87493a  and  a87486a );
 a87498a <=( (not A199)  and  (not A167) );
 a87499a <=( (not A168)  and  a87498a );
 a87502a <=( (not A201)  and  A200 );
 a87505a <=( (not A265)  and  (not A203) );
 a87506a <=( a87505a  and  a87502a );
 a87507a <=( a87506a  and  a87499a );
 a87511a <=( (not A269)  and  A268 );
 a87512a <=( (not A266)  and  a87511a );
 a87515a <=( (not A299)  and  A298 );
 a87518a <=( (not A302)  and  (not A300) );
 a87519a <=( a87518a  and  a87515a );
 a87520a <=( a87519a  and  a87512a );
 a87524a <=( (not A199)  and  (not A167) );
 a87525a <=( (not A168)  and  a87524a );
 a87528a <=( (not A201)  and  A200 );
 a87531a <=( (not A265)  and  (not A203) );
 a87532a <=( a87531a  and  a87528a );
 a87533a <=( a87532a  and  a87525a );
 a87537a <=( (not A269)  and  A268 );
 a87538a <=( (not A266)  and  a87537a );
 a87541a <=( A299  and  (not A298) );
 a87544a <=( A301  and  (not A300) );
 a87545a <=( a87544a  and  a87541a );
 a87546a <=( a87545a  and  a87538a );
 a87550a <=( (not A199)  and  (not A167) );
 a87551a <=( (not A168)  and  a87550a );
 a87554a <=( (not A201)  and  A200 );
 a87557a <=( (not A265)  and  (not A203) );
 a87558a <=( a87557a  and  a87554a );
 a87559a <=( a87558a  and  a87551a );
 a87563a <=( (not A269)  and  A268 );
 a87564a <=( (not A266)  and  a87563a );
 a87567a <=( A299  and  (not A298) );
 a87570a <=( (not A302)  and  (not A300) );
 a87571a <=( a87570a  and  a87567a );
 a87572a <=( a87571a  and  a87564a );
 a87576a <=( A199  and  (not A167) );
 a87577a <=( (not A168)  and  a87576a );
 a87580a <=( (not A202)  and  (not A200) );
 a87583a <=( A265  and  A203 );
 a87584a <=( a87583a  and  a87580a );
 a87585a <=( a87584a  and  a87577a );
 a87589a <=( (not A268)  and  (not A267) );
 a87590a <=( A266  and  a87589a );
 a87593a <=( A299  and  A298 );
 a87596a <=( (not A302)  and  A301 );
 a87597a <=( a87596a  and  a87593a );
 a87598a <=( a87597a  and  a87590a );
 a87602a <=( A199  and  (not A167) );
 a87603a <=( (not A168)  and  a87602a );
 a87606a <=( (not A202)  and  (not A200) );
 a87609a <=( A265  and  A203 );
 a87610a <=( a87609a  and  a87606a );
 a87611a <=( a87610a  and  a87603a );
 a87615a <=( (not A268)  and  (not A267) );
 a87616a <=( A266  and  a87615a );
 a87619a <=( (not A299)  and  A298 );
 a87622a <=( A302  and  (not A301) );
 a87623a <=( a87622a  and  a87619a );
 a87624a <=( a87623a  and  a87616a );
 a87628a <=( A199  and  (not A167) );
 a87629a <=( (not A168)  and  a87628a );
 a87632a <=( (not A202)  and  (not A200) );
 a87635a <=( A265  and  A203 );
 a87636a <=( a87635a  and  a87632a );
 a87637a <=( a87636a  and  a87629a );
 a87641a <=( (not A268)  and  (not A267) );
 a87642a <=( A266  and  a87641a );
 a87645a <=( A299  and  (not A298) );
 a87648a <=( A302  and  (not A301) );
 a87649a <=( a87648a  and  a87645a );
 a87650a <=( a87649a  and  a87642a );
 a87654a <=( A199  and  (not A167) );
 a87655a <=( (not A168)  and  a87654a );
 a87658a <=( (not A202)  and  (not A200) );
 a87661a <=( A265  and  A203 );
 a87662a <=( a87661a  and  a87658a );
 a87663a <=( a87662a  and  a87655a );
 a87667a <=( (not A268)  and  (not A267) );
 a87668a <=( A266  and  a87667a );
 a87671a <=( (not A299)  and  (not A298) );
 a87674a <=( (not A302)  and  A301 );
 a87675a <=( a87674a  and  a87671a );
 a87676a <=( a87675a  and  a87668a );
 a87680a <=( A199  and  (not A167) );
 a87681a <=( (not A168)  and  a87680a );
 a87684a <=( (not A202)  and  (not A200) );
 a87687a <=( A265  and  A203 );
 a87688a <=( a87687a  and  a87684a );
 a87689a <=( a87688a  and  a87681a );
 a87693a <=( A269  and  (not A267) );
 a87694a <=( A266  and  a87693a );
 a87697a <=( A299  and  A298 );
 a87700a <=( (not A302)  and  A301 );
 a87701a <=( a87700a  and  a87697a );
 a87702a <=( a87701a  and  a87694a );
 a87706a <=( A199  and  (not A167) );
 a87707a <=( (not A168)  and  a87706a );
 a87710a <=( (not A202)  and  (not A200) );
 a87713a <=( A265  and  A203 );
 a87714a <=( a87713a  and  a87710a );
 a87715a <=( a87714a  and  a87707a );
 a87719a <=( A269  and  (not A267) );
 a87720a <=( A266  and  a87719a );
 a87723a <=( (not A299)  and  A298 );
 a87726a <=( A302  and  (not A301) );
 a87727a <=( a87726a  and  a87723a );
 a87728a <=( a87727a  and  a87720a );
 a87732a <=( A199  and  (not A167) );
 a87733a <=( (not A168)  and  a87732a );
 a87736a <=( (not A202)  and  (not A200) );
 a87739a <=( A265  and  A203 );
 a87740a <=( a87739a  and  a87736a );
 a87741a <=( a87740a  and  a87733a );
 a87745a <=( A269  and  (not A267) );
 a87746a <=( A266  and  a87745a );
 a87749a <=( A299  and  (not A298) );
 a87752a <=( A302  and  (not A301) );
 a87753a <=( a87752a  and  a87749a );
 a87754a <=( a87753a  and  a87746a );
 a87758a <=( A199  and  (not A167) );
 a87759a <=( (not A168)  and  a87758a );
 a87762a <=( (not A202)  and  (not A200) );
 a87765a <=( A265  and  A203 );
 a87766a <=( a87765a  and  a87762a );
 a87767a <=( a87766a  and  a87759a );
 a87771a <=( A269  and  (not A267) );
 a87772a <=( A266  and  a87771a );
 a87775a <=( (not A299)  and  (not A298) );
 a87778a <=( (not A302)  and  A301 );
 a87779a <=( a87778a  and  a87775a );
 a87780a <=( a87779a  and  a87772a );
 a87784a <=( A199  and  (not A167) );
 a87785a <=( (not A168)  and  a87784a );
 a87788a <=( (not A202)  and  (not A200) );
 a87791a <=( (not A265)  and  A203 );
 a87792a <=( a87791a  and  a87788a );
 a87793a <=( a87792a  and  a87785a );
 a87797a <=( A268  and  (not A267) );
 a87798a <=( A266  and  a87797a );
 a87801a <=( A299  and  A298 );
 a87804a <=( (not A302)  and  A301 );
 a87805a <=( a87804a  and  a87801a );
 a87806a <=( a87805a  and  a87798a );
 a87810a <=( A199  and  (not A167) );
 a87811a <=( (not A168)  and  a87810a );
 a87814a <=( (not A202)  and  (not A200) );
 a87817a <=( (not A265)  and  A203 );
 a87818a <=( a87817a  and  a87814a );
 a87819a <=( a87818a  and  a87811a );
 a87823a <=( A268  and  (not A267) );
 a87824a <=( A266  and  a87823a );
 a87827a <=( (not A299)  and  A298 );
 a87830a <=( A302  and  (not A301) );
 a87831a <=( a87830a  and  a87827a );
 a87832a <=( a87831a  and  a87824a );
 a87836a <=( A199  and  (not A167) );
 a87837a <=( (not A168)  and  a87836a );
 a87840a <=( (not A202)  and  (not A200) );
 a87843a <=( (not A265)  and  A203 );
 a87844a <=( a87843a  and  a87840a );
 a87845a <=( a87844a  and  a87837a );
 a87849a <=( A268  and  (not A267) );
 a87850a <=( A266  and  a87849a );
 a87853a <=( A299  and  (not A298) );
 a87856a <=( A302  and  (not A301) );
 a87857a <=( a87856a  and  a87853a );
 a87858a <=( a87857a  and  a87850a );
 a87862a <=( A199  and  (not A167) );
 a87863a <=( (not A168)  and  a87862a );
 a87866a <=( (not A202)  and  (not A200) );
 a87869a <=( (not A265)  and  A203 );
 a87870a <=( a87869a  and  a87866a );
 a87871a <=( a87870a  and  a87863a );
 a87875a <=( A268  and  (not A267) );
 a87876a <=( A266  and  a87875a );
 a87879a <=( (not A299)  and  (not A298) );
 a87882a <=( (not A302)  and  A301 );
 a87883a <=( a87882a  and  a87879a );
 a87884a <=( a87883a  and  a87876a );
 a87888a <=( A199  and  (not A167) );
 a87889a <=( (not A168)  and  a87888a );
 a87892a <=( (not A202)  and  (not A200) );
 a87895a <=( (not A265)  and  A203 );
 a87896a <=( a87895a  and  a87892a );
 a87897a <=( a87896a  and  a87889a );
 a87901a <=( (not A269)  and  (not A267) );
 a87902a <=( A266  and  a87901a );
 a87905a <=( A299  and  A298 );
 a87908a <=( (not A302)  and  A301 );
 a87909a <=( a87908a  and  a87905a );
 a87910a <=( a87909a  and  a87902a );
 a87914a <=( A199  and  (not A167) );
 a87915a <=( (not A168)  and  a87914a );
 a87918a <=( (not A202)  and  (not A200) );
 a87921a <=( (not A265)  and  A203 );
 a87922a <=( a87921a  and  a87918a );
 a87923a <=( a87922a  and  a87915a );
 a87927a <=( (not A269)  and  (not A267) );
 a87928a <=( A266  and  a87927a );
 a87931a <=( (not A299)  and  A298 );
 a87934a <=( A302  and  (not A301) );
 a87935a <=( a87934a  and  a87931a );
 a87936a <=( a87935a  and  a87928a );
 a87940a <=( A199  and  (not A167) );
 a87941a <=( (not A168)  and  a87940a );
 a87944a <=( (not A202)  and  (not A200) );
 a87947a <=( (not A265)  and  A203 );
 a87948a <=( a87947a  and  a87944a );
 a87949a <=( a87948a  and  a87941a );
 a87953a <=( (not A269)  and  (not A267) );
 a87954a <=( A266  and  a87953a );
 a87957a <=( A299  and  (not A298) );
 a87960a <=( A302  and  (not A301) );
 a87961a <=( a87960a  and  a87957a );
 a87962a <=( a87961a  and  a87954a );
 a87966a <=( A199  and  (not A167) );
 a87967a <=( (not A168)  and  a87966a );
 a87970a <=( (not A202)  and  (not A200) );
 a87973a <=( (not A265)  and  A203 );
 a87974a <=( a87973a  and  a87970a );
 a87975a <=( a87974a  and  a87967a );
 a87979a <=( (not A269)  and  (not A267) );
 a87980a <=( A266  and  a87979a );
 a87983a <=( (not A299)  and  (not A298) );
 a87986a <=( (not A302)  and  A301 );
 a87987a <=( a87986a  and  a87983a );
 a87988a <=( a87987a  and  a87980a );
 a87992a <=( A199  and  (not A167) );
 a87993a <=( (not A168)  and  a87992a );
 a87996a <=( (not A202)  and  (not A200) );
 a87999a <=( A265  and  A203 );
 a88000a <=( a87999a  and  a87996a );
 a88001a <=( a88000a  and  a87993a );
 a88005a <=( A268  and  (not A267) );
 a88006a <=( (not A266)  and  a88005a );
 a88009a <=( A299  and  A298 );
 a88012a <=( (not A302)  and  A301 );
 a88013a <=( a88012a  and  a88009a );
 a88014a <=( a88013a  and  a88006a );
 a88018a <=( A199  and  (not A167) );
 a88019a <=( (not A168)  and  a88018a );
 a88022a <=( (not A202)  and  (not A200) );
 a88025a <=( A265  and  A203 );
 a88026a <=( a88025a  and  a88022a );
 a88027a <=( a88026a  and  a88019a );
 a88031a <=( A268  and  (not A267) );
 a88032a <=( (not A266)  and  a88031a );
 a88035a <=( (not A299)  and  A298 );
 a88038a <=( A302  and  (not A301) );
 a88039a <=( a88038a  and  a88035a );
 a88040a <=( a88039a  and  a88032a );
 a88044a <=( A199  and  (not A167) );
 a88045a <=( (not A168)  and  a88044a );
 a88048a <=( (not A202)  and  (not A200) );
 a88051a <=( A265  and  A203 );
 a88052a <=( a88051a  and  a88048a );
 a88053a <=( a88052a  and  a88045a );
 a88057a <=( A268  and  (not A267) );
 a88058a <=( (not A266)  and  a88057a );
 a88061a <=( A299  and  (not A298) );
 a88064a <=( A302  and  (not A301) );
 a88065a <=( a88064a  and  a88061a );
 a88066a <=( a88065a  and  a88058a );
 a88070a <=( A199  and  (not A167) );
 a88071a <=( (not A168)  and  a88070a );
 a88074a <=( (not A202)  and  (not A200) );
 a88077a <=( A265  and  A203 );
 a88078a <=( a88077a  and  a88074a );
 a88079a <=( a88078a  and  a88071a );
 a88083a <=( A268  and  (not A267) );
 a88084a <=( (not A266)  and  a88083a );
 a88087a <=( (not A299)  and  (not A298) );
 a88090a <=( (not A302)  and  A301 );
 a88091a <=( a88090a  and  a88087a );
 a88092a <=( a88091a  and  a88084a );
 a88096a <=( A199  and  (not A167) );
 a88097a <=( (not A168)  and  a88096a );
 a88100a <=( (not A202)  and  (not A200) );
 a88103a <=( A265  and  A203 );
 a88104a <=( a88103a  and  a88100a );
 a88105a <=( a88104a  and  a88097a );
 a88109a <=( (not A269)  and  (not A267) );
 a88110a <=( (not A266)  and  a88109a );
 a88113a <=( A299  and  A298 );
 a88116a <=( (not A302)  and  A301 );
 a88117a <=( a88116a  and  a88113a );
 a88118a <=( a88117a  and  a88110a );
 a88122a <=( A199  and  (not A167) );
 a88123a <=( (not A168)  and  a88122a );
 a88126a <=( (not A202)  and  (not A200) );
 a88129a <=( A265  and  A203 );
 a88130a <=( a88129a  and  a88126a );
 a88131a <=( a88130a  and  a88123a );
 a88135a <=( (not A269)  and  (not A267) );
 a88136a <=( (not A266)  and  a88135a );
 a88139a <=( (not A299)  and  A298 );
 a88142a <=( A302  and  (not A301) );
 a88143a <=( a88142a  and  a88139a );
 a88144a <=( a88143a  and  a88136a );
 a88148a <=( A199  and  (not A167) );
 a88149a <=( (not A168)  and  a88148a );
 a88152a <=( (not A202)  and  (not A200) );
 a88155a <=( A265  and  A203 );
 a88156a <=( a88155a  and  a88152a );
 a88157a <=( a88156a  and  a88149a );
 a88161a <=( (not A269)  and  (not A267) );
 a88162a <=( (not A266)  and  a88161a );
 a88165a <=( A299  and  (not A298) );
 a88168a <=( A302  and  (not A301) );
 a88169a <=( a88168a  and  a88165a );
 a88170a <=( a88169a  and  a88162a );
 a88174a <=( A199  and  (not A167) );
 a88175a <=( (not A168)  and  a88174a );
 a88178a <=( (not A202)  and  (not A200) );
 a88181a <=( A265  and  A203 );
 a88182a <=( a88181a  and  a88178a );
 a88183a <=( a88182a  and  a88175a );
 a88187a <=( (not A269)  and  (not A267) );
 a88188a <=( (not A266)  and  a88187a );
 a88191a <=( (not A299)  and  (not A298) );
 a88194a <=( (not A302)  and  A301 );
 a88195a <=( a88194a  and  a88191a );
 a88196a <=( a88195a  and  a88188a );
 a88200a <=( A199  and  (not A167) );
 a88201a <=( (not A168)  and  a88200a );
 a88204a <=( (not A201)  and  (not A200) );
 a88207a <=( A265  and  A202 );
 a88208a <=( a88207a  and  a88204a );
 a88209a <=( a88208a  and  a88201a );
 a88213a <=( (not A269)  and  A268 );
 a88214a <=( A266  and  a88213a );
 a88217a <=( A299  and  A298 );
 a88220a <=( (not A301)  and  (not A300) );
 a88221a <=( a88220a  and  a88217a );
 a88222a <=( a88221a  and  a88214a );
 a88226a <=( A199  and  (not A167) );
 a88227a <=( (not A168)  and  a88226a );
 a88230a <=( (not A201)  and  (not A200) );
 a88233a <=( A265  and  A202 );
 a88234a <=( a88233a  and  a88230a );
 a88235a <=( a88234a  and  a88227a );
 a88239a <=( (not A269)  and  A268 );
 a88240a <=( A266  and  a88239a );
 a88243a <=( A299  and  A298 );
 a88246a <=( A302  and  (not A300) );
 a88247a <=( a88246a  and  a88243a );
 a88248a <=( a88247a  and  a88240a );
 a88252a <=( A199  and  (not A167) );
 a88253a <=( (not A168)  and  a88252a );
 a88256a <=( (not A201)  and  (not A200) );
 a88259a <=( A265  and  A202 );
 a88260a <=( a88259a  and  a88256a );
 a88261a <=( a88260a  and  a88253a );
 a88265a <=( (not A269)  and  A268 );
 a88266a <=( A266  and  a88265a );
 a88269a <=( (not A299)  and  A298 );
 a88272a <=( A301  and  (not A300) );
 a88273a <=( a88272a  and  a88269a );
 a88274a <=( a88273a  and  a88266a );
 a88278a <=( A199  and  (not A167) );
 a88279a <=( (not A168)  and  a88278a );
 a88282a <=( (not A201)  and  (not A200) );
 a88285a <=( A265  and  A202 );
 a88286a <=( a88285a  and  a88282a );
 a88287a <=( a88286a  and  a88279a );
 a88291a <=( (not A269)  and  A268 );
 a88292a <=( A266  and  a88291a );
 a88295a <=( (not A299)  and  A298 );
 a88298a <=( (not A302)  and  (not A300) );
 a88299a <=( a88298a  and  a88295a );
 a88300a <=( a88299a  and  a88292a );
 a88304a <=( A199  and  (not A167) );
 a88305a <=( (not A168)  and  a88304a );
 a88308a <=( (not A201)  and  (not A200) );
 a88311a <=( A265  and  A202 );
 a88312a <=( a88311a  and  a88308a );
 a88313a <=( a88312a  and  a88305a );
 a88317a <=( (not A269)  and  A268 );
 a88318a <=( A266  and  a88317a );
 a88321a <=( A299  and  (not A298) );
 a88324a <=( A301  and  (not A300) );
 a88325a <=( a88324a  and  a88321a );
 a88326a <=( a88325a  and  a88318a );
 a88330a <=( A199  and  (not A167) );
 a88331a <=( (not A168)  and  a88330a );
 a88334a <=( (not A201)  and  (not A200) );
 a88337a <=( A265  and  A202 );
 a88338a <=( a88337a  and  a88334a );
 a88339a <=( a88338a  and  a88331a );
 a88343a <=( (not A269)  and  A268 );
 a88344a <=( A266  and  a88343a );
 a88347a <=( A299  and  (not A298) );
 a88350a <=( (not A302)  and  (not A300) );
 a88351a <=( a88350a  and  a88347a );
 a88352a <=( a88351a  and  a88344a );
 a88356a <=( A199  and  (not A167) );
 a88357a <=( (not A168)  and  a88356a );
 a88360a <=( (not A201)  and  (not A200) );
 a88363a <=( (not A265)  and  A202 );
 a88364a <=( a88363a  and  a88360a );
 a88365a <=( a88364a  and  a88357a );
 a88369a <=( A269  and  (not A268) );
 a88370a <=( A266  and  a88369a );
 a88373a <=( A299  and  A298 );
 a88376a <=( (not A301)  and  (not A300) );
 a88377a <=( a88376a  and  a88373a );
 a88378a <=( a88377a  and  a88370a );
 a88382a <=( A199  and  (not A167) );
 a88383a <=( (not A168)  and  a88382a );
 a88386a <=( (not A201)  and  (not A200) );
 a88389a <=( (not A265)  and  A202 );
 a88390a <=( a88389a  and  a88386a );
 a88391a <=( a88390a  and  a88383a );
 a88395a <=( A269  and  (not A268) );
 a88396a <=( A266  and  a88395a );
 a88399a <=( A299  and  A298 );
 a88402a <=( A302  and  (not A300) );
 a88403a <=( a88402a  and  a88399a );
 a88404a <=( a88403a  and  a88396a );
 a88408a <=( A199  and  (not A167) );
 a88409a <=( (not A168)  and  a88408a );
 a88412a <=( (not A201)  and  (not A200) );
 a88415a <=( (not A265)  and  A202 );
 a88416a <=( a88415a  and  a88412a );
 a88417a <=( a88416a  and  a88409a );
 a88421a <=( A269  and  (not A268) );
 a88422a <=( A266  and  a88421a );
 a88425a <=( (not A299)  and  A298 );
 a88428a <=( A301  and  (not A300) );
 a88429a <=( a88428a  and  a88425a );
 a88430a <=( a88429a  and  a88422a );
 a88434a <=( A199  and  (not A167) );
 a88435a <=( (not A168)  and  a88434a );
 a88438a <=( (not A201)  and  (not A200) );
 a88441a <=( (not A265)  and  A202 );
 a88442a <=( a88441a  and  a88438a );
 a88443a <=( a88442a  and  a88435a );
 a88447a <=( A269  and  (not A268) );
 a88448a <=( A266  and  a88447a );
 a88451a <=( (not A299)  and  A298 );
 a88454a <=( (not A302)  and  (not A300) );
 a88455a <=( a88454a  and  a88451a );
 a88456a <=( a88455a  and  a88448a );
 a88460a <=( A199  and  (not A167) );
 a88461a <=( (not A168)  and  a88460a );
 a88464a <=( (not A201)  and  (not A200) );
 a88467a <=( (not A265)  and  A202 );
 a88468a <=( a88467a  and  a88464a );
 a88469a <=( a88468a  and  a88461a );
 a88473a <=( A269  and  (not A268) );
 a88474a <=( A266  and  a88473a );
 a88477a <=( A299  and  (not A298) );
 a88480a <=( A301  and  (not A300) );
 a88481a <=( a88480a  and  a88477a );
 a88482a <=( a88481a  and  a88474a );
 a88486a <=( A199  and  (not A167) );
 a88487a <=( (not A168)  and  a88486a );
 a88490a <=( (not A201)  and  (not A200) );
 a88493a <=( (not A265)  and  A202 );
 a88494a <=( a88493a  and  a88490a );
 a88495a <=( a88494a  and  a88487a );
 a88499a <=( A269  and  (not A268) );
 a88500a <=( A266  and  a88499a );
 a88503a <=( A299  and  (not A298) );
 a88506a <=( (not A302)  and  (not A300) );
 a88507a <=( a88506a  and  a88503a );
 a88508a <=( a88507a  and  a88500a );
 a88512a <=( A199  and  (not A167) );
 a88513a <=( (not A168)  and  a88512a );
 a88516a <=( (not A201)  and  (not A200) );
 a88519a <=( A265  and  A202 );
 a88520a <=( a88519a  and  a88516a );
 a88521a <=( a88520a  and  a88513a );
 a88525a <=( A269  and  (not A268) );
 a88526a <=( (not A266)  and  a88525a );
 a88529a <=( A299  and  A298 );
 a88532a <=( (not A301)  and  (not A300) );
 a88533a <=( a88532a  and  a88529a );
 a88534a <=( a88533a  and  a88526a );
 a88538a <=( A199  and  (not A167) );
 a88539a <=( (not A168)  and  a88538a );
 a88542a <=( (not A201)  and  (not A200) );
 a88545a <=( A265  and  A202 );
 a88546a <=( a88545a  and  a88542a );
 a88547a <=( a88546a  and  a88539a );
 a88551a <=( A269  and  (not A268) );
 a88552a <=( (not A266)  and  a88551a );
 a88555a <=( A299  and  A298 );
 a88558a <=( A302  and  (not A300) );
 a88559a <=( a88558a  and  a88555a );
 a88560a <=( a88559a  and  a88552a );
 a88564a <=( A199  and  (not A167) );
 a88565a <=( (not A168)  and  a88564a );
 a88568a <=( (not A201)  and  (not A200) );
 a88571a <=( A265  and  A202 );
 a88572a <=( a88571a  and  a88568a );
 a88573a <=( a88572a  and  a88565a );
 a88577a <=( A269  and  (not A268) );
 a88578a <=( (not A266)  and  a88577a );
 a88581a <=( (not A299)  and  A298 );
 a88584a <=( A301  and  (not A300) );
 a88585a <=( a88584a  and  a88581a );
 a88586a <=( a88585a  and  a88578a );
 a88590a <=( A199  and  (not A167) );
 a88591a <=( (not A168)  and  a88590a );
 a88594a <=( (not A201)  and  (not A200) );
 a88597a <=( A265  and  A202 );
 a88598a <=( a88597a  and  a88594a );
 a88599a <=( a88598a  and  a88591a );
 a88603a <=( A269  and  (not A268) );
 a88604a <=( (not A266)  and  a88603a );
 a88607a <=( (not A299)  and  A298 );
 a88610a <=( (not A302)  and  (not A300) );
 a88611a <=( a88610a  and  a88607a );
 a88612a <=( a88611a  and  a88604a );
 a88616a <=( A199  and  (not A167) );
 a88617a <=( (not A168)  and  a88616a );
 a88620a <=( (not A201)  and  (not A200) );
 a88623a <=( A265  and  A202 );
 a88624a <=( a88623a  and  a88620a );
 a88625a <=( a88624a  and  a88617a );
 a88629a <=( A269  and  (not A268) );
 a88630a <=( (not A266)  and  a88629a );
 a88633a <=( A299  and  (not A298) );
 a88636a <=( A301  and  (not A300) );
 a88637a <=( a88636a  and  a88633a );
 a88638a <=( a88637a  and  a88630a );
 a88642a <=( A199  and  (not A167) );
 a88643a <=( (not A168)  and  a88642a );
 a88646a <=( (not A201)  and  (not A200) );
 a88649a <=( A265  and  A202 );
 a88650a <=( a88649a  and  a88646a );
 a88651a <=( a88650a  and  a88643a );
 a88655a <=( A269  and  (not A268) );
 a88656a <=( (not A266)  and  a88655a );
 a88659a <=( A299  and  (not A298) );
 a88662a <=( (not A302)  and  (not A300) );
 a88663a <=( a88662a  and  a88659a );
 a88664a <=( a88663a  and  a88656a );
 a88668a <=( A199  and  (not A167) );
 a88669a <=( (not A168)  and  a88668a );
 a88672a <=( (not A201)  and  (not A200) );
 a88675a <=( (not A265)  and  A202 );
 a88676a <=( a88675a  and  a88672a );
 a88677a <=( a88676a  and  a88669a );
 a88681a <=( (not A269)  and  A268 );
 a88682a <=( (not A266)  and  a88681a );
 a88685a <=( A299  and  A298 );
 a88688a <=( (not A301)  and  (not A300) );
 a88689a <=( a88688a  and  a88685a );
 a88690a <=( a88689a  and  a88682a );
 a88694a <=( A199  and  (not A167) );
 a88695a <=( (not A168)  and  a88694a );
 a88698a <=( (not A201)  and  (not A200) );
 a88701a <=( (not A265)  and  A202 );
 a88702a <=( a88701a  and  a88698a );
 a88703a <=( a88702a  and  a88695a );
 a88707a <=( (not A269)  and  A268 );
 a88708a <=( (not A266)  and  a88707a );
 a88711a <=( A299  and  A298 );
 a88714a <=( A302  and  (not A300) );
 a88715a <=( a88714a  and  a88711a );
 a88716a <=( a88715a  and  a88708a );
 a88720a <=( A199  and  (not A167) );
 a88721a <=( (not A168)  and  a88720a );
 a88724a <=( (not A201)  and  (not A200) );
 a88727a <=( (not A265)  and  A202 );
 a88728a <=( a88727a  and  a88724a );
 a88729a <=( a88728a  and  a88721a );
 a88733a <=( (not A269)  and  A268 );
 a88734a <=( (not A266)  and  a88733a );
 a88737a <=( (not A299)  and  A298 );
 a88740a <=( A301  and  (not A300) );
 a88741a <=( a88740a  and  a88737a );
 a88742a <=( a88741a  and  a88734a );
 a88746a <=( A199  and  (not A167) );
 a88747a <=( (not A168)  and  a88746a );
 a88750a <=( (not A201)  and  (not A200) );
 a88753a <=( (not A265)  and  A202 );
 a88754a <=( a88753a  and  a88750a );
 a88755a <=( a88754a  and  a88747a );
 a88759a <=( (not A269)  and  A268 );
 a88760a <=( (not A266)  and  a88759a );
 a88763a <=( (not A299)  and  A298 );
 a88766a <=( (not A302)  and  (not A300) );
 a88767a <=( a88766a  and  a88763a );
 a88768a <=( a88767a  and  a88760a );
 a88772a <=( A199  and  (not A167) );
 a88773a <=( (not A168)  and  a88772a );
 a88776a <=( (not A201)  and  (not A200) );
 a88779a <=( (not A265)  and  A202 );
 a88780a <=( a88779a  and  a88776a );
 a88781a <=( a88780a  and  a88773a );
 a88785a <=( (not A269)  and  A268 );
 a88786a <=( (not A266)  and  a88785a );
 a88789a <=( A299  and  (not A298) );
 a88792a <=( A301  and  (not A300) );
 a88793a <=( a88792a  and  a88789a );
 a88794a <=( a88793a  and  a88786a );
 a88798a <=( A199  and  (not A167) );
 a88799a <=( (not A168)  and  a88798a );
 a88802a <=( (not A201)  and  (not A200) );
 a88805a <=( (not A265)  and  A202 );
 a88806a <=( a88805a  and  a88802a );
 a88807a <=( a88806a  and  a88799a );
 a88811a <=( (not A269)  and  A268 );
 a88812a <=( (not A266)  and  a88811a );
 a88815a <=( A299  and  (not A298) );
 a88818a <=( (not A302)  and  (not A300) );
 a88819a <=( a88818a  and  a88815a );
 a88820a <=( a88819a  and  a88812a );
 a88824a <=( A199  and  (not A167) );
 a88825a <=( (not A168)  and  a88824a );
 a88828a <=( (not A201)  and  (not A200) );
 a88831a <=( A265  and  (not A203) );
 a88832a <=( a88831a  and  a88828a );
 a88833a <=( a88832a  and  a88825a );
 a88837a <=( (not A269)  and  A268 );
 a88838a <=( A266  and  a88837a );
 a88841a <=( A299  and  A298 );
 a88844a <=( (not A301)  and  (not A300) );
 a88845a <=( a88844a  and  a88841a );
 a88846a <=( a88845a  and  a88838a );
 a88850a <=( A199  and  (not A167) );
 a88851a <=( (not A168)  and  a88850a );
 a88854a <=( (not A201)  and  (not A200) );
 a88857a <=( A265  and  (not A203) );
 a88858a <=( a88857a  and  a88854a );
 a88859a <=( a88858a  and  a88851a );
 a88863a <=( (not A269)  and  A268 );
 a88864a <=( A266  and  a88863a );
 a88867a <=( A299  and  A298 );
 a88870a <=( A302  and  (not A300) );
 a88871a <=( a88870a  and  a88867a );
 a88872a <=( a88871a  and  a88864a );
 a88876a <=( A199  and  (not A167) );
 a88877a <=( (not A168)  and  a88876a );
 a88880a <=( (not A201)  and  (not A200) );
 a88883a <=( A265  and  (not A203) );
 a88884a <=( a88883a  and  a88880a );
 a88885a <=( a88884a  and  a88877a );
 a88889a <=( (not A269)  and  A268 );
 a88890a <=( A266  and  a88889a );
 a88893a <=( (not A299)  and  A298 );
 a88896a <=( A301  and  (not A300) );
 a88897a <=( a88896a  and  a88893a );
 a88898a <=( a88897a  and  a88890a );
 a88902a <=( A199  and  (not A167) );
 a88903a <=( (not A168)  and  a88902a );
 a88906a <=( (not A201)  and  (not A200) );
 a88909a <=( A265  and  (not A203) );
 a88910a <=( a88909a  and  a88906a );
 a88911a <=( a88910a  and  a88903a );
 a88915a <=( (not A269)  and  A268 );
 a88916a <=( A266  and  a88915a );
 a88919a <=( (not A299)  and  A298 );
 a88922a <=( (not A302)  and  (not A300) );
 a88923a <=( a88922a  and  a88919a );
 a88924a <=( a88923a  and  a88916a );
 a88928a <=( A199  and  (not A167) );
 a88929a <=( (not A168)  and  a88928a );
 a88932a <=( (not A201)  and  (not A200) );
 a88935a <=( A265  and  (not A203) );
 a88936a <=( a88935a  and  a88932a );
 a88937a <=( a88936a  and  a88929a );
 a88941a <=( (not A269)  and  A268 );
 a88942a <=( A266  and  a88941a );
 a88945a <=( A299  and  (not A298) );
 a88948a <=( A301  and  (not A300) );
 a88949a <=( a88948a  and  a88945a );
 a88950a <=( a88949a  and  a88942a );
 a88954a <=( A199  and  (not A167) );
 a88955a <=( (not A168)  and  a88954a );
 a88958a <=( (not A201)  and  (not A200) );
 a88961a <=( A265  and  (not A203) );
 a88962a <=( a88961a  and  a88958a );
 a88963a <=( a88962a  and  a88955a );
 a88967a <=( (not A269)  and  A268 );
 a88968a <=( A266  and  a88967a );
 a88971a <=( A299  and  (not A298) );
 a88974a <=( (not A302)  and  (not A300) );
 a88975a <=( a88974a  and  a88971a );
 a88976a <=( a88975a  and  a88968a );
 a88980a <=( A199  and  (not A167) );
 a88981a <=( (not A168)  and  a88980a );
 a88984a <=( (not A201)  and  (not A200) );
 a88987a <=( (not A265)  and  (not A203) );
 a88988a <=( a88987a  and  a88984a );
 a88989a <=( a88988a  and  a88981a );
 a88993a <=( A269  and  (not A268) );
 a88994a <=( A266  and  a88993a );
 a88997a <=( A299  and  A298 );
 a89000a <=( (not A301)  and  (not A300) );
 a89001a <=( a89000a  and  a88997a );
 a89002a <=( a89001a  and  a88994a );
 a89006a <=( A199  and  (not A167) );
 a89007a <=( (not A168)  and  a89006a );
 a89010a <=( (not A201)  and  (not A200) );
 a89013a <=( (not A265)  and  (not A203) );
 a89014a <=( a89013a  and  a89010a );
 a89015a <=( a89014a  and  a89007a );
 a89019a <=( A269  and  (not A268) );
 a89020a <=( A266  and  a89019a );
 a89023a <=( A299  and  A298 );
 a89026a <=( A302  and  (not A300) );
 a89027a <=( a89026a  and  a89023a );
 a89028a <=( a89027a  and  a89020a );
 a89032a <=( A199  and  (not A167) );
 a89033a <=( (not A168)  and  a89032a );
 a89036a <=( (not A201)  and  (not A200) );
 a89039a <=( (not A265)  and  (not A203) );
 a89040a <=( a89039a  and  a89036a );
 a89041a <=( a89040a  and  a89033a );
 a89045a <=( A269  and  (not A268) );
 a89046a <=( A266  and  a89045a );
 a89049a <=( (not A299)  and  A298 );
 a89052a <=( A301  and  (not A300) );
 a89053a <=( a89052a  and  a89049a );
 a89054a <=( a89053a  and  a89046a );
 a89058a <=( A199  and  (not A167) );
 a89059a <=( (not A168)  and  a89058a );
 a89062a <=( (not A201)  and  (not A200) );
 a89065a <=( (not A265)  and  (not A203) );
 a89066a <=( a89065a  and  a89062a );
 a89067a <=( a89066a  and  a89059a );
 a89071a <=( A269  and  (not A268) );
 a89072a <=( A266  and  a89071a );
 a89075a <=( (not A299)  and  A298 );
 a89078a <=( (not A302)  and  (not A300) );
 a89079a <=( a89078a  and  a89075a );
 a89080a <=( a89079a  and  a89072a );
 a89084a <=( A199  and  (not A167) );
 a89085a <=( (not A168)  and  a89084a );
 a89088a <=( (not A201)  and  (not A200) );
 a89091a <=( (not A265)  and  (not A203) );
 a89092a <=( a89091a  and  a89088a );
 a89093a <=( a89092a  and  a89085a );
 a89097a <=( A269  and  (not A268) );
 a89098a <=( A266  and  a89097a );
 a89101a <=( A299  and  (not A298) );
 a89104a <=( A301  and  (not A300) );
 a89105a <=( a89104a  and  a89101a );
 a89106a <=( a89105a  and  a89098a );
 a89110a <=( A199  and  (not A167) );
 a89111a <=( (not A168)  and  a89110a );
 a89114a <=( (not A201)  and  (not A200) );
 a89117a <=( (not A265)  and  (not A203) );
 a89118a <=( a89117a  and  a89114a );
 a89119a <=( a89118a  and  a89111a );
 a89123a <=( A269  and  (not A268) );
 a89124a <=( A266  and  a89123a );
 a89127a <=( A299  and  (not A298) );
 a89130a <=( (not A302)  and  (not A300) );
 a89131a <=( a89130a  and  a89127a );
 a89132a <=( a89131a  and  a89124a );
 a89136a <=( A199  and  (not A167) );
 a89137a <=( (not A168)  and  a89136a );
 a89140a <=( (not A201)  and  (not A200) );
 a89143a <=( A265  and  (not A203) );
 a89144a <=( a89143a  and  a89140a );
 a89145a <=( a89144a  and  a89137a );
 a89149a <=( A269  and  (not A268) );
 a89150a <=( (not A266)  and  a89149a );
 a89153a <=( A299  and  A298 );
 a89156a <=( (not A301)  and  (not A300) );
 a89157a <=( a89156a  and  a89153a );
 a89158a <=( a89157a  and  a89150a );
 a89162a <=( A199  and  (not A167) );
 a89163a <=( (not A168)  and  a89162a );
 a89166a <=( (not A201)  and  (not A200) );
 a89169a <=( A265  and  (not A203) );
 a89170a <=( a89169a  and  a89166a );
 a89171a <=( a89170a  and  a89163a );
 a89175a <=( A269  and  (not A268) );
 a89176a <=( (not A266)  and  a89175a );
 a89179a <=( A299  and  A298 );
 a89182a <=( A302  and  (not A300) );
 a89183a <=( a89182a  and  a89179a );
 a89184a <=( a89183a  and  a89176a );
 a89188a <=( A199  and  (not A167) );
 a89189a <=( (not A168)  and  a89188a );
 a89192a <=( (not A201)  and  (not A200) );
 a89195a <=( A265  and  (not A203) );
 a89196a <=( a89195a  and  a89192a );
 a89197a <=( a89196a  and  a89189a );
 a89201a <=( A269  and  (not A268) );
 a89202a <=( (not A266)  and  a89201a );
 a89205a <=( (not A299)  and  A298 );
 a89208a <=( A301  and  (not A300) );
 a89209a <=( a89208a  and  a89205a );
 a89210a <=( a89209a  and  a89202a );
 a89214a <=( A199  and  (not A167) );
 a89215a <=( (not A168)  and  a89214a );
 a89218a <=( (not A201)  and  (not A200) );
 a89221a <=( A265  and  (not A203) );
 a89222a <=( a89221a  and  a89218a );
 a89223a <=( a89222a  and  a89215a );
 a89227a <=( A269  and  (not A268) );
 a89228a <=( (not A266)  and  a89227a );
 a89231a <=( (not A299)  and  A298 );
 a89234a <=( (not A302)  and  (not A300) );
 a89235a <=( a89234a  and  a89231a );
 a89236a <=( a89235a  and  a89228a );
 a89240a <=( A199  and  (not A167) );
 a89241a <=( (not A168)  and  a89240a );
 a89244a <=( (not A201)  and  (not A200) );
 a89247a <=( A265  and  (not A203) );
 a89248a <=( a89247a  and  a89244a );
 a89249a <=( a89248a  and  a89241a );
 a89253a <=( A269  and  (not A268) );
 a89254a <=( (not A266)  and  a89253a );
 a89257a <=( A299  and  (not A298) );
 a89260a <=( A301  and  (not A300) );
 a89261a <=( a89260a  and  a89257a );
 a89262a <=( a89261a  and  a89254a );
 a89266a <=( A199  and  (not A167) );
 a89267a <=( (not A168)  and  a89266a );
 a89270a <=( (not A201)  and  (not A200) );
 a89273a <=( A265  and  (not A203) );
 a89274a <=( a89273a  and  a89270a );
 a89275a <=( a89274a  and  a89267a );
 a89279a <=( A269  and  (not A268) );
 a89280a <=( (not A266)  and  a89279a );
 a89283a <=( A299  and  (not A298) );
 a89286a <=( (not A302)  and  (not A300) );
 a89287a <=( a89286a  and  a89283a );
 a89288a <=( a89287a  and  a89280a );
 a89292a <=( A199  and  (not A167) );
 a89293a <=( (not A168)  and  a89292a );
 a89296a <=( (not A201)  and  (not A200) );
 a89299a <=( (not A265)  and  (not A203) );
 a89300a <=( a89299a  and  a89296a );
 a89301a <=( a89300a  and  a89293a );
 a89305a <=( (not A269)  and  A268 );
 a89306a <=( (not A266)  and  a89305a );
 a89309a <=( A299  and  A298 );
 a89312a <=( (not A301)  and  (not A300) );
 a89313a <=( a89312a  and  a89309a );
 a89314a <=( a89313a  and  a89306a );
 a89318a <=( A199  and  (not A167) );
 a89319a <=( (not A168)  and  a89318a );
 a89322a <=( (not A201)  and  (not A200) );
 a89325a <=( (not A265)  and  (not A203) );
 a89326a <=( a89325a  and  a89322a );
 a89327a <=( a89326a  and  a89319a );
 a89331a <=( (not A269)  and  A268 );
 a89332a <=( (not A266)  and  a89331a );
 a89335a <=( A299  and  A298 );
 a89338a <=( A302  and  (not A300) );
 a89339a <=( a89338a  and  a89335a );
 a89340a <=( a89339a  and  a89332a );
 a89344a <=( A199  and  (not A167) );
 a89345a <=( (not A168)  and  a89344a );
 a89348a <=( (not A201)  and  (not A200) );
 a89351a <=( (not A265)  and  (not A203) );
 a89352a <=( a89351a  and  a89348a );
 a89353a <=( a89352a  and  a89345a );
 a89357a <=( (not A269)  and  A268 );
 a89358a <=( (not A266)  and  a89357a );
 a89361a <=( (not A299)  and  A298 );
 a89364a <=( A301  and  (not A300) );
 a89365a <=( a89364a  and  a89361a );
 a89366a <=( a89365a  and  a89358a );
 a89370a <=( A199  and  (not A167) );
 a89371a <=( (not A168)  and  a89370a );
 a89374a <=( (not A201)  and  (not A200) );
 a89377a <=( (not A265)  and  (not A203) );
 a89378a <=( a89377a  and  a89374a );
 a89379a <=( a89378a  and  a89371a );
 a89383a <=( (not A269)  and  A268 );
 a89384a <=( (not A266)  and  a89383a );
 a89387a <=( (not A299)  and  A298 );
 a89390a <=( (not A302)  and  (not A300) );
 a89391a <=( a89390a  and  a89387a );
 a89392a <=( a89391a  and  a89384a );
 a89396a <=( A199  and  (not A167) );
 a89397a <=( (not A168)  and  a89396a );
 a89400a <=( (not A201)  and  (not A200) );
 a89403a <=( (not A265)  and  (not A203) );
 a89404a <=( a89403a  and  a89400a );
 a89405a <=( a89404a  and  a89397a );
 a89409a <=( (not A269)  and  A268 );
 a89410a <=( (not A266)  and  a89409a );
 a89413a <=( A299  and  (not A298) );
 a89416a <=( A301  and  (not A300) );
 a89417a <=( a89416a  and  a89413a );
 a89418a <=( a89417a  and  a89410a );
 a89422a <=( A199  and  (not A167) );
 a89423a <=( (not A168)  and  a89422a );
 a89426a <=( (not A201)  and  (not A200) );
 a89429a <=( (not A265)  and  (not A203) );
 a89430a <=( a89429a  and  a89426a );
 a89431a <=( a89430a  and  a89423a );
 a89435a <=( (not A269)  and  A268 );
 a89436a <=( (not A266)  and  a89435a );
 a89439a <=( A299  and  (not A298) );
 a89442a <=( (not A302)  and  (not A300) );
 a89443a <=( a89442a  and  a89439a );
 a89444a <=( a89443a  and  a89436a );
 a89448a <=( (not A199)  and  (not A167) );
 a89449a <=( (not A168)  and  a89448a );
 a89452a <=( A202  and  (not A200) );
 a89455a <=( A265  and  (not A203) );
 a89456a <=( a89455a  and  a89452a );
 a89457a <=( a89456a  and  a89449a );
 a89461a <=( (not A268)  and  (not A267) );
 a89462a <=( A266  and  a89461a );
 a89465a <=( A299  and  A298 );
 a89468a <=( (not A302)  and  A301 );
 a89469a <=( a89468a  and  a89465a );
 a89470a <=( a89469a  and  a89462a );
 a89474a <=( (not A199)  and  (not A167) );
 a89475a <=( (not A168)  and  a89474a );
 a89478a <=( A202  and  (not A200) );
 a89481a <=( A265  and  (not A203) );
 a89482a <=( a89481a  and  a89478a );
 a89483a <=( a89482a  and  a89475a );
 a89487a <=( (not A268)  and  (not A267) );
 a89488a <=( A266  and  a89487a );
 a89491a <=( (not A299)  and  A298 );
 a89494a <=( A302  and  (not A301) );
 a89495a <=( a89494a  and  a89491a );
 a89496a <=( a89495a  and  a89488a );
 a89500a <=( (not A199)  and  (not A167) );
 a89501a <=( (not A168)  and  a89500a );
 a89504a <=( A202  and  (not A200) );
 a89507a <=( A265  and  (not A203) );
 a89508a <=( a89507a  and  a89504a );
 a89509a <=( a89508a  and  a89501a );
 a89513a <=( (not A268)  and  (not A267) );
 a89514a <=( A266  and  a89513a );
 a89517a <=( A299  and  (not A298) );
 a89520a <=( A302  and  (not A301) );
 a89521a <=( a89520a  and  a89517a );
 a89522a <=( a89521a  and  a89514a );
 a89526a <=( (not A199)  and  (not A167) );
 a89527a <=( (not A168)  and  a89526a );
 a89530a <=( A202  and  (not A200) );
 a89533a <=( A265  and  (not A203) );
 a89534a <=( a89533a  and  a89530a );
 a89535a <=( a89534a  and  a89527a );
 a89539a <=( (not A268)  and  (not A267) );
 a89540a <=( A266  and  a89539a );
 a89543a <=( (not A299)  and  (not A298) );
 a89546a <=( (not A302)  and  A301 );
 a89547a <=( a89546a  and  a89543a );
 a89548a <=( a89547a  and  a89540a );
 a89552a <=( (not A199)  and  (not A167) );
 a89553a <=( (not A168)  and  a89552a );
 a89556a <=( A202  and  (not A200) );
 a89559a <=( A265  and  (not A203) );
 a89560a <=( a89559a  and  a89556a );
 a89561a <=( a89560a  and  a89553a );
 a89565a <=( A269  and  (not A267) );
 a89566a <=( A266  and  a89565a );
 a89569a <=( A299  and  A298 );
 a89572a <=( (not A302)  and  A301 );
 a89573a <=( a89572a  and  a89569a );
 a89574a <=( a89573a  and  a89566a );
 a89578a <=( (not A199)  and  (not A167) );
 a89579a <=( (not A168)  and  a89578a );
 a89582a <=( A202  and  (not A200) );
 a89585a <=( A265  and  (not A203) );
 a89586a <=( a89585a  and  a89582a );
 a89587a <=( a89586a  and  a89579a );
 a89591a <=( A269  and  (not A267) );
 a89592a <=( A266  and  a89591a );
 a89595a <=( (not A299)  and  A298 );
 a89598a <=( A302  and  (not A301) );
 a89599a <=( a89598a  and  a89595a );
 a89600a <=( a89599a  and  a89592a );
 a89604a <=( (not A199)  and  (not A167) );
 a89605a <=( (not A168)  and  a89604a );
 a89608a <=( A202  and  (not A200) );
 a89611a <=( A265  and  (not A203) );
 a89612a <=( a89611a  and  a89608a );
 a89613a <=( a89612a  and  a89605a );
 a89617a <=( A269  and  (not A267) );
 a89618a <=( A266  and  a89617a );
 a89621a <=( A299  and  (not A298) );
 a89624a <=( A302  and  (not A301) );
 a89625a <=( a89624a  and  a89621a );
 a89626a <=( a89625a  and  a89618a );
 a89630a <=( (not A199)  and  (not A167) );
 a89631a <=( (not A168)  and  a89630a );
 a89634a <=( A202  and  (not A200) );
 a89637a <=( A265  and  (not A203) );
 a89638a <=( a89637a  and  a89634a );
 a89639a <=( a89638a  and  a89631a );
 a89643a <=( A269  and  (not A267) );
 a89644a <=( A266  and  a89643a );
 a89647a <=( (not A299)  and  (not A298) );
 a89650a <=( (not A302)  and  A301 );
 a89651a <=( a89650a  and  a89647a );
 a89652a <=( a89651a  and  a89644a );
 a89656a <=( (not A199)  and  (not A167) );
 a89657a <=( (not A168)  and  a89656a );
 a89660a <=( A202  and  (not A200) );
 a89663a <=( (not A265)  and  (not A203) );
 a89664a <=( a89663a  and  a89660a );
 a89665a <=( a89664a  and  a89657a );
 a89669a <=( A268  and  (not A267) );
 a89670a <=( A266  and  a89669a );
 a89673a <=( A299  and  A298 );
 a89676a <=( (not A302)  and  A301 );
 a89677a <=( a89676a  and  a89673a );
 a89678a <=( a89677a  and  a89670a );
 a89682a <=( (not A199)  and  (not A167) );
 a89683a <=( (not A168)  and  a89682a );
 a89686a <=( A202  and  (not A200) );
 a89689a <=( (not A265)  and  (not A203) );
 a89690a <=( a89689a  and  a89686a );
 a89691a <=( a89690a  and  a89683a );
 a89695a <=( A268  and  (not A267) );
 a89696a <=( A266  and  a89695a );
 a89699a <=( (not A299)  and  A298 );
 a89702a <=( A302  and  (not A301) );
 a89703a <=( a89702a  and  a89699a );
 a89704a <=( a89703a  and  a89696a );
 a89708a <=( (not A199)  and  (not A167) );
 a89709a <=( (not A168)  and  a89708a );
 a89712a <=( A202  and  (not A200) );
 a89715a <=( (not A265)  and  (not A203) );
 a89716a <=( a89715a  and  a89712a );
 a89717a <=( a89716a  and  a89709a );
 a89721a <=( A268  and  (not A267) );
 a89722a <=( A266  and  a89721a );
 a89725a <=( A299  and  (not A298) );
 a89728a <=( A302  and  (not A301) );
 a89729a <=( a89728a  and  a89725a );
 a89730a <=( a89729a  and  a89722a );
 a89734a <=( (not A199)  and  (not A167) );
 a89735a <=( (not A168)  and  a89734a );
 a89738a <=( A202  and  (not A200) );
 a89741a <=( (not A265)  and  (not A203) );
 a89742a <=( a89741a  and  a89738a );
 a89743a <=( a89742a  and  a89735a );
 a89747a <=( A268  and  (not A267) );
 a89748a <=( A266  and  a89747a );
 a89751a <=( (not A299)  and  (not A298) );
 a89754a <=( (not A302)  and  A301 );
 a89755a <=( a89754a  and  a89751a );
 a89756a <=( a89755a  and  a89748a );
 a89760a <=( (not A199)  and  (not A167) );
 a89761a <=( (not A168)  and  a89760a );
 a89764a <=( A202  and  (not A200) );
 a89767a <=( (not A265)  and  (not A203) );
 a89768a <=( a89767a  and  a89764a );
 a89769a <=( a89768a  and  a89761a );
 a89773a <=( (not A269)  and  (not A267) );
 a89774a <=( A266  and  a89773a );
 a89777a <=( A299  and  A298 );
 a89780a <=( (not A302)  and  A301 );
 a89781a <=( a89780a  and  a89777a );
 a89782a <=( a89781a  and  a89774a );
 a89786a <=( (not A199)  and  (not A167) );
 a89787a <=( (not A168)  and  a89786a );
 a89790a <=( A202  and  (not A200) );
 a89793a <=( (not A265)  and  (not A203) );
 a89794a <=( a89793a  and  a89790a );
 a89795a <=( a89794a  and  a89787a );
 a89799a <=( (not A269)  and  (not A267) );
 a89800a <=( A266  and  a89799a );
 a89803a <=( (not A299)  and  A298 );
 a89806a <=( A302  and  (not A301) );
 a89807a <=( a89806a  and  a89803a );
 a89808a <=( a89807a  and  a89800a );
 a89812a <=( (not A199)  and  (not A167) );
 a89813a <=( (not A168)  and  a89812a );
 a89816a <=( A202  and  (not A200) );
 a89819a <=( (not A265)  and  (not A203) );
 a89820a <=( a89819a  and  a89816a );
 a89821a <=( a89820a  and  a89813a );
 a89825a <=( (not A269)  and  (not A267) );
 a89826a <=( A266  and  a89825a );
 a89829a <=( A299  and  (not A298) );
 a89832a <=( A302  and  (not A301) );
 a89833a <=( a89832a  and  a89829a );
 a89834a <=( a89833a  and  a89826a );
 a89838a <=( (not A199)  and  (not A167) );
 a89839a <=( (not A168)  and  a89838a );
 a89842a <=( A202  and  (not A200) );
 a89845a <=( (not A265)  and  (not A203) );
 a89846a <=( a89845a  and  a89842a );
 a89847a <=( a89846a  and  a89839a );
 a89851a <=( (not A269)  and  (not A267) );
 a89852a <=( A266  and  a89851a );
 a89855a <=( (not A299)  and  (not A298) );
 a89858a <=( (not A302)  and  A301 );
 a89859a <=( a89858a  and  a89855a );
 a89860a <=( a89859a  and  a89852a );
 a89864a <=( (not A199)  and  (not A167) );
 a89865a <=( (not A168)  and  a89864a );
 a89868a <=( A202  and  (not A200) );
 a89871a <=( A265  and  (not A203) );
 a89872a <=( a89871a  and  a89868a );
 a89873a <=( a89872a  and  a89865a );
 a89877a <=( A268  and  (not A267) );
 a89878a <=( (not A266)  and  a89877a );
 a89881a <=( A299  and  A298 );
 a89884a <=( (not A302)  and  A301 );
 a89885a <=( a89884a  and  a89881a );
 a89886a <=( a89885a  and  a89878a );
 a89890a <=( (not A199)  and  (not A167) );
 a89891a <=( (not A168)  and  a89890a );
 a89894a <=( A202  and  (not A200) );
 a89897a <=( A265  and  (not A203) );
 a89898a <=( a89897a  and  a89894a );
 a89899a <=( a89898a  and  a89891a );
 a89903a <=( A268  and  (not A267) );
 a89904a <=( (not A266)  and  a89903a );
 a89907a <=( (not A299)  and  A298 );
 a89910a <=( A302  and  (not A301) );
 a89911a <=( a89910a  and  a89907a );
 a89912a <=( a89911a  and  a89904a );
 a89916a <=( (not A199)  and  (not A167) );
 a89917a <=( (not A168)  and  a89916a );
 a89920a <=( A202  and  (not A200) );
 a89923a <=( A265  and  (not A203) );
 a89924a <=( a89923a  and  a89920a );
 a89925a <=( a89924a  and  a89917a );
 a89929a <=( A268  and  (not A267) );
 a89930a <=( (not A266)  and  a89929a );
 a89933a <=( A299  and  (not A298) );
 a89936a <=( A302  and  (not A301) );
 a89937a <=( a89936a  and  a89933a );
 a89938a <=( a89937a  and  a89930a );
 a89942a <=( (not A199)  and  (not A167) );
 a89943a <=( (not A168)  and  a89942a );
 a89946a <=( A202  and  (not A200) );
 a89949a <=( A265  and  (not A203) );
 a89950a <=( a89949a  and  a89946a );
 a89951a <=( a89950a  and  a89943a );
 a89955a <=( A268  and  (not A267) );
 a89956a <=( (not A266)  and  a89955a );
 a89959a <=( (not A299)  and  (not A298) );
 a89962a <=( (not A302)  and  A301 );
 a89963a <=( a89962a  and  a89959a );
 a89964a <=( a89963a  and  a89956a );
 a89968a <=( (not A199)  and  (not A167) );
 a89969a <=( (not A168)  and  a89968a );
 a89972a <=( A202  and  (not A200) );
 a89975a <=( A265  and  (not A203) );
 a89976a <=( a89975a  and  a89972a );
 a89977a <=( a89976a  and  a89969a );
 a89981a <=( (not A269)  and  (not A267) );
 a89982a <=( (not A266)  and  a89981a );
 a89985a <=( A299  and  A298 );
 a89988a <=( (not A302)  and  A301 );
 a89989a <=( a89988a  and  a89985a );
 a89990a <=( a89989a  and  a89982a );
 a89994a <=( (not A199)  and  (not A167) );
 a89995a <=( (not A168)  and  a89994a );
 a89998a <=( A202  and  (not A200) );
 a90001a <=( A265  and  (not A203) );
 a90002a <=( a90001a  and  a89998a );
 a90003a <=( a90002a  and  a89995a );
 a90007a <=( (not A269)  and  (not A267) );
 a90008a <=( (not A266)  and  a90007a );
 a90011a <=( (not A299)  and  A298 );
 a90014a <=( A302  and  (not A301) );
 a90015a <=( a90014a  and  a90011a );
 a90016a <=( a90015a  and  a90008a );
 a90020a <=( (not A199)  and  (not A167) );
 a90021a <=( (not A168)  and  a90020a );
 a90024a <=( A202  and  (not A200) );
 a90027a <=( A265  and  (not A203) );
 a90028a <=( a90027a  and  a90024a );
 a90029a <=( a90028a  and  a90021a );
 a90033a <=( (not A269)  and  (not A267) );
 a90034a <=( (not A266)  and  a90033a );
 a90037a <=( A299  and  (not A298) );
 a90040a <=( A302  and  (not A301) );
 a90041a <=( a90040a  and  a90037a );
 a90042a <=( a90041a  and  a90034a );
 a90046a <=( (not A199)  and  (not A167) );
 a90047a <=( (not A168)  and  a90046a );
 a90050a <=( A202  and  (not A200) );
 a90053a <=( A265  and  (not A203) );
 a90054a <=( a90053a  and  a90050a );
 a90055a <=( a90054a  and  a90047a );
 a90059a <=( (not A269)  and  (not A267) );
 a90060a <=( (not A266)  and  a90059a );
 a90063a <=( (not A299)  and  (not A298) );
 a90066a <=( (not A302)  and  A301 );
 a90067a <=( a90066a  and  a90063a );
 a90068a <=( a90067a  and  a90060a );
 a90072a <=( (not A167)  and  A168 );
 a90073a <=( A170  and  a90072a );
 a90076a <=( A199  and  A166 );
 a90079a <=( A265  and  A201 );
 a90080a <=( a90079a  and  a90076a );
 a90081a <=( a90080a  and  a90073a );
 a90085a <=( (not A269)  and  A268 );
 a90086a <=( A266  and  a90085a );
 a90089a <=( A299  and  A298 );
 a90092a <=( (not A301)  and  (not A300) );
 a90093a <=( a90092a  and  a90089a );
 a90094a <=( a90093a  and  a90086a );
 a90098a <=( (not A167)  and  A168 );
 a90099a <=( A170  and  a90098a );
 a90102a <=( A199  and  A166 );
 a90105a <=( A265  and  A201 );
 a90106a <=( a90105a  and  a90102a );
 a90107a <=( a90106a  and  a90099a );
 a90111a <=( (not A269)  and  A268 );
 a90112a <=( A266  and  a90111a );
 a90115a <=( A299  and  A298 );
 a90118a <=( A302  and  (not A300) );
 a90119a <=( a90118a  and  a90115a );
 a90120a <=( a90119a  and  a90112a );
 a90124a <=( (not A167)  and  A168 );
 a90125a <=( A170  and  a90124a );
 a90128a <=( A199  and  A166 );
 a90131a <=( A265  and  A201 );
 a90132a <=( a90131a  and  a90128a );
 a90133a <=( a90132a  and  a90125a );
 a90137a <=( (not A269)  and  A268 );
 a90138a <=( A266  and  a90137a );
 a90141a <=( (not A299)  and  A298 );
 a90144a <=( A301  and  (not A300) );
 a90145a <=( a90144a  and  a90141a );
 a90146a <=( a90145a  and  a90138a );
 a90150a <=( (not A167)  and  A168 );
 a90151a <=( A170  and  a90150a );
 a90154a <=( A199  and  A166 );
 a90157a <=( A265  and  A201 );
 a90158a <=( a90157a  and  a90154a );
 a90159a <=( a90158a  and  a90151a );
 a90163a <=( (not A269)  and  A268 );
 a90164a <=( A266  and  a90163a );
 a90167a <=( (not A299)  and  A298 );
 a90170a <=( (not A302)  and  (not A300) );
 a90171a <=( a90170a  and  a90167a );
 a90172a <=( a90171a  and  a90164a );
 a90176a <=( (not A167)  and  A168 );
 a90177a <=( A170  and  a90176a );
 a90180a <=( A199  and  A166 );
 a90183a <=( A265  and  A201 );
 a90184a <=( a90183a  and  a90180a );
 a90185a <=( a90184a  and  a90177a );
 a90189a <=( (not A269)  and  A268 );
 a90190a <=( A266  and  a90189a );
 a90193a <=( A299  and  (not A298) );
 a90196a <=( A301  and  (not A300) );
 a90197a <=( a90196a  and  a90193a );
 a90198a <=( a90197a  and  a90190a );
 a90202a <=( (not A167)  and  A168 );
 a90203a <=( A170  and  a90202a );
 a90206a <=( A199  and  A166 );
 a90209a <=( A265  and  A201 );
 a90210a <=( a90209a  and  a90206a );
 a90211a <=( a90210a  and  a90203a );
 a90215a <=( (not A269)  and  A268 );
 a90216a <=( A266  and  a90215a );
 a90219a <=( A299  and  (not A298) );
 a90222a <=( (not A302)  and  (not A300) );
 a90223a <=( a90222a  and  a90219a );
 a90224a <=( a90223a  and  a90216a );
 a90228a <=( (not A167)  and  A168 );
 a90229a <=( A170  and  a90228a );
 a90232a <=( A199  and  A166 );
 a90235a <=( (not A265)  and  A201 );
 a90236a <=( a90235a  and  a90232a );
 a90237a <=( a90236a  and  a90229a );
 a90241a <=( A269  and  (not A268) );
 a90242a <=( A266  and  a90241a );
 a90245a <=( A299  and  A298 );
 a90248a <=( (not A301)  and  (not A300) );
 a90249a <=( a90248a  and  a90245a );
 a90250a <=( a90249a  and  a90242a );
 a90254a <=( (not A167)  and  A168 );
 a90255a <=( A170  and  a90254a );
 a90258a <=( A199  and  A166 );
 a90261a <=( (not A265)  and  A201 );
 a90262a <=( a90261a  and  a90258a );
 a90263a <=( a90262a  and  a90255a );
 a90267a <=( A269  and  (not A268) );
 a90268a <=( A266  and  a90267a );
 a90271a <=( A299  and  A298 );
 a90274a <=( A302  and  (not A300) );
 a90275a <=( a90274a  and  a90271a );
 a90276a <=( a90275a  and  a90268a );
 a90280a <=( (not A167)  and  A168 );
 a90281a <=( A170  and  a90280a );
 a90284a <=( A199  and  A166 );
 a90287a <=( (not A265)  and  A201 );
 a90288a <=( a90287a  and  a90284a );
 a90289a <=( a90288a  and  a90281a );
 a90293a <=( A269  and  (not A268) );
 a90294a <=( A266  and  a90293a );
 a90297a <=( (not A299)  and  A298 );
 a90300a <=( A301  and  (not A300) );
 a90301a <=( a90300a  and  a90297a );
 a90302a <=( a90301a  and  a90294a );
 a90306a <=( (not A167)  and  A168 );
 a90307a <=( A170  and  a90306a );
 a90310a <=( A199  and  A166 );
 a90313a <=( (not A265)  and  A201 );
 a90314a <=( a90313a  and  a90310a );
 a90315a <=( a90314a  and  a90307a );
 a90319a <=( A269  and  (not A268) );
 a90320a <=( A266  and  a90319a );
 a90323a <=( (not A299)  and  A298 );
 a90326a <=( (not A302)  and  (not A300) );
 a90327a <=( a90326a  and  a90323a );
 a90328a <=( a90327a  and  a90320a );
 a90332a <=( (not A167)  and  A168 );
 a90333a <=( A170  and  a90332a );
 a90336a <=( A199  and  A166 );
 a90339a <=( (not A265)  and  A201 );
 a90340a <=( a90339a  and  a90336a );
 a90341a <=( a90340a  and  a90333a );
 a90345a <=( A269  and  (not A268) );
 a90346a <=( A266  and  a90345a );
 a90349a <=( A299  and  (not A298) );
 a90352a <=( A301  and  (not A300) );
 a90353a <=( a90352a  and  a90349a );
 a90354a <=( a90353a  and  a90346a );
 a90358a <=( (not A167)  and  A168 );
 a90359a <=( A170  and  a90358a );
 a90362a <=( A199  and  A166 );
 a90365a <=( (not A265)  and  A201 );
 a90366a <=( a90365a  and  a90362a );
 a90367a <=( a90366a  and  a90359a );
 a90371a <=( A269  and  (not A268) );
 a90372a <=( A266  and  a90371a );
 a90375a <=( A299  and  (not A298) );
 a90378a <=( (not A302)  and  (not A300) );
 a90379a <=( a90378a  and  a90375a );
 a90380a <=( a90379a  and  a90372a );
 a90384a <=( (not A167)  and  A168 );
 a90385a <=( A170  and  a90384a );
 a90388a <=( A199  and  A166 );
 a90391a <=( A265  and  A201 );
 a90392a <=( a90391a  and  a90388a );
 a90393a <=( a90392a  and  a90385a );
 a90397a <=( A269  and  (not A268) );
 a90398a <=( (not A266)  and  a90397a );
 a90401a <=( A299  and  A298 );
 a90404a <=( (not A301)  and  (not A300) );
 a90405a <=( a90404a  and  a90401a );
 a90406a <=( a90405a  and  a90398a );
 a90410a <=( (not A167)  and  A168 );
 a90411a <=( A170  and  a90410a );
 a90414a <=( A199  and  A166 );
 a90417a <=( A265  and  A201 );
 a90418a <=( a90417a  and  a90414a );
 a90419a <=( a90418a  and  a90411a );
 a90423a <=( A269  and  (not A268) );
 a90424a <=( (not A266)  and  a90423a );
 a90427a <=( A299  and  A298 );
 a90430a <=( A302  and  (not A300) );
 a90431a <=( a90430a  and  a90427a );
 a90432a <=( a90431a  and  a90424a );
 a90436a <=( (not A167)  and  A168 );
 a90437a <=( A170  and  a90436a );
 a90440a <=( A199  and  A166 );
 a90443a <=( A265  and  A201 );
 a90444a <=( a90443a  and  a90440a );
 a90445a <=( a90444a  and  a90437a );
 a90449a <=( A269  and  (not A268) );
 a90450a <=( (not A266)  and  a90449a );
 a90453a <=( (not A299)  and  A298 );
 a90456a <=( A301  and  (not A300) );
 a90457a <=( a90456a  and  a90453a );
 a90458a <=( a90457a  and  a90450a );
 a90462a <=( (not A167)  and  A168 );
 a90463a <=( A170  and  a90462a );
 a90466a <=( A199  and  A166 );
 a90469a <=( A265  and  A201 );
 a90470a <=( a90469a  and  a90466a );
 a90471a <=( a90470a  and  a90463a );
 a90475a <=( A269  and  (not A268) );
 a90476a <=( (not A266)  and  a90475a );
 a90479a <=( (not A299)  and  A298 );
 a90482a <=( (not A302)  and  (not A300) );
 a90483a <=( a90482a  and  a90479a );
 a90484a <=( a90483a  and  a90476a );
 a90488a <=( (not A167)  and  A168 );
 a90489a <=( A170  and  a90488a );
 a90492a <=( A199  and  A166 );
 a90495a <=( A265  and  A201 );
 a90496a <=( a90495a  and  a90492a );
 a90497a <=( a90496a  and  a90489a );
 a90501a <=( A269  and  (not A268) );
 a90502a <=( (not A266)  and  a90501a );
 a90505a <=( A299  and  (not A298) );
 a90508a <=( A301  and  (not A300) );
 a90509a <=( a90508a  and  a90505a );
 a90510a <=( a90509a  and  a90502a );
 a90514a <=( (not A167)  and  A168 );
 a90515a <=( A170  and  a90514a );
 a90518a <=( A199  and  A166 );
 a90521a <=( A265  and  A201 );
 a90522a <=( a90521a  and  a90518a );
 a90523a <=( a90522a  and  a90515a );
 a90527a <=( A269  and  (not A268) );
 a90528a <=( (not A266)  and  a90527a );
 a90531a <=( A299  and  (not A298) );
 a90534a <=( (not A302)  and  (not A300) );
 a90535a <=( a90534a  and  a90531a );
 a90536a <=( a90535a  and  a90528a );
 a90540a <=( (not A167)  and  A168 );
 a90541a <=( A170  and  a90540a );
 a90544a <=( A199  and  A166 );
 a90547a <=( (not A265)  and  A201 );
 a90548a <=( a90547a  and  a90544a );
 a90549a <=( a90548a  and  a90541a );
 a90553a <=( (not A269)  and  A268 );
 a90554a <=( (not A266)  and  a90553a );
 a90557a <=( A299  and  A298 );
 a90560a <=( (not A301)  and  (not A300) );
 a90561a <=( a90560a  and  a90557a );
 a90562a <=( a90561a  and  a90554a );
 a90566a <=( (not A167)  and  A168 );
 a90567a <=( A170  and  a90566a );
 a90570a <=( A199  and  A166 );
 a90573a <=( (not A265)  and  A201 );
 a90574a <=( a90573a  and  a90570a );
 a90575a <=( a90574a  and  a90567a );
 a90579a <=( (not A269)  and  A268 );
 a90580a <=( (not A266)  and  a90579a );
 a90583a <=( A299  and  A298 );
 a90586a <=( A302  and  (not A300) );
 a90587a <=( a90586a  and  a90583a );
 a90588a <=( a90587a  and  a90580a );
 a90592a <=( (not A167)  and  A168 );
 a90593a <=( A170  and  a90592a );
 a90596a <=( A199  and  A166 );
 a90599a <=( (not A265)  and  A201 );
 a90600a <=( a90599a  and  a90596a );
 a90601a <=( a90600a  and  a90593a );
 a90605a <=( (not A269)  and  A268 );
 a90606a <=( (not A266)  and  a90605a );
 a90609a <=( (not A299)  and  A298 );
 a90612a <=( A301  and  (not A300) );
 a90613a <=( a90612a  and  a90609a );
 a90614a <=( a90613a  and  a90606a );
 a90618a <=( (not A167)  and  A168 );
 a90619a <=( A170  and  a90618a );
 a90622a <=( A199  and  A166 );
 a90625a <=( (not A265)  and  A201 );
 a90626a <=( a90625a  and  a90622a );
 a90627a <=( a90626a  and  a90619a );
 a90631a <=( (not A269)  and  A268 );
 a90632a <=( (not A266)  and  a90631a );
 a90635a <=( (not A299)  and  A298 );
 a90638a <=( (not A302)  and  (not A300) );
 a90639a <=( a90638a  and  a90635a );
 a90640a <=( a90639a  and  a90632a );
 a90644a <=( (not A167)  and  A168 );
 a90645a <=( A170  and  a90644a );
 a90648a <=( A199  and  A166 );
 a90651a <=( (not A265)  and  A201 );
 a90652a <=( a90651a  and  a90648a );
 a90653a <=( a90652a  and  a90645a );
 a90657a <=( (not A269)  and  A268 );
 a90658a <=( (not A266)  and  a90657a );
 a90661a <=( A299  and  (not A298) );
 a90664a <=( A301  and  (not A300) );
 a90665a <=( a90664a  and  a90661a );
 a90666a <=( a90665a  and  a90658a );
 a90670a <=( (not A167)  and  A168 );
 a90671a <=( A170  and  a90670a );
 a90674a <=( A199  and  A166 );
 a90677a <=( (not A265)  and  A201 );
 a90678a <=( a90677a  and  a90674a );
 a90679a <=( a90678a  and  a90671a );
 a90683a <=( (not A269)  and  A268 );
 a90684a <=( (not A266)  and  a90683a );
 a90687a <=( A299  and  (not A298) );
 a90690a <=( (not A302)  and  (not A300) );
 a90691a <=( a90690a  and  a90687a );
 a90692a <=( a90691a  and  a90684a );
 a90696a <=( (not A167)  and  A168 );
 a90697a <=( A170  and  a90696a );
 a90700a <=( A200  and  A166 );
 a90703a <=( A265  and  A201 );
 a90704a <=( a90703a  and  a90700a );
 a90705a <=( a90704a  and  a90697a );
 a90709a <=( (not A269)  and  A268 );
 a90710a <=( A266  and  a90709a );
 a90713a <=( A299  and  A298 );
 a90716a <=( (not A301)  and  (not A300) );
 a90717a <=( a90716a  and  a90713a );
 a90718a <=( a90717a  and  a90710a );
 a90722a <=( (not A167)  and  A168 );
 a90723a <=( A170  and  a90722a );
 a90726a <=( A200  and  A166 );
 a90729a <=( A265  and  A201 );
 a90730a <=( a90729a  and  a90726a );
 a90731a <=( a90730a  and  a90723a );
 a90735a <=( (not A269)  and  A268 );
 a90736a <=( A266  and  a90735a );
 a90739a <=( A299  and  A298 );
 a90742a <=( A302  and  (not A300) );
 a90743a <=( a90742a  and  a90739a );
 a90744a <=( a90743a  and  a90736a );
 a90748a <=( (not A167)  and  A168 );
 a90749a <=( A170  and  a90748a );
 a90752a <=( A200  and  A166 );
 a90755a <=( A265  and  A201 );
 a90756a <=( a90755a  and  a90752a );
 a90757a <=( a90756a  and  a90749a );
 a90761a <=( (not A269)  and  A268 );
 a90762a <=( A266  and  a90761a );
 a90765a <=( (not A299)  and  A298 );
 a90768a <=( A301  and  (not A300) );
 a90769a <=( a90768a  and  a90765a );
 a90770a <=( a90769a  and  a90762a );
 a90774a <=( (not A167)  and  A168 );
 a90775a <=( A170  and  a90774a );
 a90778a <=( A200  and  A166 );
 a90781a <=( A265  and  A201 );
 a90782a <=( a90781a  and  a90778a );
 a90783a <=( a90782a  and  a90775a );
 a90787a <=( (not A269)  and  A268 );
 a90788a <=( A266  and  a90787a );
 a90791a <=( (not A299)  and  A298 );
 a90794a <=( (not A302)  and  (not A300) );
 a90795a <=( a90794a  and  a90791a );
 a90796a <=( a90795a  and  a90788a );
 a90800a <=( (not A167)  and  A168 );
 a90801a <=( A170  and  a90800a );
 a90804a <=( A200  and  A166 );
 a90807a <=( A265  and  A201 );
 a90808a <=( a90807a  and  a90804a );
 a90809a <=( a90808a  and  a90801a );
 a90813a <=( (not A269)  and  A268 );
 a90814a <=( A266  and  a90813a );
 a90817a <=( A299  and  (not A298) );
 a90820a <=( A301  and  (not A300) );
 a90821a <=( a90820a  and  a90817a );
 a90822a <=( a90821a  and  a90814a );
 a90826a <=( (not A167)  and  A168 );
 a90827a <=( A170  and  a90826a );
 a90830a <=( A200  and  A166 );
 a90833a <=( A265  and  A201 );
 a90834a <=( a90833a  and  a90830a );
 a90835a <=( a90834a  and  a90827a );
 a90839a <=( (not A269)  and  A268 );
 a90840a <=( A266  and  a90839a );
 a90843a <=( A299  and  (not A298) );
 a90846a <=( (not A302)  and  (not A300) );
 a90847a <=( a90846a  and  a90843a );
 a90848a <=( a90847a  and  a90840a );
 a90852a <=( (not A167)  and  A168 );
 a90853a <=( A170  and  a90852a );
 a90856a <=( A200  and  A166 );
 a90859a <=( (not A265)  and  A201 );
 a90860a <=( a90859a  and  a90856a );
 a90861a <=( a90860a  and  a90853a );
 a90865a <=( A269  and  (not A268) );
 a90866a <=( A266  and  a90865a );
 a90869a <=( A299  and  A298 );
 a90872a <=( (not A301)  and  (not A300) );
 a90873a <=( a90872a  and  a90869a );
 a90874a <=( a90873a  and  a90866a );
 a90878a <=( (not A167)  and  A168 );
 a90879a <=( A170  and  a90878a );
 a90882a <=( A200  and  A166 );
 a90885a <=( (not A265)  and  A201 );
 a90886a <=( a90885a  and  a90882a );
 a90887a <=( a90886a  and  a90879a );
 a90891a <=( A269  and  (not A268) );
 a90892a <=( A266  and  a90891a );
 a90895a <=( A299  and  A298 );
 a90898a <=( A302  and  (not A300) );
 a90899a <=( a90898a  and  a90895a );
 a90900a <=( a90899a  and  a90892a );
 a90904a <=( (not A167)  and  A168 );
 a90905a <=( A170  and  a90904a );
 a90908a <=( A200  and  A166 );
 a90911a <=( (not A265)  and  A201 );
 a90912a <=( a90911a  and  a90908a );
 a90913a <=( a90912a  and  a90905a );
 a90917a <=( A269  and  (not A268) );
 a90918a <=( A266  and  a90917a );
 a90921a <=( (not A299)  and  A298 );
 a90924a <=( A301  and  (not A300) );
 a90925a <=( a90924a  and  a90921a );
 a90926a <=( a90925a  and  a90918a );
 a90930a <=( (not A167)  and  A168 );
 a90931a <=( A170  and  a90930a );
 a90934a <=( A200  and  A166 );
 a90937a <=( (not A265)  and  A201 );
 a90938a <=( a90937a  and  a90934a );
 a90939a <=( a90938a  and  a90931a );
 a90943a <=( A269  and  (not A268) );
 a90944a <=( A266  and  a90943a );
 a90947a <=( (not A299)  and  A298 );
 a90950a <=( (not A302)  and  (not A300) );
 a90951a <=( a90950a  and  a90947a );
 a90952a <=( a90951a  and  a90944a );
 a90956a <=( (not A167)  and  A168 );
 a90957a <=( A170  and  a90956a );
 a90960a <=( A200  and  A166 );
 a90963a <=( (not A265)  and  A201 );
 a90964a <=( a90963a  and  a90960a );
 a90965a <=( a90964a  and  a90957a );
 a90969a <=( A269  and  (not A268) );
 a90970a <=( A266  and  a90969a );
 a90973a <=( A299  and  (not A298) );
 a90976a <=( A301  and  (not A300) );
 a90977a <=( a90976a  and  a90973a );
 a90978a <=( a90977a  and  a90970a );
 a90982a <=( (not A167)  and  A168 );
 a90983a <=( A170  and  a90982a );
 a90986a <=( A200  and  A166 );
 a90989a <=( (not A265)  and  A201 );
 a90990a <=( a90989a  and  a90986a );
 a90991a <=( a90990a  and  a90983a );
 a90995a <=( A269  and  (not A268) );
 a90996a <=( A266  and  a90995a );
 a90999a <=( A299  and  (not A298) );
 a91002a <=( (not A302)  and  (not A300) );
 a91003a <=( a91002a  and  a90999a );
 a91004a <=( a91003a  and  a90996a );
 a91008a <=( (not A167)  and  A168 );
 a91009a <=( A170  and  a91008a );
 a91012a <=( A200  and  A166 );
 a91015a <=( A265  and  A201 );
 a91016a <=( a91015a  and  a91012a );
 a91017a <=( a91016a  and  a91009a );
 a91021a <=( A269  and  (not A268) );
 a91022a <=( (not A266)  and  a91021a );
 a91025a <=( A299  and  A298 );
 a91028a <=( (not A301)  and  (not A300) );
 a91029a <=( a91028a  and  a91025a );
 a91030a <=( a91029a  and  a91022a );
 a91034a <=( (not A167)  and  A168 );
 a91035a <=( A170  and  a91034a );
 a91038a <=( A200  and  A166 );
 a91041a <=( A265  and  A201 );
 a91042a <=( a91041a  and  a91038a );
 a91043a <=( a91042a  and  a91035a );
 a91047a <=( A269  and  (not A268) );
 a91048a <=( (not A266)  and  a91047a );
 a91051a <=( A299  and  A298 );
 a91054a <=( A302  and  (not A300) );
 a91055a <=( a91054a  and  a91051a );
 a91056a <=( a91055a  and  a91048a );
 a91060a <=( (not A167)  and  A168 );
 a91061a <=( A170  and  a91060a );
 a91064a <=( A200  and  A166 );
 a91067a <=( A265  and  A201 );
 a91068a <=( a91067a  and  a91064a );
 a91069a <=( a91068a  and  a91061a );
 a91073a <=( A269  and  (not A268) );
 a91074a <=( (not A266)  and  a91073a );
 a91077a <=( (not A299)  and  A298 );
 a91080a <=( A301  and  (not A300) );
 a91081a <=( a91080a  and  a91077a );
 a91082a <=( a91081a  and  a91074a );
 a91086a <=( (not A167)  and  A168 );
 a91087a <=( A170  and  a91086a );
 a91090a <=( A200  and  A166 );
 a91093a <=( A265  and  A201 );
 a91094a <=( a91093a  and  a91090a );
 a91095a <=( a91094a  and  a91087a );
 a91099a <=( A269  and  (not A268) );
 a91100a <=( (not A266)  and  a91099a );
 a91103a <=( (not A299)  and  A298 );
 a91106a <=( (not A302)  and  (not A300) );
 a91107a <=( a91106a  and  a91103a );
 a91108a <=( a91107a  and  a91100a );
 a91112a <=( (not A167)  and  A168 );
 a91113a <=( A170  and  a91112a );
 a91116a <=( A200  and  A166 );
 a91119a <=( A265  and  A201 );
 a91120a <=( a91119a  and  a91116a );
 a91121a <=( a91120a  and  a91113a );
 a91125a <=( A269  and  (not A268) );
 a91126a <=( (not A266)  and  a91125a );
 a91129a <=( A299  and  (not A298) );
 a91132a <=( A301  and  (not A300) );
 a91133a <=( a91132a  and  a91129a );
 a91134a <=( a91133a  and  a91126a );
 a91138a <=( (not A167)  and  A168 );
 a91139a <=( A170  and  a91138a );
 a91142a <=( A200  and  A166 );
 a91145a <=( A265  and  A201 );
 a91146a <=( a91145a  and  a91142a );
 a91147a <=( a91146a  and  a91139a );
 a91151a <=( A269  and  (not A268) );
 a91152a <=( (not A266)  and  a91151a );
 a91155a <=( A299  and  (not A298) );
 a91158a <=( (not A302)  and  (not A300) );
 a91159a <=( a91158a  and  a91155a );
 a91160a <=( a91159a  and  a91152a );
 a91164a <=( (not A167)  and  A168 );
 a91165a <=( A170  and  a91164a );
 a91168a <=( A200  and  A166 );
 a91171a <=( (not A265)  and  A201 );
 a91172a <=( a91171a  and  a91168a );
 a91173a <=( a91172a  and  a91165a );
 a91177a <=( (not A269)  and  A268 );
 a91178a <=( (not A266)  and  a91177a );
 a91181a <=( A299  and  A298 );
 a91184a <=( (not A301)  and  (not A300) );
 a91185a <=( a91184a  and  a91181a );
 a91186a <=( a91185a  and  a91178a );
 a91190a <=( (not A167)  and  A168 );
 a91191a <=( A170  and  a91190a );
 a91194a <=( A200  and  A166 );
 a91197a <=( (not A265)  and  A201 );
 a91198a <=( a91197a  and  a91194a );
 a91199a <=( a91198a  and  a91191a );
 a91203a <=( (not A269)  and  A268 );
 a91204a <=( (not A266)  and  a91203a );
 a91207a <=( A299  and  A298 );
 a91210a <=( A302  and  (not A300) );
 a91211a <=( a91210a  and  a91207a );
 a91212a <=( a91211a  and  a91204a );
 a91216a <=( (not A167)  and  A168 );
 a91217a <=( A170  and  a91216a );
 a91220a <=( A200  and  A166 );
 a91223a <=( (not A265)  and  A201 );
 a91224a <=( a91223a  and  a91220a );
 a91225a <=( a91224a  and  a91217a );
 a91229a <=( (not A269)  and  A268 );
 a91230a <=( (not A266)  and  a91229a );
 a91233a <=( (not A299)  and  A298 );
 a91236a <=( A301  and  (not A300) );
 a91237a <=( a91236a  and  a91233a );
 a91238a <=( a91237a  and  a91230a );
 a91242a <=( (not A167)  and  A168 );
 a91243a <=( A170  and  a91242a );
 a91246a <=( A200  and  A166 );
 a91249a <=( (not A265)  and  A201 );
 a91250a <=( a91249a  and  a91246a );
 a91251a <=( a91250a  and  a91243a );
 a91255a <=( (not A269)  and  A268 );
 a91256a <=( (not A266)  and  a91255a );
 a91259a <=( (not A299)  and  A298 );
 a91262a <=( (not A302)  and  (not A300) );
 a91263a <=( a91262a  and  a91259a );
 a91264a <=( a91263a  and  a91256a );
 a91268a <=( (not A167)  and  A168 );
 a91269a <=( A170  and  a91268a );
 a91272a <=( A200  and  A166 );
 a91275a <=( (not A265)  and  A201 );
 a91276a <=( a91275a  and  a91272a );
 a91277a <=( a91276a  and  a91269a );
 a91281a <=( (not A269)  and  A268 );
 a91282a <=( (not A266)  and  a91281a );
 a91285a <=( A299  and  (not A298) );
 a91288a <=( A301  and  (not A300) );
 a91289a <=( a91288a  and  a91285a );
 a91290a <=( a91289a  and  a91282a );
 a91294a <=( (not A167)  and  A168 );
 a91295a <=( A170  and  a91294a );
 a91298a <=( A200  and  A166 );
 a91301a <=( (not A265)  and  A201 );
 a91302a <=( a91301a  and  a91298a );
 a91303a <=( a91302a  and  a91295a );
 a91307a <=( (not A269)  and  A268 );
 a91308a <=( (not A266)  and  a91307a );
 a91311a <=( A299  and  (not A298) );
 a91314a <=( (not A302)  and  (not A300) );
 a91315a <=( a91314a  and  a91311a );
 a91316a <=( a91315a  and  a91308a );
 a91320a <=( (not A167)  and  A168 );
 a91321a <=( A170  and  a91320a );
 a91324a <=( A199  and  A166 );
 a91327a <=( A202  and  A200 );
 a91328a <=( a91327a  and  a91324a );
 a91329a <=( a91328a  and  a91321a );
 a91333a <=( A267  and  A265 );
 a91334a <=( (not A203)  and  a91333a );
 a91337a <=( A299  and  A298 );
 a91340a <=( (not A301)  and  (not A300) );
 a91341a <=( a91340a  and  a91337a );
 a91342a <=( a91341a  and  a91334a );
 a91346a <=( (not A167)  and  A168 );
 a91347a <=( A170  and  a91346a );
 a91350a <=( A199  and  A166 );
 a91353a <=( A202  and  A200 );
 a91354a <=( a91353a  and  a91350a );
 a91355a <=( a91354a  and  a91347a );
 a91359a <=( A267  and  A265 );
 a91360a <=( (not A203)  and  a91359a );
 a91363a <=( A299  and  A298 );
 a91366a <=( A302  and  (not A300) );
 a91367a <=( a91366a  and  a91363a );
 a91368a <=( a91367a  and  a91360a );
 a91372a <=( (not A167)  and  A168 );
 a91373a <=( A170  and  a91372a );
 a91376a <=( A199  and  A166 );
 a91379a <=( A202  and  A200 );
 a91380a <=( a91379a  and  a91376a );
 a91381a <=( a91380a  and  a91373a );
 a91385a <=( A267  and  A265 );
 a91386a <=( (not A203)  and  a91385a );
 a91389a <=( (not A299)  and  A298 );
 a91392a <=( A301  and  (not A300) );
 a91393a <=( a91392a  and  a91389a );
 a91394a <=( a91393a  and  a91386a );
 a91398a <=( (not A167)  and  A168 );
 a91399a <=( A170  and  a91398a );
 a91402a <=( A199  and  A166 );
 a91405a <=( A202  and  A200 );
 a91406a <=( a91405a  and  a91402a );
 a91407a <=( a91406a  and  a91399a );
 a91411a <=( A267  and  A265 );
 a91412a <=( (not A203)  and  a91411a );
 a91415a <=( (not A299)  and  A298 );
 a91418a <=( (not A302)  and  (not A300) );
 a91419a <=( a91418a  and  a91415a );
 a91420a <=( a91419a  and  a91412a );
 a91424a <=( (not A167)  and  A168 );
 a91425a <=( A170  and  a91424a );
 a91428a <=( A199  and  A166 );
 a91431a <=( A202  and  A200 );
 a91432a <=( a91431a  and  a91428a );
 a91433a <=( a91432a  and  a91425a );
 a91437a <=( A267  and  A265 );
 a91438a <=( (not A203)  and  a91437a );
 a91441a <=( A299  and  (not A298) );
 a91444a <=( A301  and  (not A300) );
 a91445a <=( a91444a  and  a91441a );
 a91446a <=( a91445a  and  a91438a );
 a91450a <=( (not A167)  and  A168 );
 a91451a <=( A170  and  a91450a );
 a91454a <=( A199  and  A166 );
 a91457a <=( A202  and  A200 );
 a91458a <=( a91457a  and  a91454a );
 a91459a <=( a91458a  and  a91451a );
 a91463a <=( A267  and  A265 );
 a91464a <=( (not A203)  and  a91463a );
 a91467a <=( A299  and  (not A298) );
 a91470a <=( (not A302)  and  (not A300) );
 a91471a <=( a91470a  and  a91467a );
 a91472a <=( a91471a  and  a91464a );
 a91476a <=( (not A167)  and  A168 );
 a91477a <=( A170  and  a91476a );
 a91480a <=( A199  and  A166 );
 a91483a <=( A202  and  A200 );
 a91484a <=( a91483a  and  a91480a );
 a91485a <=( a91484a  and  a91477a );
 a91489a <=( A267  and  A266 );
 a91490a <=( (not A203)  and  a91489a );
 a91493a <=( A299  and  A298 );
 a91496a <=( (not A301)  and  (not A300) );
 a91497a <=( a91496a  and  a91493a );
 a91498a <=( a91497a  and  a91490a );
 a91502a <=( (not A167)  and  A168 );
 a91503a <=( A170  and  a91502a );
 a91506a <=( A199  and  A166 );
 a91509a <=( A202  and  A200 );
 a91510a <=( a91509a  and  a91506a );
 a91511a <=( a91510a  and  a91503a );
 a91515a <=( A267  and  A266 );
 a91516a <=( (not A203)  and  a91515a );
 a91519a <=( A299  and  A298 );
 a91522a <=( A302  and  (not A300) );
 a91523a <=( a91522a  and  a91519a );
 a91524a <=( a91523a  and  a91516a );
 a91528a <=( (not A167)  and  A168 );
 a91529a <=( A170  and  a91528a );
 a91532a <=( A199  and  A166 );
 a91535a <=( A202  and  A200 );
 a91536a <=( a91535a  and  a91532a );
 a91537a <=( a91536a  and  a91529a );
 a91541a <=( A267  and  A266 );
 a91542a <=( (not A203)  and  a91541a );
 a91545a <=( (not A299)  and  A298 );
 a91548a <=( A301  and  (not A300) );
 a91549a <=( a91548a  and  a91545a );
 a91550a <=( a91549a  and  a91542a );
 a91554a <=( (not A167)  and  A168 );
 a91555a <=( A170  and  a91554a );
 a91558a <=( A199  and  A166 );
 a91561a <=( A202  and  A200 );
 a91562a <=( a91561a  and  a91558a );
 a91563a <=( a91562a  and  a91555a );
 a91567a <=( A267  and  A266 );
 a91568a <=( (not A203)  and  a91567a );
 a91571a <=( (not A299)  and  A298 );
 a91574a <=( (not A302)  and  (not A300) );
 a91575a <=( a91574a  and  a91571a );
 a91576a <=( a91575a  and  a91568a );
 a91580a <=( (not A167)  and  A168 );
 a91581a <=( A170  and  a91580a );
 a91584a <=( A199  and  A166 );
 a91587a <=( A202  and  A200 );
 a91588a <=( a91587a  and  a91584a );
 a91589a <=( a91588a  and  a91581a );
 a91593a <=( A267  and  A266 );
 a91594a <=( (not A203)  and  a91593a );
 a91597a <=( A299  and  (not A298) );
 a91600a <=( A301  and  (not A300) );
 a91601a <=( a91600a  and  a91597a );
 a91602a <=( a91601a  and  a91594a );
 a91606a <=( (not A167)  and  A168 );
 a91607a <=( A170  and  a91606a );
 a91610a <=( A199  and  A166 );
 a91613a <=( A202  and  A200 );
 a91614a <=( a91613a  and  a91610a );
 a91615a <=( a91614a  and  a91607a );
 a91619a <=( A267  and  A266 );
 a91620a <=( (not A203)  and  a91619a );
 a91623a <=( A299  and  (not A298) );
 a91626a <=( (not A302)  and  (not A300) );
 a91627a <=( a91626a  and  a91623a );
 a91628a <=( a91627a  and  a91620a );
 a91632a <=( (not A167)  and  A168 );
 a91633a <=( A170  and  a91632a );
 a91636a <=( A199  and  A166 );
 a91639a <=( (not A201)  and  A200 );
 a91640a <=( a91639a  and  a91636a );
 a91641a <=( a91640a  and  a91633a );
 a91645a <=( A266  and  A265 );
 a91646a <=( (not A202)  and  a91645a );
 a91649a <=( (not A268)  and  (not A267) );
 a91652a <=( A300  and  A299 );
 a91653a <=( a91652a  and  a91649a );
 a91654a <=( a91653a  and  a91646a );
 a91658a <=( (not A167)  and  A168 );
 a91659a <=( A170  and  a91658a );
 a91662a <=( A199  and  A166 );
 a91665a <=( (not A201)  and  A200 );
 a91666a <=( a91665a  and  a91662a );
 a91667a <=( a91666a  and  a91659a );
 a91671a <=( A266  and  A265 );
 a91672a <=( (not A202)  and  a91671a );
 a91675a <=( (not A268)  and  (not A267) );
 a91678a <=( A300  and  A298 );
 a91679a <=( a91678a  and  a91675a );
 a91680a <=( a91679a  and  a91672a );
 a91684a <=( (not A167)  and  A168 );
 a91685a <=( A170  and  a91684a );
 a91688a <=( A199  and  A166 );
 a91691a <=( (not A201)  and  A200 );
 a91692a <=( a91691a  and  a91688a );
 a91693a <=( a91692a  and  a91685a );
 a91697a <=( A266  and  A265 );
 a91698a <=( (not A202)  and  a91697a );
 a91701a <=( A269  and  (not A267) );
 a91704a <=( A300  and  A299 );
 a91705a <=( a91704a  and  a91701a );
 a91706a <=( a91705a  and  a91698a );
 a91710a <=( (not A167)  and  A168 );
 a91711a <=( A170  and  a91710a );
 a91714a <=( A199  and  A166 );
 a91717a <=( (not A201)  and  A200 );
 a91718a <=( a91717a  and  a91714a );
 a91719a <=( a91718a  and  a91711a );
 a91723a <=( A266  and  A265 );
 a91724a <=( (not A202)  and  a91723a );
 a91727a <=( A269  and  (not A267) );
 a91730a <=( A300  and  A298 );
 a91731a <=( a91730a  and  a91727a );
 a91732a <=( a91731a  and  a91724a );
 a91736a <=( (not A167)  and  A168 );
 a91737a <=( A170  and  a91736a );
 a91740a <=( A199  and  A166 );
 a91743a <=( (not A201)  and  A200 );
 a91744a <=( a91743a  and  a91740a );
 a91745a <=( a91744a  and  a91737a );
 a91749a <=( A266  and  (not A265) );
 a91750a <=( (not A202)  and  a91749a );
 a91753a <=( A268  and  (not A267) );
 a91756a <=( A300  and  A299 );
 a91757a <=( a91756a  and  a91753a );
 a91758a <=( a91757a  and  a91750a );
 a91762a <=( (not A167)  and  A168 );
 a91763a <=( A170  and  a91762a );
 a91766a <=( A199  and  A166 );
 a91769a <=( (not A201)  and  A200 );
 a91770a <=( a91769a  and  a91766a );
 a91771a <=( a91770a  and  a91763a );
 a91775a <=( A266  and  (not A265) );
 a91776a <=( (not A202)  and  a91775a );
 a91779a <=( A268  and  (not A267) );
 a91782a <=( A300  and  A298 );
 a91783a <=( a91782a  and  a91779a );
 a91784a <=( a91783a  and  a91776a );
 a91788a <=( (not A167)  and  A168 );
 a91789a <=( A170  and  a91788a );
 a91792a <=( A199  and  A166 );
 a91795a <=( (not A201)  and  A200 );
 a91796a <=( a91795a  and  a91792a );
 a91797a <=( a91796a  and  a91789a );
 a91801a <=( A266  and  (not A265) );
 a91802a <=( (not A202)  and  a91801a );
 a91805a <=( (not A269)  and  (not A267) );
 a91808a <=( A300  and  A299 );
 a91809a <=( a91808a  and  a91805a );
 a91810a <=( a91809a  and  a91802a );
 a91814a <=( (not A167)  and  A168 );
 a91815a <=( A170  and  a91814a );
 a91818a <=( A199  and  A166 );
 a91821a <=( (not A201)  and  A200 );
 a91822a <=( a91821a  and  a91818a );
 a91823a <=( a91822a  and  a91815a );
 a91827a <=( A266  and  (not A265) );
 a91828a <=( (not A202)  and  a91827a );
 a91831a <=( (not A269)  and  (not A267) );
 a91834a <=( A300  and  A298 );
 a91835a <=( a91834a  and  a91831a );
 a91836a <=( a91835a  and  a91828a );
 a91840a <=( (not A167)  and  A168 );
 a91841a <=( A170  and  a91840a );
 a91844a <=( A199  and  A166 );
 a91847a <=( (not A201)  and  A200 );
 a91848a <=( a91847a  and  a91844a );
 a91849a <=( a91848a  and  a91841a );
 a91853a <=( (not A266)  and  A265 );
 a91854a <=( (not A202)  and  a91853a );
 a91857a <=( A268  and  (not A267) );
 a91860a <=( A300  and  A299 );
 a91861a <=( a91860a  and  a91857a );
 a91862a <=( a91861a  and  a91854a );
 a91866a <=( (not A167)  and  A168 );
 a91867a <=( A170  and  a91866a );
 a91870a <=( A199  and  A166 );
 a91873a <=( (not A201)  and  A200 );
 a91874a <=( a91873a  and  a91870a );
 a91875a <=( a91874a  and  a91867a );
 a91879a <=( (not A266)  and  A265 );
 a91880a <=( (not A202)  and  a91879a );
 a91883a <=( A268  and  (not A267) );
 a91886a <=( A300  and  A298 );
 a91887a <=( a91886a  and  a91883a );
 a91888a <=( a91887a  and  a91880a );
 a91892a <=( (not A167)  and  A168 );
 a91893a <=( A170  and  a91892a );
 a91896a <=( A199  and  A166 );
 a91899a <=( (not A201)  and  A200 );
 a91900a <=( a91899a  and  a91896a );
 a91901a <=( a91900a  and  a91893a );
 a91905a <=( (not A266)  and  A265 );
 a91906a <=( (not A202)  and  a91905a );
 a91909a <=( (not A269)  and  (not A267) );
 a91912a <=( A300  and  A299 );
 a91913a <=( a91912a  and  a91909a );
 a91914a <=( a91913a  and  a91906a );
 a91918a <=( (not A167)  and  A168 );
 a91919a <=( A170  and  a91918a );
 a91922a <=( A199  and  A166 );
 a91925a <=( (not A201)  and  A200 );
 a91926a <=( a91925a  and  a91922a );
 a91927a <=( a91926a  and  a91919a );
 a91931a <=( (not A266)  and  A265 );
 a91932a <=( (not A202)  and  a91931a );
 a91935a <=( (not A269)  and  (not A267) );
 a91938a <=( A300  and  A298 );
 a91939a <=( a91938a  and  a91935a );
 a91940a <=( a91939a  and  a91932a );
 a91944a <=( (not A167)  and  A168 );
 a91945a <=( A170  and  a91944a );
 a91948a <=( A199  and  A166 );
 a91951a <=( (not A201)  and  A200 );
 a91952a <=( a91951a  and  a91948a );
 a91953a <=( a91952a  and  a91945a );
 a91957a <=( A266  and  A265 );
 a91958a <=( A203  and  a91957a );
 a91961a <=( (not A268)  and  (not A267) );
 a91964a <=( A300  and  A299 );
 a91965a <=( a91964a  and  a91961a );
 a91966a <=( a91965a  and  a91958a );
 a91970a <=( (not A167)  and  A168 );
 a91971a <=( A170  and  a91970a );
 a91974a <=( A199  and  A166 );
 a91977a <=( (not A201)  and  A200 );
 a91978a <=( a91977a  and  a91974a );
 a91979a <=( a91978a  and  a91971a );
 a91983a <=( A266  and  A265 );
 a91984a <=( A203  and  a91983a );
 a91987a <=( (not A268)  and  (not A267) );
 a91990a <=( A300  and  A298 );
 a91991a <=( a91990a  and  a91987a );
 a91992a <=( a91991a  and  a91984a );
 a91996a <=( (not A167)  and  A168 );
 a91997a <=( A170  and  a91996a );
 a92000a <=( A199  and  A166 );
 a92003a <=( (not A201)  and  A200 );
 a92004a <=( a92003a  and  a92000a );
 a92005a <=( a92004a  and  a91997a );
 a92009a <=( A266  and  A265 );
 a92010a <=( A203  and  a92009a );
 a92013a <=( A269  and  (not A267) );
 a92016a <=( A300  and  A299 );
 a92017a <=( a92016a  and  a92013a );
 a92018a <=( a92017a  and  a92010a );
 a92022a <=( (not A167)  and  A168 );
 a92023a <=( A170  and  a92022a );
 a92026a <=( A199  and  A166 );
 a92029a <=( (not A201)  and  A200 );
 a92030a <=( a92029a  and  a92026a );
 a92031a <=( a92030a  and  a92023a );
 a92035a <=( A266  and  A265 );
 a92036a <=( A203  and  a92035a );
 a92039a <=( A269  and  (not A267) );
 a92042a <=( A300  and  A298 );
 a92043a <=( a92042a  and  a92039a );
 a92044a <=( a92043a  and  a92036a );
 a92048a <=( (not A167)  and  A168 );
 a92049a <=( A170  and  a92048a );
 a92052a <=( A199  and  A166 );
 a92055a <=( (not A201)  and  A200 );
 a92056a <=( a92055a  and  a92052a );
 a92057a <=( a92056a  and  a92049a );
 a92061a <=( A266  and  (not A265) );
 a92062a <=( A203  and  a92061a );
 a92065a <=( A268  and  (not A267) );
 a92068a <=( A300  and  A299 );
 a92069a <=( a92068a  and  a92065a );
 a92070a <=( a92069a  and  a92062a );
 a92074a <=( (not A167)  and  A168 );
 a92075a <=( A170  and  a92074a );
 a92078a <=( A199  and  A166 );
 a92081a <=( (not A201)  and  A200 );
 a92082a <=( a92081a  and  a92078a );
 a92083a <=( a92082a  and  a92075a );
 a92087a <=( A266  and  (not A265) );
 a92088a <=( A203  and  a92087a );
 a92091a <=( A268  and  (not A267) );
 a92094a <=( A300  and  A298 );
 a92095a <=( a92094a  and  a92091a );
 a92096a <=( a92095a  and  a92088a );
 a92100a <=( (not A167)  and  A168 );
 a92101a <=( A170  and  a92100a );
 a92104a <=( A199  and  A166 );
 a92107a <=( (not A201)  and  A200 );
 a92108a <=( a92107a  and  a92104a );
 a92109a <=( a92108a  and  a92101a );
 a92113a <=( A266  and  (not A265) );
 a92114a <=( A203  and  a92113a );
 a92117a <=( (not A269)  and  (not A267) );
 a92120a <=( A300  and  A299 );
 a92121a <=( a92120a  and  a92117a );
 a92122a <=( a92121a  and  a92114a );
 a92126a <=( (not A167)  and  A168 );
 a92127a <=( A170  and  a92126a );
 a92130a <=( A199  and  A166 );
 a92133a <=( (not A201)  and  A200 );
 a92134a <=( a92133a  and  a92130a );
 a92135a <=( a92134a  and  a92127a );
 a92139a <=( A266  and  (not A265) );
 a92140a <=( A203  and  a92139a );
 a92143a <=( (not A269)  and  (not A267) );
 a92146a <=( A300  and  A298 );
 a92147a <=( a92146a  and  a92143a );
 a92148a <=( a92147a  and  a92140a );
 a92152a <=( (not A167)  and  A168 );
 a92153a <=( A170  and  a92152a );
 a92156a <=( A199  and  A166 );
 a92159a <=( (not A201)  and  A200 );
 a92160a <=( a92159a  and  a92156a );
 a92161a <=( a92160a  and  a92153a );
 a92165a <=( (not A266)  and  A265 );
 a92166a <=( A203  and  a92165a );
 a92169a <=( A268  and  (not A267) );
 a92172a <=( A300  and  A299 );
 a92173a <=( a92172a  and  a92169a );
 a92174a <=( a92173a  and  a92166a );
 a92178a <=( (not A167)  and  A168 );
 a92179a <=( A170  and  a92178a );
 a92182a <=( A199  and  A166 );
 a92185a <=( (not A201)  and  A200 );
 a92186a <=( a92185a  and  a92182a );
 a92187a <=( a92186a  and  a92179a );
 a92191a <=( (not A266)  and  A265 );
 a92192a <=( A203  and  a92191a );
 a92195a <=( A268  and  (not A267) );
 a92198a <=( A300  and  A298 );
 a92199a <=( a92198a  and  a92195a );
 a92200a <=( a92199a  and  a92192a );
 a92204a <=( (not A167)  and  A168 );
 a92205a <=( A170  and  a92204a );
 a92208a <=( A199  and  A166 );
 a92211a <=( (not A201)  and  A200 );
 a92212a <=( a92211a  and  a92208a );
 a92213a <=( a92212a  and  a92205a );
 a92217a <=( (not A266)  and  A265 );
 a92218a <=( A203  and  a92217a );
 a92221a <=( (not A269)  and  (not A267) );
 a92224a <=( A300  and  A299 );
 a92225a <=( a92224a  and  a92221a );
 a92226a <=( a92225a  and  a92218a );
 a92230a <=( (not A167)  and  A168 );
 a92231a <=( A170  and  a92230a );
 a92234a <=( A199  and  A166 );
 a92237a <=( (not A201)  and  A200 );
 a92238a <=( a92237a  and  a92234a );
 a92239a <=( a92238a  and  a92231a );
 a92243a <=( (not A266)  and  A265 );
 a92244a <=( A203  and  a92243a );
 a92247a <=( (not A269)  and  (not A267) );
 a92250a <=( A300  and  A298 );
 a92251a <=( a92250a  and  a92247a );
 a92252a <=( a92251a  and  a92244a );
 a92256a <=( (not A167)  and  A168 );
 a92257a <=( A170  and  a92256a );
 a92260a <=( (not A199)  and  A166 );
 a92263a <=( (not A202)  and  A200 );
 a92264a <=( a92263a  and  a92260a );
 a92265a <=( a92264a  and  a92257a );
 a92269a <=( A267  and  A265 );
 a92270a <=( A203  and  a92269a );
 a92273a <=( A299  and  A298 );
 a92276a <=( (not A301)  and  (not A300) );
 a92277a <=( a92276a  and  a92273a );
 a92278a <=( a92277a  and  a92270a );
 a92282a <=( (not A167)  and  A168 );
 a92283a <=( A170  and  a92282a );
 a92286a <=( (not A199)  and  A166 );
 a92289a <=( (not A202)  and  A200 );
 a92290a <=( a92289a  and  a92286a );
 a92291a <=( a92290a  and  a92283a );
 a92295a <=( A267  and  A265 );
 a92296a <=( A203  and  a92295a );
 a92299a <=( A299  and  A298 );
 a92302a <=( A302  and  (not A300) );
 a92303a <=( a92302a  and  a92299a );
 a92304a <=( a92303a  and  a92296a );
 a92308a <=( (not A167)  and  A168 );
 a92309a <=( A170  and  a92308a );
 a92312a <=( (not A199)  and  A166 );
 a92315a <=( (not A202)  and  A200 );
 a92316a <=( a92315a  and  a92312a );
 a92317a <=( a92316a  and  a92309a );
 a92321a <=( A267  and  A265 );
 a92322a <=( A203  and  a92321a );
 a92325a <=( (not A299)  and  A298 );
 a92328a <=( A301  and  (not A300) );
 a92329a <=( a92328a  and  a92325a );
 a92330a <=( a92329a  and  a92322a );
 a92334a <=( (not A167)  and  A168 );
 a92335a <=( A170  and  a92334a );
 a92338a <=( (not A199)  and  A166 );
 a92341a <=( (not A202)  and  A200 );
 a92342a <=( a92341a  and  a92338a );
 a92343a <=( a92342a  and  a92335a );
 a92347a <=( A267  and  A265 );
 a92348a <=( A203  and  a92347a );
 a92351a <=( (not A299)  and  A298 );
 a92354a <=( (not A302)  and  (not A300) );
 a92355a <=( a92354a  and  a92351a );
 a92356a <=( a92355a  and  a92348a );
 a92360a <=( (not A167)  and  A168 );
 a92361a <=( A170  and  a92360a );
 a92364a <=( (not A199)  and  A166 );
 a92367a <=( (not A202)  and  A200 );
 a92368a <=( a92367a  and  a92364a );
 a92369a <=( a92368a  and  a92361a );
 a92373a <=( A267  and  A265 );
 a92374a <=( A203  and  a92373a );
 a92377a <=( A299  and  (not A298) );
 a92380a <=( A301  and  (not A300) );
 a92381a <=( a92380a  and  a92377a );
 a92382a <=( a92381a  and  a92374a );
 a92386a <=( (not A167)  and  A168 );
 a92387a <=( A170  and  a92386a );
 a92390a <=( (not A199)  and  A166 );
 a92393a <=( (not A202)  and  A200 );
 a92394a <=( a92393a  and  a92390a );
 a92395a <=( a92394a  and  a92387a );
 a92399a <=( A267  and  A265 );
 a92400a <=( A203  and  a92399a );
 a92403a <=( A299  and  (not A298) );
 a92406a <=( (not A302)  and  (not A300) );
 a92407a <=( a92406a  and  a92403a );
 a92408a <=( a92407a  and  a92400a );
 a92412a <=( (not A167)  and  A168 );
 a92413a <=( A170  and  a92412a );
 a92416a <=( (not A199)  and  A166 );
 a92419a <=( (not A202)  and  A200 );
 a92420a <=( a92419a  and  a92416a );
 a92421a <=( a92420a  and  a92413a );
 a92425a <=( A267  and  A266 );
 a92426a <=( A203  and  a92425a );
 a92429a <=( A299  and  A298 );
 a92432a <=( (not A301)  and  (not A300) );
 a92433a <=( a92432a  and  a92429a );
 a92434a <=( a92433a  and  a92426a );
 a92438a <=( (not A167)  and  A168 );
 a92439a <=( A170  and  a92438a );
 a92442a <=( (not A199)  and  A166 );
 a92445a <=( (not A202)  and  A200 );
 a92446a <=( a92445a  and  a92442a );
 a92447a <=( a92446a  and  a92439a );
 a92451a <=( A267  and  A266 );
 a92452a <=( A203  and  a92451a );
 a92455a <=( A299  and  A298 );
 a92458a <=( A302  and  (not A300) );
 a92459a <=( a92458a  and  a92455a );
 a92460a <=( a92459a  and  a92452a );
 a92464a <=( (not A167)  and  A168 );
 a92465a <=( A170  and  a92464a );
 a92468a <=( (not A199)  and  A166 );
 a92471a <=( (not A202)  and  A200 );
 a92472a <=( a92471a  and  a92468a );
 a92473a <=( a92472a  and  a92465a );
 a92477a <=( A267  and  A266 );
 a92478a <=( A203  and  a92477a );
 a92481a <=( (not A299)  and  A298 );
 a92484a <=( A301  and  (not A300) );
 a92485a <=( a92484a  and  a92481a );
 a92486a <=( a92485a  and  a92478a );
 a92490a <=( (not A167)  and  A168 );
 a92491a <=( A170  and  a92490a );
 a92494a <=( (not A199)  and  A166 );
 a92497a <=( (not A202)  and  A200 );
 a92498a <=( a92497a  and  a92494a );
 a92499a <=( a92498a  and  a92491a );
 a92503a <=( A267  and  A266 );
 a92504a <=( A203  and  a92503a );
 a92507a <=( (not A299)  and  A298 );
 a92510a <=( (not A302)  and  (not A300) );
 a92511a <=( a92510a  and  a92507a );
 a92512a <=( a92511a  and  a92504a );
 a92516a <=( (not A167)  and  A168 );
 a92517a <=( A170  and  a92516a );
 a92520a <=( (not A199)  and  A166 );
 a92523a <=( (not A202)  and  A200 );
 a92524a <=( a92523a  and  a92520a );
 a92525a <=( a92524a  and  a92517a );
 a92529a <=( A267  and  A266 );
 a92530a <=( A203  and  a92529a );
 a92533a <=( A299  and  (not A298) );
 a92536a <=( A301  and  (not A300) );
 a92537a <=( a92536a  and  a92533a );
 a92538a <=( a92537a  and  a92530a );
 a92542a <=( (not A167)  and  A168 );
 a92543a <=( A170  and  a92542a );
 a92546a <=( (not A199)  and  A166 );
 a92549a <=( (not A202)  and  A200 );
 a92550a <=( a92549a  and  a92546a );
 a92551a <=( a92550a  and  a92543a );
 a92555a <=( A267  and  A266 );
 a92556a <=( A203  and  a92555a );
 a92559a <=( A299  and  (not A298) );
 a92562a <=( (not A302)  and  (not A300) );
 a92563a <=( a92562a  and  a92559a );
 a92564a <=( a92563a  and  a92556a );
 a92568a <=( (not A167)  and  A168 );
 a92569a <=( A170  and  a92568a );
 a92572a <=( (not A199)  and  A166 );
 a92575a <=( (not A201)  and  A200 );
 a92576a <=( a92575a  and  a92572a );
 a92577a <=( a92576a  and  a92569a );
 a92581a <=( A266  and  A265 );
 a92582a <=( A202  and  a92581a );
 a92585a <=( (not A268)  and  (not A267) );
 a92588a <=( A300  and  A299 );
 a92589a <=( a92588a  and  a92585a );
 a92590a <=( a92589a  and  a92582a );
 a92594a <=( (not A167)  and  A168 );
 a92595a <=( A170  and  a92594a );
 a92598a <=( (not A199)  and  A166 );
 a92601a <=( (not A201)  and  A200 );
 a92602a <=( a92601a  and  a92598a );
 a92603a <=( a92602a  and  a92595a );
 a92607a <=( A266  and  A265 );
 a92608a <=( A202  and  a92607a );
 a92611a <=( (not A268)  and  (not A267) );
 a92614a <=( A300  and  A298 );
 a92615a <=( a92614a  and  a92611a );
 a92616a <=( a92615a  and  a92608a );
 a92620a <=( (not A167)  and  A168 );
 a92621a <=( A170  and  a92620a );
 a92624a <=( (not A199)  and  A166 );
 a92627a <=( (not A201)  and  A200 );
 a92628a <=( a92627a  and  a92624a );
 a92629a <=( a92628a  and  a92621a );
 a92633a <=( A266  and  A265 );
 a92634a <=( A202  and  a92633a );
 a92637a <=( A269  and  (not A267) );
 a92640a <=( A300  and  A299 );
 a92641a <=( a92640a  and  a92637a );
 a92642a <=( a92641a  and  a92634a );
 a92646a <=( (not A167)  and  A168 );
 a92647a <=( A170  and  a92646a );
 a92650a <=( (not A199)  and  A166 );
 a92653a <=( (not A201)  and  A200 );
 a92654a <=( a92653a  and  a92650a );
 a92655a <=( a92654a  and  a92647a );
 a92659a <=( A266  and  A265 );
 a92660a <=( A202  and  a92659a );
 a92663a <=( A269  and  (not A267) );
 a92666a <=( A300  and  A298 );
 a92667a <=( a92666a  and  a92663a );
 a92668a <=( a92667a  and  a92660a );
 a92672a <=( (not A167)  and  A168 );
 a92673a <=( A170  and  a92672a );
 a92676a <=( (not A199)  and  A166 );
 a92679a <=( (not A201)  and  A200 );
 a92680a <=( a92679a  and  a92676a );
 a92681a <=( a92680a  and  a92673a );
 a92685a <=( A266  and  (not A265) );
 a92686a <=( A202  and  a92685a );
 a92689a <=( A268  and  (not A267) );
 a92692a <=( A300  and  A299 );
 a92693a <=( a92692a  and  a92689a );
 a92694a <=( a92693a  and  a92686a );
 a92698a <=( (not A167)  and  A168 );
 a92699a <=( A170  and  a92698a );
 a92702a <=( (not A199)  and  A166 );
 a92705a <=( (not A201)  and  A200 );
 a92706a <=( a92705a  and  a92702a );
 a92707a <=( a92706a  and  a92699a );
 a92711a <=( A266  and  (not A265) );
 a92712a <=( A202  and  a92711a );
 a92715a <=( A268  and  (not A267) );
 a92718a <=( A300  and  A298 );
 a92719a <=( a92718a  and  a92715a );
 a92720a <=( a92719a  and  a92712a );
 a92724a <=( (not A167)  and  A168 );
 a92725a <=( A170  and  a92724a );
 a92728a <=( (not A199)  and  A166 );
 a92731a <=( (not A201)  and  A200 );
 a92732a <=( a92731a  and  a92728a );
 a92733a <=( a92732a  and  a92725a );
 a92737a <=( A266  and  (not A265) );
 a92738a <=( A202  and  a92737a );
 a92741a <=( (not A269)  and  (not A267) );
 a92744a <=( A300  and  A299 );
 a92745a <=( a92744a  and  a92741a );
 a92746a <=( a92745a  and  a92738a );
 a92750a <=( (not A167)  and  A168 );
 a92751a <=( A170  and  a92750a );
 a92754a <=( (not A199)  and  A166 );
 a92757a <=( (not A201)  and  A200 );
 a92758a <=( a92757a  and  a92754a );
 a92759a <=( a92758a  and  a92751a );
 a92763a <=( A266  and  (not A265) );
 a92764a <=( A202  and  a92763a );
 a92767a <=( (not A269)  and  (not A267) );
 a92770a <=( A300  and  A298 );
 a92771a <=( a92770a  and  a92767a );
 a92772a <=( a92771a  and  a92764a );
 a92776a <=( (not A167)  and  A168 );
 a92777a <=( A170  and  a92776a );
 a92780a <=( (not A199)  and  A166 );
 a92783a <=( (not A201)  and  A200 );
 a92784a <=( a92783a  and  a92780a );
 a92785a <=( a92784a  and  a92777a );
 a92789a <=( (not A266)  and  A265 );
 a92790a <=( A202  and  a92789a );
 a92793a <=( A268  and  (not A267) );
 a92796a <=( A300  and  A299 );
 a92797a <=( a92796a  and  a92793a );
 a92798a <=( a92797a  and  a92790a );
 a92802a <=( (not A167)  and  A168 );
 a92803a <=( A170  and  a92802a );
 a92806a <=( (not A199)  and  A166 );
 a92809a <=( (not A201)  and  A200 );
 a92810a <=( a92809a  and  a92806a );
 a92811a <=( a92810a  and  a92803a );
 a92815a <=( (not A266)  and  A265 );
 a92816a <=( A202  and  a92815a );
 a92819a <=( A268  and  (not A267) );
 a92822a <=( A300  and  A298 );
 a92823a <=( a92822a  and  a92819a );
 a92824a <=( a92823a  and  a92816a );
 a92828a <=( (not A167)  and  A168 );
 a92829a <=( A170  and  a92828a );
 a92832a <=( (not A199)  and  A166 );
 a92835a <=( (not A201)  and  A200 );
 a92836a <=( a92835a  and  a92832a );
 a92837a <=( a92836a  and  a92829a );
 a92841a <=( (not A266)  and  A265 );
 a92842a <=( A202  and  a92841a );
 a92845a <=( (not A269)  and  (not A267) );
 a92848a <=( A300  and  A299 );
 a92849a <=( a92848a  and  a92845a );
 a92850a <=( a92849a  and  a92842a );
 a92854a <=( (not A167)  and  A168 );
 a92855a <=( A170  and  a92854a );
 a92858a <=( (not A199)  and  A166 );
 a92861a <=( (not A201)  and  A200 );
 a92862a <=( a92861a  and  a92858a );
 a92863a <=( a92862a  and  a92855a );
 a92867a <=( (not A266)  and  A265 );
 a92868a <=( A202  and  a92867a );
 a92871a <=( (not A269)  and  (not A267) );
 a92874a <=( A300  and  A298 );
 a92875a <=( a92874a  and  a92871a );
 a92876a <=( a92875a  and  a92868a );
 a92880a <=( (not A167)  and  A168 );
 a92881a <=( A170  and  a92880a );
 a92884a <=( (not A199)  and  A166 );
 a92887a <=( (not A201)  and  A200 );
 a92888a <=( a92887a  and  a92884a );
 a92889a <=( a92888a  and  a92881a );
 a92893a <=( A266  and  A265 );
 a92894a <=( (not A203)  and  a92893a );
 a92897a <=( (not A268)  and  (not A267) );
 a92900a <=( A300  and  A299 );
 a92901a <=( a92900a  and  a92897a );
 a92902a <=( a92901a  and  a92894a );
 a92906a <=( (not A167)  and  A168 );
 a92907a <=( A170  and  a92906a );
 a92910a <=( (not A199)  and  A166 );
 a92913a <=( (not A201)  and  A200 );
 a92914a <=( a92913a  and  a92910a );
 a92915a <=( a92914a  and  a92907a );
 a92919a <=( A266  and  A265 );
 a92920a <=( (not A203)  and  a92919a );
 a92923a <=( (not A268)  and  (not A267) );
 a92926a <=( A300  and  A298 );
 a92927a <=( a92926a  and  a92923a );
 a92928a <=( a92927a  and  a92920a );
 a92932a <=( (not A167)  and  A168 );
 a92933a <=( A170  and  a92932a );
 a92936a <=( (not A199)  and  A166 );
 a92939a <=( (not A201)  and  A200 );
 a92940a <=( a92939a  and  a92936a );
 a92941a <=( a92940a  and  a92933a );
 a92945a <=( A266  and  A265 );
 a92946a <=( (not A203)  and  a92945a );
 a92949a <=( A269  and  (not A267) );
 a92952a <=( A300  and  A299 );
 a92953a <=( a92952a  and  a92949a );
 a92954a <=( a92953a  and  a92946a );
 a92958a <=( (not A167)  and  A168 );
 a92959a <=( A170  and  a92958a );
 a92962a <=( (not A199)  and  A166 );
 a92965a <=( (not A201)  and  A200 );
 a92966a <=( a92965a  and  a92962a );
 a92967a <=( a92966a  and  a92959a );
 a92971a <=( A266  and  A265 );
 a92972a <=( (not A203)  and  a92971a );
 a92975a <=( A269  and  (not A267) );
 a92978a <=( A300  and  A298 );
 a92979a <=( a92978a  and  a92975a );
 a92980a <=( a92979a  and  a92972a );
 a92984a <=( (not A167)  and  A168 );
 a92985a <=( A170  and  a92984a );
 a92988a <=( (not A199)  and  A166 );
 a92991a <=( (not A201)  and  A200 );
 a92992a <=( a92991a  and  a92988a );
 a92993a <=( a92992a  and  a92985a );
 a92997a <=( A266  and  (not A265) );
 a92998a <=( (not A203)  and  a92997a );
 a93001a <=( A268  and  (not A267) );
 a93004a <=( A300  and  A299 );
 a93005a <=( a93004a  and  a93001a );
 a93006a <=( a93005a  and  a92998a );
 a93010a <=( (not A167)  and  A168 );
 a93011a <=( A170  and  a93010a );
 a93014a <=( (not A199)  and  A166 );
 a93017a <=( (not A201)  and  A200 );
 a93018a <=( a93017a  and  a93014a );
 a93019a <=( a93018a  and  a93011a );
 a93023a <=( A266  and  (not A265) );
 a93024a <=( (not A203)  and  a93023a );
 a93027a <=( A268  and  (not A267) );
 a93030a <=( A300  and  A298 );
 a93031a <=( a93030a  and  a93027a );
 a93032a <=( a93031a  and  a93024a );
 a93036a <=( (not A167)  and  A168 );
 a93037a <=( A170  and  a93036a );
 a93040a <=( (not A199)  and  A166 );
 a93043a <=( (not A201)  and  A200 );
 a93044a <=( a93043a  and  a93040a );
 a93045a <=( a93044a  and  a93037a );
 a93049a <=( A266  and  (not A265) );
 a93050a <=( (not A203)  and  a93049a );
 a93053a <=( (not A269)  and  (not A267) );
 a93056a <=( A300  and  A299 );
 a93057a <=( a93056a  and  a93053a );
 a93058a <=( a93057a  and  a93050a );
 a93062a <=( (not A167)  and  A168 );
 a93063a <=( A170  and  a93062a );
 a93066a <=( (not A199)  and  A166 );
 a93069a <=( (not A201)  and  A200 );
 a93070a <=( a93069a  and  a93066a );
 a93071a <=( a93070a  and  a93063a );
 a93075a <=( A266  and  (not A265) );
 a93076a <=( (not A203)  and  a93075a );
 a93079a <=( (not A269)  and  (not A267) );
 a93082a <=( A300  and  A298 );
 a93083a <=( a93082a  and  a93079a );
 a93084a <=( a93083a  and  a93076a );
 a93088a <=( (not A167)  and  A168 );
 a93089a <=( A170  and  a93088a );
 a93092a <=( (not A199)  and  A166 );
 a93095a <=( (not A201)  and  A200 );
 a93096a <=( a93095a  and  a93092a );
 a93097a <=( a93096a  and  a93089a );
 a93101a <=( (not A266)  and  A265 );
 a93102a <=( (not A203)  and  a93101a );
 a93105a <=( A268  and  (not A267) );
 a93108a <=( A300  and  A299 );
 a93109a <=( a93108a  and  a93105a );
 a93110a <=( a93109a  and  a93102a );
 a93114a <=( (not A167)  and  A168 );
 a93115a <=( A170  and  a93114a );
 a93118a <=( (not A199)  and  A166 );
 a93121a <=( (not A201)  and  A200 );
 a93122a <=( a93121a  and  a93118a );
 a93123a <=( a93122a  and  a93115a );
 a93127a <=( (not A266)  and  A265 );
 a93128a <=( (not A203)  and  a93127a );
 a93131a <=( A268  and  (not A267) );
 a93134a <=( A300  and  A298 );
 a93135a <=( a93134a  and  a93131a );
 a93136a <=( a93135a  and  a93128a );
 a93140a <=( (not A167)  and  A168 );
 a93141a <=( A170  and  a93140a );
 a93144a <=( (not A199)  and  A166 );
 a93147a <=( (not A201)  and  A200 );
 a93148a <=( a93147a  and  a93144a );
 a93149a <=( a93148a  and  a93141a );
 a93153a <=( (not A266)  and  A265 );
 a93154a <=( (not A203)  and  a93153a );
 a93157a <=( (not A269)  and  (not A267) );
 a93160a <=( A300  and  A299 );
 a93161a <=( a93160a  and  a93157a );
 a93162a <=( a93161a  and  a93154a );
 a93166a <=( (not A167)  and  A168 );
 a93167a <=( A170  and  a93166a );
 a93170a <=( (not A199)  and  A166 );
 a93173a <=( (not A201)  and  A200 );
 a93174a <=( a93173a  and  a93170a );
 a93175a <=( a93174a  and  a93167a );
 a93179a <=( (not A266)  and  A265 );
 a93180a <=( (not A203)  and  a93179a );
 a93183a <=( (not A269)  and  (not A267) );
 a93186a <=( A300  and  A298 );
 a93187a <=( a93186a  and  a93183a );
 a93188a <=( a93187a  and  a93180a );
 a93192a <=( (not A167)  and  A168 );
 a93193a <=( A170  and  a93192a );
 a93196a <=( A199  and  A166 );
 a93199a <=( (not A202)  and  (not A200) );
 a93200a <=( a93199a  and  a93196a );
 a93201a <=( a93200a  and  a93193a );
 a93205a <=( A267  and  A265 );
 a93206a <=( A203  and  a93205a );
 a93209a <=( A299  and  A298 );
 a93212a <=( (not A301)  and  (not A300) );
 a93213a <=( a93212a  and  a93209a );
 a93214a <=( a93213a  and  a93206a );
 a93218a <=( (not A167)  and  A168 );
 a93219a <=( A170  and  a93218a );
 a93222a <=( A199  and  A166 );
 a93225a <=( (not A202)  and  (not A200) );
 a93226a <=( a93225a  and  a93222a );
 a93227a <=( a93226a  and  a93219a );
 a93231a <=( A267  and  A265 );
 a93232a <=( A203  and  a93231a );
 a93235a <=( A299  and  A298 );
 a93238a <=( A302  and  (not A300) );
 a93239a <=( a93238a  and  a93235a );
 a93240a <=( a93239a  and  a93232a );
 a93244a <=( (not A167)  and  A168 );
 a93245a <=( A170  and  a93244a );
 a93248a <=( A199  and  A166 );
 a93251a <=( (not A202)  and  (not A200) );
 a93252a <=( a93251a  and  a93248a );
 a93253a <=( a93252a  and  a93245a );
 a93257a <=( A267  and  A265 );
 a93258a <=( A203  and  a93257a );
 a93261a <=( (not A299)  and  A298 );
 a93264a <=( A301  and  (not A300) );
 a93265a <=( a93264a  and  a93261a );
 a93266a <=( a93265a  and  a93258a );
 a93270a <=( (not A167)  and  A168 );
 a93271a <=( A170  and  a93270a );
 a93274a <=( A199  and  A166 );
 a93277a <=( (not A202)  and  (not A200) );
 a93278a <=( a93277a  and  a93274a );
 a93279a <=( a93278a  and  a93271a );
 a93283a <=( A267  and  A265 );
 a93284a <=( A203  and  a93283a );
 a93287a <=( (not A299)  and  A298 );
 a93290a <=( (not A302)  and  (not A300) );
 a93291a <=( a93290a  and  a93287a );
 a93292a <=( a93291a  and  a93284a );
 a93296a <=( (not A167)  and  A168 );
 a93297a <=( A170  and  a93296a );
 a93300a <=( A199  and  A166 );
 a93303a <=( (not A202)  and  (not A200) );
 a93304a <=( a93303a  and  a93300a );
 a93305a <=( a93304a  and  a93297a );
 a93309a <=( A267  and  A265 );
 a93310a <=( A203  and  a93309a );
 a93313a <=( A299  and  (not A298) );
 a93316a <=( A301  and  (not A300) );
 a93317a <=( a93316a  and  a93313a );
 a93318a <=( a93317a  and  a93310a );
 a93322a <=( (not A167)  and  A168 );
 a93323a <=( A170  and  a93322a );
 a93326a <=( A199  and  A166 );
 a93329a <=( (not A202)  and  (not A200) );
 a93330a <=( a93329a  and  a93326a );
 a93331a <=( a93330a  and  a93323a );
 a93335a <=( A267  and  A265 );
 a93336a <=( A203  and  a93335a );
 a93339a <=( A299  and  (not A298) );
 a93342a <=( (not A302)  and  (not A300) );
 a93343a <=( a93342a  and  a93339a );
 a93344a <=( a93343a  and  a93336a );
 a93348a <=( (not A167)  and  A168 );
 a93349a <=( A170  and  a93348a );
 a93352a <=( A199  and  A166 );
 a93355a <=( (not A202)  and  (not A200) );
 a93356a <=( a93355a  and  a93352a );
 a93357a <=( a93356a  and  a93349a );
 a93361a <=( A267  and  A266 );
 a93362a <=( A203  and  a93361a );
 a93365a <=( A299  and  A298 );
 a93368a <=( (not A301)  and  (not A300) );
 a93369a <=( a93368a  and  a93365a );
 a93370a <=( a93369a  and  a93362a );
 a93374a <=( (not A167)  and  A168 );
 a93375a <=( A170  and  a93374a );
 a93378a <=( A199  and  A166 );
 a93381a <=( (not A202)  and  (not A200) );
 a93382a <=( a93381a  and  a93378a );
 a93383a <=( a93382a  and  a93375a );
 a93387a <=( A267  and  A266 );
 a93388a <=( A203  and  a93387a );
 a93391a <=( A299  and  A298 );
 a93394a <=( A302  and  (not A300) );
 a93395a <=( a93394a  and  a93391a );
 a93396a <=( a93395a  and  a93388a );
 a93400a <=( (not A167)  and  A168 );
 a93401a <=( A170  and  a93400a );
 a93404a <=( A199  and  A166 );
 a93407a <=( (not A202)  and  (not A200) );
 a93408a <=( a93407a  and  a93404a );
 a93409a <=( a93408a  and  a93401a );
 a93413a <=( A267  and  A266 );
 a93414a <=( A203  and  a93413a );
 a93417a <=( (not A299)  and  A298 );
 a93420a <=( A301  and  (not A300) );
 a93421a <=( a93420a  and  a93417a );
 a93422a <=( a93421a  and  a93414a );
 a93426a <=( (not A167)  and  A168 );
 a93427a <=( A170  and  a93426a );
 a93430a <=( A199  and  A166 );
 a93433a <=( (not A202)  and  (not A200) );
 a93434a <=( a93433a  and  a93430a );
 a93435a <=( a93434a  and  a93427a );
 a93439a <=( A267  and  A266 );
 a93440a <=( A203  and  a93439a );
 a93443a <=( (not A299)  and  A298 );
 a93446a <=( (not A302)  and  (not A300) );
 a93447a <=( a93446a  and  a93443a );
 a93448a <=( a93447a  and  a93440a );
 a93452a <=( (not A167)  and  A168 );
 a93453a <=( A170  and  a93452a );
 a93456a <=( A199  and  A166 );
 a93459a <=( (not A202)  and  (not A200) );
 a93460a <=( a93459a  and  a93456a );
 a93461a <=( a93460a  and  a93453a );
 a93465a <=( A267  and  A266 );
 a93466a <=( A203  and  a93465a );
 a93469a <=( A299  and  (not A298) );
 a93472a <=( A301  and  (not A300) );
 a93473a <=( a93472a  and  a93469a );
 a93474a <=( a93473a  and  a93466a );
 a93478a <=( (not A167)  and  A168 );
 a93479a <=( A170  and  a93478a );
 a93482a <=( A199  and  A166 );
 a93485a <=( (not A202)  and  (not A200) );
 a93486a <=( a93485a  and  a93482a );
 a93487a <=( a93486a  and  a93479a );
 a93491a <=( A267  and  A266 );
 a93492a <=( A203  and  a93491a );
 a93495a <=( A299  and  (not A298) );
 a93498a <=( (not A302)  and  (not A300) );
 a93499a <=( a93498a  and  a93495a );
 a93500a <=( a93499a  and  a93492a );
 a93504a <=( (not A167)  and  A168 );
 a93505a <=( A170  and  a93504a );
 a93508a <=( A199  and  A166 );
 a93511a <=( (not A201)  and  (not A200) );
 a93512a <=( a93511a  and  a93508a );
 a93513a <=( a93512a  and  a93505a );
 a93517a <=( A266  and  A265 );
 a93518a <=( A202  and  a93517a );
 a93521a <=( (not A268)  and  (not A267) );
 a93524a <=( A300  and  A299 );
 a93525a <=( a93524a  and  a93521a );
 a93526a <=( a93525a  and  a93518a );
 a93530a <=( (not A167)  and  A168 );
 a93531a <=( A170  and  a93530a );
 a93534a <=( A199  and  A166 );
 a93537a <=( (not A201)  and  (not A200) );
 a93538a <=( a93537a  and  a93534a );
 a93539a <=( a93538a  and  a93531a );
 a93543a <=( A266  and  A265 );
 a93544a <=( A202  and  a93543a );
 a93547a <=( (not A268)  and  (not A267) );
 a93550a <=( A300  and  A298 );
 a93551a <=( a93550a  and  a93547a );
 a93552a <=( a93551a  and  a93544a );
 a93556a <=( (not A167)  and  A168 );
 a93557a <=( A170  and  a93556a );
 a93560a <=( A199  and  A166 );
 a93563a <=( (not A201)  and  (not A200) );
 a93564a <=( a93563a  and  a93560a );
 a93565a <=( a93564a  and  a93557a );
 a93569a <=( A266  and  A265 );
 a93570a <=( A202  and  a93569a );
 a93573a <=( A269  and  (not A267) );
 a93576a <=( A300  and  A299 );
 a93577a <=( a93576a  and  a93573a );
 a93578a <=( a93577a  and  a93570a );
 a93582a <=( (not A167)  and  A168 );
 a93583a <=( A170  and  a93582a );
 a93586a <=( A199  and  A166 );
 a93589a <=( (not A201)  and  (not A200) );
 a93590a <=( a93589a  and  a93586a );
 a93591a <=( a93590a  and  a93583a );
 a93595a <=( A266  and  A265 );
 a93596a <=( A202  and  a93595a );
 a93599a <=( A269  and  (not A267) );
 a93602a <=( A300  and  A298 );
 a93603a <=( a93602a  and  a93599a );
 a93604a <=( a93603a  and  a93596a );
 a93608a <=( (not A167)  and  A168 );
 a93609a <=( A170  and  a93608a );
 a93612a <=( A199  and  A166 );
 a93615a <=( (not A201)  and  (not A200) );
 a93616a <=( a93615a  and  a93612a );
 a93617a <=( a93616a  and  a93609a );
 a93621a <=( A266  and  (not A265) );
 a93622a <=( A202  and  a93621a );
 a93625a <=( A268  and  (not A267) );
 a93628a <=( A300  and  A299 );
 a93629a <=( a93628a  and  a93625a );
 a93630a <=( a93629a  and  a93622a );
 a93634a <=( (not A167)  and  A168 );
 a93635a <=( A170  and  a93634a );
 a93638a <=( A199  and  A166 );
 a93641a <=( (not A201)  and  (not A200) );
 a93642a <=( a93641a  and  a93638a );
 a93643a <=( a93642a  and  a93635a );
 a93647a <=( A266  and  (not A265) );
 a93648a <=( A202  and  a93647a );
 a93651a <=( A268  and  (not A267) );
 a93654a <=( A300  and  A298 );
 a93655a <=( a93654a  and  a93651a );
 a93656a <=( a93655a  and  a93648a );
 a93660a <=( (not A167)  and  A168 );
 a93661a <=( A170  and  a93660a );
 a93664a <=( A199  and  A166 );
 a93667a <=( (not A201)  and  (not A200) );
 a93668a <=( a93667a  and  a93664a );
 a93669a <=( a93668a  and  a93661a );
 a93673a <=( A266  and  (not A265) );
 a93674a <=( A202  and  a93673a );
 a93677a <=( (not A269)  and  (not A267) );
 a93680a <=( A300  and  A299 );
 a93681a <=( a93680a  and  a93677a );
 a93682a <=( a93681a  and  a93674a );
 a93686a <=( (not A167)  and  A168 );
 a93687a <=( A170  and  a93686a );
 a93690a <=( A199  and  A166 );
 a93693a <=( (not A201)  and  (not A200) );
 a93694a <=( a93693a  and  a93690a );
 a93695a <=( a93694a  and  a93687a );
 a93699a <=( A266  and  (not A265) );
 a93700a <=( A202  and  a93699a );
 a93703a <=( (not A269)  and  (not A267) );
 a93706a <=( A300  and  A298 );
 a93707a <=( a93706a  and  a93703a );
 a93708a <=( a93707a  and  a93700a );
 a93712a <=( (not A167)  and  A168 );
 a93713a <=( A170  and  a93712a );
 a93716a <=( A199  and  A166 );
 a93719a <=( (not A201)  and  (not A200) );
 a93720a <=( a93719a  and  a93716a );
 a93721a <=( a93720a  and  a93713a );
 a93725a <=( (not A266)  and  A265 );
 a93726a <=( A202  and  a93725a );
 a93729a <=( A268  and  (not A267) );
 a93732a <=( A300  and  A299 );
 a93733a <=( a93732a  and  a93729a );
 a93734a <=( a93733a  and  a93726a );
 a93738a <=( (not A167)  and  A168 );
 a93739a <=( A170  and  a93738a );
 a93742a <=( A199  and  A166 );
 a93745a <=( (not A201)  and  (not A200) );
 a93746a <=( a93745a  and  a93742a );
 a93747a <=( a93746a  and  a93739a );
 a93751a <=( (not A266)  and  A265 );
 a93752a <=( A202  and  a93751a );
 a93755a <=( A268  and  (not A267) );
 a93758a <=( A300  and  A298 );
 a93759a <=( a93758a  and  a93755a );
 a93760a <=( a93759a  and  a93752a );
 a93764a <=( (not A167)  and  A168 );
 a93765a <=( A170  and  a93764a );
 a93768a <=( A199  and  A166 );
 a93771a <=( (not A201)  and  (not A200) );
 a93772a <=( a93771a  and  a93768a );
 a93773a <=( a93772a  and  a93765a );
 a93777a <=( (not A266)  and  A265 );
 a93778a <=( A202  and  a93777a );
 a93781a <=( (not A269)  and  (not A267) );
 a93784a <=( A300  and  A299 );
 a93785a <=( a93784a  and  a93781a );
 a93786a <=( a93785a  and  a93778a );
 a93790a <=( (not A167)  and  A168 );
 a93791a <=( A170  and  a93790a );
 a93794a <=( A199  and  A166 );
 a93797a <=( (not A201)  and  (not A200) );
 a93798a <=( a93797a  and  a93794a );
 a93799a <=( a93798a  and  a93791a );
 a93803a <=( (not A266)  and  A265 );
 a93804a <=( A202  and  a93803a );
 a93807a <=( (not A269)  and  (not A267) );
 a93810a <=( A300  and  A298 );
 a93811a <=( a93810a  and  a93807a );
 a93812a <=( a93811a  and  a93804a );
 a93816a <=( (not A167)  and  A168 );
 a93817a <=( A170  and  a93816a );
 a93820a <=( A199  and  A166 );
 a93823a <=( (not A201)  and  (not A200) );
 a93824a <=( a93823a  and  a93820a );
 a93825a <=( a93824a  and  a93817a );
 a93829a <=( A266  and  A265 );
 a93830a <=( (not A203)  and  a93829a );
 a93833a <=( (not A268)  and  (not A267) );
 a93836a <=( A300  and  A299 );
 a93837a <=( a93836a  and  a93833a );
 a93838a <=( a93837a  and  a93830a );
 a93842a <=( (not A167)  and  A168 );
 a93843a <=( A170  and  a93842a );
 a93846a <=( A199  and  A166 );
 a93849a <=( (not A201)  and  (not A200) );
 a93850a <=( a93849a  and  a93846a );
 a93851a <=( a93850a  and  a93843a );
 a93855a <=( A266  and  A265 );
 a93856a <=( (not A203)  and  a93855a );
 a93859a <=( (not A268)  and  (not A267) );
 a93862a <=( A300  and  A298 );
 a93863a <=( a93862a  and  a93859a );
 a93864a <=( a93863a  and  a93856a );
 a93868a <=( (not A167)  and  A168 );
 a93869a <=( A170  and  a93868a );
 a93872a <=( A199  and  A166 );
 a93875a <=( (not A201)  and  (not A200) );
 a93876a <=( a93875a  and  a93872a );
 a93877a <=( a93876a  and  a93869a );
 a93881a <=( A266  and  A265 );
 a93882a <=( (not A203)  and  a93881a );
 a93885a <=( A269  and  (not A267) );
 a93888a <=( A300  and  A299 );
 a93889a <=( a93888a  and  a93885a );
 a93890a <=( a93889a  and  a93882a );
 a93894a <=( (not A167)  and  A168 );
 a93895a <=( A170  and  a93894a );
 a93898a <=( A199  and  A166 );
 a93901a <=( (not A201)  and  (not A200) );
 a93902a <=( a93901a  and  a93898a );
 a93903a <=( a93902a  and  a93895a );
 a93907a <=( A266  and  A265 );
 a93908a <=( (not A203)  and  a93907a );
 a93911a <=( A269  and  (not A267) );
 a93914a <=( A300  and  A298 );
 a93915a <=( a93914a  and  a93911a );
 a93916a <=( a93915a  and  a93908a );
 a93920a <=( (not A167)  and  A168 );
 a93921a <=( A170  and  a93920a );
 a93924a <=( A199  and  A166 );
 a93927a <=( (not A201)  and  (not A200) );
 a93928a <=( a93927a  and  a93924a );
 a93929a <=( a93928a  and  a93921a );
 a93933a <=( A266  and  (not A265) );
 a93934a <=( (not A203)  and  a93933a );
 a93937a <=( A268  and  (not A267) );
 a93940a <=( A300  and  A299 );
 a93941a <=( a93940a  and  a93937a );
 a93942a <=( a93941a  and  a93934a );
 a93946a <=( (not A167)  and  A168 );
 a93947a <=( A170  and  a93946a );
 a93950a <=( A199  and  A166 );
 a93953a <=( (not A201)  and  (not A200) );
 a93954a <=( a93953a  and  a93950a );
 a93955a <=( a93954a  and  a93947a );
 a93959a <=( A266  and  (not A265) );
 a93960a <=( (not A203)  and  a93959a );
 a93963a <=( A268  and  (not A267) );
 a93966a <=( A300  and  A298 );
 a93967a <=( a93966a  and  a93963a );
 a93968a <=( a93967a  and  a93960a );
 a93972a <=( (not A167)  and  A168 );
 a93973a <=( A170  and  a93972a );
 a93976a <=( A199  and  A166 );
 a93979a <=( (not A201)  and  (not A200) );
 a93980a <=( a93979a  and  a93976a );
 a93981a <=( a93980a  and  a93973a );
 a93985a <=( A266  and  (not A265) );
 a93986a <=( (not A203)  and  a93985a );
 a93989a <=( (not A269)  and  (not A267) );
 a93992a <=( A300  and  A299 );
 a93993a <=( a93992a  and  a93989a );
 a93994a <=( a93993a  and  a93986a );
 a93998a <=( (not A167)  and  A168 );
 a93999a <=( A170  and  a93998a );
 a94002a <=( A199  and  A166 );
 a94005a <=( (not A201)  and  (not A200) );
 a94006a <=( a94005a  and  a94002a );
 a94007a <=( a94006a  and  a93999a );
 a94011a <=( A266  and  (not A265) );
 a94012a <=( (not A203)  and  a94011a );
 a94015a <=( (not A269)  and  (not A267) );
 a94018a <=( A300  and  A298 );
 a94019a <=( a94018a  and  a94015a );
 a94020a <=( a94019a  and  a94012a );
 a94024a <=( (not A167)  and  A168 );
 a94025a <=( A170  and  a94024a );
 a94028a <=( A199  and  A166 );
 a94031a <=( (not A201)  and  (not A200) );
 a94032a <=( a94031a  and  a94028a );
 a94033a <=( a94032a  and  a94025a );
 a94037a <=( (not A266)  and  A265 );
 a94038a <=( (not A203)  and  a94037a );
 a94041a <=( A268  and  (not A267) );
 a94044a <=( A300  and  A299 );
 a94045a <=( a94044a  and  a94041a );
 a94046a <=( a94045a  and  a94038a );
 a94050a <=( (not A167)  and  A168 );
 a94051a <=( A170  and  a94050a );
 a94054a <=( A199  and  A166 );
 a94057a <=( (not A201)  and  (not A200) );
 a94058a <=( a94057a  and  a94054a );
 a94059a <=( a94058a  and  a94051a );
 a94063a <=( (not A266)  and  A265 );
 a94064a <=( (not A203)  and  a94063a );
 a94067a <=( A268  and  (not A267) );
 a94070a <=( A300  and  A298 );
 a94071a <=( a94070a  and  a94067a );
 a94072a <=( a94071a  and  a94064a );
 a94076a <=( (not A167)  and  A168 );
 a94077a <=( A170  and  a94076a );
 a94080a <=( A199  and  A166 );
 a94083a <=( (not A201)  and  (not A200) );
 a94084a <=( a94083a  and  a94080a );
 a94085a <=( a94084a  and  a94077a );
 a94089a <=( (not A266)  and  A265 );
 a94090a <=( (not A203)  and  a94089a );
 a94093a <=( (not A269)  and  (not A267) );
 a94096a <=( A300  and  A299 );
 a94097a <=( a94096a  and  a94093a );
 a94098a <=( a94097a  and  a94090a );
 a94102a <=( (not A167)  and  A168 );
 a94103a <=( A170  and  a94102a );
 a94106a <=( A199  and  A166 );
 a94109a <=( (not A201)  and  (not A200) );
 a94110a <=( a94109a  and  a94106a );
 a94111a <=( a94110a  and  a94103a );
 a94115a <=( (not A266)  and  A265 );
 a94116a <=( (not A203)  and  a94115a );
 a94119a <=( (not A269)  and  (not A267) );
 a94122a <=( A300  and  A298 );
 a94123a <=( a94122a  and  a94119a );
 a94124a <=( a94123a  and  a94116a );
 a94128a <=( (not A167)  and  A168 );
 a94129a <=( A170  and  a94128a );
 a94132a <=( (not A199)  and  A166 );
 a94135a <=( (not A202)  and  (not A200) );
 a94136a <=( a94135a  and  a94132a );
 a94137a <=( a94136a  and  a94129a );
 a94141a <=( (not A268)  and  (not A266) );
 a94142a <=( (not A265)  and  a94141a );
 a94145a <=( A299  and  A298 );
 a94148a <=( (not A302)  and  A301 );
 a94149a <=( a94148a  and  a94145a );
 a94150a <=( a94149a  and  a94142a );
 a94154a <=( (not A167)  and  A168 );
 a94155a <=( A170  and  a94154a );
 a94158a <=( (not A199)  and  A166 );
 a94161a <=( (not A202)  and  (not A200) );
 a94162a <=( a94161a  and  a94158a );
 a94163a <=( a94162a  and  a94155a );
 a94167a <=( (not A268)  and  (not A266) );
 a94168a <=( (not A265)  and  a94167a );
 a94171a <=( (not A299)  and  A298 );
 a94174a <=( A302  and  (not A301) );
 a94175a <=( a94174a  and  a94171a );
 a94176a <=( a94175a  and  a94168a );
 a94180a <=( (not A167)  and  A168 );
 a94181a <=( A170  and  a94180a );
 a94184a <=( (not A199)  and  A166 );
 a94187a <=( (not A202)  and  (not A200) );
 a94188a <=( a94187a  and  a94184a );
 a94189a <=( a94188a  and  a94181a );
 a94193a <=( (not A268)  and  (not A266) );
 a94194a <=( (not A265)  and  a94193a );
 a94197a <=( A299  and  (not A298) );
 a94200a <=( A302  and  (not A301) );
 a94201a <=( a94200a  and  a94197a );
 a94202a <=( a94201a  and  a94194a );
 a94206a <=( (not A167)  and  A168 );
 a94207a <=( A170  and  a94206a );
 a94210a <=( (not A199)  and  A166 );
 a94213a <=( (not A202)  and  (not A200) );
 a94214a <=( a94213a  and  a94210a );
 a94215a <=( a94214a  and  a94207a );
 a94219a <=( (not A268)  and  (not A266) );
 a94220a <=( (not A265)  and  a94219a );
 a94223a <=( (not A299)  and  (not A298) );
 a94226a <=( (not A302)  and  A301 );
 a94227a <=( a94226a  and  a94223a );
 a94228a <=( a94227a  and  a94220a );
 a94232a <=( (not A167)  and  A168 );
 a94233a <=( A170  and  a94232a );
 a94236a <=( (not A199)  and  A166 );
 a94239a <=( (not A202)  and  (not A200) );
 a94240a <=( a94239a  and  a94236a );
 a94241a <=( a94240a  and  a94233a );
 a94245a <=( A269  and  (not A266) );
 a94246a <=( (not A265)  and  a94245a );
 a94249a <=( A299  and  A298 );
 a94252a <=( (not A302)  and  A301 );
 a94253a <=( a94252a  and  a94249a );
 a94254a <=( a94253a  and  a94246a );
 a94258a <=( (not A167)  and  A168 );
 a94259a <=( A170  and  a94258a );
 a94262a <=( (not A199)  and  A166 );
 a94265a <=( (not A202)  and  (not A200) );
 a94266a <=( a94265a  and  a94262a );
 a94267a <=( a94266a  and  a94259a );
 a94271a <=( A269  and  (not A266) );
 a94272a <=( (not A265)  and  a94271a );
 a94275a <=( (not A299)  and  A298 );
 a94278a <=( A302  and  (not A301) );
 a94279a <=( a94278a  and  a94275a );
 a94280a <=( a94279a  and  a94272a );
 a94284a <=( (not A167)  and  A168 );
 a94285a <=( A170  and  a94284a );
 a94288a <=( (not A199)  and  A166 );
 a94291a <=( (not A202)  and  (not A200) );
 a94292a <=( a94291a  and  a94288a );
 a94293a <=( a94292a  and  a94285a );
 a94297a <=( A269  and  (not A266) );
 a94298a <=( (not A265)  and  a94297a );
 a94301a <=( A299  and  (not A298) );
 a94304a <=( A302  and  (not A301) );
 a94305a <=( a94304a  and  a94301a );
 a94306a <=( a94305a  and  a94298a );
 a94310a <=( (not A167)  and  A168 );
 a94311a <=( A170  and  a94310a );
 a94314a <=( (not A199)  and  A166 );
 a94317a <=( (not A202)  and  (not A200) );
 a94318a <=( a94317a  and  a94314a );
 a94319a <=( a94318a  and  a94311a );
 a94323a <=( A269  and  (not A266) );
 a94324a <=( (not A265)  and  a94323a );
 a94327a <=( (not A299)  and  (not A298) );
 a94330a <=( (not A302)  and  A301 );
 a94331a <=( a94330a  and  a94327a );
 a94332a <=( a94331a  and  a94324a );
 a94336a <=( (not A167)  and  A168 );
 a94337a <=( A170  and  a94336a );
 a94340a <=( (not A199)  and  A166 );
 a94343a <=( A203  and  (not A200) );
 a94344a <=( a94343a  and  a94340a );
 a94345a <=( a94344a  and  a94337a );
 a94349a <=( (not A268)  and  (not A266) );
 a94350a <=( (not A265)  and  a94349a );
 a94353a <=( A299  and  A298 );
 a94356a <=( (not A302)  and  A301 );
 a94357a <=( a94356a  and  a94353a );
 a94358a <=( a94357a  and  a94350a );
 a94362a <=( (not A167)  and  A168 );
 a94363a <=( A170  and  a94362a );
 a94366a <=( (not A199)  and  A166 );
 a94369a <=( A203  and  (not A200) );
 a94370a <=( a94369a  and  a94366a );
 a94371a <=( a94370a  and  a94363a );
 a94375a <=( (not A268)  and  (not A266) );
 a94376a <=( (not A265)  and  a94375a );
 a94379a <=( (not A299)  and  A298 );
 a94382a <=( A302  and  (not A301) );
 a94383a <=( a94382a  and  a94379a );
 a94384a <=( a94383a  and  a94376a );
 a94388a <=( (not A167)  and  A168 );
 a94389a <=( A170  and  a94388a );
 a94392a <=( (not A199)  and  A166 );
 a94395a <=( A203  and  (not A200) );
 a94396a <=( a94395a  and  a94392a );
 a94397a <=( a94396a  and  a94389a );
 a94401a <=( (not A268)  and  (not A266) );
 a94402a <=( (not A265)  and  a94401a );
 a94405a <=( A299  and  (not A298) );
 a94408a <=( A302  and  (not A301) );
 a94409a <=( a94408a  and  a94405a );
 a94410a <=( a94409a  and  a94402a );
 a94414a <=( (not A167)  and  A168 );
 a94415a <=( A170  and  a94414a );
 a94418a <=( (not A199)  and  A166 );
 a94421a <=( A203  and  (not A200) );
 a94422a <=( a94421a  and  a94418a );
 a94423a <=( a94422a  and  a94415a );
 a94427a <=( (not A268)  and  (not A266) );
 a94428a <=( (not A265)  and  a94427a );
 a94431a <=( (not A299)  and  (not A298) );
 a94434a <=( (not A302)  and  A301 );
 a94435a <=( a94434a  and  a94431a );
 a94436a <=( a94435a  and  a94428a );
 a94440a <=( (not A167)  and  A168 );
 a94441a <=( A170  and  a94440a );
 a94444a <=( (not A199)  and  A166 );
 a94447a <=( A203  and  (not A200) );
 a94448a <=( a94447a  and  a94444a );
 a94449a <=( a94448a  and  a94441a );
 a94453a <=( A269  and  (not A266) );
 a94454a <=( (not A265)  and  a94453a );
 a94457a <=( A299  and  A298 );
 a94460a <=( (not A302)  and  A301 );
 a94461a <=( a94460a  and  a94457a );
 a94462a <=( a94461a  and  a94454a );
 a94466a <=( (not A167)  and  A168 );
 a94467a <=( A170  and  a94466a );
 a94470a <=( (not A199)  and  A166 );
 a94473a <=( A203  and  (not A200) );
 a94474a <=( a94473a  and  a94470a );
 a94475a <=( a94474a  and  a94467a );
 a94479a <=( A269  and  (not A266) );
 a94480a <=( (not A265)  and  a94479a );
 a94483a <=( (not A299)  and  A298 );
 a94486a <=( A302  and  (not A301) );
 a94487a <=( a94486a  and  a94483a );
 a94488a <=( a94487a  and  a94480a );
 a94492a <=( (not A167)  and  A168 );
 a94493a <=( A170  and  a94492a );
 a94496a <=( (not A199)  and  A166 );
 a94499a <=( A203  and  (not A200) );
 a94500a <=( a94499a  and  a94496a );
 a94501a <=( a94500a  and  a94493a );
 a94505a <=( A269  and  (not A266) );
 a94506a <=( (not A265)  and  a94505a );
 a94509a <=( A299  and  (not A298) );
 a94512a <=( A302  and  (not A301) );
 a94513a <=( a94512a  and  a94509a );
 a94514a <=( a94513a  and  a94506a );
 a94518a <=( (not A167)  and  A168 );
 a94519a <=( A170  and  a94518a );
 a94522a <=( (not A199)  and  A166 );
 a94525a <=( A203  and  (not A200) );
 a94526a <=( a94525a  and  a94522a );
 a94527a <=( a94526a  and  a94519a );
 a94531a <=( A269  and  (not A266) );
 a94532a <=( (not A265)  and  a94531a );
 a94535a <=( (not A299)  and  (not A298) );
 a94538a <=( (not A302)  and  A301 );
 a94539a <=( a94538a  and  a94535a );
 a94540a <=( a94539a  and  a94532a );
 a94544a <=( (not A167)  and  A168 );
 a94545a <=( A170  and  a94544a );
 a94548a <=( (not A199)  and  A166 );
 a94551a <=( A202  and  (not A200) );
 a94552a <=( a94551a  and  a94548a );
 a94553a <=( a94552a  and  a94545a );
 a94557a <=( A267  and  A265 );
 a94558a <=( (not A203)  and  a94557a );
 a94561a <=( A299  and  A298 );
 a94564a <=( (not A301)  and  (not A300) );
 a94565a <=( a94564a  and  a94561a );
 a94566a <=( a94565a  and  a94558a );
 a94570a <=( (not A167)  and  A168 );
 a94571a <=( A170  and  a94570a );
 a94574a <=( (not A199)  and  A166 );
 a94577a <=( A202  and  (not A200) );
 a94578a <=( a94577a  and  a94574a );
 a94579a <=( a94578a  and  a94571a );
 a94583a <=( A267  and  A265 );
 a94584a <=( (not A203)  and  a94583a );
 a94587a <=( A299  and  A298 );
 a94590a <=( A302  and  (not A300) );
 a94591a <=( a94590a  and  a94587a );
 a94592a <=( a94591a  and  a94584a );
 a94596a <=( (not A167)  and  A168 );
 a94597a <=( A170  and  a94596a );
 a94600a <=( (not A199)  and  A166 );
 a94603a <=( A202  and  (not A200) );
 a94604a <=( a94603a  and  a94600a );
 a94605a <=( a94604a  and  a94597a );
 a94609a <=( A267  and  A265 );
 a94610a <=( (not A203)  and  a94609a );
 a94613a <=( (not A299)  and  A298 );
 a94616a <=( A301  and  (not A300) );
 a94617a <=( a94616a  and  a94613a );
 a94618a <=( a94617a  and  a94610a );
 a94622a <=( (not A167)  and  A168 );
 a94623a <=( A170  and  a94622a );
 a94626a <=( (not A199)  and  A166 );
 a94629a <=( A202  and  (not A200) );
 a94630a <=( a94629a  and  a94626a );
 a94631a <=( a94630a  and  a94623a );
 a94635a <=( A267  and  A265 );
 a94636a <=( (not A203)  and  a94635a );
 a94639a <=( (not A299)  and  A298 );
 a94642a <=( (not A302)  and  (not A300) );
 a94643a <=( a94642a  and  a94639a );
 a94644a <=( a94643a  and  a94636a );
 a94648a <=( (not A167)  and  A168 );
 a94649a <=( A170  and  a94648a );
 a94652a <=( (not A199)  and  A166 );
 a94655a <=( A202  and  (not A200) );
 a94656a <=( a94655a  and  a94652a );
 a94657a <=( a94656a  and  a94649a );
 a94661a <=( A267  and  A265 );
 a94662a <=( (not A203)  and  a94661a );
 a94665a <=( A299  and  (not A298) );
 a94668a <=( A301  and  (not A300) );
 a94669a <=( a94668a  and  a94665a );
 a94670a <=( a94669a  and  a94662a );
 a94674a <=( (not A167)  and  A168 );
 a94675a <=( A170  and  a94674a );
 a94678a <=( (not A199)  and  A166 );
 a94681a <=( A202  and  (not A200) );
 a94682a <=( a94681a  and  a94678a );
 a94683a <=( a94682a  and  a94675a );
 a94687a <=( A267  and  A265 );
 a94688a <=( (not A203)  and  a94687a );
 a94691a <=( A299  and  (not A298) );
 a94694a <=( (not A302)  and  (not A300) );
 a94695a <=( a94694a  and  a94691a );
 a94696a <=( a94695a  and  a94688a );
 a94700a <=( (not A167)  and  A168 );
 a94701a <=( A170  and  a94700a );
 a94704a <=( (not A199)  and  A166 );
 a94707a <=( A202  and  (not A200) );
 a94708a <=( a94707a  and  a94704a );
 a94709a <=( a94708a  and  a94701a );
 a94713a <=( A267  and  A266 );
 a94714a <=( (not A203)  and  a94713a );
 a94717a <=( A299  and  A298 );
 a94720a <=( (not A301)  and  (not A300) );
 a94721a <=( a94720a  and  a94717a );
 a94722a <=( a94721a  and  a94714a );
 a94726a <=( (not A167)  and  A168 );
 a94727a <=( A170  and  a94726a );
 a94730a <=( (not A199)  and  A166 );
 a94733a <=( A202  and  (not A200) );
 a94734a <=( a94733a  and  a94730a );
 a94735a <=( a94734a  and  a94727a );
 a94739a <=( A267  and  A266 );
 a94740a <=( (not A203)  and  a94739a );
 a94743a <=( A299  and  A298 );
 a94746a <=( A302  and  (not A300) );
 a94747a <=( a94746a  and  a94743a );
 a94748a <=( a94747a  and  a94740a );
 a94752a <=( (not A167)  and  A168 );
 a94753a <=( A170  and  a94752a );
 a94756a <=( (not A199)  and  A166 );
 a94759a <=( A202  and  (not A200) );
 a94760a <=( a94759a  and  a94756a );
 a94761a <=( a94760a  and  a94753a );
 a94765a <=( A267  and  A266 );
 a94766a <=( (not A203)  and  a94765a );
 a94769a <=( (not A299)  and  A298 );
 a94772a <=( A301  and  (not A300) );
 a94773a <=( a94772a  and  a94769a );
 a94774a <=( a94773a  and  a94766a );
 a94778a <=( (not A167)  and  A168 );
 a94779a <=( A170  and  a94778a );
 a94782a <=( (not A199)  and  A166 );
 a94785a <=( A202  and  (not A200) );
 a94786a <=( a94785a  and  a94782a );
 a94787a <=( a94786a  and  a94779a );
 a94791a <=( A267  and  A266 );
 a94792a <=( (not A203)  and  a94791a );
 a94795a <=( (not A299)  and  A298 );
 a94798a <=( (not A302)  and  (not A300) );
 a94799a <=( a94798a  and  a94795a );
 a94800a <=( a94799a  and  a94792a );
 a94804a <=( (not A167)  and  A168 );
 a94805a <=( A170  and  a94804a );
 a94808a <=( (not A199)  and  A166 );
 a94811a <=( A202  and  (not A200) );
 a94812a <=( a94811a  and  a94808a );
 a94813a <=( a94812a  and  a94805a );
 a94817a <=( A267  and  A266 );
 a94818a <=( (not A203)  and  a94817a );
 a94821a <=( A299  and  (not A298) );
 a94824a <=( A301  and  (not A300) );
 a94825a <=( a94824a  and  a94821a );
 a94826a <=( a94825a  and  a94818a );
 a94830a <=( (not A167)  and  A168 );
 a94831a <=( A170  and  a94830a );
 a94834a <=( (not A199)  and  A166 );
 a94837a <=( A202  and  (not A200) );
 a94838a <=( a94837a  and  a94834a );
 a94839a <=( a94838a  and  a94831a );
 a94843a <=( A267  and  A266 );
 a94844a <=( (not A203)  and  a94843a );
 a94847a <=( A299  and  (not A298) );
 a94850a <=( (not A302)  and  (not A300) );
 a94851a <=( a94850a  and  a94847a );
 a94852a <=( a94851a  and  a94844a );
 a94856a <=( (not A167)  and  A168 );
 a94857a <=( A169  and  a94856a );
 a94860a <=( A199  and  A166 );
 a94863a <=( A265  and  A201 );
 a94864a <=( a94863a  and  a94860a );
 a94865a <=( a94864a  and  a94857a );
 a94869a <=( (not A269)  and  A268 );
 a94870a <=( A266  and  a94869a );
 a94873a <=( A299  and  A298 );
 a94876a <=( (not A301)  and  (not A300) );
 a94877a <=( a94876a  and  a94873a );
 a94878a <=( a94877a  and  a94870a );
 a94882a <=( (not A167)  and  A168 );
 a94883a <=( A169  and  a94882a );
 a94886a <=( A199  and  A166 );
 a94889a <=( A265  and  A201 );
 a94890a <=( a94889a  and  a94886a );
 a94891a <=( a94890a  and  a94883a );
 a94895a <=( (not A269)  and  A268 );
 a94896a <=( A266  and  a94895a );
 a94899a <=( A299  and  A298 );
 a94902a <=( A302  and  (not A300) );
 a94903a <=( a94902a  and  a94899a );
 a94904a <=( a94903a  and  a94896a );
 a94908a <=( (not A167)  and  A168 );
 a94909a <=( A169  and  a94908a );
 a94912a <=( A199  and  A166 );
 a94915a <=( A265  and  A201 );
 a94916a <=( a94915a  and  a94912a );
 a94917a <=( a94916a  and  a94909a );
 a94921a <=( (not A269)  and  A268 );
 a94922a <=( A266  and  a94921a );
 a94925a <=( (not A299)  and  A298 );
 a94928a <=( A301  and  (not A300) );
 a94929a <=( a94928a  and  a94925a );
 a94930a <=( a94929a  and  a94922a );
 a94934a <=( (not A167)  and  A168 );
 a94935a <=( A169  and  a94934a );
 a94938a <=( A199  and  A166 );
 a94941a <=( A265  and  A201 );
 a94942a <=( a94941a  and  a94938a );
 a94943a <=( a94942a  and  a94935a );
 a94947a <=( (not A269)  and  A268 );
 a94948a <=( A266  and  a94947a );
 a94951a <=( (not A299)  and  A298 );
 a94954a <=( (not A302)  and  (not A300) );
 a94955a <=( a94954a  and  a94951a );
 a94956a <=( a94955a  and  a94948a );
 a94960a <=( (not A167)  and  A168 );
 a94961a <=( A169  and  a94960a );
 a94964a <=( A199  and  A166 );
 a94967a <=( A265  and  A201 );
 a94968a <=( a94967a  and  a94964a );
 a94969a <=( a94968a  and  a94961a );
 a94973a <=( (not A269)  and  A268 );
 a94974a <=( A266  and  a94973a );
 a94977a <=( A299  and  (not A298) );
 a94980a <=( A301  and  (not A300) );
 a94981a <=( a94980a  and  a94977a );
 a94982a <=( a94981a  and  a94974a );
 a94986a <=( (not A167)  and  A168 );
 a94987a <=( A169  and  a94986a );
 a94990a <=( A199  and  A166 );
 a94993a <=( A265  and  A201 );
 a94994a <=( a94993a  and  a94990a );
 a94995a <=( a94994a  and  a94987a );
 a94999a <=( (not A269)  and  A268 );
 a95000a <=( A266  and  a94999a );
 a95003a <=( A299  and  (not A298) );
 a95006a <=( (not A302)  and  (not A300) );
 a95007a <=( a95006a  and  a95003a );
 a95008a <=( a95007a  and  a95000a );
 a95012a <=( (not A167)  and  A168 );
 a95013a <=( A169  and  a95012a );
 a95016a <=( A199  and  A166 );
 a95019a <=( (not A265)  and  A201 );
 a95020a <=( a95019a  and  a95016a );
 a95021a <=( a95020a  and  a95013a );
 a95025a <=( A269  and  (not A268) );
 a95026a <=( A266  and  a95025a );
 a95029a <=( A299  and  A298 );
 a95032a <=( (not A301)  and  (not A300) );
 a95033a <=( a95032a  and  a95029a );
 a95034a <=( a95033a  and  a95026a );
 a95038a <=( (not A167)  and  A168 );
 a95039a <=( A169  and  a95038a );
 a95042a <=( A199  and  A166 );
 a95045a <=( (not A265)  and  A201 );
 a95046a <=( a95045a  and  a95042a );
 a95047a <=( a95046a  and  a95039a );
 a95051a <=( A269  and  (not A268) );
 a95052a <=( A266  and  a95051a );
 a95055a <=( A299  and  A298 );
 a95058a <=( A302  and  (not A300) );
 a95059a <=( a95058a  and  a95055a );
 a95060a <=( a95059a  and  a95052a );
 a95064a <=( (not A167)  and  A168 );
 a95065a <=( A169  and  a95064a );
 a95068a <=( A199  and  A166 );
 a95071a <=( (not A265)  and  A201 );
 a95072a <=( a95071a  and  a95068a );
 a95073a <=( a95072a  and  a95065a );
 a95077a <=( A269  and  (not A268) );
 a95078a <=( A266  and  a95077a );
 a95081a <=( (not A299)  and  A298 );
 a95084a <=( A301  and  (not A300) );
 a95085a <=( a95084a  and  a95081a );
 a95086a <=( a95085a  and  a95078a );
 a95090a <=( (not A167)  and  A168 );
 a95091a <=( A169  and  a95090a );
 a95094a <=( A199  and  A166 );
 a95097a <=( (not A265)  and  A201 );
 a95098a <=( a95097a  and  a95094a );
 a95099a <=( a95098a  and  a95091a );
 a95103a <=( A269  and  (not A268) );
 a95104a <=( A266  and  a95103a );
 a95107a <=( (not A299)  and  A298 );
 a95110a <=( (not A302)  and  (not A300) );
 a95111a <=( a95110a  and  a95107a );
 a95112a <=( a95111a  and  a95104a );
 a95116a <=( (not A167)  and  A168 );
 a95117a <=( A169  and  a95116a );
 a95120a <=( A199  and  A166 );
 a95123a <=( (not A265)  and  A201 );
 a95124a <=( a95123a  and  a95120a );
 a95125a <=( a95124a  and  a95117a );
 a95129a <=( A269  and  (not A268) );
 a95130a <=( A266  and  a95129a );
 a95133a <=( A299  and  (not A298) );
 a95136a <=( A301  and  (not A300) );
 a95137a <=( a95136a  and  a95133a );
 a95138a <=( a95137a  and  a95130a );
 a95142a <=( (not A167)  and  A168 );
 a95143a <=( A169  and  a95142a );
 a95146a <=( A199  and  A166 );
 a95149a <=( (not A265)  and  A201 );
 a95150a <=( a95149a  and  a95146a );
 a95151a <=( a95150a  and  a95143a );
 a95155a <=( A269  and  (not A268) );
 a95156a <=( A266  and  a95155a );
 a95159a <=( A299  and  (not A298) );
 a95162a <=( (not A302)  and  (not A300) );
 a95163a <=( a95162a  and  a95159a );
 a95164a <=( a95163a  and  a95156a );
 a95168a <=( (not A167)  and  A168 );
 a95169a <=( A169  and  a95168a );
 a95172a <=( A199  and  A166 );
 a95175a <=( A265  and  A201 );
 a95176a <=( a95175a  and  a95172a );
 a95177a <=( a95176a  and  a95169a );
 a95181a <=( A269  and  (not A268) );
 a95182a <=( (not A266)  and  a95181a );
 a95185a <=( A299  and  A298 );
 a95188a <=( (not A301)  and  (not A300) );
 a95189a <=( a95188a  and  a95185a );
 a95190a <=( a95189a  and  a95182a );
 a95194a <=( (not A167)  and  A168 );
 a95195a <=( A169  and  a95194a );
 a95198a <=( A199  and  A166 );
 a95201a <=( A265  and  A201 );
 a95202a <=( a95201a  and  a95198a );
 a95203a <=( a95202a  and  a95195a );
 a95207a <=( A269  and  (not A268) );
 a95208a <=( (not A266)  and  a95207a );
 a95211a <=( A299  and  A298 );
 a95214a <=( A302  and  (not A300) );
 a95215a <=( a95214a  and  a95211a );
 a95216a <=( a95215a  and  a95208a );
 a95220a <=( (not A167)  and  A168 );
 a95221a <=( A169  and  a95220a );
 a95224a <=( A199  and  A166 );
 a95227a <=( A265  and  A201 );
 a95228a <=( a95227a  and  a95224a );
 a95229a <=( a95228a  and  a95221a );
 a95233a <=( A269  and  (not A268) );
 a95234a <=( (not A266)  and  a95233a );
 a95237a <=( (not A299)  and  A298 );
 a95240a <=( A301  and  (not A300) );
 a95241a <=( a95240a  and  a95237a );
 a95242a <=( a95241a  and  a95234a );
 a95246a <=( (not A167)  and  A168 );
 a95247a <=( A169  and  a95246a );
 a95250a <=( A199  and  A166 );
 a95253a <=( A265  and  A201 );
 a95254a <=( a95253a  and  a95250a );
 a95255a <=( a95254a  and  a95247a );
 a95259a <=( A269  and  (not A268) );
 a95260a <=( (not A266)  and  a95259a );
 a95263a <=( (not A299)  and  A298 );
 a95266a <=( (not A302)  and  (not A300) );
 a95267a <=( a95266a  and  a95263a );
 a95268a <=( a95267a  and  a95260a );
 a95272a <=( (not A167)  and  A168 );
 a95273a <=( A169  and  a95272a );
 a95276a <=( A199  and  A166 );
 a95279a <=( A265  and  A201 );
 a95280a <=( a95279a  and  a95276a );
 a95281a <=( a95280a  and  a95273a );
 a95285a <=( A269  and  (not A268) );
 a95286a <=( (not A266)  and  a95285a );
 a95289a <=( A299  and  (not A298) );
 a95292a <=( A301  and  (not A300) );
 a95293a <=( a95292a  and  a95289a );
 a95294a <=( a95293a  and  a95286a );
 a95298a <=( (not A167)  and  A168 );
 a95299a <=( A169  and  a95298a );
 a95302a <=( A199  and  A166 );
 a95305a <=( A265  and  A201 );
 a95306a <=( a95305a  and  a95302a );
 a95307a <=( a95306a  and  a95299a );
 a95311a <=( A269  and  (not A268) );
 a95312a <=( (not A266)  and  a95311a );
 a95315a <=( A299  and  (not A298) );
 a95318a <=( (not A302)  and  (not A300) );
 a95319a <=( a95318a  and  a95315a );
 a95320a <=( a95319a  and  a95312a );
 a95324a <=( (not A167)  and  A168 );
 a95325a <=( A169  and  a95324a );
 a95328a <=( A199  and  A166 );
 a95331a <=( (not A265)  and  A201 );
 a95332a <=( a95331a  and  a95328a );
 a95333a <=( a95332a  and  a95325a );
 a95337a <=( (not A269)  and  A268 );
 a95338a <=( (not A266)  and  a95337a );
 a95341a <=( A299  and  A298 );
 a95344a <=( (not A301)  and  (not A300) );
 a95345a <=( a95344a  and  a95341a );
 a95346a <=( a95345a  and  a95338a );
 a95350a <=( (not A167)  and  A168 );
 a95351a <=( A169  and  a95350a );
 a95354a <=( A199  and  A166 );
 a95357a <=( (not A265)  and  A201 );
 a95358a <=( a95357a  and  a95354a );
 a95359a <=( a95358a  and  a95351a );
 a95363a <=( (not A269)  and  A268 );
 a95364a <=( (not A266)  and  a95363a );
 a95367a <=( A299  and  A298 );
 a95370a <=( A302  and  (not A300) );
 a95371a <=( a95370a  and  a95367a );
 a95372a <=( a95371a  and  a95364a );
 a95376a <=( (not A167)  and  A168 );
 a95377a <=( A169  and  a95376a );
 a95380a <=( A199  and  A166 );
 a95383a <=( (not A265)  and  A201 );
 a95384a <=( a95383a  and  a95380a );
 a95385a <=( a95384a  and  a95377a );
 a95389a <=( (not A269)  and  A268 );
 a95390a <=( (not A266)  and  a95389a );
 a95393a <=( (not A299)  and  A298 );
 a95396a <=( A301  and  (not A300) );
 a95397a <=( a95396a  and  a95393a );
 a95398a <=( a95397a  and  a95390a );
 a95402a <=( (not A167)  and  A168 );
 a95403a <=( A169  and  a95402a );
 a95406a <=( A199  and  A166 );
 a95409a <=( (not A265)  and  A201 );
 a95410a <=( a95409a  and  a95406a );
 a95411a <=( a95410a  and  a95403a );
 a95415a <=( (not A269)  and  A268 );
 a95416a <=( (not A266)  and  a95415a );
 a95419a <=( (not A299)  and  A298 );
 a95422a <=( (not A302)  and  (not A300) );
 a95423a <=( a95422a  and  a95419a );
 a95424a <=( a95423a  and  a95416a );
 a95428a <=( (not A167)  and  A168 );
 a95429a <=( A169  and  a95428a );
 a95432a <=( A199  and  A166 );
 a95435a <=( (not A265)  and  A201 );
 a95436a <=( a95435a  and  a95432a );
 a95437a <=( a95436a  and  a95429a );
 a95441a <=( (not A269)  and  A268 );
 a95442a <=( (not A266)  and  a95441a );
 a95445a <=( A299  and  (not A298) );
 a95448a <=( A301  and  (not A300) );
 a95449a <=( a95448a  and  a95445a );
 a95450a <=( a95449a  and  a95442a );
 a95454a <=( (not A167)  and  A168 );
 a95455a <=( A169  and  a95454a );
 a95458a <=( A199  and  A166 );
 a95461a <=( (not A265)  and  A201 );
 a95462a <=( a95461a  and  a95458a );
 a95463a <=( a95462a  and  a95455a );
 a95467a <=( (not A269)  and  A268 );
 a95468a <=( (not A266)  and  a95467a );
 a95471a <=( A299  and  (not A298) );
 a95474a <=( (not A302)  and  (not A300) );
 a95475a <=( a95474a  and  a95471a );
 a95476a <=( a95475a  and  a95468a );
 a95480a <=( (not A167)  and  A168 );
 a95481a <=( A169  and  a95480a );
 a95484a <=( A200  and  A166 );
 a95487a <=( A265  and  A201 );
 a95488a <=( a95487a  and  a95484a );
 a95489a <=( a95488a  and  a95481a );
 a95493a <=( (not A269)  and  A268 );
 a95494a <=( A266  and  a95493a );
 a95497a <=( A299  and  A298 );
 a95500a <=( (not A301)  and  (not A300) );
 a95501a <=( a95500a  and  a95497a );
 a95502a <=( a95501a  and  a95494a );
 a95506a <=( (not A167)  and  A168 );
 a95507a <=( A169  and  a95506a );
 a95510a <=( A200  and  A166 );
 a95513a <=( A265  and  A201 );
 a95514a <=( a95513a  and  a95510a );
 a95515a <=( a95514a  and  a95507a );
 a95519a <=( (not A269)  and  A268 );
 a95520a <=( A266  and  a95519a );
 a95523a <=( A299  and  A298 );
 a95526a <=( A302  and  (not A300) );
 a95527a <=( a95526a  and  a95523a );
 a95528a <=( a95527a  and  a95520a );
 a95532a <=( (not A167)  and  A168 );
 a95533a <=( A169  and  a95532a );
 a95536a <=( A200  and  A166 );
 a95539a <=( A265  and  A201 );
 a95540a <=( a95539a  and  a95536a );
 a95541a <=( a95540a  and  a95533a );
 a95545a <=( (not A269)  and  A268 );
 a95546a <=( A266  and  a95545a );
 a95549a <=( (not A299)  and  A298 );
 a95552a <=( A301  and  (not A300) );
 a95553a <=( a95552a  and  a95549a );
 a95554a <=( a95553a  and  a95546a );
 a95558a <=( (not A167)  and  A168 );
 a95559a <=( A169  and  a95558a );
 a95562a <=( A200  and  A166 );
 a95565a <=( A265  and  A201 );
 a95566a <=( a95565a  and  a95562a );
 a95567a <=( a95566a  and  a95559a );
 a95571a <=( (not A269)  and  A268 );
 a95572a <=( A266  and  a95571a );
 a95575a <=( (not A299)  and  A298 );
 a95578a <=( (not A302)  and  (not A300) );
 a95579a <=( a95578a  and  a95575a );
 a95580a <=( a95579a  and  a95572a );
 a95584a <=( (not A167)  and  A168 );
 a95585a <=( A169  and  a95584a );
 a95588a <=( A200  and  A166 );
 a95591a <=( A265  and  A201 );
 a95592a <=( a95591a  and  a95588a );
 a95593a <=( a95592a  and  a95585a );
 a95597a <=( (not A269)  and  A268 );
 a95598a <=( A266  and  a95597a );
 a95601a <=( A299  and  (not A298) );
 a95604a <=( A301  and  (not A300) );
 a95605a <=( a95604a  and  a95601a );
 a95606a <=( a95605a  and  a95598a );
 a95610a <=( (not A167)  and  A168 );
 a95611a <=( A169  and  a95610a );
 a95614a <=( A200  and  A166 );
 a95617a <=( A265  and  A201 );
 a95618a <=( a95617a  and  a95614a );
 a95619a <=( a95618a  and  a95611a );
 a95623a <=( (not A269)  and  A268 );
 a95624a <=( A266  and  a95623a );
 a95627a <=( A299  and  (not A298) );
 a95630a <=( (not A302)  and  (not A300) );
 a95631a <=( a95630a  and  a95627a );
 a95632a <=( a95631a  and  a95624a );
 a95636a <=( (not A167)  and  A168 );
 a95637a <=( A169  and  a95636a );
 a95640a <=( A200  and  A166 );
 a95643a <=( (not A265)  and  A201 );
 a95644a <=( a95643a  and  a95640a );
 a95645a <=( a95644a  and  a95637a );
 a95649a <=( A269  and  (not A268) );
 a95650a <=( A266  and  a95649a );
 a95653a <=( A299  and  A298 );
 a95656a <=( (not A301)  and  (not A300) );
 a95657a <=( a95656a  and  a95653a );
 a95658a <=( a95657a  and  a95650a );
 a95662a <=( (not A167)  and  A168 );
 a95663a <=( A169  and  a95662a );
 a95666a <=( A200  and  A166 );
 a95669a <=( (not A265)  and  A201 );
 a95670a <=( a95669a  and  a95666a );
 a95671a <=( a95670a  and  a95663a );
 a95675a <=( A269  and  (not A268) );
 a95676a <=( A266  and  a95675a );
 a95679a <=( A299  and  A298 );
 a95682a <=( A302  and  (not A300) );
 a95683a <=( a95682a  and  a95679a );
 a95684a <=( a95683a  and  a95676a );
 a95688a <=( (not A167)  and  A168 );
 a95689a <=( A169  and  a95688a );
 a95692a <=( A200  and  A166 );
 a95695a <=( (not A265)  and  A201 );
 a95696a <=( a95695a  and  a95692a );
 a95697a <=( a95696a  and  a95689a );
 a95701a <=( A269  and  (not A268) );
 a95702a <=( A266  and  a95701a );
 a95705a <=( (not A299)  and  A298 );
 a95708a <=( A301  and  (not A300) );
 a95709a <=( a95708a  and  a95705a );
 a95710a <=( a95709a  and  a95702a );
 a95714a <=( (not A167)  and  A168 );
 a95715a <=( A169  and  a95714a );
 a95718a <=( A200  and  A166 );
 a95721a <=( (not A265)  and  A201 );
 a95722a <=( a95721a  and  a95718a );
 a95723a <=( a95722a  and  a95715a );
 a95727a <=( A269  and  (not A268) );
 a95728a <=( A266  and  a95727a );
 a95731a <=( (not A299)  and  A298 );
 a95734a <=( (not A302)  and  (not A300) );
 a95735a <=( a95734a  and  a95731a );
 a95736a <=( a95735a  and  a95728a );
 a95740a <=( (not A167)  and  A168 );
 a95741a <=( A169  and  a95740a );
 a95744a <=( A200  and  A166 );
 a95747a <=( (not A265)  and  A201 );
 a95748a <=( a95747a  and  a95744a );
 a95749a <=( a95748a  and  a95741a );
 a95753a <=( A269  and  (not A268) );
 a95754a <=( A266  and  a95753a );
 a95757a <=( A299  and  (not A298) );
 a95760a <=( A301  and  (not A300) );
 a95761a <=( a95760a  and  a95757a );
 a95762a <=( a95761a  and  a95754a );
 a95766a <=( (not A167)  and  A168 );
 a95767a <=( A169  and  a95766a );
 a95770a <=( A200  and  A166 );
 a95773a <=( (not A265)  and  A201 );
 a95774a <=( a95773a  and  a95770a );
 a95775a <=( a95774a  and  a95767a );
 a95779a <=( A269  and  (not A268) );
 a95780a <=( A266  and  a95779a );
 a95783a <=( A299  and  (not A298) );
 a95786a <=( (not A302)  and  (not A300) );
 a95787a <=( a95786a  and  a95783a );
 a95788a <=( a95787a  and  a95780a );
 a95792a <=( (not A167)  and  A168 );
 a95793a <=( A169  and  a95792a );
 a95796a <=( A200  and  A166 );
 a95799a <=( A265  and  A201 );
 a95800a <=( a95799a  and  a95796a );
 a95801a <=( a95800a  and  a95793a );
 a95805a <=( A269  and  (not A268) );
 a95806a <=( (not A266)  and  a95805a );
 a95809a <=( A299  and  A298 );
 a95812a <=( (not A301)  and  (not A300) );
 a95813a <=( a95812a  and  a95809a );
 a95814a <=( a95813a  and  a95806a );
 a95818a <=( (not A167)  and  A168 );
 a95819a <=( A169  and  a95818a );
 a95822a <=( A200  and  A166 );
 a95825a <=( A265  and  A201 );
 a95826a <=( a95825a  and  a95822a );
 a95827a <=( a95826a  and  a95819a );
 a95831a <=( A269  and  (not A268) );
 a95832a <=( (not A266)  and  a95831a );
 a95835a <=( A299  and  A298 );
 a95838a <=( A302  and  (not A300) );
 a95839a <=( a95838a  and  a95835a );
 a95840a <=( a95839a  and  a95832a );
 a95844a <=( (not A167)  and  A168 );
 a95845a <=( A169  and  a95844a );
 a95848a <=( A200  and  A166 );
 a95851a <=( A265  and  A201 );
 a95852a <=( a95851a  and  a95848a );
 a95853a <=( a95852a  and  a95845a );
 a95857a <=( A269  and  (not A268) );
 a95858a <=( (not A266)  and  a95857a );
 a95861a <=( (not A299)  and  A298 );
 a95864a <=( A301  and  (not A300) );
 a95865a <=( a95864a  and  a95861a );
 a95866a <=( a95865a  and  a95858a );
 a95870a <=( (not A167)  and  A168 );
 a95871a <=( A169  and  a95870a );
 a95874a <=( A200  and  A166 );
 a95877a <=( A265  and  A201 );
 a95878a <=( a95877a  and  a95874a );
 a95879a <=( a95878a  and  a95871a );
 a95883a <=( A269  and  (not A268) );
 a95884a <=( (not A266)  and  a95883a );
 a95887a <=( (not A299)  and  A298 );
 a95890a <=( (not A302)  and  (not A300) );
 a95891a <=( a95890a  and  a95887a );
 a95892a <=( a95891a  and  a95884a );
 a95896a <=( (not A167)  and  A168 );
 a95897a <=( A169  and  a95896a );
 a95900a <=( A200  and  A166 );
 a95903a <=( A265  and  A201 );
 a95904a <=( a95903a  and  a95900a );
 a95905a <=( a95904a  and  a95897a );
 a95909a <=( A269  and  (not A268) );
 a95910a <=( (not A266)  and  a95909a );
 a95913a <=( A299  and  (not A298) );
 a95916a <=( A301  and  (not A300) );
 a95917a <=( a95916a  and  a95913a );
 a95918a <=( a95917a  and  a95910a );
 a95922a <=( (not A167)  and  A168 );
 a95923a <=( A169  and  a95922a );
 a95926a <=( A200  and  A166 );
 a95929a <=( A265  and  A201 );
 a95930a <=( a95929a  and  a95926a );
 a95931a <=( a95930a  and  a95923a );
 a95935a <=( A269  and  (not A268) );
 a95936a <=( (not A266)  and  a95935a );
 a95939a <=( A299  and  (not A298) );
 a95942a <=( (not A302)  and  (not A300) );
 a95943a <=( a95942a  and  a95939a );
 a95944a <=( a95943a  and  a95936a );
 a95948a <=( (not A167)  and  A168 );
 a95949a <=( A169  and  a95948a );
 a95952a <=( A200  and  A166 );
 a95955a <=( (not A265)  and  A201 );
 a95956a <=( a95955a  and  a95952a );
 a95957a <=( a95956a  and  a95949a );
 a95961a <=( (not A269)  and  A268 );
 a95962a <=( (not A266)  and  a95961a );
 a95965a <=( A299  and  A298 );
 a95968a <=( (not A301)  and  (not A300) );
 a95969a <=( a95968a  and  a95965a );
 a95970a <=( a95969a  and  a95962a );
 a95974a <=( (not A167)  and  A168 );
 a95975a <=( A169  and  a95974a );
 a95978a <=( A200  and  A166 );
 a95981a <=( (not A265)  and  A201 );
 a95982a <=( a95981a  and  a95978a );
 a95983a <=( a95982a  and  a95975a );
 a95987a <=( (not A269)  and  A268 );
 a95988a <=( (not A266)  and  a95987a );
 a95991a <=( A299  and  A298 );
 a95994a <=( A302  and  (not A300) );
 a95995a <=( a95994a  and  a95991a );
 a95996a <=( a95995a  and  a95988a );
 a96000a <=( (not A167)  and  A168 );
 a96001a <=( A169  and  a96000a );
 a96004a <=( A200  and  A166 );
 a96007a <=( (not A265)  and  A201 );
 a96008a <=( a96007a  and  a96004a );
 a96009a <=( a96008a  and  a96001a );
 a96013a <=( (not A269)  and  A268 );
 a96014a <=( (not A266)  and  a96013a );
 a96017a <=( (not A299)  and  A298 );
 a96020a <=( A301  and  (not A300) );
 a96021a <=( a96020a  and  a96017a );
 a96022a <=( a96021a  and  a96014a );
 a96026a <=( (not A167)  and  A168 );
 a96027a <=( A169  and  a96026a );
 a96030a <=( A200  and  A166 );
 a96033a <=( (not A265)  and  A201 );
 a96034a <=( a96033a  and  a96030a );
 a96035a <=( a96034a  and  a96027a );
 a96039a <=( (not A269)  and  A268 );
 a96040a <=( (not A266)  and  a96039a );
 a96043a <=( (not A299)  and  A298 );
 a96046a <=( (not A302)  and  (not A300) );
 a96047a <=( a96046a  and  a96043a );
 a96048a <=( a96047a  and  a96040a );
 a96052a <=( (not A167)  and  A168 );
 a96053a <=( A169  and  a96052a );
 a96056a <=( A200  and  A166 );
 a96059a <=( (not A265)  and  A201 );
 a96060a <=( a96059a  and  a96056a );
 a96061a <=( a96060a  and  a96053a );
 a96065a <=( (not A269)  and  A268 );
 a96066a <=( (not A266)  and  a96065a );
 a96069a <=( A299  and  (not A298) );
 a96072a <=( A301  and  (not A300) );
 a96073a <=( a96072a  and  a96069a );
 a96074a <=( a96073a  and  a96066a );
 a96078a <=( (not A167)  and  A168 );
 a96079a <=( A169  and  a96078a );
 a96082a <=( A200  and  A166 );
 a96085a <=( (not A265)  and  A201 );
 a96086a <=( a96085a  and  a96082a );
 a96087a <=( a96086a  and  a96079a );
 a96091a <=( (not A269)  and  A268 );
 a96092a <=( (not A266)  and  a96091a );
 a96095a <=( A299  and  (not A298) );
 a96098a <=( (not A302)  and  (not A300) );
 a96099a <=( a96098a  and  a96095a );
 a96100a <=( a96099a  and  a96092a );
 a96104a <=( (not A167)  and  A168 );
 a96105a <=( A169  and  a96104a );
 a96108a <=( A199  and  A166 );
 a96111a <=( A202  and  A200 );
 a96112a <=( a96111a  and  a96108a );
 a96113a <=( a96112a  and  a96105a );
 a96117a <=( A267  and  A265 );
 a96118a <=( (not A203)  and  a96117a );
 a96121a <=( A299  and  A298 );
 a96124a <=( (not A301)  and  (not A300) );
 a96125a <=( a96124a  and  a96121a );
 a96126a <=( a96125a  and  a96118a );
 a96130a <=( (not A167)  and  A168 );
 a96131a <=( A169  and  a96130a );
 a96134a <=( A199  and  A166 );
 a96137a <=( A202  and  A200 );
 a96138a <=( a96137a  and  a96134a );
 a96139a <=( a96138a  and  a96131a );
 a96143a <=( A267  and  A265 );
 a96144a <=( (not A203)  and  a96143a );
 a96147a <=( A299  and  A298 );
 a96150a <=( A302  and  (not A300) );
 a96151a <=( a96150a  and  a96147a );
 a96152a <=( a96151a  and  a96144a );
 a96156a <=( (not A167)  and  A168 );
 a96157a <=( A169  and  a96156a );
 a96160a <=( A199  and  A166 );
 a96163a <=( A202  and  A200 );
 a96164a <=( a96163a  and  a96160a );
 a96165a <=( a96164a  and  a96157a );
 a96169a <=( A267  and  A265 );
 a96170a <=( (not A203)  and  a96169a );
 a96173a <=( (not A299)  and  A298 );
 a96176a <=( A301  and  (not A300) );
 a96177a <=( a96176a  and  a96173a );
 a96178a <=( a96177a  and  a96170a );
 a96182a <=( (not A167)  and  A168 );
 a96183a <=( A169  and  a96182a );
 a96186a <=( A199  and  A166 );
 a96189a <=( A202  and  A200 );
 a96190a <=( a96189a  and  a96186a );
 a96191a <=( a96190a  and  a96183a );
 a96195a <=( A267  and  A265 );
 a96196a <=( (not A203)  and  a96195a );
 a96199a <=( (not A299)  and  A298 );
 a96202a <=( (not A302)  and  (not A300) );
 a96203a <=( a96202a  and  a96199a );
 a96204a <=( a96203a  and  a96196a );
 a96208a <=( (not A167)  and  A168 );
 a96209a <=( A169  and  a96208a );
 a96212a <=( A199  and  A166 );
 a96215a <=( A202  and  A200 );
 a96216a <=( a96215a  and  a96212a );
 a96217a <=( a96216a  and  a96209a );
 a96221a <=( A267  and  A265 );
 a96222a <=( (not A203)  and  a96221a );
 a96225a <=( A299  and  (not A298) );
 a96228a <=( A301  and  (not A300) );
 a96229a <=( a96228a  and  a96225a );
 a96230a <=( a96229a  and  a96222a );
 a96234a <=( (not A167)  and  A168 );
 a96235a <=( A169  and  a96234a );
 a96238a <=( A199  and  A166 );
 a96241a <=( A202  and  A200 );
 a96242a <=( a96241a  and  a96238a );
 a96243a <=( a96242a  and  a96235a );
 a96247a <=( A267  and  A265 );
 a96248a <=( (not A203)  and  a96247a );
 a96251a <=( A299  and  (not A298) );
 a96254a <=( (not A302)  and  (not A300) );
 a96255a <=( a96254a  and  a96251a );
 a96256a <=( a96255a  and  a96248a );
 a96260a <=( (not A167)  and  A168 );
 a96261a <=( A169  and  a96260a );
 a96264a <=( A199  and  A166 );
 a96267a <=( A202  and  A200 );
 a96268a <=( a96267a  and  a96264a );
 a96269a <=( a96268a  and  a96261a );
 a96273a <=( A267  and  A266 );
 a96274a <=( (not A203)  and  a96273a );
 a96277a <=( A299  and  A298 );
 a96280a <=( (not A301)  and  (not A300) );
 a96281a <=( a96280a  and  a96277a );
 a96282a <=( a96281a  and  a96274a );
 a96286a <=( (not A167)  and  A168 );
 a96287a <=( A169  and  a96286a );
 a96290a <=( A199  and  A166 );
 a96293a <=( A202  and  A200 );
 a96294a <=( a96293a  and  a96290a );
 a96295a <=( a96294a  and  a96287a );
 a96299a <=( A267  and  A266 );
 a96300a <=( (not A203)  and  a96299a );
 a96303a <=( A299  and  A298 );
 a96306a <=( A302  and  (not A300) );
 a96307a <=( a96306a  and  a96303a );
 a96308a <=( a96307a  and  a96300a );
 a96312a <=( (not A167)  and  A168 );
 a96313a <=( A169  and  a96312a );
 a96316a <=( A199  and  A166 );
 a96319a <=( A202  and  A200 );
 a96320a <=( a96319a  and  a96316a );
 a96321a <=( a96320a  and  a96313a );
 a96325a <=( A267  and  A266 );
 a96326a <=( (not A203)  and  a96325a );
 a96329a <=( (not A299)  and  A298 );
 a96332a <=( A301  and  (not A300) );
 a96333a <=( a96332a  and  a96329a );
 a96334a <=( a96333a  and  a96326a );
 a96338a <=( (not A167)  and  A168 );
 a96339a <=( A169  and  a96338a );
 a96342a <=( A199  and  A166 );
 a96345a <=( A202  and  A200 );
 a96346a <=( a96345a  and  a96342a );
 a96347a <=( a96346a  and  a96339a );
 a96351a <=( A267  and  A266 );
 a96352a <=( (not A203)  and  a96351a );
 a96355a <=( (not A299)  and  A298 );
 a96358a <=( (not A302)  and  (not A300) );
 a96359a <=( a96358a  and  a96355a );
 a96360a <=( a96359a  and  a96352a );
 a96364a <=( (not A167)  and  A168 );
 a96365a <=( A169  and  a96364a );
 a96368a <=( A199  and  A166 );
 a96371a <=( A202  and  A200 );
 a96372a <=( a96371a  and  a96368a );
 a96373a <=( a96372a  and  a96365a );
 a96377a <=( A267  and  A266 );
 a96378a <=( (not A203)  and  a96377a );
 a96381a <=( A299  and  (not A298) );
 a96384a <=( A301  and  (not A300) );
 a96385a <=( a96384a  and  a96381a );
 a96386a <=( a96385a  and  a96378a );
 a96390a <=( (not A167)  and  A168 );
 a96391a <=( A169  and  a96390a );
 a96394a <=( A199  and  A166 );
 a96397a <=( A202  and  A200 );
 a96398a <=( a96397a  and  a96394a );
 a96399a <=( a96398a  and  a96391a );
 a96403a <=( A267  and  A266 );
 a96404a <=( (not A203)  and  a96403a );
 a96407a <=( A299  and  (not A298) );
 a96410a <=( (not A302)  and  (not A300) );
 a96411a <=( a96410a  and  a96407a );
 a96412a <=( a96411a  and  a96404a );
 a96416a <=( (not A167)  and  A168 );
 a96417a <=( A169  and  a96416a );
 a96420a <=( A199  and  A166 );
 a96423a <=( (not A201)  and  A200 );
 a96424a <=( a96423a  and  a96420a );
 a96425a <=( a96424a  and  a96417a );
 a96429a <=( A266  and  A265 );
 a96430a <=( (not A202)  and  a96429a );
 a96433a <=( (not A268)  and  (not A267) );
 a96436a <=( A300  and  A299 );
 a96437a <=( a96436a  and  a96433a );
 a96438a <=( a96437a  and  a96430a );
 a96442a <=( (not A167)  and  A168 );
 a96443a <=( A169  and  a96442a );
 a96446a <=( A199  and  A166 );
 a96449a <=( (not A201)  and  A200 );
 a96450a <=( a96449a  and  a96446a );
 a96451a <=( a96450a  and  a96443a );
 a96455a <=( A266  and  A265 );
 a96456a <=( (not A202)  and  a96455a );
 a96459a <=( (not A268)  and  (not A267) );
 a96462a <=( A300  and  A298 );
 a96463a <=( a96462a  and  a96459a );
 a96464a <=( a96463a  and  a96456a );
 a96468a <=( (not A167)  and  A168 );
 a96469a <=( A169  and  a96468a );
 a96472a <=( A199  and  A166 );
 a96475a <=( (not A201)  and  A200 );
 a96476a <=( a96475a  and  a96472a );
 a96477a <=( a96476a  and  a96469a );
 a96481a <=( A266  and  A265 );
 a96482a <=( (not A202)  and  a96481a );
 a96485a <=( A269  and  (not A267) );
 a96488a <=( A300  and  A299 );
 a96489a <=( a96488a  and  a96485a );
 a96490a <=( a96489a  and  a96482a );
 a96494a <=( (not A167)  and  A168 );
 a96495a <=( A169  and  a96494a );
 a96498a <=( A199  and  A166 );
 a96501a <=( (not A201)  and  A200 );
 a96502a <=( a96501a  and  a96498a );
 a96503a <=( a96502a  and  a96495a );
 a96507a <=( A266  and  A265 );
 a96508a <=( (not A202)  and  a96507a );
 a96511a <=( A269  and  (not A267) );
 a96514a <=( A300  and  A298 );
 a96515a <=( a96514a  and  a96511a );
 a96516a <=( a96515a  and  a96508a );
 a96520a <=( (not A167)  and  A168 );
 a96521a <=( A169  and  a96520a );
 a96524a <=( A199  and  A166 );
 a96527a <=( (not A201)  and  A200 );
 a96528a <=( a96527a  and  a96524a );
 a96529a <=( a96528a  and  a96521a );
 a96533a <=( A266  and  (not A265) );
 a96534a <=( (not A202)  and  a96533a );
 a96537a <=( A268  and  (not A267) );
 a96540a <=( A300  and  A299 );
 a96541a <=( a96540a  and  a96537a );
 a96542a <=( a96541a  and  a96534a );
 a96546a <=( (not A167)  and  A168 );
 a96547a <=( A169  and  a96546a );
 a96550a <=( A199  and  A166 );
 a96553a <=( (not A201)  and  A200 );
 a96554a <=( a96553a  and  a96550a );
 a96555a <=( a96554a  and  a96547a );
 a96559a <=( A266  and  (not A265) );
 a96560a <=( (not A202)  and  a96559a );
 a96563a <=( A268  and  (not A267) );
 a96566a <=( A300  and  A298 );
 a96567a <=( a96566a  and  a96563a );
 a96568a <=( a96567a  and  a96560a );
 a96572a <=( (not A167)  and  A168 );
 a96573a <=( A169  and  a96572a );
 a96576a <=( A199  and  A166 );
 a96579a <=( (not A201)  and  A200 );
 a96580a <=( a96579a  and  a96576a );
 a96581a <=( a96580a  and  a96573a );
 a96585a <=( A266  and  (not A265) );
 a96586a <=( (not A202)  and  a96585a );
 a96589a <=( (not A269)  and  (not A267) );
 a96592a <=( A300  and  A299 );
 a96593a <=( a96592a  and  a96589a );
 a96594a <=( a96593a  and  a96586a );
 a96598a <=( (not A167)  and  A168 );
 a96599a <=( A169  and  a96598a );
 a96602a <=( A199  and  A166 );
 a96605a <=( (not A201)  and  A200 );
 a96606a <=( a96605a  and  a96602a );
 a96607a <=( a96606a  and  a96599a );
 a96611a <=( A266  and  (not A265) );
 a96612a <=( (not A202)  and  a96611a );
 a96615a <=( (not A269)  and  (not A267) );
 a96618a <=( A300  and  A298 );
 a96619a <=( a96618a  and  a96615a );
 a96620a <=( a96619a  and  a96612a );
 a96624a <=( (not A167)  and  A168 );
 a96625a <=( A169  and  a96624a );
 a96628a <=( A199  and  A166 );
 a96631a <=( (not A201)  and  A200 );
 a96632a <=( a96631a  and  a96628a );
 a96633a <=( a96632a  and  a96625a );
 a96637a <=( (not A266)  and  A265 );
 a96638a <=( (not A202)  and  a96637a );
 a96641a <=( A268  and  (not A267) );
 a96644a <=( A300  and  A299 );
 a96645a <=( a96644a  and  a96641a );
 a96646a <=( a96645a  and  a96638a );
 a96650a <=( (not A167)  and  A168 );
 a96651a <=( A169  and  a96650a );
 a96654a <=( A199  and  A166 );
 a96657a <=( (not A201)  and  A200 );
 a96658a <=( a96657a  and  a96654a );
 a96659a <=( a96658a  and  a96651a );
 a96663a <=( (not A266)  and  A265 );
 a96664a <=( (not A202)  and  a96663a );
 a96667a <=( A268  and  (not A267) );
 a96670a <=( A300  and  A298 );
 a96671a <=( a96670a  and  a96667a );
 a96672a <=( a96671a  and  a96664a );
 a96676a <=( (not A167)  and  A168 );
 a96677a <=( A169  and  a96676a );
 a96680a <=( A199  and  A166 );
 a96683a <=( (not A201)  and  A200 );
 a96684a <=( a96683a  and  a96680a );
 a96685a <=( a96684a  and  a96677a );
 a96689a <=( (not A266)  and  A265 );
 a96690a <=( (not A202)  and  a96689a );
 a96693a <=( (not A269)  and  (not A267) );
 a96696a <=( A300  and  A299 );
 a96697a <=( a96696a  and  a96693a );
 a96698a <=( a96697a  and  a96690a );
 a96702a <=( (not A167)  and  A168 );
 a96703a <=( A169  and  a96702a );
 a96706a <=( A199  and  A166 );
 a96709a <=( (not A201)  and  A200 );
 a96710a <=( a96709a  and  a96706a );
 a96711a <=( a96710a  and  a96703a );
 a96715a <=( (not A266)  and  A265 );
 a96716a <=( (not A202)  and  a96715a );
 a96719a <=( (not A269)  and  (not A267) );
 a96722a <=( A300  and  A298 );
 a96723a <=( a96722a  and  a96719a );
 a96724a <=( a96723a  and  a96716a );
 a96728a <=( (not A167)  and  A168 );
 a96729a <=( A169  and  a96728a );
 a96732a <=( A199  and  A166 );
 a96735a <=( (not A201)  and  A200 );
 a96736a <=( a96735a  and  a96732a );
 a96737a <=( a96736a  and  a96729a );
 a96741a <=( A266  and  A265 );
 a96742a <=( A203  and  a96741a );
 a96745a <=( (not A268)  and  (not A267) );
 a96748a <=( A300  and  A299 );
 a96749a <=( a96748a  and  a96745a );
 a96750a <=( a96749a  and  a96742a );
 a96754a <=( (not A167)  and  A168 );
 a96755a <=( A169  and  a96754a );
 a96758a <=( A199  and  A166 );
 a96761a <=( (not A201)  and  A200 );
 a96762a <=( a96761a  and  a96758a );
 a96763a <=( a96762a  and  a96755a );
 a96767a <=( A266  and  A265 );
 a96768a <=( A203  and  a96767a );
 a96771a <=( (not A268)  and  (not A267) );
 a96774a <=( A300  and  A298 );
 a96775a <=( a96774a  and  a96771a );
 a96776a <=( a96775a  and  a96768a );
 a96780a <=( (not A167)  and  A168 );
 a96781a <=( A169  and  a96780a );
 a96784a <=( A199  and  A166 );
 a96787a <=( (not A201)  and  A200 );
 a96788a <=( a96787a  and  a96784a );
 a96789a <=( a96788a  and  a96781a );
 a96793a <=( A266  and  A265 );
 a96794a <=( A203  and  a96793a );
 a96797a <=( A269  and  (not A267) );
 a96800a <=( A300  and  A299 );
 a96801a <=( a96800a  and  a96797a );
 a96802a <=( a96801a  and  a96794a );
 a96806a <=( (not A167)  and  A168 );
 a96807a <=( A169  and  a96806a );
 a96810a <=( A199  and  A166 );
 a96813a <=( (not A201)  and  A200 );
 a96814a <=( a96813a  and  a96810a );
 a96815a <=( a96814a  and  a96807a );
 a96819a <=( A266  and  A265 );
 a96820a <=( A203  and  a96819a );
 a96823a <=( A269  and  (not A267) );
 a96826a <=( A300  and  A298 );
 a96827a <=( a96826a  and  a96823a );
 a96828a <=( a96827a  and  a96820a );
 a96832a <=( (not A167)  and  A168 );
 a96833a <=( A169  and  a96832a );
 a96836a <=( A199  and  A166 );
 a96839a <=( (not A201)  and  A200 );
 a96840a <=( a96839a  and  a96836a );
 a96841a <=( a96840a  and  a96833a );
 a96845a <=( A266  and  (not A265) );
 a96846a <=( A203  and  a96845a );
 a96849a <=( A268  and  (not A267) );
 a96852a <=( A300  and  A299 );
 a96853a <=( a96852a  and  a96849a );
 a96854a <=( a96853a  and  a96846a );
 a96858a <=( (not A167)  and  A168 );
 a96859a <=( A169  and  a96858a );
 a96862a <=( A199  and  A166 );
 a96865a <=( (not A201)  and  A200 );
 a96866a <=( a96865a  and  a96862a );
 a96867a <=( a96866a  and  a96859a );
 a96871a <=( A266  and  (not A265) );
 a96872a <=( A203  and  a96871a );
 a96875a <=( A268  and  (not A267) );
 a96878a <=( A300  and  A298 );
 a96879a <=( a96878a  and  a96875a );
 a96880a <=( a96879a  and  a96872a );
 a96884a <=( (not A167)  and  A168 );
 a96885a <=( A169  and  a96884a );
 a96888a <=( A199  and  A166 );
 a96891a <=( (not A201)  and  A200 );
 a96892a <=( a96891a  and  a96888a );
 a96893a <=( a96892a  and  a96885a );
 a96897a <=( A266  and  (not A265) );
 a96898a <=( A203  and  a96897a );
 a96901a <=( (not A269)  and  (not A267) );
 a96904a <=( A300  and  A299 );
 a96905a <=( a96904a  and  a96901a );
 a96906a <=( a96905a  and  a96898a );
 a96910a <=( (not A167)  and  A168 );
 a96911a <=( A169  and  a96910a );
 a96914a <=( A199  and  A166 );
 a96917a <=( (not A201)  and  A200 );
 a96918a <=( a96917a  and  a96914a );
 a96919a <=( a96918a  and  a96911a );
 a96923a <=( A266  and  (not A265) );
 a96924a <=( A203  and  a96923a );
 a96927a <=( (not A269)  and  (not A267) );
 a96930a <=( A300  and  A298 );
 a96931a <=( a96930a  and  a96927a );
 a96932a <=( a96931a  and  a96924a );
 a96936a <=( (not A167)  and  A168 );
 a96937a <=( A169  and  a96936a );
 a96940a <=( A199  and  A166 );
 a96943a <=( (not A201)  and  A200 );
 a96944a <=( a96943a  and  a96940a );
 a96945a <=( a96944a  and  a96937a );
 a96949a <=( (not A266)  and  A265 );
 a96950a <=( A203  and  a96949a );
 a96953a <=( A268  and  (not A267) );
 a96956a <=( A300  and  A299 );
 a96957a <=( a96956a  and  a96953a );
 a96958a <=( a96957a  and  a96950a );
 a96962a <=( (not A167)  and  A168 );
 a96963a <=( A169  and  a96962a );
 a96966a <=( A199  and  A166 );
 a96969a <=( (not A201)  and  A200 );
 a96970a <=( a96969a  and  a96966a );
 a96971a <=( a96970a  and  a96963a );
 a96975a <=( (not A266)  and  A265 );
 a96976a <=( A203  and  a96975a );
 a96979a <=( A268  and  (not A267) );
 a96982a <=( A300  and  A298 );
 a96983a <=( a96982a  and  a96979a );
 a96984a <=( a96983a  and  a96976a );
 a96988a <=( (not A167)  and  A168 );
 a96989a <=( A169  and  a96988a );
 a96992a <=( A199  and  A166 );
 a96995a <=( (not A201)  and  A200 );
 a96996a <=( a96995a  and  a96992a );
 a96997a <=( a96996a  and  a96989a );
 a97001a <=( (not A266)  and  A265 );
 a97002a <=( A203  and  a97001a );
 a97005a <=( (not A269)  and  (not A267) );
 a97008a <=( A300  and  A299 );
 a97009a <=( a97008a  and  a97005a );
 a97010a <=( a97009a  and  a97002a );
 a97014a <=( (not A167)  and  A168 );
 a97015a <=( A169  and  a97014a );
 a97018a <=( A199  and  A166 );
 a97021a <=( (not A201)  and  A200 );
 a97022a <=( a97021a  and  a97018a );
 a97023a <=( a97022a  and  a97015a );
 a97027a <=( (not A266)  and  A265 );
 a97028a <=( A203  and  a97027a );
 a97031a <=( (not A269)  and  (not A267) );
 a97034a <=( A300  and  A298 );
 a97035a <=( a97034a  and  a97031a );
 a97036a <=( a97035a  and  a97028a );
 a97040a <=( (not A167)  and  A168 );
 a97041a <=( A169  and  a97040a );
 a97044a <=( (not A199)  and  A166 );
 a97047a <=( (not A202)  and  A200 );
 a97048a <=( a97047a  and  a97044a );
 a97049a <=( a97048a  and  a97041a );
 a97053a <=( A267  and  A265 );
 a97054a <=( A203  and  a97053a );
 a97057a <=( A299  and  A298 );
 a97060a <=( (not A301)  and  (not A300) );
 a97061a <=( a97060a  and  a97057a );
 a97062a <=( a97061a  and  a97054a );
 a97066a <=( (not A167)  and  A168 );
 a97067a <=( A169  and  a97066a );
 a97070a <=( (not A199)  and  A166 );
 a97073a <=( (not A202)  and  A200 );
 a97074a <=( a97073a  and  a97070a );
 a97075a <=( a97074a  and  a97067a );
 a97079a <=( A267  and  A265 );
 a97080a <=( A203  and  a97079a );
 a97083a <=( A299  and  A298 );
 a97086a <=( A302  and  (not A300) );
 a97087a <=( a97086a  and  a97083a );
 a97088a <=( a97087a  and  a97080a );
 a97092a <=( (not A167)  and  A168 );
 a97093a <=( A169  and  a97092a );
 a97096a <=( (not A199)  and  A166 );
 a97099a <=( (not A202)  and  A200 );
 a97100a <=( a97099a  and  a97096a );
 a97101a <=( a97100a  and  a97093a );
 a97105a <=( A267  and  A265 );
 a97106a <=( A203  and  a97105a );
 a97109a <=( (not A299)  and  A298 );
 a97112a <=( A301  and  (not A300) );
 a97113a <=( a97112a  and  a97109a );
 a97114a <=( a97113a  and  a97106a );
 a97118a <=( (not A167)  and  A168 );
 a97119a <=( A169  and  a97118a );
 a97122a <=( (not A199)  and  A166 );
 a97125a <=( (not A202)  and  A200 );
 a97126a <=( a97125a  and  a97122a );
 a97127a <=( a97126a  and  a97119a );
 a97131a <=( A267  and  A265 );
 a97132a <=( A203  and  a97131a );
 a97135a <=( (not A299)  and  A298 );
 a97138a <=( (not A302)  and  (not A300) );
 a97139a <=( a97138a  and  a97135a );
 a97140a <=( a97139a  and  a97132a );
 a97144a <=( (not A167)  and  A168 );
 a97145a <=( A169  and  a97144a );
 a97148a <=( (not A199)  and  A166 );
 a97151a <=( (not A202)  and  A200 );
 a97152a <=( a97151a  and  a97148a );
 a97153a <=( a97152a  and  a97145a );
 a97157a <=( A267  and  A265 );
 a97158a <=( A203  and  a97157a );
 a97161a <=( A299  and  (not A298) );
 a97164a <=( A301  and  (not A300) );
 a97165a <=( a97164a  and  a97161a );
 a97166a <=( a97165a  and  a97158a );
 a97170a <=( (not A167)  and  A168 );
 a97171a <=( A169  and  a97170a );
 a97174a <=( (not A199)  and  A166 );
 a97177a <=( (not A202)  and  A200 );
 a97178a <=( a97177a  and  a97174a );
 a97179a <=( a97178a  and  a97171a );
 a97183a <=( A267  and  A265 );
 a97184a <=( A203  and  a97183a );
 a97187a <=( A299  and  (not A298) );
 a97190a <=( (not A302)  and  (not A300) );
 a97191a <=( a97190a  and  a97187a );
 a97192a <=( a97191a  and  a97184a );
 a97196a <=( (not A167)  and  A168 );
 a97197a <=( A169  and  a97196a );
 a97200a <=( (not A199)  and  A166 );
 a97203a <=( (not A202)  and  A200 );
 a97204a <=( a97203a  and  a97200a );
 a97205a <=( a97204a  and  a97197a );
 a97209a <=( A267  and  A266 );
 a97210a <=( A203  and  a97209a );
 a97213a <=( A299  and  A298 );
 a97216a <=( (not A301)  and  (not A300) );
 a97217a <=( a97216a  and  a97213a );
 a97218a <=( a97217a  and  a97210a );
 a97222a <=( (not A167)  and  A168 );
 a97223a <=( A169  and  a97222a );
 a97226a <=( (not A199)  and  A166 );
 a97229a <=( (not A202)  and  A200 );
 a97230a <=( a97229a  and  a97226a );
 a97231a <=( a97230a  and  a97223a );
 a97235a <=( A267  and  A266 );
 a97236a <=( A203  and  a97235a );
 a97239a <=( A299  and  A298 );
 a97242a <=( A302  and  (not A300) );
 a97243a <=( a97242a  and  a97239a );
 a97244a <=( a97243a  and  a97236a );
 a97248a <=( (not A167)  and  A168 );
 a97249a <=( A169  and  a97248a );
 a97252a <=( (not A199)  and  A166 );
 a97255a <=( (not A202)  and  A200 );
 a97256a <=( a97255a  and  a97252a );
 a97257a <=( a97256a  and  a97249a );
 a97261a <=( A267  and  A266 );
 a97262a <=( A203  and  a97261a );
 a97265a <=( (not A299)  and  A298 );
 a97268a <=( A301  and  (not A300) );
 a97269a <=( a97268a  and  a97265a );
 a97270a <=( a97269a  and  a97262a );
 a97274a <=( (not A167)  and  A168 );
 a97275a <=( A169  and  a97274a );
 a97278a <=( (not A199)  and  A166 );
 a97281a <=( (not A202)  and  A200 );
 a97282a <=( a97281a  and  a97278a );
 a97283a <=( a97282a  and  a97275a );
 a97287a <=( A267  and  A266 );
 a97288a <=( A203  and  a97287a );
 a97291a <=( (not A299)  and  A298 );
 a97294a <=( (not A302)  and  (not A300) );
 a97295a <=( a97294a  and  a97291a );
 a97296a <=( a97295a  and  a97288a );
 a97300a <=( (not A167)  and  A168 );
 a97301a <=( A169  and  a97300a );
 a97304a <=( (not A199)  and  A166 );
 a97307a <=( (not A202)  and  A200 );
 a97308a <=( a97307a  and  a97304a );
 a97309a <=( a97308a  and  a97301a );
 a97313a <=( A267  and  A266 );
 a97314a <=( A203  and  a97313a );
 a97317a <=( A299  and  (not A298) );
 a97320a <=( A301  and  (not A300) );
 a97321a <=( a97320a  and  a97317a );
 a97322a <=( a97321a  and  a97314a );
 a97326a <=( (not A167)  and  A168 );
 a97327a <=( A169  and  a97326a );
 a97330a <=( (not A199)  and  A166 );
 a97333a <=( (not A202)  and  A200 );
 a97334a <=( a97333a  and  a97330a );
 a97335a <=( a97334a  and  a97327a );
 a97339a <=( A267  and  A266 );
 a97340a <=( A203  and  a97339a );
 a97343a <=( A299  and  (not A298) );
 a97346a <=( (not A302)  and  (not A300) );
 a97347a <=( a97346a  and  a97343a );
 a97348a <=( a97347a  and  a97340a );
 a97352a <=( (not A167)  and  A168 );
 a97353a <=( A169  and  a97352a );
 a97356a <=( (not A199)  and  A166 );
 a97359a <=( (not A201)  and  A200 );
 a97360a <=( a97359a  and  a97356a );
 a97361a <=( a97360a  and  a97353a );
 a97365a <=( A266  and  A265 );
 a97366a <=( A202  and  a97365a );
 a97369a <=( (not A268)  and  (not A267) );
 a97372a <=( A300  and  A299 );
 a97373a <=( a97372a  and  a97369a );
 a97374a <=( a97373a  and  a97366a );
 a97378a <=( (not A167)  and  A168 );
 a97379a <=( A169  and  a97378a );
 a97382a <=( (not A199)  and  A166 );
 a97385a <=( (not A201)  and  A200 );
 a97386a <=( a97385a  and  a97382a );
 a97387a <=( a97386a  and  a97379a );
 a97391a <=( A266  and  A265 );
 a97392a <=( A202  and  a97391a );
 a97395a <=( (not A268)  and  (not A267) );
 a97398a <=( A300  and  A298 );
 a97399a <=( a97398a  and  a97395a );
 a97400a <=( a97399a  and  a97392a );
 a97404a <=( (not A167)  and  A168 );
 a97405a <=( A169  and  a97404a );
 a97408a <=( (not A199)  and  A166 );
 a97411a <=( (not A201)  and  A200 );
 a97412a <=( a97411a  and  a97408a );
 a97413a <=( a97412a  and  a97405a );
 a97417a <=( A266  and  A265 );
 a97418a <=( A202  and  a97417a );
 a97421a <=( A269  and  (not A267) );
 a97424a <=( A300  and  A299 );
 a97425a <=( a97424a  and  a97421a );
 a97426a <=( a97425a  and  a97418a );
 a97430a <=( (not A167)  and  A168 );
 a97431a <=( A169  and  a97430a );
 a97434a <=( (not A199)  and  A166 );
 a97437a <=( (not A201)  and  A200 );
 a97438a <=( a97437a  and  a97434a );
 a97439a <=( a97438a  and  a97431a );
 a97443a <=( A266  and  A265 );
 a97444a <=( A202  and  a97443a );
 a97447a <=( A269  and  (not A267) );
 a97450a <=( A300  and  A298 );
 a97451a <=( a97450a  and  a97447a );
 a97452a <=( a97451a  and  a97444a );
 a97456a <=( (not A167)  and  A168 );
 a97457a <=( A169  and  a97456a );
 a97460a <=( (not A199)  and  A166 );
 a97463a <=( (not A201)  and  A200 );
 a97464a <=( a97463a  and  a97460a );
 a97465a <=( a97464a  and  a97457a );
 a97469a <=( A266  and  (not A265) );
 a97470a <=( A202  and  a97469a );
 a97473a <=( A268  and  (not A267) );
 a97476a <=( A300  and  A299 );
 a97477a <=( a97476a  and  a97473a );
 a97478a <=( a97477a  and  a97470a );
 a97482a <=( (not A167)  and  A168 );
 a97483a <=( A169  and  a97482a );
 a97486a <=( (not A199)  and  A166 );
 a97489a <=( (not A201)  and  A200 );
 a97490a <=( a97489a  and  a97486a );
 a97491a <=( a97490a  and  a97483a );
 a97495a <=( A266  and  (not A265) );
 a97496a <=( A202  and  a97495a );
 a97499a <=( A268  and  (not A267) );
 a97502a <=( A300  and  A298 );
 a97503a <=( a97502a  and  a97499a );
 a97504a <=( a97503a  and  a97496a );
 a97508a <=( (not A167)  and  A168 );
 a97509a <=( A169  and  a97508a );
 a97512a <=( (not A199)  and  A166 );
 a97515a <=( (not A201)  and  A200 );
 a97516a <=( a97515a  and  a97512a );
 a97517a <=( a97516a  and  a97509a );
 a97521a <=( A266  and  (not A265) );
 a97522a <=( A202  and  a97521a );
 a97525a <=( (not A269)  and  (not A267) );
 a97528a <=( A300  and  A299 );
 a97529a <=( a97528a  and  a97525a );
 a97530a <=( a97529a  and  a97522a );
 a97534a <=( (not A167)  and  A168 );
 a97535a <=( A169  and  a97534a );
 a97538a <=( (not A199)  and  A166 );
 a97541a <=( (not A201)  and  A200 );
 a97542a <=( a97541a  and  a97538a );
 a97543a <=( a97542a  and  a97535a );
 a97547a <=( A266  and  (not A265) );
 a97548a <=( A202  and  a97547a );
 a97551a <=( (not A269)  and  (not A267) );
 a97554a <=( A300  and  A298 );
 a97555a <=( a97554a  and  a97551a );
 a97556a <=( a97555a  and  a97548a );
 a97560a <=( (not A167)  and  A168 );
 a97561a <=( A169  and  a97560a );
 a97564a <=( (not A199)  and  A166 );
 a97567a <=( (not A201)  and  A200 );
 a97568a <=( a97567a  and  a97564a );
 a97569a <=( a97568a  and  a97561a );
 a97573a <=( (not A266)  and  A265 );
 a97574a <=( A202  and  a97573a );
 a97577a <=( A268  and  (not A267) );
 a97580a <=( A300  and  A299 );
 a97581a <=( a97580a  and  a97577a );
 a97582a <=( a97581a  and  a97574a );
 a97586a <=( (not A167)  and  A168 );
 a97587a <=( A169  and  a97586a );
 a97590a <=( (not A199)  and  A166 );
 a97593a <=( (not A201)  and  A200 );
 a97594a <=( a97593a  and  a97590a );
 a97595a <=( a97594a  and  a97587a );
 a97599a <=( (not A266)  and  A265 );
 a97600a <=( A202  and  a97599a );
 a97603a <=( A268  and  (not A267) );
 a97606a <=( A300  and  A298 );
 a97607a <=( a97606a  and  a97603a );
 a97608a <=( a97607a  and  a97600a );
 a97612a <=( (not A167)  and  A168 );
 a97613a <=( A169  and  a97612a );
 a97616a <=( (not A199)  and  A166 );
 a97619a <=( (not A201)  and  A200 );
 a97620a <=( a97619a  and  a97616a );
 a97621a <=( a97620a  and  a97613a );
 a97625a <=( (not A266)  and  A265 );
 a97626a <=( A202  and  a97625a );
 a97629a <=( (not A269)  and  (not A267) );
 a97632a <=( A300  and  A299 );
 a97633a <=( a97632a  and  a97629a );
 a97634a <=( a97633a  and  a97626a );
 a97638a <=( (not A167)  and  A168 );
 a97639a <=( A169  and  a97638a );
 a97642a <=( (not A199)  and  A166 );
 a97645a <=( (not A201)  and  A200 );
 a97646a <=( a97645a  and  a97642a );
 a97647a <=( a97646a  and  a97639a );
 a97651a <=( (not A266)  and  A265 );
 a97652a <=( A202  and  a97651a );
 a97655a <=( (not A269)  and  (not A267) );
 a97658a <=( A300  and  A298 );
 a97659a <=( a97658a  and  a97655a );
 a97660a <=( a97659a  and  a97652a );
 a97664a <=( (not A167)  and  A168 );
 a97665a <=( A169  and  a97664a );
 a97668a <=( (not A199)  and  A166 );
 a97671a <=( (not A201)  and  A200 );
 a97672a <=( a97671a  and  a97668a );
 a97673a <=( a97672a  and  a97665a );
 a97677a <=( A266  and  A265 );
 a97678a <=( (not A203)  and  a97677a );
 a97681a <=( (not A268)  and  (not A267) );
 a97684a <=( A300  and  A299 );
 a97685a <=( a97684a  and  a97681a );
 a97686a <=( a97685a  and  a97678a );
 a97690a <=( (not A167)  and  A168 );
 a97691a <=( A169  and  a97690a );
 a97694a <=( (not A199)  and  A166 );
 a97697a <=( (not A201)  and  A200 );
 a97698a <=( a97697a  and  a97694a );
 a97699a <=( a97698a  and  a97691a );
 a97703a <=( A266  and  A265 );
 a97704a <=( (not A203)  and  a97703a );
 a97707a <=( (not A268)  and  (not A267) );
 a97710a <=( A300  and  A298 );
 a97711a <=( a97710a  and  a97707a );
 a97712a <=( a97711a  and  a97704a );
 a97716a <=( (not A167)  and  A168 );
 a97717a <=( A169  and  a97716a );
 a97720a <=( (not A199)  and  A166 );
 a97723a <=( (not A201)  and  A200 );
 a97724a <=( a97723a  and  a97720a );
 a97725a <=( a97724a  and  a97717a );
 a97729a <=( A266  and  A265 );
 a97730a <=( (not A203)  and  a97729a );
 a97733a <=( A269  and  (not A267) );
 a97736a <=( A300  and  A299 );
 a97737a <=( a97736a  and  a97733a );
 a97738a <=( a97737a  and  a97730a );
 a97742a <=( (not A167)  and  A168 );
 a97743a <=( A169  and  a97742a );
 a97746a <=( (not A199)  and  A166 );
 a97749a <=( (not A201)  and  A200 );
 a97750a <=( a97749a  and  a97746a );
 a97751a <=( a97750a  and  a97743a );
 a97755a <=( A266  and  A265 );
 a97756a <=( (not A203)  and  a97755a );
 a97759a <=( A269  and  (not A267) );
 a97762a <=( A300  and  A298 );
 a97763a <=( a97762a  and  a97759a );
 a97764a <=( a97763a  and  a97756a );
 a97768a <=( (not A167)  and  A168 );
 a97769a <=( A169  and  a97768a );
 a97772a <=( (not A199)  and  A166 );
 a97775a <=( (not A201)  and  A200 );
 a97776a <=( a97775a  and  a97772a );
 a97777a <=( a97776a  and  a97769a );
 a97781a <=( A266  and  (not A265) );
 a97782a <=( (not A203)  and  a97781a );
 a97785a <=( A268  and  (not A267) );
 a97788a <=( A300  and  A299 );
 a97789a <=( a97788a  and  a97785a );
 a97790a <=( a97789a  and  a97782a );
 a97794a <=( (not A167)  and  A168 );
 a97795a <=( A169  and  a97794a );
 a97798a <=( (not A199)  and  A166 );
 a97801a <=( (not A201)  and  A200 );
 a97802a <=( a97801a  and  a97798a );
 a97803a <=( a97802a  and  a97795a );
 a97807a <=( A266  and  (not A265) );
 a97808a <=( (not A203)  and  a97807a );
 a97811a <=( A268  and  (not A267) );
 a97814a <=( A300  and  A298 );
 a97815a <=( a97814a  and  a97811a );
 a97816a <=( a97815a  and  a97808a );
 a97820a <=( (not A167)  and  A168 );
 a97821a <=( A169  and  a97820a );
 a97824a <=( (not A199)  and  A166 );
 a97827a <=( (not A201)  and  A200 );
 a97828a <=( a97827a  and  a97824a );
 a97829a <=( a97828a  and  a97821a );
 a97833a <=( A266  and  (not A265) );
 a97834a <=( (not A203)  and  a97833a );
 a97837a <=( (not A269)  and  (not A267) );
 a97840a <=( A300  and  A299 );
 a97841a <=( a97840a  and  a97837a );
 a97842a <=( a97841a  and  a97834a );
 a97846a <=( (not A167)  and  A168 );
 a97847a <=( A169  and  a97846a );
 a97850a <=( (not A199)  and  A166 );
 a97853a <=( (not A201)  and  A200 );
 a97854a <=( a97853a  and  a97850a );
 a97855a <=( a97854a  and  a97847a );
 a97859a <=( A266  and  (not A265) );
 a97860a <=( (not A203)  and  a97859a );
 a97863a <=( (not A269)  and  (not A267) );
 a97866a <=( A300  and  A298 );
 a97867a <=( a97866a  and  a97863a );
 a97868a <=( a97867a  and  a97860a );
 a97872a <=( (not A167)  and  A168 );
 a97873a <=( A169  and  a97872a );
 a97876a <=( (not A199)  and  A166 );
 a97879a <=( (not A201)  and  A200 );
 a97880a <=( a97879a  and  a97876a );
 a97881a <=( a97880a  and  a97873a );
 a97885a <=( (not A266)  and  A265 );
 a97886a <=( (not A203)  and  a97885a );
 a97889a <=( A268  and  (not A267) );
 a97892a <=( A300  and  A299 );
 a97893a <=( a97892a  and  a97889a );
 a97894a <=( a97893a  and  a97886a );
 a97898a <=( (not A167)  and  A168 );
 a97899a <=( A169  and  a97898a );
 a97902a <=( (not A199)  and  A166 );
 a97905a <=( (not A201)  and  A200 );
 a97906a <=( a97905a  and  a97902a );
 a97907a <=( a97906a  and  a97899a );
 a97911a <=( (not A266)  and  A265 );
 a97912a <=( (not A203)  and  a97911a );
 a97915a <=( A268  and  (not A267) );
 a97918a <=( A300  and  A298 );
 a97919a <=( a97918a  and  a97915a );
 a97920a <=( a97919a  and  a97912a );
 a97924a <=( (not A167)  and  A168 );
 a97925a <=( A169  and  a97924a );
 a97928a <=( (not A199)  and  A166 );
 a97931a <=( (not A201)  and  A200 );
 a97932a <=( a97931a  and  a97928a );
 a97933a <=( a97932a  and  a97925a );
 a97937a <=( (not A266)  and  A265 );
 a97938a <=( (not A203)  and  a97937a );
 a97941a <=( (not A269)  and  (not A267) );
 a97944a <=( A300  and  A299 );
 a97945a <=( a97944a  and  a97941a );
 a97946a <=( a97945a  and  a97938a );
 a97950a <=( (not A167)  and  A168 );
 a97951a <=( A169  and  a97950a );
 a97954a <=( (not A199)  and  A166 );
 a97957a <=( (not A201)  and  A200 );
 a97958a <=( a97957a  and  a97954a );
 a97959a <=( a97958a  and  a97951a );
 a97963a <=( (not A266)  and  A265 );
 a97964a <=( (not A203)  and  a97963a );
 a97967a <=( (not A269)  and  (not A267) );
 a97970a <=( A300  and  A298 );
 a97971a <=( a97970a  and  a97967a );
 a97972a <=( a97971a  and  a97964a );
 a97976a <=( (not A167)  and  A168 );
 a97977a <=( A169  and  a97976a );
 a97980a <=( A199  and  A166 );
 a97983a <=( (not A202)  and  (not A200) );
 a97984a <=( a97983a  and  a97980a );
 a97985a <=( a97984a  and  a97977a );
 a97989a <=( A267  and  A265 );
 a97990a <=( A203  and  a97989a );
 a97993a <=( A299  and  A298 );
 a97996a <=( (not A301)  and  (not A300) );
 a97997a <=( a97996a  and  a97993a );
 a97998a <=( a97997a  and  a97990a );
 a98002a <=( (not A167)  and  A168 );
 a98003a <=( A169  and  a98002a );
 a98006a <=( A199  and  A166 );
 a98009a <=( (not A202)  and  (not A200) );
 a98010a <=( a98009a  and  a98006a );
 a98011a <=( a98010a  and  a98003a );
 a98015a <=( A267  and  A265 );
 a98016a <=( A203  and  a98015a );
 a98019a <=( A299  and  A298 );
 a98022a <=( A302  and  (not A300) );
 a98023a <=( a98022a  and  a98019a );
 a98024a <=( a98023a  and  a98016a );
 a98028a <=( (not A167)  and  A168 );
 a98029a <=( A169  and  a98028a );
 a98032a <=( A199  and  A166 );
 a98035a <=( (not A202)  and  (not A200) );
 a98036a <=( a98035a  and  a98032a );
 a98037a <=( a98036a  and  a98029a );
 a98041a <=( A267  and  A265 );
 a98042a <=( A203  and  a98041a );
 a98045a <=( (not A299)  and  A298 );
 a98048a <=( A301  and  (not A300) );
 a98049a <=( a98048a  and  a98045a );
 a98050a <=( a98049a  and  a98042a );
 a98054a <=( (not A167)  and  A168 );
 a98055a <=( A169  and  a98054a );
 a98058a <=( A199  and  A166 );
 a98061a <=( (not A202)  and  (not A200) );
 a98062a <=( a98061a  and  a98058a );
 a98063a <=( a98062a  and  a98055a );
 a98067a <=( A267  and  A265 );
 a98068a <=( A203  and  a98067a );
 a98071a <=( (not A299)  and  A298 );
 a98074a <=( (not A302)  and  (not A300) );
 a98075a <=( a98074a  and  a98071a );
 a98076a <=( a98075a  and  a98068a );
 a98080a <=( (not A167)  and  A168 );
 a98081a <=( A169  and  a98080a );
 a98084a <=( A199  and  A166 );
 a98087a <=( (not A202)  and  (not A200) );
 a98088a <=( a98087a  and  a98084a );
 a98089a <=( a98088a  and  a98081a );
 a98093a <=( A267  and  A265 );
 a98094a <=( A203  and  a98093a );
 a98097a <=( A299  and  (not A298) );
 a98100a <=( A301  and  (not A300) );
 a98101a <=( a98100a  and  a98097a );
 a98102a <=( a98101a  and  a98094a );
 a98106a <=( (not A167)  and  A168 );
 a98107a <=( A169  and  a98106a );
 a98110a <=( A199  and  A166 );
 a98113a <=( (not A202)  and  (not A200) );
 a98114a <=( a98113a  and  a98110a );
 a98115a <=( a98114a  and  a98107a );
 a98119a <=( A267  and  A265 );
 a98120a <=( A203  and  a98119a );
 a98123a <=( A299  and  (not A298) );
 a98126a <=( (not A302)  and  (not A300) );
 a98127a <=( a98126a  and  a98123a );
 a98128a <=( a98127a  and  a98120a );
 a98132a <=( (not A167)  and  A168 );
 a98133a <=( A169  and  a98132a );
 a98136a <=( A199  and  A166 );
 a98139a <=( (not A202)  and  (not A200) );
 a98140a <=( a98139a  and  a98136a );
 a98141a <=( a98140a  and  a98133a );
 a98145a <=( A267  and  A266 );
 a98146a <=( A203  and  a98145a );
 a98149a <=( A299  and  A298 );
 a98152a <=( (not A301)  and  (not A300) );
 a98153a <=( a98152a  and  a98149a );
 a98154a <=( a98153a  and  a98146a );
 a98158a <=( (not A167)  and  A168 );
 a98159a <=( A169  and  a98158a );
 a98162a <=( A199  and  A166 );
 a98165a <=( (not A202)  and  (not A200) );
 a98166a <=( a98165a  and  a98162a );
 a98167a <=( a98166a  and  a98159a );
 a98171a <=( A267  and  A266 );
 a98172a <=( A203  and  a98171a );
 a98175a <=( A299  and  A298 );
 a98178a <=( A302  and  (not A300) );
 a98179a <=( a98178a  and  a98175a );
 a98180a <=( a98179a  and  a98172a );
 a98184a <=( (not A167)  and  A168 );
 a98185a <=( A169  and  a98184a );
 a98188a <=( A199  and  A166 );
 a98191a <=( (not A202)  and  (not A200) );
 a98192a <=( a98191a  and  a98188a );
 a98193a <=( a98192a  and  a98185a );
 a98197a <=( A267  and  A266 );
 a98198a <=( A203  and  a98197a );
 a98201a <=( (not A299)  and  A298 );
 a98204a <=( A301  and  (not A300) );
 a98205a <=( a98204a  and  a98201a );
 a98206a <=( a98205a  and  a98198a );
 a98210a <=( (not A167)  and  A168 );
 a98211a <=( A169  and  a98210a );
 a98214a <=( A199  and  A166 );
 a98217a <=( (not A202)  and  (not A200) );
 a98218a <=( a98217a  and  a98214a );
 a98219a <=( a98218a  and  a98211a );
 a98223a <=( A267  and  A266 );
 a98224a <=( A203  and  a98223a );
 a98227a <=( (not A299)  and  A298 );
 a98230a <=( (not A302)  and  (not A300) );
 a98231a <=( a98230a  and  a98227a );
 a98232a <=( a98231a  and  a98224a );
 a98236a <=( (not A167)  and  A168 );
 a98237a <=( A169  and  a98236a );
 a98240a <=( A199  and  A166 );
 a98243a <=( (not A202)  and  (not A200) );
 a98244a <=( a98243a  and  a98240a );
 a98245a <=( a98244a  and  a98237a );
 a98249a <=( A267  and  A266 );
 a98250a <=( A203  and  a98249a );
 a98253a <=( A299  and  (not A298) );
 a98256a <=( A301  and  (not A300) );
 a98257a <=( a98256a  and  a98253a );
 a98258a <=( a98257a  and  a98250a );
 a98262a <=( (not A167)  and  A168 );
 a98263a <=( A169  and  a98262a );
 a98266a <=( A199  and  A166 );
 a98269a <=( (not A202)  and  (not A200) );
 a98270a <=( a98269a  and  a98266a );
 a98271a <=( a98270a  and  a98263a );
 a98275a <=( A267  and  A266 );
 a98276a <=( A203  and  a98275a );
 a98279a <=( A299  and  (not A298) );
 a98282a <=( (not A302)  and  (not A300) );
 a98283a <=( a98282a  and  a98279a );
 a98284a <=( a98283a  and  a98276a );
 a98288a <=( (not A167)  and  A168 );
 a98289a <=( A169  and  a98288a );
 a98292a <=( A199  and  A166 );
 a98295a <=( (not A201)  and  (not A200) );
 a98296a <=( a98295a  and  a98292a );
 a98297a <=( a98296a  and  a98289a );
 a98301a <=( A266  and  A265 );
 a98302a <=( A202  and  a98301a );
 a98305a <=( (not A268)  and  (not A267) );
 a98308a <=( A300  and  A299 );
 a98309a <=( a98308a  and  a98305a );
 a98310a <=( a98309a  and  a98302a );
 a98314a <=( (not A167)  and  A168 );
 a98315a <=( A169  and  a98314a );
 a98318a <=( A199  and  A166 );
 a98321a <=( (not A201)  and  (not A200) );
 a98322a <=( a98321a  and  a98318a );
 a98323a <=( a98322a  and  a98315a );
 a98327a <=( A266  and  A265 );
 a98328a <=( A202  and  a98327a );
 a98331a <=( (not A268)  and  (not A267) );
 a98334a <=( A300  and  A298 );
 a98335a <=( a98334a  and  a98331a );
 a98336a <=( a98335a  and  a98328a );
 a98340a <=( (not A167)  and  A168 );
 a98341a <=( A169  and  a98340a );
 a98344a <=( A199  and  A166 );
 a98347a <=( (not A201)  and  (not A200) );
 a98348a <=( a98347a  and  a98344a );
 a98349a <=( a98348a  and  a98341a );
 a98353a <=( A266  and  A265 );
 a98354a <=( A202  and  a98353a );
 a98357a <=( A269  and  (not A267) );
 a98360a <=( A300  and  A299 );
 a98361a <=( a98360a  and  a98357a );
 a98362a <=( a98361a  and  a98354a );
 a98366a <=( (not A167)  and  A168 );
 a98367a <=( A169  and  a98366a );
 a98370a <=( A199  and  A166 );
 a98373a <=( (not A201)  and  (not A200) );
 a98374a <=( a98373a  and  a98370a );
 a98375a <=( a98374a  and  a98367a );
 a98379a <=( A266  and  A265 );
 a98380a <=( A202  and  a98379a );
 a98383a <=( A269  and  (not A267) );
 a98386a <=( A300  and  A298 );
 a98387a <=( a98386a  and  a98383a );
 a98388a <=( a98387a  and  a98380a );
 a98392a <=( (not A167)  and  A168 );
 a98393a <=( A169  and  a98392a );
 a98396a <=( A199  and  A166 );
 a98399a <=( (not A201)  and  (not A200) );
 a98400a <=( a98399a  and  a98396a );
 a98401a <=( a98400a  and  a98393a );
 a98405a <=( A266  and  (not A265) );
 a98406a <=( A202  and  a98405a );
 a98409a <=( A268  and  (not A267) );
 a98412a <=( A300  and  A299 );
 a98413a <=( a98412a  and  a98409a );
 a98414a <=( a98413a  and  a98406a );
 a98418a <=( (not A167)  and  A168 );
 a98419a <=( A169  and  a98418a );
 a98422a <=( A199  and  A166 );
 a98425a <=( (not A201)  and  (not A200) );
 a98426a <=( a98425a  and  a98422a );
 a98427a <=( a98426a  and  a98419a );
 a98431a <=( A266  and  (not A265) );
 a98432a <=( A202  and  a98431a );
 a98435a <=( A268  and  (not A267) );
 a98438a <=( A300  and  A298 );
 a98439a <=( a98438a  and  a98435a );
 a98440a <=( a98439a  and  a98432a );
 a98444a <=( (not A167)  and  A168 );
 a98445a <=( A169  and  a98444a );
 a98448a <=( A199  and  A166 );
 a98451a <=( (not A201)  and  (not A200) );
 a98452a <=( a98451a  and  a98448a );
 a98453a <=( a98452a  and  a98445a );
 a98457a <=( A266  and  (not A265) );
 a98458a <=( A202  and  a98457a );
 a98461a <=( (not A269)  and  (not A267) );
 a98464a <=( A300  and  A299 );
 a98465a <=( a98464a  and  a98461a );
 a98466a <=( a98465a  and  a98458a );
 a98470a <=( (not A167)  and  A168 );
 a98471a <=( A169  and  a98470a );
 a98474a <=( A199  and  A166 );
 a98477a <=( (not A201)  and  (not A200) );
 a98478a <=( a98477a  and  a98474a );
 a98479a <=( a98478a  and  a98471a );
 a98483a <=( A266  and  (not A265) );
 a98484a <=( A202  and  a98483a );
 a98487a <=( (not A269)  and  (not A267) );
 a98490a <=( A300  and  A298 );
 a98491a <=( a98490a  and  a98487a );
 a98492a <=( a98491a  and  a98484a );
 a98496a <=( (not A167)  and  A168 );
 a98497a <=( A169  and  a98496a );
 a98500a <=( A199  and  A166 );
 a98503a <=( (not A201)  and  (not A200) );
 a98504a <=( a98503a  and  a98500a );
 a98505a <=( a98504a  and  a98497a );
 a98509a <=( (not A266)  and  A265 );
 a98510a <=( A202  and  a98509a );
 a98513a <=( A268  and  (not A267) );
 a98516a <=( A300  and  A299 );
 a98517a <=( a98516a  and  a98513a );
 a98518a <=( a98517a  and  a98510a );
 a98522a <=( (not A167)  and  A168 );
 a98523a <=( A169  and  a98522a );
 a98526a <=( A199  and  A166 );
 a98529a <=( (not A201)  and  (not A200) );
 a98530a <=( a98529a  and  a98526a );
 a98531a <=( a98530a  and  a98523a );
 a98535a <=( (not A266)  and  A265 );
 a98536a <=( A202  and  a98535a );
 a98539a <=( A268  and  (not A267) );
 a98542a <=( A300  and  A298 );
 a98543a <=( a98542a  and  a98539a );
 a98544a <=( a98543a  and  a98536a );
 a98548a <=( (not A167)  and  A168 );
 a98549a <=( A169  and  a98548a );
 a98552a <=( A199  and  A166 );
 a98555a <=( (not A201)  and  (not A200) );
 a98556a <=( a98555a  and  a98552a );
 a98557a <=( a98556a  and  a98549a );
 a98561a <=( (not A266)  and  A265 );
 a98562a <=( A202  and  a98561a );
 a98565a <=( (not A269)  and  (not A267) );
 a98568a <=( A300  and  A299 );
 a98569a <=( a98568a  and  a98565a );
 a98570a <=( a98569a  and  a98562a );
 a98574a <=( (not A167)  and  A168 );
 a98575a <=( A169  and  a98574a );
 a98578a <=( A199  and  A166 );
 a98581a <=( (not A201)  and  (not A200) );
 a98582a <=( a98581a  and  a98578a );
 a98583a <=( a98582a  and  a98575a );
 a98587a <=( (not A266)  and  A265 );
 a98588a <=( A202  and  a98587a );
 a98591a <=( (not A269)  and  (not A267) );
 a98594a <=( A300  and  A298 );
 a98595a <=( a98594a  and  a98591a );
 a98596a <=( a98595a  and  a98588a );
 a98600a <=( (not A167)  and  A168 );
 a98601a <=( A169  and  a98600a );
 a98604a <=( A199  and  A166 );
 a98607a <=( (not A201)  and  (not A200) );
 a98608a <=( a98607a  and  a98604a );
 a98609a <=( a98608a  and  a98601a );
 a98613a <=( A266  and  A265 );
 a98614a <=( (not A203)  and  a98613a );
 a98617a <=( (not A268)  and  (not A267) );
 a98620a <=( A300  and  A299 );
 a98621a <=( a98620a  and  a98617a );
 a98622a <=( a98621a  and  a98614a );
 a98626a <=( (not A167)  and  A168 );
 a98627a <=( A169  and  a98626a );
 a98630a <=( A199  and  A166 );
 a98633a <=( (not A201)  and  (not A200) );
 a98634a <=( a98633a  and  a98630a );
 a98635a <=( a98634a  and  a98627a );
 a98639a <=( A266  and  A265 );
 a98640a <=( (not A203)  and  a98639a );
 a98643a <=( (not A268)  and  (not A267) );
 a98646a <=( A300  and  A298 );
 a98647a <=( a98646a  and  a98643a );
 a98648a <=( a98647a  and  a98640a );
 a98652a <=( (not A167)  and  A168 );
 a98653a <=( A169  and  a98652a );
 a98656a <=( A199  and  A166 );
 a98659a <=( (not A201)  and  (not A200) );
 a98660a <=( a98659a  and  a98656a );
 a98661a <=( a98660a  and  a98653a );
 a98665a <=( A266  and  A265 );
 a98666a <=( (not A203)  and  a98665a );
 a98669a <=( A269  and  (not A267) );
 a98672a <=( A300  and  A299 );
 a98673a <=( a98672a  and  a98669a );
 a98674a <=( a98673a  and  a98666a );
 a98678a <=( (not A167)  and  A168 );
 a98679a <=( A169  and  a98678a );
 a98682a <=( A199  and  A166 );
 a98685a <=( (not A201)  and  (not A200) );
 a98686a <=( a98685a  and  a98682a );
 a98687a <=( a98686a  and  a98679a );
 a98691a <=( A266  and  A265 );
 a98692a <=( (not A203)  and  a98691a );
 a98695a <=( A269  and  (not A267) );
 a98698a <=( A300  and  A298 );
 a98699a <=( a98698a  and  a98695a );
 a98700a <=( a98699a  and  a98692a );
 a98704a <=( (not A167)  and  A168 );
 a98705a <=( A169  and  a98704a );
 a98708a <=( A199  and  A166 );
 a98711a <=( (not A201)  and  (not A200) );
 a98712a <=( a98711a  and  a98708a );
 a98713a <=( a98712a  and  a98705a );
 a98717a <=( A266  and  (not A265) );
 a98718a <=( (not A203)  and  a98717a );
 a98721a <=( A268  and  (not A267) );
 a98724a <=( A300  and  A299 );
 a98725a <=( a98724a  and  a98721a );
 a98726a <=( a98725a  and  a98718a );
 a98730a <=( (not A167)  and  A168 );
 a98731a <=( A169  and  a98730a );
 a98734a <=( A199  and  A166 );
 a98737a <=( (not A201)  and  (not A200) );
 a98738a <=( a98737a  and  a98734a );
 a98739a <=( a98738a  and  a98731a );
 a98743a <=( A266  and  (not A265) );
 a98744a <=( (not A203)  and  a98743a );
 a98747a <=( A268  and  (not A267) );
 a98750a <=( A300  and  A298 );
 a98751a <=( a98750a  and  a98747a );
 a98752a <=( a98751a  and  a98744a );
 a98756a <=( (not A167)  and  A168 );
 a98757a <=( A169  and  a98756a );
 a98760a <=( A199  and  A166 );
 a98763a <=( (not A201)  and  (not A200) );
 a98764a <=( a98763a  and  a98760a );
 a98765a <=( a98764a  and  a98757a );
 a98769a <=( A266  and  (not A265) );
 a98770a <=( (not A203)  and  a98769a );
 a98773a <=( (not A269)  and  (not A267) );
 a98776a <=( A300  and  A299 );
 a98777a <=( a98776a  and  a98773a );
 a98778a <=( a98777a  and  a98770a );
 a98782a <=( (not A167)  and  A168 );
 a98783a <=( A169  and  a98782a );
 a98786a <=( A199  and  A166 );
 a98789a <=( (not A201)  and  (not A200) );
 a98790a <=( a98789a  and  a98786a );
 a98791a <=( a98790a  and  a98783a );
 a98795a <=( A266  and  (not A265) );
 a98796a <=( (not A203)  and  a98795a );
 a98799a <=( (not A269)  and  (not A267) );
 a98802a <=( A300  and  A298 );
 a98803a <=( a98802a  and  a98799a );
 a98804a <=( a98803a  and  a98796a );
 a98808a <=( (not A167)  and  A168 );
 a98809a <=( A169  and  a98808a );
 a98812a <=( A199  and  A166 );
 a98815a <=( (not A201)  and  (not A200) );
 a98816a <=( a98815a  and  a98812a );
 a98817a <=( a98816a  and  a98809a );
 a98821a <=( (not A266)  and  A265 );
 a98822a <=( (not A203)  and  a98821a );
 a98825a <=( A268  and  (not A267) );
 a98828a <=( A300  and  A299 );
 a98829a <=( a98828a  and  a98825a );
 a98830a <=( a98829a  and  a98822a );
 a98834a <=( (not A167)  and  A168 );
 a98835a <=( A169  and  a98834a );
 a98838a <=( A199  and  A166 );
 a98841a <=( (not A201)  and  (not A200) );
 a98842a <=( a98841a  and  a98838a );
 a98843a <=( a98842a  and  a98835a );
 a98847a <=( (not A266)  and  A265 );
 a98848a <=( (not A203)  and  a98847a );
 a98851a <=( A268  and  (not A267) );
 a98854a <=( A300  and  A298 );
 a98855a <=( a98854a  and  a98851a );
 a98856a <=( a98855a  and  a98848a );
 a98860a <=( (not A167)  and  A168 );
 a98861a <=( A169  and  a98860a );
 a98864a <=( A199  and  A166 );
 a98867a <=( (not A201)  and  (not A200) );
 a98868a <=( a98867a  and  a98864a );
 a98869a <=( a98868a  and  a98861a );
 a98873a <=( (not A266)  and  A265 );
 a98874a <=( (not A203)  and  a98873a );
 a98877a <=( (not A269)  and  (not A267) );
 a98880a <=( A300  and  A299 );
 a98881a <=( a98880a  and  a98877a );
 a98882a <=( a98881a  and  a98874a );
 a98886a <=( (not A167)  and  A168 );
 a98887a <=( A169  and  a98886a );
 a98890a <=( A199  and  A166 );
 a98893a <=( (not A201)  and  (not A200) );
 a98894a <=( a98893a  and  a98890a );
 a98895a <=( a98894a  and  a98887a );
 a98899a <=( (not A266)  and  A265 );
 a98900a <=( (not A203)  and  a98899a );
 a98903a <=( (not A269)  and  (not A267) );
 a98906a <=( A300  and  A298 );
 a98907a <=( a98906a  and  a98903a );
 a98908a <=( a98907a  and  a98900a );
 a98912a <=( (not A167)  and  A168 );
 a98913a <=( A169  and  a98912a );
 a98916a <=( (not A199)  and  A166 );
 a98919a <=( (not A202)  and  (not A200) );
 a98920a <=( a98919a  and  a98916a );
 a98921a <=( a98920a  and  a98913a );
 a98925a <=( (not A268)  and  (not A266) );
 a98926a <=( (not A265)  and  a98925a );
 a98929a <=( A299  and  A298 );
 a98932a <=( (not A302)  and  A301 );
 a98933a <=( a98932a  and  a98929a );
 a98934a <=( a98933a  and  a98926a );
 a98938a <=( (not A167)  and  A168 );
 a98939a <=( A169  and  a98938a );
 a98942a <=( (not A199)  and  A166 );
 a98945a <=( (not A202)  and  (not A200) );
 a98946a <=( a98945a  and  a98942a );
 a98947a <=( a98946a  and  a98939a );
 a98951a <=( (not A268)  and  (not A266) );
 a98952a <=( (not A265)  and  a98951a );
 a98955a <=( (not A299)  and  A298 );
 a98958a <=( A302  and  (not A301) );
 a98959a <=( a98958a  and  a98955a );
 a98960a <=( a98959a  and  a98952a );
 a98964a <=( (not A167)  and  A168 );
 a98965a <=( A169  and  a98964a );
 a98968a <=( (not A199)  and  A166 );
 a98971a <=( (not A202)  and  (not A200) );
 a98972a <=( a98971a  and  a98968a );
 a98973a <=( a98972a  and  a98965a );
 a98977a <=( (not A268)  and  (not A266) );
 a98978a <=( (not A265)  and  a98977a );
 a98981a <=( A299  and  (not A298) );
 a98984a <=( A302  and  (not A301) );
 a98985a <=( a98984a  and  a98981a );
 a98986a <=( a98985a  and  a98978a );
 a98990a <=( (not A167)  and  A168 );
 a98991a <=( A169  and  a98990a );
 a98994a <=( (not A199)  and  A166 );
 a98997a <=( (not A202)  and  (not A200) );
 a98998a <=( a98997a  and  a98994a );
 a98999a <=( a98998a  and  a98991a );
 a99003a <=( (not A268)  and  (not A266) );
 a99004a <=( (not A265)  and  a99003a );
 a99007a <=( (not A299)  and  (not A298) );
 a99010a <=( (not A302)  and  A301 );
 a99011a <=( a99010a  and  a99007a );
 a99012a <=( a99011a  and  a99004a );
 a99016a <=( (not A167)  and  A168 );
 a99017a <=( A169  and  a99016a );
 a99020a <=( (not A199)  and  A166 );
 a99023a <=( (not A202)  and  (not A200) );
 a99024a <=( a99023a  and  a99020a );
 a99025a <=( a99024a  and  a99017a );
 a99029a <=( A269  and  (not A266) );
 a99030a <=( (not A265)  and  a99029a );
 a99033a <=( A299  and  A298 );
 a99036a <=( (not A302)  and  A301 );
 a99037a <=( a99036a  and  a99033a );
 a99038a <=( a99037a  and  a99030a );
 a99042a <=( (not A167)  and  A168 );
 a99043a <=( A169  and  a99042a );
 a99046a <=( (not A199)  and  A166 );
 a99049a <=( (not A202)  and  (not A200) );
 a99050a <=( a99049a  and  a99046a );
 a99051a <=( a99050a  and  a99043a );
 a99055a <=( A269  and  (not A266) );
 a99056a <=( (not A265)  and  a99055a );
 a99059a <=( (not A299)  and  A298 );
 a99062a <=( A302  and  (not A301) );
 a99063a <=( a99062a  and  a99059a );
 a99064a <=( a99063a  and  a99056a );
 a99068a <=( (not A167)  and  A168 );
 a99069a <=( A169  and  a99068a );
 a99072a <=( (not A199)  and  A166 );
 a99075a <=( (not A202)  and  (not A200) );
 a99076a <=( a99075a  and  a99072a );
 a99077a <=( a99076a  and  a99069a );
 a99081a <=( A269  and  (not A266) );
 a99082a <=( (not A265)  and  a99081a );
 a99085a <=( A299  and  (not A298) );
 a99088a <=( A302  and  (not A301) );
 a99089a <=( a99088a  and  a99085a );
 a99090a <=( a99089a  and  a99082a );
 a99094a <=( (not A167)  and  A168 );
 a99095a <=( A169  and  a99094a );
 a99098a <=( (not A199)  and  A166 );
 a99101a <=( (not A202)  and  (not A200) );
 a99102a <=( a99101a  and  a99098a );
 a99103a <=( a99102a  and  a99095a );
 a99107a <=( A269  and  (not A266) );
 a99108a <=( (not A265)  and  a99107a );
 a99111a <=( (not A299)  and  (not A298) );
 a99114a <=( (not A302)  and  A301 );
 a99115a <=( a99114a  and  a99111a );
 a99116a <=( a99115a  and  a99108a );
 a99120a <=( (not A167)  and  A168 );
 a99121a <=( A169  and  a99120a );
 a99124a <=( (not A199)  and  A166 );
 a99127a <=( A203  and  (not A200) );
 a99128a <=( a99127a  and  a99124a );
 a99129a <=( a99128a  and  a99121a );
 a99133a <=( (not A268)  and  (not A266) );
 a99134a <=( (not A265)  and  a99133a );
 a99137a <=( A299  and  A298 );
 a99140a <=( (not A302)  and  A301 );
 a99141a <=( a99140a  and  a99137a );
 a99142a <=( a99141a  and  a99134a );
 a99146a <=( (not A167)  and  A168 );
 a99147a <=( A169  and  a99146a );
 a99150a <=( (not A199)  and  A166 );
 a99153a <=( A203  and  (not A200) );
 a99154a <=( a99153a  and  a99150a );
 a99155a <=( a99154a  and  a99147a );
 a99159a <=( (not A268)  and  (not A266) );
 a99160a <=( (not A265)  and  a99159a );
 a99163a <=( (not A299)  and  A298 );
 a99166a <=( A302  and  (not A301) );
 a99167a <=( a99166a  and  a99163a );
 a99168a <=( a99167a  and  a99160a );
 a99172a <=( (not A167)  and  A168 );
 a99173a <=( A169  and  a99172a );
 a99176a <=( (not A199)  and  A166 );
 a99179a <=( A203  and  (not A200) );
 a99180a <=( a99179a  and  a99176a );
 a99181a <=( a99180a  and  a99173a );
 a99185a <=( (not A268)  and  (not A266) );
 a99186a <=( (not A265)  and  a99185a );
 a99189a <=( A299  and  (not A298) );
 a99192a <=( A302  and  (not A301) );
 a99193a <=( a99192a  and  a99189a );
 a99194a <=( a99193a  and  a99186a );
 a99198a <=( (not A167)  and  A168 );
 a99199a <=( A169  and  a99198a );
 a99202a <=( (not A199)  and  A166 );
 a99205a <=( A203  and  (not A200) );
 a99206a <=( a99205a  and  a99202a );
 a99207a <=( a99206a  and  a99199a );
 a99211a <=( (not A268)  and  (not A266) );
 a99212a <=( (not A265)  and  a99211a );
 a99215a <=( (not A299)  and  (not A298) );
 a99218a <=( (not A302)  and  A301 );
 a99219a <=( a99218a  and  a99215a );
 a99220a <=( a99219a  and  a99212a );
 a99224a <=( (not A167)  and  A168 );
 a99225a <=( A169  and  a99224a );
 a99228a <=( (not A199)  and  A166 );
 a99231a <=( A203  and  (not A200) );
 a99232a <=( a99231a  and  a99228a );
 a99233a <=( a99232a  and  a99225a );
 a99237a <=( A269  and  (not A266) );
 a99238a <=( (not A265)  and  a99237a );
 a99241a <=( A299  and  A298 );
 a99244a <=( (not A302)  and  A301 );
 a99245a <=( a99244a  and  a99241a );
 a99246a <=( a99245a  and  a99238a );
 a99250a <=( (not A167)  and  A168 );
 a99251a <=( A169  and  a99250a );
 a99254a <=( (not A199)  and  A166 );
 a99257a <=( A203  and  (not A200) );
 a99258a <=( a99257a  and  a99254a );
 a99259a <=( a99258a  and  a99251a );
 a99263a <=( A269  and  (not A266) );
 a99264a <=( (not A265)  and  a99263a );
 a99267a <=( (not A299)  and  A298 );
 a99270a <=( A302  and  (not A301) );
 a99271a <=( a99270a  and  a99267a );
 a99272a <=( a99271a  and  a99264a );
 a99276a <=( (not A167)  and  A168 );
 a99277a <=( A169  and  a99276a );
 a99280a <=( (not A199)  and  A166 );
 a99283a <=( A203  and  (not A200) );
 a99284a <=( a99283a  and  a99280a );
 a99285a <=( a99284a  and  a99277a );
 a99289a <=( A269  and  (not A266) );
 a99290a <=( (not A265)  and  a99289a );
 a99293a <=( A299  and  (not A298) );
 a99296a <=( A302  and  (not A301) );
 a99297a <=( a99296a  and  a99293a );
 a99298a <=( a99297a  and  a99290a );
 a99302a <=( (not A167)  and  A168 );
 a99303a <=( A169  and  a99302a );
 a99306a <=( (not A199)  and  A166 );
 a99309a <=( A203  and  (not A200) );
 a99310a <=( a99309a  and  a99306a );
 a99311a <=( a99310a  and  a99303a );
 a99315a <=( A269  and  (not A266) );
 a99316a <=( (not A265)  and  a99315a );
 a99319a <=( (not A299)  and  (not A298) );
 a99322a <=( (not A302)  and  A301 );
 a99323a <=( a99322a  and  a99319a );
 a99324a <=( a99323a  and  a99316a );
 a99328a <=( (not A167)  and  A168 );
 a99329a <=( A169  and  a99328a );
 a99332a <=( (not A199)  and  A166 );
 a99335a <=( A202  and  (not A200) );
 a99336a <=( a99335a  and  a99332a );
 a99337a <=( a99336a  and  a99329a );
 a99341a <=( A267  and  A265 );
 a99342a <=( (not A203)  and  a99341a );
 a99345a <=( A299  and  A298 );
 a99348a <=( (not A301)  and  (not A300) );
 a99349a <=( a99348a  and  a99345a );
 a99350a <=( a99349a  and  a99342a );
 a99354a <=( (not A167)  and  A168 );
 a99355a <=( A169  and  a99354a );
 a99358a <=( (not A199)  and  A166 );
 a99361a <=( A202  and  (not A200) );
 a99362a <=( a99361a  and  a99358a );
 a99363a <=( a99362a  and  a99355a );
 a99367a <=( A267  and  A265 );
 a99368a <=( (not A203)  and  a99367a );
 a99371a <=( A299  and  A298 );
 a99374a <=( A302  and  (not A300) );
 a99375a <=( a99374a  and  a99371a );
 a99376a <=( a99375a  and  a99368a );
 a99380a <=( (not A167)  and  A168 );
 a99381a <=( A169  and  a99380a );
 a99384a <=( (not A199)  and  A166 );
 a99387a <=( A202  and  (not A200) );
 a99388a <=( a99387a  and  a99384a );
 a99389a <=( a99388a  and  a99381a );
 a99393a <=( A267  and  A265 );
 a99394a <=( (not A203)  and  a99393a );
 a99397a <=( (not A299)  and  A298 );
 a99400a <=( A301  and  (not A300) );
 a99401a <=( a99400a  and  a99397a );
 a99402a <=( a99401a  and  a99394a );
 a99406a <=( (not A167)  and  A168 );
 a99407a <=( A169  and  a99406a );
 a99410a <=( (not A199)  and  A166 );
 a99413a <=( A202  and  (not A200) );
 a99414a <=( a99413a  and  a99410a );
 a99415a <=( a99414a  and  a99407a );
 a99419a <=( A267  and  A265 );
 a99420a <=( (not A203)  and  a99419a );
 a99423a <=( (not A299)  and  A298 );
 a99426a <=( (not A302)  and  (not A300) );
 a99427a <=( a99426a  and  a99423a );
 a99428a <=( a99427a  and  a99420a );
 a99432a <=( (not A167)  and  A168 );
 a99433a <=( A169  and  a99432a );
 a99436a <=( (not A199)  and  A166 );
 a99439a <=( A202  and  (not A200) );
 a99440a <=( a99439a  and  a99436a );
 a99441a <=( a99440a  and  a99433a );
 a99445a <=( A267  and  A265 );
 a99446a <=( (not A203)  and  a99445a );
 a99449a <=( A299  and  (not A298) );
 a99452a <=( A301  and  (not A300) );
 a99453a <=( a99452a  and  a99449a );
 a99454a <=( a99453a  and  a99446a );
 a99458a <=( (not A167)  and  A168 );
 a99459a <=( A169  and  a99458a );
 a99462a <=( (not A199)  and  A166 );
 a99465a <=( A202  and  (not A200) );
 a99466a <=( a99465a  and  a99462a );
 a99467a <=( a99466a  and  a99459a );
 a99471a <=( A267  and  A265 );
 a99472a <=( (not A203)  and  a99471a );
 a99475a <=( A299  and  (not A298) );
 a99478a <=( (not A302)  and  (not A300) );
 a99479a <=( a99478a  and  a99475a );
 a99480a <=( a99479a  and  a99472a );
 a99484a <=( (not A167)  and  A168 );
 a99485a <=( A169  and  a99484a );
 a99488a <=( (not A199)  and  A166 );
 a99491a <=( A202  and  (not A200) );
 a99492a <=( a99491a  and  a99488a );
 a99493a <=( a99492a  and  a99485a );
 a99497a <=( A267  and  A266 );
 a99498a <=( (not A203)  and  a99497a );
 a99501a <=( A299  and  A298 );
 a99504a <=( (not A301)  and  (not A300) );
 a99505a <=( a99504a  and  a99501a );
 a99506a <=( a99505a  and  a99498a );
 a99510a <=( (not A167)  and  A168 );
 a99511a <=( A169  and  a99510a );
 a99514a <=( (not A199)  and  A166 );
 a99517a <=( A202  and  (not A200) );
 a99518a <=( a99517a  and  a99514a );
 a99519a <=( a99518a  and  a99511a );
 a99523a <=( A267  and  A266 );
 a99524a <=( (not A203)  and  a99523a );
 a99527a <=( A299  and  A298 );
 a99530a <=( A302  and  (not A300) );
 a99531a <=( a99530a  and  a99527a );
 a99532a <=( a99531a  and  a99524a );
 a99536a <=( (not A167)  and  A168 );
 a99537a <=( A169  and  a99536a );
 a99540a <=( (not A199)  and  A166 );
 a99543a <=( A202  and  (not A200) );
 a99544a <=( a99543a  and  a99540a );
 a99545a <=( a99544a  and  a99537a );
 a99549a <=( A267  and  A266 );
 a99550a <=( (not A203)  and  a99549a );
 a99553a <=( (not A299)  and  A298 );
 a99556a <=( A301  and  (not A300) );
 a99557a <=( a99556a  and  a99553a );
 a99558a <=( a99557a  and  a99550a );
 a99562a <=( (not A167)  and  A168 );
 a99563a <=( A169  and  a99562a );
 a99566a <=( (not A199)  and  A166 );
 a99569a <=( A202  and  (not A200) );
 a99570a <=( a99569a  and  a99566a );
 a99571a <=( a99570a  and  a99563a );
 a99575a <=( A267  and  A266 );
 a99576a <=( (not A203)  and  a99575a );
 a99579a <=( (not A299)  and  A298 );
 a99582a <=( (not A302)  and  (not A300) );
 a99583a <=( a99582a  and  a99579a );
 a99584a <=( a99583a  and  a99576a );
 a99588a <=( (not A167)  and  A168 );
 a99589a <=( A169  and  a99588a );
 a99592a <=( (not A199)  and  A166 );
 a99595a <=( A202  and  (not A200) );
 a99596a <=( a99595a  and  a99592a );
 a99597a <=( a99596a  and  a99589a );
 a99601a <=( A267  and  A266 );
 a99602a <=( (not A203)  and  a99601a );
 a99605a <=( A299  and  (not A298) );
 a99608a <=( A301  and  (not A300) );
 a99609a <=( a99608a  and  a99605a );
 a99610a <=( a99609a  and  a99602a );
 a99614a <=( (not A167)  and  A168 );
 a99615a <=( A169  and  a99614a );
 a99618a <=( (not A199)  and  A166 );
 a99621a <=( A202  and  (not A200) );
 a99622a <=( a99621a  and  a99618a );
 a99623a <=( a99622a  and  a99615a );
 a99627a <=( A267  and  A266 );
 a99628a <=( (not A203)  and  a99627a );
 a99631a <=( A299  and  (not A298) );
 a99634a <=( (not A302)  and  (not A300) );
 a99635a <=( a99634a  and  a99631a );
 a99636a <=( a99635a  and  a99628a );
 a99640a <=( (not A167)  and  (not A169) );
 a99641a <=( (not A170)  and  a99640a );
 a99644a <=( A200  and  A199 );
 a99647a <=( (not A203)  and  A202 );
 a99648a <=( a99647a  and  a99644a );
 a99649a <=( a99648a  and  a99641a );
 a99653a <=( (not A268)  and  (not A266) );
 a99654a <=( (not A265)  and  a99653a );
 a99657a <=( A299  and  A298 );
 a99660a <=( (not A302)  and  A301 );
 a99661a <=( a99660a  and  a99657a );
 a99662a <=( a99661a  and  a99654a );
 a99666a <=( (not A167)  and  (not A169) );
 a99667a <=( (not A170)  and  a99666a );
 a99670a <=( A200  and  A199 );
 a99673a <=( (not A203)  and  A202 );
 a99674a <=( a99673a  and  a99670a );
 a99675a <=( a99674a  and  a99667a );
 a99679a <=( (not A268)  and  (not A266) );
 a99680a <=( (not A265)  and  a99679a );
 a99683a <=( (not A299)  and  A298 );
 a99686a <=( A302  and  (not A301) );
 a99687a <=( a99686a  and  a99683a );
 a99688a <=( a99687a  and  a99680a );
 a99692a <=( (not A167)  and  (not A169) );
 a99693a <=( (not A170)  and  a99692a );
 a99696a <=( A200  and  A199 );
 a99699a <=( (not A203)  and  A202 );
 a99700a <=( a99699a  and  a99696a );
 a99701a <=( a99700a  and  a99693a );
 a99705a <=( (not A268)  and  (not A266) );
 a99706a <=( (not A265)  and  a99705a );
 a99709a <=( A299  and  (not A298) );
 a99712a <=( A302  and  (not A301) );
 a99713a <=( a99712a  and  a99709a );
 a99714a <=( a99713a  and  a99706a );
 a99718a <=( (not A167)  and  (not A169) );
 a99719a <=( (not A170)  and  a99718a );
 a99722a <=( A200  and  A199 );
 a99725a <=( (not A203)  and  A202 );
 a99726a <=( a99725a  and  a99722a );
 a99727a <=( a99726a  and  a99719a );
 a99731a <=( (not A268)  and  (not A266) );
 a99732a <=( (not A265)  and  a99731a );
 a99735a <=( (not A299)  and  (not A298) );
 a99738a <=( (not A302)  and  A301 );
 a99739a <=( a99738a  and  a99735a );
 a99740a <=( a99739a  and  a99732a );
 a99744a <=( (not A167)  and  (not A169) );
 a99745a <=( (not A170)  and  a99744a );
 a99748a <=( A200  and  A199 );
 a99751a <=( (not A203)  and  A202 );
 a99752a <=( a99751a  and  a99748a );
 a99753a <=( a99752a  and  a99745a );
 a99757a <=( A269  and  (not A266) );
 a99758a <=( (not A265)  and  a99757a );
 a99761a <=( A299  and  A298 );
 a99764a <=( (not A302)  and  A301 );
 a99765a <=( a99764a  and  a99761a );
 a99766a <=( a99765a  and  a99758a );
 a99770a <=( (not A167)  and  (not A169) );
 a99771a <=( (not A170)  and  a99770a );
 a99774a <=( A200  and  A199 );
 a99777a <=( (not A203)  and  A202 );
 a99778a <=( a99777a  and  a99774a );
 a99779a <=( a99778a  and  a99771a );
 a99783a <=( A269  and  (not A266) );
 a99784a <=( (not A265)  and  a99783a );
 a99787a <=( (not A299)  and  A298 );
 a99790a <=( A302  and  (not A301) );
 a99791a <=( a99790a  and  a99787a );
 a99792a <=( a99791a  and  a99784a );
 a99796a <=( (not A167)  and  (not A169) );
 a99797a <=( (not A170)  and  a99796a );
 a99800a <=( A200  and  A199 );
 a99803a <=( (not A203)  and  A202 );
 a99804a <=( a99803a  and  a99800a );
 a99805a <=( a99804a  and  a99797a );
 a99809a <=( A269  and  (not A266) );
 a99810a <=( (not A265)  and  a99809a );
 a99813a <=( A299  and  (not A298) );
 a99816a <=( A302  and  (not A301) );
 a99817a <=( a99816a  and  a99813a );
 a99818a <=( a99817a  and  a99810a );
 a99822a <=( (not A167)  and  (not A169) );
 a99823a <=( (not A170)  and  a99822a );
 a99826a <=( A200  and  A199 );
 a99829a <=( (not A203)  and  A202 );
 a99830a <=( a99829a  and  a99826a );
 a99831a <=( a99830a  and  a99823a );
 a99835a <=( A269  and  (not A266) );
 a99836a <=( (not A265)  and  a99835a );
 a99839a <=( (not A299)  and  (not A298) );
 a99842a <=( (not A302)  and  A301 );
 a99843a <=( a99842a  and  a99839a );
 a99844a <=( a99843a  and  a99836a );
 a99848a <=( (not A167)  and  (not A169) );
 a99849a <=( (not A170)  and  a99848a );
 a99852a <=( A200  and  A199 );
 a99855a <=( (not A202)  and  (not A201) );
 a99856a <=( a99855a  and  a99852a );
 a99857a <=( a99856a  and  a99849a );
 a99861a <=( A268  and  A266 );
 a99862a <=( A265  and  a99861a );
 a99865a <=( (not A298)  and  (not A269) );
 a99868a <=( (not A301)  and  (not A299) );
 a99869a <=( a99868a  and  a99865a );
 a99870a <=( a99869a  and  a99862a );
 a99874a <=( (not A167)  and  (not A169) );
 a99875a <=( (not A170)  and  a99874a );
 a99878a <=( A200  and  A199 );
 a99881a <=( (not A202)  and  (not A201) );
 a99882a <=( a99881a  and  a99878a );
 a99883a <=( a99882a  and  a99875a );
 a99887a <=( A268  and  A266 );
 a99888a <=( A265  and  a99887a );
 a99891a <=( (not A298)  and  (not A269) );
 a99894a <=( A302  and  (not A299) );
 a99895a <=( a99894a  and  a99891a );
 a99896a <=( a99895a  and  a99888a );
 a99900a <=( (not A167)  and  (not A169) );
 a99901a <=( (not A170)  and  a99900a );
 a99904a <=( A200  and  A199 );
 a99907a <=( (not A202)  and  (not A201) );
 a99908a <=( a99907a  and  a99904a );
 a99909a <=( a99908a  and  a99901a );
 a99913a <=( (not A268)  and  A266 );
 a99914a <=( (not A265)  and  a99913a );
 a99917a <=( (not A298)  and  A269 );
 a99920a <=( (not A301)  and  (not A299) );
 a99921a <=( a99920a  and  a99917a );
 a99922a <=( a99921a  and  a99914a );
 a99926a <=( (not A167)  and  (not A169) );
 a99927a <=( (not A170)  and  a99926a );
 a99930a <=( A200  and  A199 );
 a99933a <=( (not A202)  and  (not A201) );
 a99934a <=( a99933a  and  a99930a );
 a99935a <=( a99934a  and  a99927a );
 a99939a <=( (not A268)  and  A266 );
 a99940a <=( (not A265)  and  a99939a );
 a99943a <=( (not A298)  and  A269 );
 a99946a <=( A302  and  (not A299) );
 a99947a <=( a99946a  and  a99943a );
 a99948a <=( a99947a  and  a99940a );
 a99952a <=( (not A167)  and  (not A169) );
 a99953a <=( (not A170)  and  a99952a );
 a99956a <=( A200  and  A199 );
 a99959a <=( (not A202)  and  (not A201) );
 a99960a <=( a99959a  and  a99956a );
 a99961a <=( a99960a  and  a99953a );
 a99965a <=( (not A268)  and  (not A266) );
 a99966a <=( A265  and  a99965a );
 a99969a <=( (not A298)  and  A269 );
 a99972a <=( (not A301)  and  (not A299) );
 a99973a <=( a99972a  and  a99969a );
 a99974a <=( a99973a  and  a99966a );
 a99978a <=( (not A167)  and  (not A169) );
 a99979a <=( (not A170)  and  a99978a );
 a99982a <=( A200  and  A199 );
 a99985a <=( (not A202)  and  (not A201) );
 a99986a <=( a99985a  and  a99982a );
 a99987a <=( a99986a  and  a99979a );
 a99991a <=( (not A268)  and  (not A266) );
 a99992a <=( A265  and  a99991a );
 a99995a <=( (not A298)  and  A269 );
 a99998a <=( A302  and  (not A299) );
 a99999a <=( a99998a  and  a99995a );
 a100000a <=( a99999a  and  a99992a );
 a100004a <=( (not A167)  and  (not A169) );
 a100005a <=( (not A170)  and  a100004a );
 a100008a <=( A200  and  A199 );
 a100011a <=( (not A202)  and  (not A201) );
 a100012a <=( a100011a  and  a100008a );
 a100013a <=( a100012a  and  a100005a );
 a100017a <=( A268  and  (not A266) );
 a100018a <=( (not A265)  and  a100017a );
 a100021a <=( (not A298)  and  (not A269) );
 a100024a <=( (not A301)  and  (not A299) );
 a100025a <=( a100024a  and  a100021a );
 a100026a <=( a100025a  and  a100018a );
 a100030a <=( (not A167)  and  (not A169) );
 a100031a <=( (not A170)  and  a100030a );
 a100034a <=( A200  and  A199 );
 a100037a <=( (not A202)  and  (not A201) );
 a100038a <=( a100037a  and  a100034a );
 a100039a <=( a100038a  and  a100031a );
 a100043a <=( A268  and  (not A266) );
 a100044a <=( (not A265)  and  a100043a );
 a100047a <=( (not A298)  and  (not A269) );
 a100050a <=( A302  and  (not A299) );
 a100051a <=( a100050a  and  a100047a );
 a100052a <=( a100051a  and  a100044a );
 a100056a <=( (not A167)  and  (not A169) );
 a100057a <=( (not A170)  and  a100056a );
 a100060a <=( A200  and  A199 );
 a100063a <=( A203  and  (not A201) );
 a100064a <=( a100063a  and  a100060a );
 a100065a <=( a100064a  and  a100057a );
 a100069a <=( A268  and  A266 );
 a100070a <=( A265  and  a100069a );
 a100073a <=( (not A298)  and  (not A269) );
 a100076a <=( (not A301)  and  (not A299) );
 a100077a <=( a100076a  and  a100073a );
 a100078a <=( a100077a  and  a100070a );
 a100082a <=( (not A167)  and  (not A169) );
 a100083a <=( (not A170)  and  a100082a );
 a100086a <=( A200  and  A199 );
 a100089a <=( A203  and  (not A201) );
 a100090a <=( a100089a  and  a100086a );
 a100091a <=( a100090a  and  a100083a );
 a100095a <=( A268  and  A266 );
 a100096a <=( A265  and  a100095a );
 a100099a <=( (not A298)  and  (not A269) );
 a100102a <=( A302  and  (not A299) );
 a100103a <=( a100102a  and  a100099a );
 a100104a <=( a100103a  and  a100096a );
 a100108a <=( (not A167)  and  (not A169) );
 a100109a <=( (not A170)  and  a100108a );
 a100112a <=( A200  and  A199 );
 a100115a <=( A203  and  (not A201) );
 a100116a <=( a100115a  and  a100112a );
 a100117a <=( a100116a  and  a100109a );
 a100121a <=( (not A268)  and  A266 );
 a100122a <=( (not A265)  and  a100121a );
 a100125a <=( (not A298)  and  A269 );
 a100128a <=( (not A301)  and  (not A299) );
 a100129a <=( a100128a  and  a100125a );
 a100130a <=( a100129a  and  a100122a );
 a100134a <=( (not A167)  and  (not A169) );
 a100135a <=( (not A170)  and  a100134a );
 a100138a <=( A200  and  A199 );
 a100141a <=( A203  and  (not A201) );
 a100142a <=( a100141a  and  a100138a );
 a100143a <=( a100142a  and  a100135a );
 a100147a <=( (not A268)  and  A266 );
 a100148a <=( (not A265)  and  a100147a );
 a100151a <=( (not A298)  and  A269 );
 a100154a <=( A302  and  (not A299) );
 a100155a <=( a100154a  and  a100151a );
 a100156a <=( a100155a  and  a100148a );
 a100160a <=( (not A167)  and  (not A169) );
 a100161a <=( (not A170)  and  a100160a );
 a100164a <=( A200  and  A199 );
 a100167a <=( A203  and  (not A201) );
 a100168a <=( a100167a  and  a100164a );
 a100169a <=( a100168a  and  a100161a );
 a100173a <=( (not A268)  and  (not A266) );
 a100174a <=( A265  and  a100173a );
 a100177a <=( (not A298)  and  A269 );
 a100180a <=( (not A301)  and  (not A299) );
 a100181a <=( a100180a  and  a100177a );
 a100182a <=( a100181a  and  a100174a );
 a100186a <=( (not A167)  and  (not A169) );
 a100187a <=( (not A170)  and  a100186a );
 a100190a <=( A200  and  A199 );
 a100193a <=( A203  and  (not A201) );
 a100194a <=( a100193a  and  a100190a );
 a100195a <=( a100194a  and  a100187a );
 a100199a <=( (not A268)  and  (not A266) );
 a100200a <=( A265  and  a100199a );
 a100203a <=( (not A298)  and  A269 );
 a100206a <=( A302  and  (not A299) );
 a100207a <=( a100206a  and  a100203a );
 a100208a <=( a100207a  and  a100200a );
 a100212a <=( (not A167)  and  (not A169) );
 a100213a <=( (not A170)  and  a100212a );
 a100216a <=( A200  and  A199 );
 a100219a <=( A203  and  (not A201) );
 a100220a <=( a100219a  and  a100216a );
 a100221a <=( a100220a  and  a100213a );
 a100225a <=( A268  and  (not A266) );
 a100226a <=( (not A265)  and  a100225a );
 a100229a <=( (not A298)  and  (not A269) );
 a100232a <=( (not A301)  and  (not A299) );
 a100233a <=( a100232a  and  a100229a );
 a100234a <=( a100233a  and  a100226a );
 a100238a <=( (not A167)  and  (not A169) );
 a100239a <=( (not A170)  and  a100238a );
 a100242a <=( A200  and  A199 );
 a100245a <=( A203  and  (not A201) );
 a100246a <=( a100245a  and  a100242a );
 a100247a <=( a100246a  and  a100239a );
 a100251a <=( A268  and  (not A266) );
 a100252a <=( (not A265)  and  a100251a );
 a100255a <=( (not A298)  and  (not A269) );
 a100258a <=( A302  and  (not A299) );
 a100259a <=( a100258a  and  a100255a );
 a100260a <=( a100259a  and  a100252a );
 a100264a <=( (not A167)  and  (not A169) );
 a100265a <=( (not A170)  and  a100264a );
 a100268a <=( A200  and  (not A199) );
 a100271a <=( A203  and  (not A202) );
 a100272a <=( a100271a  and  a100268a );
 a100273a <=( a100272a  and  a100265a );
 a100277a <=( (not A268)  and  (not A266) );
 a100278a <=( (not A265)  and  a100277a );
 a100281a <=( A299  and  A298 );
 a100284a <=( (not A302)  and  A301 );
 a100285a <=( a100284a  and  a100281a );
 a100286a <=( a100285a  and  a100278a );
 a100290a <=( (not A167)  and  (not A169) );
 a100291a <=( (not A170)  and  a100290a );
 a100294a <=( A200  and  (not A199) );
 a100297a <=( A203  and  (not A202) );
 a100298a <=( a100297a  and  a100294a );
 a100299a <=( a100298a  and  a100291a );
 a100303a <=( (not A268)  and  (not A266) );
 a100304a <=( (not A265)  and  a100303a );
 a100307a <=( (not A299)  and  A298 );
 a100310a <=( A302  and  (not A301) );
 a100311a <=( a100310a  and  a100307a );
 a100312a <=( a100311a  and  a100304a );
 a100316a <=( (not A167)  and  (not A169) );
 a100317a <=( (not A170)  and  a100316a );
 a100320a <=( A200  and  (not A199) );
 a100323a <=( A203  and  (not A202) );
 a100324a <=( a100323a  and  a100320a );
 a100325a <=( a100324a  and  a100317a );
 a100329a <=( (not A268)  and  (not A266) );
 a100330a <=( (not A265)  and  a100329a );
 a100333a <=( A299  and  (not A298) );
 a100336a <=( A302  and  (not A301) );
 a100337a <=( a100336a  and  a100333a );
 a100338a <=( a100337a  and  a100330a );
 a100342a <=( (not A167)  and  (not A169) );
 a100343a <=( (not A170)  and  a100342a );
 a100346a <=( A200  and  (not A199) );
 a100349a <=( A203  and  (not A202) );
 a100350a <=( a100349a  and  a100346a );
 a100351a <=( a100350a  and  a100343a );
 a100355a <=( (not A268)  and  (not A266) );
 a100356a <=( (not A265)  and  a100355a );
 a100359a <=( (not A299)  and  (not A298) );
 a100362a <=( (not A302)  and  A301 );
 a100363a <=( a100362a  and  a100359a );
 a100364a <=( a100363a  and  a100356a );
 a100368a <=( (not A167)  and  (not A169) );
 a100369a <=( (not A170)  and  a100368a );
 a100372a <=( A200  and  (not A199) );
 a100375a <=( A203  and  (not A202) );
 a100376a <=( a100375a  and  a100372a );
 a100377a <=( a100376a  and  a100369a );
 a100381a <=( A269  and  (not A266) );
 a100382a <=( (not A265)  and  a100381a );
 a100385a <=( A299  and  A298 );
 a100388a <=( (not A302)  and  A301 );
 a100389a <=( a100388a  and  a100385a );
 a100390a <=( a100389a  and  a100382a );
 a100394a <=( (not A167)  and  (not A169) );
 a100395a <=( (not A170)  and  a100394a );
 a100398a <=( A200  and  (not A199) );
 a100401a <=( A203  and  (not A202) );
 a100402a <=( a100401a  and  a100398a );
 a100403a <=( a100402a  and  a100395a );
 a100407a <=( A269  and  (not A266) );
 a100408a <=( (not A265)  and  a100407a );
 a100411a <=( (not A299)  and  A298 );
 a100414a <=( A302  and  (not A301) );
 a100415a <=( a100414a  and  a100411a );
 a100416a <=( a100415a  and  a100408a );
 a100420a <=( (not A167)  and  (not A169) );
 a100421a <=( (not A170)  and  a100420a );
 a100424a <=( A200  and  (not A199) );
 a100427a <=( A203  and  (not A202) );
 a100428a <=( a100427a  and  a100424a );
 a100429a <=( a100428a  and  a100421a );
 a100433a <=( A269  and  (not A266) );
 a100434a <=( (not A265)  and  a100433a );
 a100437a <=( A299  and  (not A298) );
 a100440a <=( A302  and  (not A301) );
 a100441a <=( a100440a  and  a100437a );
 a100442a <=( a100441a  and  a100434a );
 a100446a <=( (not A167)  and  (not A169) );
 a100447a <=( (not A170)  and  a100446a );
 a100450a <=( A200  and  (not A199) );
 a100453a <=( A203  and  (not A202) );
 a100454a <=( a100453a  and  a100450a );
 a100455a <=( a100454a  and  a100447a );
 a100459a <=( A269  and  (not A266) );
 a100460a <=( (not A265)  and  a100459a );
 a100463a <=( (not A299)  and  (not A298) );
 a100466a <=( (not A302)  and  A301 );
 a100467a <=( a100466a  and  a100463a );
 a100468a <=( a100467a  and  a100460a );
 a100472a <=( (not A167)  and  (not A169) );
 a100473a <=( (not A170)  and  a100472a );
 a100476a <=( A200  and  (not A199) );
 a100479a <=( A202  and  (not A201) );
 a100480a <=( a100479a  and  a100476a );
 a100481a <=( a100480a  and  a100473a );
 a100485a <=( A268  and  A266 );
 a100486a <=( A265  and  a100485a );
 a100489a <=( (not A298)  and  (not A269) );
 a100492a <=( (not A301)  and  (not A299) );
 a100493a <=( a100492a  and  a100489a );
 a100494a <=( a100493a  and  a100486a );
 a100498a <=( (not A167)  and  (not A169) );
 a100499a <=( (not A170)  and  a100498a );
 a100502a <=( A200  and  (not A199) );
 a100505a <=( A202  and  (not A201) );
 a100506a <=( a100505a  and  a100502a );
 a100507a <=( a100506a  and  a100499a );
 a100511a <=( A268  and  A266 );
 a100512a <=( A265  and  a100511a );
 a100515a <=( (not A298)  and  (not A269) );
 a100518a <=( A302  and  (not A299) );
 a100519a <=( a100518a  and  a100515a );
 a100520a <=( a100519a  and  a100512a );
 a100524a <=( (not A167)  and  (not A169) );
 a100525a <=( (not A170)  and  a100524a );
 a100528a <=( A200  and  (not A199) );
 a100531a <=( A202  and  (not A201) );
 a100532a <=( a100531a  and  a100528a );
 a100533a <=( a100532a  and  a100525a );
 a100537a <=( (not A268)  and  A266 );
 a100538a <=( (not A265)  and  a100537a );
 a100541a <=( (not A298)  and  A269 );
 a100544a <=( (not A301)  and  (not A299) );
 a100545a <=( a100544a  and  a100541a );
 a100546a <=( a100545a  and  a100538a );
 a100550a <=( (not A167)  and  (not A169) );
 a100551a <=( (not A170)  and  a100550a );
 a100554a <=( A200  and  (not A199) );
 a100557a <=( A202  and  (not A201) );
 a100558a <=( a100557a  and  a100554a );
 a100559a <=( a100558a  and  a100551a );
 a100563a <=( (not A268)  and  A266 );
 a100564a <=( (not A265)  and  a100563a );
 a100567a <=( (not A298)  and  A269 );
 a100570a <=( A302  and  (not A299) );
 a100571a <=( a100570a  and  a100567a );
 a100572a <=( a100571a  and  a100564a );
 a100576a <=( (not A167)  and  (not A169) );
 a100577a <=( (not A170)  and  a100576a );
 a100580a <=( A200  and  (not A199) );
 a100583a <=( A202  and  (not A201) );
 a100584a <=( a100583a  and  a100580a );
 a100585a <=( a100584a  and  a100577a );
 a100589a <=( (not A268)  and  (not A266) );
 a100590a <=( A265  and  a100589a );
 a100593a <=( (not A298)  and  A269 );
 a100596a <=( (not A301)  and  (not A299) );
 a100597a <=( a100596a  and  a100593a );
 a100598a <=( a100597a  and  a100590a );
 a100602a <=( (not A167)  and  (not A169) );
 a100603a <=( (not A170)  and  a100602a );
 a100606a <=( A200  and  (not A199) );
 a100609a <=( A202  and  (not A201) );
 a100610a <=( a100609a  and  a100606a );
 a100611a <=( a100610a  and  a100603a );
 a100615a <=( (not A268)  and  (not A266) );
 a100616a <=( A265  and  a100615a );
 a100619a <=( (not A298)  and  A269 );
 a100622a <=( A302  and  (not A299) );
 a100623a <=( a100622a  and  a100619a );
 a100624a <=( a100623a  and  a100616a );
 a100628a <=( (not A167)  and  (not A169) );
 a100629a <=( (not A170)  and  a100628a );
 a100632a <=( A200  and  (not A199) );
 a100635a <=( A202  and  (not A201) );
 a100636a <=( a100635a  and  a100632a );
 a100637a <=( a100636a  and  a100629a );
 a100641a <=( A268  and  (not A266) );
 a100642a <=( (not A265)  and  a100641a );
 a100645a <=( (not A298)  and  (not A269) );
 a100648a <=( (not A301)  and  (not A299) );
 a100649a <=( a100648a  and  a100645a );
 a100650a <=( a100649a  and  a100642a );
 a100654a <=( (not A167)  and  (not A169) );
 a100655a <=( (not A170)  and  a100654a );
 a100658a <=( A200  and  (not A199) );
 a100661a <=( A202  and  (not A201) );
 a100662a <=( a100661a  and  a100658a );
 a100663a <=( a100662a  and  a100655a );
 a100667a <=( A268  and  (not A266) );
 a100668a <=( (not A265)  and  a100667a );
 a100671a <=( (not A298)  and  (not A269) );
 a100674a <=( A302  and  (not A299) );
 a100675a <=( a100674a  and  a100671a );
 a100676a <=( a100675a  and  a100668a );
 a100680a <=( (not A167)  and  (not A169) );
 a100681a <=( (not A170)  and  a100680a );
 a100684a <=( A200  and  (not A199) );
 a100687a <=( (not A203)  and  (not A201) );
 a100688a <=( a100687a  and  a100684a );
 a100689a <=( a100688a  and  a100681a );
 a100693a <=( A268  and  A266 );
 a100694a <=( A265  and  a100693a );
 a100697a <=( (not A298)  and  (not A269) );
 a100700a <=( (not A301)  and  (not A299) );
 a100701a <=( a100700a  and  a100697a );
 a100702a <=( a100701a  and  a100694a );
 a100706a <=( (not A167)  and  (not A169) );
 a100707a <=( (not A170)  and  a100706a );
 a100710a <=( A200  and  (not A199) );
 a100713a <=( (not A203)  and  (not A201) );
 a100714a <=( a100713a  and  a100710a );
 a100715a <=( a100714a  and  a100707a );
 a100719a <=( A268  and  A266 );
 a100720a <=( A265  and  a100719a );
 a100723a <=( (not A298)  and  (not A269) );
 a100726a <=( A302  and  (not A299) );
 a100727a <=( a100726a  and  a100723a );
 a100728a <=( a100727a  and  a100720a );
 a100732a <=( (not A167)  and  (not A169) );
 a100733a <=( (not A170)  and  a100732a );
 a100736a <=( A200  and  (not A199) );
 a100739a <=( (not A203)  and  (not A201) );
 a100740a <=( a100739a  and  a100736a );
 a100741a <=( a100740a  and  a100733a );
 a100745a <=( (not A268)  and  A266 );
 a100746a <=( (not A265)  and  a100745a );
 a100749a <=( (not A298)  and  A269 );
 a100752a <=( (not A301)  and  (not A299) );
 a100753a <=( a100752a  and  a100749a );
 a100754a <=( a100753a  and  a100746a );
 a100758a <=( (not A167)  and  (not A169) );
 a100759a <=( (not A170)  and  a100758a );
 a100762a <=( A200  and  (not A199) );
 a100765a <=( (not A203)  and  (not A201) );
 a100766a <=( a100765a  and  a100762a );
 a100767a <=( a100766a  and  a100759a );
 a100771a <=( (not A268)  and  A266 );
 a100772a <=( (not A265)  and  a100771a );
 a100775a <=( (not A298)  and  A269 );
 a100778a <=( A302  and  (not A299) );
 a100779a <=( a100778a  and  a100775a );
 a100780a <=( a100779a  and  a100772a );
 a100784a <=( (not A167)  and  (not A169) );
 a100785a <=( (not A170)  and  a100784a );
 a100788a <=( A200  and  (not A199) );
 a100791a <=( (not A203)  and  (not A201) );
 a100792a <=( a100791a  and  a100788a );
 a100793a <=( a100792a  and  a100785a );
 a100797a <=( (not A268)  and  (not A266) );
 a100798a <=( A265  and  a100797a );
 a100801a <=( (not A298)  and  A269 );
 a100804a <=( (not A301)  and  (not A299) );
 a100805a <=( a100804a  and  a100801a );
 a100806a <=( a100805a  and  a100798a );
 a100810a <=( (not A167)  and  (not A169) );
 a100811a <=( (not A170)  and  a100810a );
 a100814a <=( A200  and  (not A199) );
 a100817a <=( (not A203)  and  (not A201) );
 a100818a <=( a100817a  and  a100814a );
 a100819a <=( a100818a  and  a100811a );
 a100823a <=( (not A268)  and  (not A266) );
 a100824a <=( A265  and  a100823a );
 a100827a <=( (not A298)  and  A269 );
 a100830a <=( A302  and  (not A299) );
 a100831a <=( a100830a  and  a100827a );
 a100832a <=( a100831a  and  a100824a );
 a100836a <=( (not A167)  and  (not A169) );
 a100837a <=( (not A170)  and  a100836a );
 a100840a <=( A200  and  (not A199) );
 a100843a <=( (not A203)  and  (not A201) );
 a100844a <=( a100843a  and  a100840a );
 a100845a <=( a100844a  and  a100837a );
 a100849a <=( A268  and  (not A266) );
 a100850a <=( (not A265)  and  a100849a );
 a100853a <=( (not A298)  and  (not A269) );
 a100856a <=( (not A301)  and  (not A299) );
 a100857a <=( a100856a  and  a100853a );
 a100858a <=( a100857a  and  a100850a );
 a100862a <=( (not A167)  and  (not A169) );
 a100863a <=( (not A170)  and  a100862a );
 a100866a <=( A200  and  (not A199) );
 a100869a <=( (not A203)  and  (not A201) );
 a100870a <=( a100869a  and  a100866a );
 a100871a <=( a100870a  and  a100863a );
 a100875a <=( A268  and  (not A266) );
 a100876a <=( (not A265)  and  a100875a );
 a100879a <=( (not A298)  and  (not A269) );
 a100882a <=( A302  and  (not A299) );
 a100883a <=( a100882a  and  a100879a );
 a100884a <=( a100883a  and  a100876a );
 a100888a <=( (not A167)  and  (not A169) );
 a100889a <=( (not A170)  and  a100888a );
 a100892a <=( (not A200)  and  A199 );
 a100895a <=( A203  and  (not A202) );
 a100896a <=( a100895a  and  a100892a );
 a100897a <=( a100896a  and  a100889a );
 a100901a <=( (not A268)  and  (not A266) );
 a100902a <=( (not A265)  and  a100901a );
 a100905a <=( A299  and  A298 );
 a100908a <=( (not A302)  and  A301 );
 a100909a <=( a100908a  and  a100905a );
 a100910a <=( a100909a  and  a100902a );
 a100914a <=( (not A167)  and  (not A169) );
 a100915a <=( (not A170)  and  a100914a );
 a100918a <=( (not A200)  and  A199 );
 a100921a <=( A203  and  (not A202) );
 a100922a <=( a100921a  and  a100918a );
 a100923a <=( a100922a  and  a100915a );
 a100927a <=( (not A268)  and  (not A266) );
 a100928a <=( (not A265)  and  a100927a );
 a100931a <=( (not A299)  and  A298 );
 a100934a <=( A302  and  (not A301) );
 a100935a <=( a100934a  and  a100931a );
 a100936a <=( a100935a  and  a100928a );
 a100940a <=( (not A167)  and  (not A169) );
 a100941a <=( (not A170)  and  a100940a );
 a100944a <=( (not A200)  and  A199 );
 a100947a <=( A203  and  (not A202) );
 a100948a <=( a100947a  and  a100944a );
 a100949a <=( a100948a  and  a100941a );
 a100953a <=( (not A268)  and  (not A266) );
 a100954a <=( (not A265)  and  a100953a );
 a100957a <=( A299  and  (not A298) );
 a100960a <=( A302  and  (not A301) );
 a100961a <=( a100960a  and  a100957a );
 a100962a <=( a100961a  and  a100954a );
 a100966a <=( (not A167)  and  (not A169) );
 a100967a <=( (not A170)  and  a100966a );
 a100970a <=( (not A200)  and  A199 );
 a100973a <=( A203  and  (not A202) );
 a100974a <=( a100973a  and  a100970a );
 a100975a <=( a100974a  and  a100967a );
 a100979a <=( (not A268)  and  (not A266) );
 a100980a <=( (not A265)  and  a100979a );
 a100983a <=( (not A299)  and  (not A298) );
 a100986a <=( (not A302)  and  A301 );
 a100987a <=( a100986a  and  a100983a );
 a100988a <=( a100987a  and  a100980a );
 a100992a <=( (not A167)  and  (not A169) );
 a100993a <=( (not A170)  and  a100992a );
 a100996a <=( (not A200)  and  A199 );
 a100999a <=( A203  and  (not A202) );
 a101000a <=( a100999a  and  a100996a );
 a101001a <=( a101000a  and  a100993a );
 a101005a <=( A269  and  (not A266) );
 a101006a <=( (not A265)  and  a101005a );
 a101009a <=( A299  and  A298 );
 a101012a <=( (not A302)  and  A301 );
 a101013a <=( a101012a  and  a101009a );
 a101014a <=( a101013a  and  a101006a );
 a101018a <=( (not A167)  and  (not A169) );
 a101019a <=( (not A170)  and  a101018a );
 a101022a <=( (not A200)  and  A199 );
 a101025a <=( A203  and  (not A202) );
 a101026a <=( a101025a  and  a101022a );
 a101027a <=( a101026a  and  a101019a );
 a101031a <=( A269  and  (not A266) );
 a101032a <=( (not A265)  and  a101031a );
 a101035a <=( (not A299)  and  A298 );
 a101038a <=( A302  and  (not A301) );
 a101039a <=( a101038a  and  a101035a );
 a101040a <=( a101039a  and  a101032a );
 a101044a <=( (not A167)  and  (not A169) );
 a101045a <=( (not A170)  and  a101044a );
 a101048a <=( (not A200)  and  A199 );
 a101051a <=( A203  and  (not A202) );
 a101052a <=( a101051a  and  a101048a );
 a101053a <=( a101052a  and  a101045a );
 a101057a <=( A269  and  (not A266) );
 a101058a <=( (not A265)  and  a101057a );
 a101061a <=( A299  and  (not A298) );
 a101064a <=( A302  and  (not A301) );
 a101065a <=( a101064a  and  a101061a );
 a101066a <=( a101065a  and  a101058a );
 a101070a <=( (not A167)  and  (not A169) );
 a101071a <=( (not A170)  and  a101070a );
 a101074a <=( (not A200)  and  A199 );
 a101077a <=( A203  and  (not A202) );
 a101078a <=( a101077a  and  a101074a );
 a101079a <=( a101078a  and  a101071a );
 a101083a <=( A269  and  (not A266) );
 a101084a <=( (not A265)  and  a101083a );
 a101087a <=( (not A299)  and  (not A298) );
 a101090a <=( (not A302)  and  A301 );
 a101091a <=( a101090a  and  a101087a );
 a101092a <=( a101091a  and  a101084a );
 a101096a <=( (not A167)  and  (not A169) );
 a101097a <=( (not A170)  and  a101096a );
 a101100a <=( (not A200)  and  A199 );
 a101103a <=( A202  and  (not A201) );
 a101104a <=( a101103a  and  a101100a );
 a101105a <=( a101104a  and  a101097a );
 a101109a <=( A268  and  A266 );
 a101110a <=( A265  and  a101109a );
 a101113a <=( (not A298)  and  (not A269) );
 a101116a <=( (not A301)  and  (not A299) );
 a101117a <=( a101116a  and  a101113a );
 a101118a <=( a101117a  and  a101110a );
 a101122a <=( (not A167)  and  (not A169) );
 a101123a <=( (not A170)  and  a101122a );
 a101126a <=( (not A200)  and  A199 );
 a101129a <=( A202  and  (not A201) );
 a101130a <=( a101129a  and  a101126a );
 a101131a <=( a101130a  and  a101123a );
 a101135a <=( A268  and  A266 );
 a101136a <=( A265  and  a101135a );
 a101139a <=( (not A298)  and  (not A269) );
 a101142a <=( A302  and  (not A299) );
 a101143a <=( a101142a  and  a101139a );
 a101144a <=( a101143a  and  a101136a );
 a101148a <=( (not A167)  and  (not A169) );
 a101149a <=( (not A170)  and  a101148a );
 a101152a <=( (not A200)  and  A199 );
 a101155a <=( A202  and  (not A201) );
 a101156a <=( a101155a  and  a101152a );
 a101157a <=( a101156a  and  a101149a );
 a101161a <=( (not A268)  and  A266 );
 a101162a <=( (not A265)  and  a101161a );
 a101165a <=( (not A298)  and  A269 );
 a101168a <=( (not A301)  and  (not A299) );
 a101169a <=( a101168a  and  a101165a );
 a101170a <=( a101169a  and  a101162a );
 a101174a <=( (not A167)  and  (not A169) );
 a101175a <=( (not A170)  and  a101174a );
 a101178a <=( (not A200)  and  A199 );
 a101181a <=( A202  and  (not A201) );
 a101182a <=( a101181a  and  a101178a );
 a101183a <=( a101182a  and  a101175a );
 a101187a <=( (not A268)  and  A266 );
 a101188a <=( (not A265)  and  a101187a );
 a101191a <=( (not A298)  and  A269 );
 a101194a <=( A302  and  (not A299) );
 a101195a <=( a101194a  and  a101191a );
 a101196a <=( a101195a  and  a101188a );
 a101200a <=( (not A167)  and  (not A169) );
 a101201a <=( (not A170)  and  a101200a );
 a101204a <=( (not A200)  and  A199 );
 a101207a <=( A202  and  (not A201) );
 a101208a <=( a101207a  and  a101204a );
 a101209a <=( a101208a  and  a101201a );
 a101213a <=( (not A268)  and  (not A266) );
 a101214a <=( A265  and  a101213a );
 a101217a <=( (not A298)  and  A269 );
 a101220a <=( (not A301)  and  (not A299) );
 a101221a <=( a101220a  and  a101217a );
 a101222a <=( a101221a  and  a101214a );
 a101226a <=( (not A167)  and  (not A169) );
 a101227a <=( (not A170)  and  a101226a );
 a101230a <=( (not A200)  and  A199 );
 a101233a <=( A202  and  (not A201) );
 a101234a <=( a101233a  and  a101230a );
 a101235a <=( a101234a  and  a101227a );
 a101239a <=( (not A268)  and  (not A266) );
 a101240a <=( A265  and  a101239a );
 a101243a <=( (not A298)  and  A269 );
 a101246a <=( A302  and  (not A299) );
 a101247a <=( a101246a  and  a101243a );
 a101248a <=( a101247a  and  a101240a );
 a101252a <=( (not A167)  and  (not A169) );
 a101253a <=( (not A170)  and  a101252a );
 a101256a <=( (not A200)  and  A199 );
 a101259a <=( A202  and  (not A201) );
 a101260a <=( a101259a  and  a101256a );
 a101261a <=( a101260a  and  a101253a );
 a101265a <=( A268  and  (not A266) );
 a101266a <=( (not A265)  and  a101265a );
 a101269a <=( (not A298)  and  (not A269) );
 a101272a <=( (not A301)  and  (not A299) );
 a101273a <=( a101272a  and  a101269a );
 a101274a <=( a101273a  and  a101266a );
 a101278a <=( (not A167)  and  (not A169) );
 a101279a <=( (not A170)  and  a101278a );
 a101282a <=( (not A200)  and  A199 );
 a101285a <=( A202  and  (not A201) );
 a101286a <=( a101285a  and  a101282a );
 a101287a <=( a101286a  and  a101279a );
 a101291a <=( A268  and  (not A266) );
 a101292a <=( (not A265)  and  a101291a );
 a101295a <=( (not A298)  and  (not A269) );
 a101298a <=( A302  and  (not A299) );
 a101299a <=( a101298a  and  a101295a );
 a101300a <=( a101299a  and  a101292a );
 a101304a <=( (not A167)  and  (not A169) );
 a101305a <=( (not A170)  and  a101304a );
 a101308a <=( (not A200)  and  A199 );
 a101311a <=( (not A203)  and  (not A201) );
 a101312a <=( a101311a  and  a101308a );
 a101313a <=( a101312a  and  a101305a );
 a101317a <=( A268  and  A266 );
 a101318a <=( A265  and  a101317a );
 a101321a <=( (not A298)  and  (not A269) );
 a101324a <=( (not A301)  and  (not A299) );
 a101325a <=( a101324a  and  a101321a );
 a101326a <=( a101325a  and  a101318a );
 a101330a <=( (not A167)  and  (not A169) );
 a101331a <=( (not A170)  and  a101330a );
 a101334a <=( (not A200)  and  A199 );
 a101337a <=( (not A203)  and  (not A201) );
 a101338a <=( a101337a  and  a101334a );
 a101339a <=( a101338a  and  a101331a );
 a101343a <=( A268  and  A266 );
 a101344a <=( A265  and  a101343a );
 a101347a <=( (not A298)  and  (not A269) );
 a101350a <=( A302  and  (not A299) );
 a101351a <=( a101350a  and  a101347a );
 a101352a <=( a101351a  and  a101344a );
 a101356a <=( (not A167)  and  (not A169) );
 a101357a <=( (not A170)  and  a101356a );
 a101360a <=( (not A200)  and  A199 );
 a101363a <=( (not A203)  and  (not A201) );
 a101364a <=( a101363a  and  a101360a );
 a101365a <=( a101364a  and  a101357a );
 a101369a <=( (not A268)  and  A266 );
 a101370a <=( (not A265)  and  a101369a );
 a101373a <=( (not A298)  and  A269 );
 a101376a <=( (not A301)  and  (not A299) );
 a101377a <=( a101376a  and  a101373a );
 a101378a <=( a101377a  and  a101370a );
 a101382a <=( (not A167)  and  (not A169) );
 a101383a <=( (not A170)  and  a101382a );
 a101386a <=( (not A200)  and  A199 );
 a101389a <=( (not A203)  and  (not A201) );
 a101390a <=( a101389a  and  a101386a );
 a101391a <=( a101390a  and  a101383a );
 a101395a <=( (not A268)  and  A266 );
 a101396a <=( (not A265)  and  a101395a );
 a101399a <=( (not A298)  and  A269 );
 a101402a <=( A302  and  (not A299) );
 a101403a <=( a101402a  and  a101399a );
 a101404a <=( a101403a  and  a101396a );
 a101408a <=( (not A167)  and  (not A169) );
 a101409a <=( (not A170)  and  a101408a );
 a101412a <=( (not A200)  and  A199 );
 a101415a <=( (not A203)  and  (not A201) );
 a101416a <=( a101415a  and  a101412a );
 a101417a <=( a101416a  and  a101409a );
 a101421a <=( (not A268)  and  (not A266) );
 a101422a <=( A265  and  a101421a );
 a101425a <=( (not A298)  and  A269 );
 a101428a <=( (not A301)  and  (not A299) );
 a101429a <=( a101428a  and  a101425a );
 a101430a <=( a101429a  and  a101422a );
 a101434a <=( (not A167)  and  (not A169) );
 a101435a <=( (not A170)  and  a101434a );
 a101438a <=( (not A200)  and  A199 );
 a101441a <=( (not A203)  and  (not A201) );
 a101442a <=( a101441a  and  a101438a );
 a101443a <=( a101442a  and  a101435a );
 a101447a <=( (not A268)  and  (not A266) );
 a101448a <=( A265  and  a101447a );
 a101451a <=( (not A298)  and  A269 );
 a101454a <=( A302  and  (not A299) );
 a101455a <=( a101454a  and  a101451a );
 a101456a <=( a101455a  and  a101448a );
 a101460a <=( (not A167)  and  (not A169) );
 a101461a <=( (not A170)  and  a101460a );
 a101464a <=( (not A200)  and  A199 );
 a101467a <=( (not A203)  and  (not A201) );
 a101468a <=( a101467a  and  a101464a );
 a101469a <=( a101468a  and  a101461a );
 a101473a <=( A268  and  (not A266) );
 a101474a <=( (not A265)  and  a101473a );
 a101477a <=( (not A298)  and  (not A269) );
 a101480a <=( (not A301)  and  (not A299) );
 a101481a <=( a101480a  and  a101477a );
 a101482a <=( a101481a  and  a101474a );
 a101486a <=( (not A167)  and  (not A169) );
 a101487a <=( (not A170)  and  a101486a );
 a101490a <=( (not A200)  and  A199 );
 a101493a <=( (not A203)  and  (not A201) );
 a101494a <=( a101493a  and  a101490a );
 a101495a <=( a101494a  and  a101487a );
 a101499a <=( A268  and  (not A266) );
 a101500a <=( (not A265)  and  a101499a );
 a101503a <=( (not A298)  and  (not A269) );
 a101506a <=( A302  and  (not A299) );
 a101507a <=( a101506a  and  a101503a );
 a101508a <=( a101507a  and  a101500a );
 a101512a <=( (not A167)  and  (not A169) );
 a101513a <=( (not A170)  and  a101512a );
 a101516a <=( (not A200)  and  (not A199) );
 a101519a <=( A265  and  (not A202) );
 a101520a <=( a101519a  and  a101516a );
 a101521a <=( a101520a  and  a101513a );
 a101525a <=( (not A269)  and  A268 );
 a101526a <=( A266  and  a101525a );
 a101529a <=( A299  and  A298 );
 a101532a <=( (not A301)  and  (not A300) );
 a101533a <=( a101532a  and  a101529a );
 a101534a <=( a101533a  and  a101526a );
 a101538a <=( (not A167)  and  (not A169) );
 a101539a <=( (not A170)  and  a101538a );
 a101542a <=( (not A200)  and  (not A199) );
 a101545a <=( A265  and  (not A202) );
 a101546a <=( a101545a  and  a101542a );
 a101547a <=( a101546a  and  a101539a );
 a101551a <=( (not A269)  and  A268 );
 a101552a <=( A266  and  a101551a );
 a101555a <=( A299  and  A298 );
 a101558a <=( A302  and  (not A300) );
 a101559a <=( a101558a  and  a101555a );
 a101560a <=( a101559a  and  a101552a );
 a101564a <=( (not A167)  and  (not A169) );
 a101565a <=( (not A170)  and  a101564a );
 a101568a <=( (not A200)  and  (not A199) );
 a101571a <=( A265  and  (not A202) );
 a101572a <=( a101571a  and  a101568a );
 a101573a <=( a101572a  and  a101565a );
 a101577a <=( (not A269)  and  A268 );
 a101578a <=( A266  and  a101577a );
 a101581a <=( (not A299)  and  A298 );
 a101584a <=( A301  and  (not A300) );
 a101585a <=( a101584a  and  a101581a );
 a101586a <=( a101585a  and  a101578a );
 a101590a <=( (not A167)  and  (not A169) );
 a101591a <=( (not A170)  and  a101590a );
 a101594a <=( (not A200)  and  (not A199) );
 a101597a <=( A265  and  (not A202) );
 a101598a <=( a101597a  and  a101594a );
 a101599a <=( a101598a  and  a101591a );
 a101603a <=( (not A269)  and  A268 );
 a101604a <=( A266  and  a101603a );
 a101607a <=( (not A299)  and  A298 );
 a101610a <=( (not A302)  and  (not A300) );
 a101611a <=( a101610a  and  a101607a );
 a101612a <=( a101611a  and  a101604a );
 a101616a <=( (not A167)  and  (not A169) );
 a101617a <=( (not A170)  and  a101616a );
 a101620a <=( (not A200)  and  (not A199) );
 a101623a <=( A265  and  (not A202) );
 a101624a <=( a101623a  and  a101620a );
 a101625a <=( a101624a  and  a101617a );
 a101629a <=( (not A269)  and  A268 );
 a101630a <=( A266  and  a101629a );
 a101633a <=( A299  and  (not A298) );
 a101636a <=( A301  and  (not A300) );
 a101637a <=( a101636a  and  a101633a );
 a101638a <=( a101637a  and  a101630a );
 a101642a <=( (not A167)  and  (not A169) );
 a101643a <=( (not A170)  and  a101642a );
 a101646a <=( (not A200)  and  (not A199) );
 a101649a <=( A265  and  (not A202) );
 a101650a <=( a101649a  and  a101646a );
 a101651a <=( a101650a  and  a101643a );
 a101655a <=( (not A269)  and  A268 );
 a101656a <=( A266  and  a101655a );
 a101659a <=( A299  and  (not A298) );
 a101662a <=( (not A302)  and  (not A300) );
 a101663a <=( a101662a  and  a101659a );
 a101664a <=( a101663a  and  a101656a );
 a101668a <=( (not A167)  and  (not A169) );
 a101669a <=( (not A170)  and  a101668a );
 a101672a <=( (not A200)  and  (not A199) );
 a101675a <=( (not A265)  and  (not A202) );
 a101676a <=( a101675a  and  a101672a );
 a101677a <=( a101676a  and  a101669a );
 a101681a <=( A269  and  (not A268) );
 a101682a <=( A266  and  a101681a );
 a101685a <=( A299  and  A298 );
 a101688a <=( (not A301)  and  (not A300) );
 a101689a <=( a101688a  and  a101685a );
 a101690a <=( a101689a  and  a101682a );
 a101694a <=( (not A167)  and  (not A169) );
 a101695a <=( (not A170)  and  a101694a );
 a101698a <=( (not A200)  and  (not A199) );
 a101701a <=( (not A265)  and  (not A202) );
 a101702a <=( a101701a  and  a101698a );
 a101703a <=( a101702a  and  a101695a );
 a101707a <=( A269  and  (not A268) );
 a101708a <=( A266  and  a101707a );
 a101711a <=( A299  and  A298 );
 a101714a <=( A302  and  (not A300) );
 a101715a <=( a101714a  and  a101711a );
 a101716a <=( a101715a  and  a101708a );
 a101720a <=( (not A167)  and  (not A169) );
 a101721a <=( (not A170)  and  a101720a );
 a101724a <=( (not A200)  and  (not A199) );
 a101727a <=( (not A265)  and  (not A202) );
 a101728a <=( a101727a  and  a101724a );
 a101729a <=( a101728a  and  a101721a );
 a101733a <=( A269  and  (not A268) );
 a101734a <=( A266  and  a101733a );
 a101737a <=( (not A299)  and  A298 );
 a101740a <=( A301  and  (not A300) );
 a101741a <=( a101740a  and  a101737a );
 a101742a <=( a101741a  and  a101734a );
 a101746a <=( (not A167)  and  (not A169) );
 a101747a <=( (not A170)  and  a101746a );
 a101750a <=( (not A200)  and  (not A199) );
 a101753a <=( (not A265)  and  (not A202) );
 a101754a <=( a101753a  and  a101750a );
 a101755a <=( a101754a  and  a101747a );
 a101759a <=( A269  and  (not A268) );
 a101760a <=( A266  and  a101759a );
 a101763a <=( (not A299)  and  A298 );
 a101766a <=( (not A302)  and  (not A300) );
 a101767a <=( a101766a  and  a101763a );
 a101768a <=( a101767a  and  a101760a );
 a101772a <=( (not A167)  and  (not A169) );
 a101773a <=( (not A170)  and  a101772a );
 a101776a <=( (not A200)  and  (not A199) );
 a101779a <=( (not A265)  and  (not A202) );
 a101780a <=( a101779a  and  a101776a );
 a101781a <=( a101780a  and  a101773a );
 a101785a <=( A269  and  (not A268) );
 a101786a <=( A266  and  a101785a );
 a101789a <=( A299  and  (not A298) );
 a101792a <=( A301  and  (not A300) );
 a101793a <=( a101792a  and  a101789a );
 a101794a <=( a101793a  and  a101786a );
 a101798a <=( (not A167)  and  (not A169) );
 a101799a <=( (not A170)  and  a101798a );
 a101802a <=( (not A200)  and  (not A199) );
 a101805a <=( (not A265)  and  (not A202) );
 a101806a <=( a101805a  and  a101802a );
 a101807a <=( a101806a  and  a101799a );
 a101811a <=( A269  and  (not A268) );
 a101812a <=( A266  and  a101811a );
 a101815a <=( A299  and  (not A298) );
 a101818a <=( (not A302)  and  (not A300) );
 a101819a <=( a101818a  and  a101815a );
 a101820a <=( a101819a  and  a101812a );
 a101824a <=( (not A167)  and  (not A169) );
 a101825a <=( (not A170)  and  a101824a );
 a101828a <=( (not A200)  and  (not A199) );
 a101831a <=( A265  and  (not A202) );
 a101832a <=( a101831a  and  a101828a );
 a101833a <=( a101832a  and  a101825a );
 a101837a <=( A269  and  (not A268) );
 a101838a <=( (not A266)  and  a101837a );
 a101841a <=( A299  and  A298 );
 a101844a <=( (not A301)  and  (not A300) );
 a101845a <=( a101844a  and  a101841a );
 a101846a <=( a101845a  and  a101838a );
 a101850a <=( (not A167)  and  (not A169) );
 a101851a <=( (not A170)  and  a101850a );
 a101854a <=( (not A200)  and  (not A199) );
 a101857a <=( A265  and  (not A202) );
 a101858a <=( a101857a  and  a101854a );
 a101859a <=( a101858a  and  a101851a );
 a101863a <=( A269  and  (not A268) );
 a101864a <=( (not A266)  and  a101863a );
 a101867a <=( A299  and  A298 );
 a101870a <=( A302  and  (not A300) );
 a101871a <=( a101870a  and  a101867a );
 a101872a <=( a101871a  and  a101864a );
 a101876a <=( (not A167)  and  (not A169) );
 a101877a <=( (not A170)  and  a101876a );
 a101880a <=( (not A200)  and  (not A199) );
 a101883a <=( A265  and  (not A202) );
 a101884a <=( a101883a  and  a101880a );
 a101885a <=( a101884a  and  a101877a );
 a101889a <=( A269  and  (not A268) );
 a101890a <=( (not A266)  and  a101889a );
 a101893a <=( (not A299)  and  A298 );
 a101896a <=( A301  and  (not A300) );
 a101897a <=( a101896a  and  a101893a );
 a101898a <=( a101897a  and  a101890a );
 a101902a <=( (not A167)  and  (not A169) );
 a101903a <=( (not A170)  and  a101902a );
 a101906a <=( (not A200)  and  (not A199) );
 a101909a <=( A265  and  (not A202) );
 a101910a <=( a101909a  and  a101906a );
 a101911a <=( a101910a  and  a101903a );
 a101915a <=( A269  and  (not A268) );
 a101916a <=( (not A266)  and  a101915a );
 a101919a <=( (not A299)  and  A298 );
 a101922a <=( (not A302)  and  (not A300) );
 a101923a <=( a101922a  and  a101919a );
 a101924a <=( a101923a  and  a101916a );
 a101928a <=( (not A167)  and  (not A169) );
 a101929a <=( (not A170)  and  a101928a );
 a101932a <=( (not A200)  and  (not A199) );
 a101935a <=( A265  and  (not A202) );
 a101936a <=( a101935a  and  a101932a );
 a101937a <=( a101936a  and  a101929a );
 a101941a <=( A269  and  (not A268) );
 a101942a <=( (not A266)  and  a101941a );
 a101945a <=( A299  and  (not A298) );
 a101948a <=( A301  and  (not A300) );
 a101949a <=( a101948a  and  a101945a );
 a101950a <=( a101949a  and  a101942a );
 a101954a <=( (not A167)  and  (not A169) );
 a101955a <=( (not A170)  and  a101954a );
 a101958a <=( (not A200)  and  (not A199) );
 a101961a <=( A265  and  (not A202) );
 a101962a <=( a101961a  and  a101958a );
 a101963a <=( a101962a  and  a101955a );
 a101967a <=( A269  and  (not A268) );
 a101968a <=( (not A266)  and  a101967a );
 a101971a <=( A299  and  (not A298) );
 a101974a <=( (not A302)  and  (not A300) );
 a101975a <=( a101974a  and  a101971a );
 a101976a <=( a101975a  and  a101968a );
 a101980a <=( (not A167)  and  (not A169) );
 a101981a <=( (not A170)  and  a101980a );
 a101984a <=( (not A200)  and  (not A199) );
 a101987a <=( (not A265)  and  (not A202) );
 a101988a <=( a101987a  and  a101984a );
 a101989a <=( a101988a  and  a101981a );
 a101993a <=( (not A269)  and  A268 );
 a101994a <=( (not A266)  and  a101993a );
 a101997a <=( A299  and  A298 );
 a102000a <=( (not A301)  and  (not A300) );
 a102001a <=( a102000a  and  a101997a );
 a102002a <=( a102001a  and  a101994a );
 a102006a <=( (not A167)  and  (not A169) );
 a102007a <=( (not A170)  and  a102006a );
 a102010a <=( (not A200)  and  (not A199) );
 a102013a <=( (not A265)  and  (not A202) );
 a102014a <=( a102013a  and  a102010a );
 a102015a <=( a102014a  and  a102007a );
 a102019a <=( (not A269)  and  A268 );
 a102020a <=( (not A266)  and  a102019a );
 a102023a <=( A299  and  A298 );
 a102026a <=( A302  and  (not A300) );
 a102027a <=( a102026a  and  a102023a );
 a102028a <=( a102027a  and  a102020a );
 a102032a <=( (not A167)  and  (not A169) );
 a102033a <=( (not A170)  and  a102032a );
 a102036a <=( (not A200)  and  (not A199) );
 a102039a <=( (not A265)  and  (not A202) );
 a102040a <=( a102039a  and  a102036a );
 a102041a <=( a102040a  and  a102033a );
 a102045a <=( (not A269)  and  A268 );
 a102046a <=( (not A266)  and  a102045a );
 a102049a <=( (not A299)  and  A298 );
 a102052a <=( A301  and  (not A300) );
 a102053a <=( a102052a  and  a102049a );
 a102054a <=( a102053a  and  a102046a );
 a102058a <=( (not A167)  and  (not A169) );
 a102059a <=( (not A170)  and  a102058a );
 a102062a <=( (not A200)  and  (not A199) );
 a102065a <=( (not A265)  and  (not A202) );
 a102066a <=( a102065a  and  a102062a );
 a102067a <=( a102066a  and  a102059a );
 a102071a <=( (not A269)  and  A268 );
 a102072a <=( (not A266)  and  a102071a );
 a102075a <=( (not A299)  and  A298 );
 a102078a <=( (not A302)  and  (not A300) );
 a102079a <=( a102078a  and  a102075a );
 a102080a <=( a102079a  and  a102072a );
 a102084a <=( (not A167)  and  (not A169) );
 a102085a <=( (not A170)  and  a102084a );
 a102088a <=( (not A200)  and  (not A199) );
 a102091a <=( (not A265)  and  (not A202) );
 a102092a <=( a102091a  and  a102088a );
 a102093a <=( a102092a  and  a102085a );
 a102097a <=( (not A269)  and  A268 );
 a102098a <=( (not A266)  and  a102097a );
 a102101a <=( A299  and  (not A298) );
 a102104a <=( A301  and  (not A300) );
 a102105a <=( a102104a  and  a102101a );
 a102106a <=( a102105a  and  a102098a );
 a102110a <=( (not A167)  and  (not A169) );
 a102111a <=( (not A170)  and  a102110a );
 a102114a <=( (not A200)  and  (not A199) );
 a102117a <=( (not A265)  and  (not A202) );
 a102118a <=( a102117a  and  a102114a );
 a102119a <=( a102118a  and  a102111a );
 a102123a <=( (not A269)  and  A268 );
 a102124a <=( (not A266)  and  a102123a );
 a102127a <=( A299  and  (not A298) );
 a102130a <=( (not A302)  and  (not A300) );
 a102131a <=( a102130a  and  a102127a );
 a102132a <=( a102131a  and  a102124a );
 a102136a <=( (not A167)  and  (not A169) );
 a102137a <=( (not A170)  and  a102136a );
 a102140a <=( (not A200)  and  (not A199) );
 a102143a <=( A265  and  A203 );
 a102144a <=( a102143a  and  a102140a );
 a102145a <=( a102144a  and  a102137a );
 a102149a <=( (not A269)  and  A268 );
 a102150a <=( A266  and  a102149a );
 a102153a <=( A299  and  A298 );
 a102156a <=( (not A301)  and  (not A300) );
 a102157a <=( a102156a  and  a102153a );
 a102158a <=( a102157a  and  a102150a );
 a102162a <=( (not A167)  and  (not A169) );
 a102163a <=( (not A170)  and  a102162a );
 a102166a <=( (not A200)  and  (not A199) );
 a102169a <=( A265  and  A203 );
 a102170a <=( a102169a  and  a102166a );
 a102171a <=( a102170a  and  a102163a );
 a102175a <=( (not A269)  and  A268 );
 a102176a <=( A266  and  a102175a );
 a102179a <=( A299  and  A298 );
 a102182a <=( A302  and  (not A300) );
 a102183a <=( a102182a  and  a102179a );
 a102184a <=( a102183a  and  a102176a );
 a102188a <=( (not A167)  and  (not A169) );
 a102189a <=( (not A170)  and  a102188a );
 a102192a <=( (not A200)  and  (not A199) );
 a102195a <=( A265  and  A203 );
 a102196a <=( a102195a  and  a102192a );
 a102197a <=( a102196a  and  a102189a );
 a102201a <=( (not A269)  and  A268 );
 a102202a <=( A266  and  a102201a );
 a102205a <=( (not A299)  and  A298 );
 a102208a <=( A301  and  (not A300) );
 a102209a <=( a102208a  and  a102205a );
 a102210a <=( a102209a  and  a102202a );
 a102214a <=( (not A167)  and  (not A169) );
 a102215a <=( (not A170)  and  a102214a );
 a102218a <=( (not A200)  and  (not A199) );
 a102221a <=( A265  and  A203 );
 a102222a <=( a102221a  and  a102218a );
 a102223a <=( a102222a  and  a102215a );
 a102227a <=( (not A269)  and  A268 );
 a102228a <=( A266  and  a102227a );
 a102231a <=( (not A299)  and  A298 );
 a102234a <=( (not A302)  and  (not A300) );
 a102235a <=( a102234a  and  a102231a );
 a102236a <=( a102235a  and  a102228a );
 a102240a <=( (not A167)  and  (not A169) );
 a102241a <=( (not A170)  and  a102240a );
 a102244a <=( (not A200)  and  (not A199) );
 a102247a <=( A265  and  A203 );
 a102248a <=( a102247a  and  a102244a );
 a102249a <=( a102248a  and  a102241a );
 a102253a <=( (not A269)  and  A268 );
 a102254a <=( A266  and  a102253a );
 a102257a <=( A299  and  (not A298) );
 a102260a <=( A301  and  (not A300) );
 a102261a <=( a102260a  and  a102257a );
 a102262a <=( a102261a  and  a102254a );
 a102266a <=( (not A167)  and  (not A169) );
 a102267a <=( (not A170)  and  a102266a );
 a102270a <=( (not A200)  and  (not A199) );
 a102273a <=( A265  and  A203 );
 a102274a <=( a102273a  and  a102270a );
 a102275a <=( a102274a  and  a102267a );
 a102279a <=( (not A269)  and  A268 );
 a102280a <=( A266  and  a102279a );
 a102283a <=( A299  and  (not A298) );
 a102286a <=( (not A302)  and  (not A300) );
 a102287a <=( a102286a  and  a102283a );
 a102288a <=( a102287a  and  a102280a );
 a102292a <=( (not A167)  and  (not A169) );
 a102293a <=( (not A170)  and  a102292a );
 a102296a <=( (not A200)  and  (not A199) );
 a102299a <=( (not A265)  and  A203 );
 a102300a <=( a102299a  and  a102296a );
 a102301a <=( a102300a  and  a102293a );
 a102305a <=( A269  and  (not A268) );
 a102306a <=( A266  and  a102305a );
 a102309a <=( A299  and  A298 );
 a102312a <=( (not A301)  and  (not A300) );
 a102313a <=( a102312a  and  a102309a );
 a102314a <=( a102313a  and  a102306a );
 a102318a <=( (not A167)  and  (not A169) );
 a102319a <=( (not A170)  and  a102318a );
 a102322a <=( (not A200)  and  (not A199) );
 a102325a <=( (not A265)  and  A203 );
 a102326a <=( a102325a  and  a102322a );
 a102327a <=( a102326a  and  a102319a );
 a102331a <=( A269  and  (not A268) );
 a102332a <=( A266  and  a102331a );
 a102335a <=( A299  and  A298 );
 a102338a <=( A302  and  (not A300) );
 a102339a <=( a102338a  and  a102335a );
 a102340a <=( a102339a  and  a102332a );
 a102344a <=( (not A167)  and  (not A169) );
 a102345a <=( (not A170)  and  a102344a );
 a102348a <=( (not A200)  and  (not A199) );
 a102351a <=( (not A265)  and  A203 );
 a102352a <=( a102351a  and  a102348a );
 a102353a <=( a102352a  and  a102345a );
 a102357a <=( A269  and  (not A268) );
 a102358a <=( A266  and  a102357a );
 a102361a <=( (not A299)  and  A298 );
 a102364a <=( A301  and  (not A300) );
 a102365a <=( a102364a  and  a102361a );
 a102366a <=( a102365a  and  a102358a );
 a102370a <=( (not A167)  and  (not A169) );
 a102371a <=( (not A170)  and  a102370a );
 a102374a <=( (not A200)  and  (not A199) );
 a102377a <=( (not A265)  and  A203 );
 a102378a <=( a102377a  and  a102374a );
 a102379a <=( a102378a  and  a102371a );
 a102383a <=( A269  and  (not A268) );
 a102384a <=( A266  and  a102383a );
 a102387a <=( (not A299)  and  A298 );
 a102390a <=( (not A302)  and  (not A300) );
 a102391a <=( a102390a  and  a102387a );
 a102392a <=( a102391a  and  a102384a );
 a102396a <=( (not A167)  and  (not A169) );
 a102397a <=( (not A170)  and  a102396a );
 a102400a <=( (not A200)  and  (not A199) );
 a102403a <=( (not A265)  and  A203 );
 a102404a <=( a102403a  and  a102400a );
 a102405a <=( a102404a  and  a102397a );
 a102409a <=( A269  and  (not A268) );
 a102410a <=( A266  and  a102409a );
 a102413a <=( A299  and  (not A298) );
 a102416a <=( A301  and  (not A300) );
 a102417a <=( a102416a  and  a102413a );
 a102418a <=( a102417a  and  a102410a );
 a102422a <=( (not A167)  and  (not A169) );
 a102423a <=( (not A170)  and  a102422a );
 a102426a <=( (not A200)  and  (not A199) );
 a102429a <=( (not A265)  and  A203 );
 a102430a <=( a102429a  and  a102426a );
 a102431a <=( a102430a  and  a102423a );
 a102435a <=( A269  and  (not A268) );
 a102436a <=( A266  and  a102435a );
 a102439a <=( A299  and  (not A298) );
 a102442a <=( (not A302)  and  (not A300) );
 a102443a <=( a102442a  and  a102439a );
 a102444a <=( a102443a  and  a102436a );
 a102448a <=( (not A167)  and  (not A169) );
 a102449a <=( (not A170)  and  a102448a );
 a102452a <=( (not A200)  and  (not A199) );
 a102455a <=( A265  and  A203 );
 a102456a <=( a102455a  and  a102452a );
 a102457a <=( a102456a  and  a102449a );
 a102461a <=( A269  and  (not A268) );
 a102462a <=( (not A266)  and  a102461a );
 a102465a <=( A299  and  A298 );
 a102468a <=( (not A301)  and  (not A300) );
 a102469a <=( a102468a  and  a102465a );
 a102470a <=( a102469a  and  a102462a );
 a102474a <=( (not A167)  and  (not A169) );
 a102475a <=( (not A170)  and  a102474a );
 a102478a <=( (not A200)  and  (not A199) );
 a102481a <=( A265  and  A203 );
 a102482a <=( a102481a  and  a102478a );
 a102483a <=( a102482a  and  a102475a );
 a102487a <=( A269  and  (not A268) );
 a102488a <=( (not A266)  and  a102487a );
 a102491a <=( A299  and  A298 );
 a102494a <=( A302  and  (not A300) );
 a102495a <=( a102494a  and  a102491a );
 a102496a <=( a102495a  and  a102488a );
 a102500a <=( (not A167)  and  (not A169) );
 a102501a <=( (not A170)  and  a102500a );
 a102504a <=( (not A200)  and  (not A199) );
 a102507a <=( A265  and  A203 );
 a102508a <=( a102507a  and  a102504a );
 a102509a <=( a102508a  and  a102501a );
 a102513a <=( A269  and  (not A268) );
 a102514a <=( (not A266)  and  a102513a );
 a102517a <=( (not A299)  and  A298 );
 a102520a <=( A301  and  (not A300) );
 a102521a <=( a102520a  and  a102517a );
 a102522a <=( a102521a  and  a102514a );
 a102526a <=( (not A167)  and  (not A169) );
 a102527a <=( (not A170)  and  a102526a );
 a102530a <=( (not A200)  and  (not A199) );
 a102533a <=( A265  and  A203 );
 a102534a <=( a102533a  and  a102530a );
 a102535a <=( a102534a  and  a102527a );
 a102539a <=( A269  and  (not A268) );
 a102540a <=( (not A266)  and  a102539a );
 a102543a <=( (not A299)  and  A298 );
 a102546a <=( (not A302)  and  (not A300) );
 a102547a <=( a102546a  and  a102543a );
 a102548a <=( a102547a  and  a102540a );
 a102552a <=( (not A167)  and  (not A169) );
 a102553a <=( (not A170)  and  a102552a );
 a102556a <=( (not A200)  and  (not A199) );
 a102559a <=( A265  and  A203 );
 a102560a <=( a102559a  and  a102556a );
 a102561a <=( a102560a  and  a102553a );
 a102565a <=( A269  and  (not A268) );
 a102566a <=( (not A266)  and  a102565a );
 a102569a <=( A299  and  (not A298) );
 a102572a <=( A301  and  (not A300) );
 a102573a <=( a102572a  and  a102569a );
 a102574a <=( a102573a  and  a102566a );
 a102578a <=( (not A167)  and  (not A169) );
 a102579a <=( (not A170)  and  a102578a );
 a102582a <=( (not A200)  and  (not A199) );
 a102585a <=( A265  and  A203 );
 a102586a <=( a102585a  and  a102582a );
 a102587a <=( a102586a  and  a102579a );
 a102591a <=( A269  and  (not A268) );
 a102592a <=( (not A266)  and  a102591a );
 a102595a <=( A299  and  (not A298) );
 a102598a <=( (not A302)  and  (not A300) );
 a102599a <=( a102598a  and  a102595a );
 a102600a <=( a102599a  and  a102592a );
 a102604a <=( (not A167)  and  (not A169) );
 a102605a <=( (not A170)  and  a102604a );
 a102608a <=( (not A200)  and  (not A199) );
 a102611a <=( (not A265)  and  A203 );
 a102612a <=( a102611a  and  a102608a );
 a102613a <=( a102612a  and  a102605a );
 a102617a <=( (not A269)  and  A268 );
 a102618a <=( (not A266)  and  a102617a );
 a102621a <=( A299  and  A298 );
 a102624a <=( (not A301)  and  (not A300) );
 a102625a <=( a102624a  and  a102621a );
 a102626a <=( a102625a  and  a102618a );
 a102630a <=( (not A167)  and  (not A169) );
 a102631a <=( (not A170)  and  a102630a );
 a102634a <=( (not A200)  and  (not A199) );
 a102637a <=( (not A265)  and  A203 );
 a102638a <=( a102637a  and  a102634a );
 a102639a <=( a102638a  and  a102631a );
 a102643a <=( (not A269)  and  A268 );
 a102644a <=( (not A266)  and  a102643a );
 a102647a <=( A299  and  A298 );
 a102650a <=( A302  and  (not A300) );
 a102651a <=( a102650a  and  a102647a );
 a102652a <=( a102651a  and  a102644a );
 a102656a <=( (not A167)  and  (not A169) );
 a102657a <=( (not A170)  and  a102656a );
 a102660a <=( (not A200)  and  (not A199) );
 a102663a <=( (not A265)  and  A203 );
 a102664a <=( a102663a  and  a102660a );
 a102665a <=( a102664a  and  a102657a );
 a102669a <=( (not A269)  and  A268 );
 a102670a <=( (not A266)  and  a102669a );
 a102673a <=( (not A299)  and  A298 );
 a102676a <=( A301  and  (not A300) );
 a102677a <=( a102676a  and  a102673a );
 a102678a <=( a102677a  and  a102670a );
 a102682a <=( (not A167)  and  (not A169) );
 a102683a <=( (not A170)  and  a102682a );
 a102686a <=( (not A200)  and  (not A199) );
 a102689a <=( (not A265)  and  A203 );
 a102690a <=( a102689a  and  a102686a );
 a102691a <=( a102690a  and  a102683a );
 a102695a <=( (not A269)  and  A268 );
 a102696a <=( (not A266)  and  a102695a );
 a102699a <=( (not A299)  and  A298 );
 a102702a <=( (not A302)  and  (not A300) );
 a102703a <=( a102702a  and  a102699a );
 a102704a <=( a102703a  and  a102696a );
 a102708a <=( (not A167)  and  (not A169) );
 a102709a <=( (not A170)  and  a102708a );
 a102712a <=( (not A200)  and  (not A199) );
 a102715a <=( (not A265)  and  A203 );
 a102716a <=( a102715a  and  a102712a );
 a102717a <=( a102716a  and  a102709a );
 a102721a <=( (not A269)  and  A268 );
 a102722a <=( (not A266)  and  a102721a );
 a102725a <=( A299  and  (not A298) );
 a102728a <=( A301  and  (not A300) );
 a102729a <=( a102728a  and  a102725a );
 a102730a <=( a102729a  and  a102722a );
 a102734a <=( (not A167)  and  (not A169) );
 a102735a <=( (not A170)  and  a102734a );
 a102738a <=( (not A200)  and  (not A199) );
 a102741a <=( (not A265)  and  A203 );
 a102742a <=( a102741a  and  a102738a );
 a102743a <=( a102742a  and  a102735a );
 a102747a <=( (not A269)  and  A268 );
 a102748a <=( (not A266)  and  a102747a );
 a102751a <=( A299  and  (not A298) );
 a102754a <=( (not A302)  and  (not A300) );
 a102755a <=( a102754a  and  a102751a );
 a102756a <=( a102755a  and  a102748a );
 a102760a <=( (not A167)  and  (not A169) );
 a102761a <=( (not A170)  and  a102760a );
 a102764a <=( (not A200)  and  (not A199) );
 a102767a <=( (not A203)  and  A202 );
 a102768a <=( a102767a  and  a102764a );
 a102769a <=( a102768a  and  a102761a );
 a102773a <=( (not A268)  and  (not A266) );
 a102774a <=( (not A265)  and  a102773a );
 a102777a <=( A299  and  A298 );
 a102780a <=( (not A302)  and  A301 );
 a102781a <=( a102780a  and  a102777a );
 a102782a <=( a102781a  and  a102774a );
 a102786a <=( (not A167)  and  (not A169) );
 a102787a <=( (not A170)  and  a102786a );
 a102790a <=( (not A200)  and  (not A199) );
 a102793a <=( (not A203)  and  A202 );
 a102794a <=( a102793a  and  a102790a );
 a102795a <=( a102794a  and  a102787a );
 a102799a <=( (not A268)  and  (not A266) );
 a102800a <=( (not A265)  and  a102799a );
 a102803a <=( (not A299)  and  A298 );
 a102806a <=( A302  and  (not A301) );
 a102807a <=( a102806a  and  a102803a );
 a102808a <=( a102807a  and  a102800a );
 a102812a <=( (not A167)  and  (not A169) );
 a102813a <=( (not A170)  and  a102812a );
 a102816a <=( (not A200)  and  (not A199) );
 a102819a <=( (not A203)  and  A202 );
 a102820a <=( a102819a  and  a102816a );
 a102821a <=( a102820a  and  a102813a );
 a102825a <=( (not A268)  and  (not A266) );
 a102826a <=( (not A265)  and  a102825a );
 a102829a <=( A299  and  (not A298) );
 a102832a <=( A302  and  (not A301) );
 a102833a <=( a102832a  and  a102829a );
 a102834a <=( a102833a  and  a102826a );
 a102838a <=( (not A167)  and  (not A169) );
 a102839a <=( (not A170)  and  a102838a );
 a102842a <=( (not A200)  and  (not A199) );
 a102845a <=( (not A203)  and  A202 );
 a102846a <=( a102845a  and  a102842a );
 a102847a <=( a102846a  and  a102839a );
 a102851a <=( (not A268)  and  (not A266) );
 a102852a <=( (not A265)  and  a102851a );
 a102855a <=( (not A299)  and  (not A298) );
 a102858a <=( (not A302)  and  A301 );
 a102859a <=( a102858a  and  a102855a );
 a102860a <=( a102859a  and  a102852a );
 a102864a <=( (not A167)  and  (not A169) );
 a102865a <=( (not A170)  and  a102864a );
 a102868a <=( (not A200)  and  (not A199) );
 a102871a <=( (not A203)  and  A202 );
 a102872a <=( a102871a  and  a102868a );
 a102873a <=( a102872a  and  a102865a );
 a102877a <=( A269  and  (not A266) );
 a102878a <=( (not A265)  and  a102877a );
 a102881a <=( A299  and  A298 );
 a102884a <=( (not A302)  and  A301 );
 a102885a <=( a102884a  and  a102881a );
 a102886a <=( a102885a  and  a102878a );
 a102890a <=( (not A167)  and  (not A169) );
 a102891a <=( (not A170)  and  a102890a );
 a102894a <=( (not A200)  and  (not A199) );
 a102897a <=( (not A203)  and  A202 );
 a102898a <=( a102897a  and  a102894a );
 a102899a <=( a102898a  and  a102891a );
 a102903a <=( A269  and  (not A266) );
 a102904a <=( (not A265)  and  a102903a );
 a102907a <=( (not A299)  and  A298 );
 a102910a <=( A302  and  (not A301) );
 a102911a <=( a102910a  and  a102907a );
 a102912a <=( a102911a  and  a102904a );
 a102916a <=( (not A167)  and  (not A169) );
 a102917a <=( (not A170)  and  a102916a );
 a102920a <=( (not A200)  and  (not A199) );
 a102923a <=( (not A203)  and  A202 );
 a102924a <=( a102923a  and  a102920a );
 a102925a <=( a102924a  and  a102917a );
 a102929a <=( A269  and  (not A266) );
 a102930a <=( (not A265)  and  a102929a );
 a102933a <=( A299  and  (not A298) );
 a102936a <=( A302  and  (not A301) );
 a102937a <=( a102936a  and  a102933a );
 a102938a <=( a102937a  and  a102930a );
 a102942a <=( (not A167)  and  (not A169) );
 a102943a <=( (not A170)  and  a102942a );
 a102946a <=( (not A200)  and  (not A199) );
 a102949a <=( (not A203)  and  A202 );
 a102950a <=( a102949a  and  a102946a );
 a102951a <=( a102950a  and  a102943a );
 a102955a <=( A269  and  (not A266) );
 a102956a <=( (not A265)  and  a102955a );
 a102959a <=( (not A299)  and  (not A298) );
 a102962a <=( (not A302)  and  A301 );
 a102963a <=( a102962a  and  a102959a );
 a102964a <=( a102963a  and  a102956a );
 a102968a <=( (not A167)  and  A168 );
 a102969a <=( A170  and  a102968a );
 a102972a <=( A199  and  A166 );
 a102975a <=( A202  and  A200 );
 a102976a <=( a102975a  and  a102972a );
 a102977a <=( a102976a  and  a102969a );
 a102980a <=( A265  and  (not A203) );
 a102983a <=( A268  and  A266 );
 a102984a <=( a102983a  and  a102980a );
 a102987a <=( (not A298)  and  (not A269) );
 a102990a <=( (not A301)  and  (not A299) );
 a102991a <=( a102990a  and  a102987a );
 a102992a <=( a102991a  and  a102984a );
 a102996a <=( (not A167)  and  A168 );
 a102997a <=( A170  and  a102996a );
 a103000a <=( A199  and  A166 );
 a103003a <=( A202  and  A200 );
 a103004a <=( a103003a  and  a103000a );
 a103005a <=( a103004a  and  a102997a );
 a103008a <=( A265  and  (not A203) );
 a103011a <=( A268  and  A266 );
 a103012a <=( a103011a  and  a103008a );
 a103015a <=( (not A298)  and  (not A269) );
 a103018a <=( A302  and  (not A299) );
 a103019a <=( a103018a  and  a103015a );
 a103020a <=( a103019a  and  a103012a );
 a103024a <=( (not A167)  and  A168 );
 a103025a <=( A170  and  a103024a );
 a103028a <=( A199  and  A166 );
 a103031a <=( A202  and  A200 );
 a103032a <=( a103031a  and  a103028a );
 a103033a <=( a103032a  and  a103025a );
 a103036a <=( (not A265)  and  (not A203) );
 a103039a <=( (not A268)  and  A266 );
 a103040a <=( a103039a  and  a103036a );
 a103043a <=( (not A298)  and  A269 );
 a103046a <=( (not A301)  and  (not A299) );
 a103047a <=( a103046a  and  a103043a );
 a103048a <=( a103047a  and  a103040a );
 a103052a <=( (not A167)  and  A168 );
 a103053a <=( A170  and  a103052a );
 a103056a <=( A199  and  A166 );
 a103059a <=( A202  and  A200 );
 a103060a <=( a103059a  and  a103056a );
 a103061a <=( a103060a  and  a103053a );
 a103064a <=( (not A265)  and  (not A203) );
 a103067a <=( (not A268)  and  A266 );
 a103068a <=( a103067a  and  a103064a );
 a103071a <=( (not A298)  and  A269 );
 a103074a <=( A302  and  (not A299) );
 a103075a <=( a103074a  and  a103071a );
 a103076a <=( a103075a  and  a103068a );
 a103080a <=( (not A167)  and  A168 );
 a103081a <=( A170  and  a103080a );
 a103084a <=( A199  and  A166 );
 a103087a <=( A202  and  A200 );
 a103088a <=( a103087a  and  a103084a );
 a103089a <=( a103088a  and  a103081a );
 a103092a <=( A265  and  (not A203) );
 a103095a <=( (not A268)  and  (not A266) );
 a103096a <=( a103095a  and  a103092a );
 a103099a <=( (not A298)  and  A269 );
 a103102a <=( (not A301)  and  (not A299) );
 a103103a <=( a103102a  and  a103099a );
 a103104a <=( a103103a  and  a103096a );
 a103108a <=( (not A167)  and  A168 );
 a103109a <=( A170  and  a103108a );
 a103112a <=( A199  and  A166 );
 a103115a <=( A202  and  A200 );
 a103116a <=( a103115a  and  a103112a );
 a103117a <=( a103116a  and  a103109a );
 a103120a <=( A265  and  (not A203) );
 a103123a <=( (not A268)  and  (not A266) );
 a103124a <=( a103123a  and  a103120a );
 a103127a <=( (not A298)  and  A269 );
 a103130a <=( A302  and  (not A299) );
 a103131a <=( a103130a  and  a103127a );
 a103132a <=( a103131a  and  a103124a );
 a103136a <=( (not A167)  and  A168 );
 a103137a <=( A170  and  a103136a );
 a103140a <=( A199  and  A166 );
 a103143a <=( A202  and  A200 );
 a103144a <=( a103143a  and  a103140a );
 a103145a <=( a103144a  and  a103137a );
 a103148a <=( (not A265)  and  (not A203) );
 a103151a <=( A268  and  (not A266) );
 a103152a <=( a103151a  and  a103148a );
 a103155a <=( (not A298)  and  (not A269) );
 a103158a <=( (not A301)  and  (not A299) );
 a103159a <=( a103158a  and  a103155a );
 a103160a <=( a103159a  and  a103152a );
 a103164a <=( (not A167)  and  A168 );
 a103165a <=( A170  and  a103164a );
 a103168a <=( A199  and  A166 );
 a103171a <=( A202  and  A200 );
 a103172a <=( a103171a  and  a103168a );
 a103173a <=( a103172a  and  a103165a );
 a103176a <=( (not A265)  and  (not A203) );
 a103179a <=( A268  and  (not A266) );
 a103180a <=( a103179a  and  a103176a );
 a103183a <=( (not A298)  and  (not A269) );
 a103186a <=( A302  and  (not A299) );
 a103187a <=( a103186a  and  a103183a );
 a103188a <=( a103187a  and  a103180a );
 a103192a <=( (not A167)  and  A168 );
 a103193a <=( A170  and  a103192a );
 a103196a <=( A199  and  A166 );
 a103199a <=( (not A201)  and  A200 );
 a103200a <=( a103199a  and  a103196a );
 a103201a <=( a103200a  and  a103193a );
 a103204a <=( (not A265)  and  (not A202) );
 a103207a <=( (not A268)  and  (not A266) );
 a103208a <=( a103207a  and  a103204a );
 a103211a <=( A299  and  A298 );
 a103214a <=( (not A302)  and  A301 );
 a103215a <=( a103214a  and  a103211a );
 a103216a <=( a103215a  and  a103208a );
 a103220a <=( (not A167)  and  A168 );
 a103221a <=( A170  and  a103220a );
 a103224a <=( A199  and  A166 );
 a103227a <=( (not A201)  and  A200 );
 a103228a <=( a103227a  and  a103224a );
 a103229a <=( a103228a  and  a103221a );
 a103232a <=( (not A265)  and  (not A202) );
 a103235a <=( (not A268)  and  (not A266) );
 a103236a <=( a103235a  and  a103232a );
 a103239a <=( (not A299)  and  A298 );
 a103242a <=( A302  and  (not A301) );
 a103243a <=( a103242a  and  a103239a );
 a103244a <=( a103243a  and  a103236a );
 a103248a <=( (not A167)  and  A168 );
 a103249a <=( A170  and  a103248a );
 a103252a <=( A199  and  A166 );
 a103255a <=( (not A201)  and  A200 );
 a103256a <=( a103255a  and  a103252a );
 a103257a <=( a103256a  and  a103249a );
 a103260a <=( (not A265)  and  (not A202) );
 a103263a <=( (not A268)  and  (not A266) );
 a103264a <=( a103263a  and  a103260a );
 a103267a <=( A299  and  (not A298) );
 a103270a <=( A302  and  (not A301) );
 a103271a <=( a103270a  and  a103267a );
 a103272a <=( a103271a  and  a103264a );
 a103276a <=( (not A167)  and  A168 );
 a103277a <=( A170  and  a103276a );
 a103280a <=( A199  and  A166 );
 a103283a <=( (not A201)  and  A200 );
 a103284a <=( a103283a  and  a103280a );
 a103285a <=( a103284a  and  a103277a );
 a103288a <=( (not A265)  and  (not A202) );
 a103291a <=( (not A268)  and  (not A266) );
 a103292a <=( a103291a  and  a103288a );
 a103295a <=( (not A299)  and  (not A298) );
 a103298a <=( (not A302)  and  A301 );
 a103299a <=( a103298a  and  a103295a );
 a103300a <=( a103299a  and  a103292a );
 a103304a <=( (not A167)  and  A168 );
 a103305a <=( A170  and  a103304a );
 a103308a <=( A199  and  A166 );
 a103311a <=( (not A201)  and  A200 );
 a103312a <=( a103311a  and  a103308a );
 a103313a <=( a103312a  and  a103305a );
 a103316a <=( (not A265)  and  (not A202) );
 a103319a <=( A269  and  (not A266) );
 a103320a <=( a103319a  and  a103316a );
 a103323a <=( A299  and  A298 );
 a103326a <=( (not A302)  and  A301 );
 a103327a <=( a103326a  and  a103323a );
 a103328a <=( a103327a  and  a103320a );
 a103332a <=( (not A167)  and  A168 );
 a103333a <=( A170  and  a103332a );
 a103336a <=( A199  and  A166 );
 a103339a <=( (not A201)  and  A200 );
 a103340a <=( a103339a  and  a103336a );
 a103341a <=( a103340a  and  a103333a );
 a103344a <=( (not A265)  and  (not A202) );
 a103347a <=( A269  and  (not A266) );
 a103348a <=( a103347a  and  a103344a );
 a103351a <=( (not A299)  and  A298 );
 a103354a <=( A302  and  (not A301) );
 a103355a <=( a103354a  and  a103351a );
 a103356a <=( a103355a  and  a103348a );
 a103360a <=( (not A167)  and  A168 );
 a103361a <=( A170  and  a103360a );
 a103364a <=( A199  and  A166 );
 a103367a <=( (not A201)  and  A200 );
 a103368a <=( a103367a  and  a103364a );
 a103369a <=( a103368a  and  a103361a );
 a103372a <=( (not A265)  and  (not A202) );
 a103375a <=( A269  and  (not A266) );
 a103376a <=( a103375a  and  a103372a );
 a103379a <=( A299  and  (not A298) );
 a103382a <=( A302  and  (not A301) );
 a103383a <=( a103382a  and  a103379a );
 a103384a <=( a103383a  and  a103376a );
 a103388a <=( (not A167)  and  A168 );
 a103389a <=( A170  and  a103388a );
 a103392a <=( A199  and  A166 );
 a103395a <=( (not A201)  and  A200 );
 a103396a <=( a103395a  and  a103392a );
 a103397a <=( a103396a  and  a103389a );
 a103400a <=( (not A265)  and  (not A202) );
 a103403a <=( A269  and  (not A266) );
 a103404a <=( a103403a  and  a103400a );
 a103407a <=( (not A299)  and  (not A298) );
 a103410a <=( (not A302)  and  A301 );
 a103411a <=( a103410a  and  a103407a );
 a103412a <=( a103411a  and  a103404a );
 a103416a <=( (not A167)  and  A168 );
 a103417a <=( A170  and  a103416a );
 a103420a <=( A199  and  A166 );
 a103423a <=( (not A201)  and  A200 );
 a103424a <=( a103423a  and  a103420a );
 a103425a <=( a103424a  and  a103417a );
 a103428a <=( (not A265)  and  A203 );
 a103431a <=( (not A268)  and  (not A266) );
 a103432a <=( a103431a  and  a103428a );
 a103435a <=( A299  and  A298 );
 a103438a <=( (not A302)  and  A301 );
 a103439a <=( a103438a  and  a103435a );
 a103440a <=( a103439a  and  a103432a );
 a103444a <=( (not A167)  and  A168 );
 a103445a <=( A170  and  a103444a );
 a103448a <=( A199  and  A166 );
 a103451a <=( (not A201)  and  A200 );
 a103452a <=( a103451a  and  a103448a );
 a103453a <=( a103452a  and  a103445a );
 a103456a <=( (not A265)  and  A203 );
 a103459a <=( (not A268)  and  (not A266) );
 a103460a <=( a103459a  and  a103456a );
 a103463a <=( (not A299)  and  A298 );
 a103466a <=( A302  and  (not A301) );
 a103467a <=( a103466a  and  a103463a );
 a103468a <=( a103467a  and  a103460a );
 a103472a <=( (not A167)  and  A168 );
 a103473a <=( A170  and  a103472a );
 a103476a <=( A199  and  A166 );
 a103479a <=( (not A201)  and  A200 );
 a103480a <=( a103479a  and  a103476a );
 a103481a <=( a103480a  and  a103473a );
 a103484a <=( (not A265)  and  A203 );
 a103487a <=( (not A268)  and  (not A266) );
 a103488a <=( a103487a  and  a103484a );
 a103491a <=( A299  and  (not A298) );
 a103494a <=( A302  and  (not A301) );
 a103495a <=( a103494a  and  a103491a );
 a103496a <=( a103495a  and  a103488a );
 a103500a <=( (not A167)  and  A168 );
 a103501a <=( A170  and  a103500a );
 a103504a <=( A199  and  A166 );
 a103507a <=( (not A201)  and  A200 );
 a103508a <=( a103507a  and  a103504a );
 a103509a <=( a103508a  and  a103501a );
 a103512a <=( (not A265)  and  A203 );
 a103515a <=( (not A268)  and  (not A266) );
 a103516a <=( a103515a  and  a103512a );
 a103519a <=( (not A299)  and  (not A298) );
 a103522a <=( (not A302)  and  A301 );
 a103523a <=( a103522a  and  a103519a );
 a103524a <=( a103523a  and  a103516a );
 a103528a <=( (not A167)  and  A168 );
 a103529a <=( A170  and  a103528a );
 a103532a <=( A199  and  A166 );
 a103535a <=( (not A201)  and  A200 );
 a103536a <=( a103535a  and  a103532a );
 a103537a <=( a103536a  and  a103529a );
 a103540a <=( (not A265)  and  A203 );
 a103543a <=( A269  and  (not A266) );
 a103544a <=( a103543a  and  a103540a );
 a103547a <=( A299  and  A298 );
 a103550a <=( (not A302)  and  A301 );
 a103551a <=( a103550a  and  a103547a );
 a103552a <=( a103551a  and  a103544a );
 a103556a <=( (not A167)  and  A168 );
 a103557a <=( A170  and  a103556a );
 a103560a <=( A199  and  A166 );
 a103563a <=( (not A201)  and  A200 );
 a103564a <=( a103563a  and  a103560a );
 a103565a <=( a103564a  and  a103557a );
 a103568a <=( (not A265)  and  A203 );
 a103571a <=( A269  and  (not A266) );
 a103572a <=( a103571a  and  a103568a );
 a103575a <=( (not A299)  and  A298 );
 a103578a <=( A302  and  (not A301) );
 a103579a <=( a103578a  and  a103575a );
 a103580a <=( a103579a  and  a103572a );
 a103584a <=( (not A167)  and  A168 );
 a103585a <=( A170  and  a103584a );
 a103588a <=( A199  and  A166 );
 a103591a <=( (not A201)  and  A200 );
 a103592a <=( a103591a  and  a103588a );
 a103593a <=( a103592a  and  a103585a );
 a103596a <=( (not A265)  and  A203 );
 a103599a <=( A269  and  (not A266) );
 a103600a <=( a103599a  and  a103596a );
 a103603a <=( A299  and  (not A298) );
 a103606a <=( A302  and  (not A301) );
 a103607a <=( a103606a  and  a103603a );
 a103608a <=( a103607a  and  a103600a );
 a103612a <=( (not A167)  and  A168 );
 a103613a <=( A170  and  a103612a );
 a103616a <=( A199  and  A166 );
 a103619a <=( (not A201)  and  A200 );
 a103620a <=( a103619a  and  a103616a );
 a103621a <=( a103620a  and  a103613a );
 a103624a <=( (not A265)  and  A203 );
 a103627a <=( A269  and  (not A266) );
 a103628a <=( a103627a  and  a103624a );
 a103631a <=( (not A299)  and  (not A298) );
 a103634a <=( (not A302)  and  A301 );
 a103635a <=( a103634a  and  a103631a );
 a103636a <=( a103635a  and  a103628a );
 a103640a <=( (not A167)  and  A168 );
 a103641a <=( A170  and  a103640a );
 a103644a <=( (not A199)  and  A166 );
 a103647a <=( (not A202)  and  A200 );
 a103648a <=( a103647a  and  a103644a );
 a103649a <=( a103648a  and  a103641a );
 a103652a <=( A265  and  A203 );
 a103655a <=( A268  and  A266 );
 a103656a <=( a103655a  and  a103652a );
 a103659a <=( (not A298)  and  (not A269) );
 a103662a <=( (not A301)  and  (not A299) );
 a103663a <=( a103662a  and  a103659a );
 a103664a <=( a103663a  and  a103656a );
 a103668a <=( (not A167)  and  A168 );
 a103669a <=( A170  and  a103668a );
 a103672a <=( (not A199)  and  A166 );
 a103675a <=( (not A202)  and  A200 );
 a103676a <=( a103675a  and  a103672a );
 a103677a <=( a103676a  and  a103669a );
 a103680a <=( A265  and  A203 );
 a103683a <=( A268  and  A266 );
 a103684a <=( a103683a  and  a103680a );
 a103687a <=( (not A298)  and  (not A269) );
 a103690a <=( A302  and  (not A299) );
 a103691a <=( a103690a  and  a103687a );
 a103692a <=( a103691a  and  a103684a );
 a103696a <=( (not A167)  and  A168 );
 a103697a <=( A170  and  a103696a );
 a103700a <=( (not A199)  and  A166 );
 a103703a <=( (not A202)  and  A200 );
 a103704a <=( a103703a  and  a103700a );
 a103705a <=( a103704a  and  a103697a );
 a103708a <=( (not A265)  and  A203 );
 a103711a <=( (not A268)  and  A266 );
 a103712a <=( a103711a  and  a103708a );
 a103715a <=( (not A298)  and  A269 );
 a103718a <=( (not A301)  and  (not A299) );
 a103719a <=( a103718a  and  a103715a );
 a103720a <=( a103719a  and  a103712a );
 a103724a <=( (not A167)  and  A168 );
 a103725a <=( A170  and  a103724a );
 a103728a <=( (not A199)  and  A166 );
 a103731a <=( (not A202)  and  A200 );
 a103732a <=( a103731a  and  a103728a );
 a103733a <=( a103732a  and  a103725a );
 a103736a <=( (not A265)  and  A203 );
 a103739a <=( (not A268)  and  A266 );
 a103740a <=( a103739a  and  a103736a );
 a103743a <=( (not A298)  and  A269 );
 a103746a <=( A302  and  (not A299) );
 a103747a <=( a103746a  and  a103743a );
 a103748a <=( a103747a  and  a103740a );
 a103752a <=( (not A167)  and  A168 );
 a103753a <=( A170  and  a103752a );
 a103756a <=( (not A199)  and  A166 );
 a103759a <=( (not A202)  and  A200 );
 a103760a <=( a103759a  and  a103756a );
 a103761a <=( a103760a  and  a103753a );
 a103764a <=( A265  and  A203 );
 a103767a <=( (not A268)  and  (not A266) );
 a103768a <=( a103767a  and  a103764a );
 a103771a <=( (not A298)  and  A269 );
 a103774a <=( (not A301)  and  (not A299) );
 a103775a <=( a103774a  and  a103771a );
 a103776a <=( a103775a  and  a103768a );
 a103780a <=( (not A167)  and  A168 );
 a103781a <=( A170  and  a103780a );
 a103784a <=( (not A199)  and  A166 );
 a103787a <=( (not A202)  and  A200 );
 a103788a <=( a103787a  and  a103784a );
 a103789a <=( a103788a  and  a103781a );
 a103792a <=( A265  and  A203 );
 a103795a <=( (not A268)  and  (not A266) );
 a103796a <=( a103795a  and  a103792a );
 a103799a <=( (not A298)  and  A269 );
 a103802a <=( A302  and  (not A299) );
 a103803a <=( a103802a  and  a103799a );
 a103804a <=( a103803a  and  a103796a );
 a103808a <=( (not A167)  and  A168 );
 a103809a <=( A170  and  a103808a );
 a103812a <=( (not A199)  and  A166 );
 a103815a <=( (not A202)  and  A200 );
 a103816a <=( a103815a  and  a103812a );
 a103817a <=( a103816a  and  a103809a );
 a103820a <=( (not A265)  and  A203 );
 a103823a <=( A268  and  (not A266) );
 a103824a <=( a103823a  and  a103820a );
 a103827a <=( (not A298)  and  (not A269) );
 a103830a <=( (not A301)  and  (not A299) );
 a103831a <=( a103830a  and  a103827a );
 a103832a <=( a103831a  and  a103824a );
 a103836a <=( (not A167)  and  A168 );
 a103837a <=( A170  and  a103836a );
 a103840a <=( (not A199)  and  A166 );
 a103843a <=( (not A202)  and  A200 );
 a103844a <=( a103843a  and  a103840a );
 a103845a <=( a103844a  and  a103837a );
 a103848a <=( (not A265)  and  A203 );
 a103851a <=( A268  and  (not A266) );
 a103852a <=( a103851a  and  a103848a );
 a103855a <=( (not A298)  and  (not A269) );
 a103858a <=( A302  and  (not A299) );
 a103859a <=( a103858a  and  a103855a );
 a103860a <=( a103859a  and  a103852a );
 a103864a <=( (not A167)  and  A168 );
 a103865a <=( A170  and  a103864a );
 a103868a <=( (not A199)  and  A166 );
 a103871a <=( (not A201)  and  A200 );
 a103872a <=( a103871a  and  a103868a );
 a103873a <=( a103872a  and  a103865a );
 a103876a <=( (not A265)  and  A202 );
 a103879a <=( (not A268)  and  (not A266) );
 a103880a <=( a103879a  and  a103876a );
 a103883a <=( A299  and  A298 );
 a103886a <=( (not A302)  and  A301 );
 a103887a <=( a103886a  and  a103883a );
 a103888a <=( a103887a  and  a103880a );
 a103892a <=( (not A167)  and  A168 );
 a103893a <=( A170  and  a103892a );
 a103896a <=( (not A199)  and  A166 );
 a103899a <=( (not A201)  and  A200 );
 a103900a <=( a103899a  and  a103896a );
 a103901a <=( a103900a  and  a103893a );
 a103904a <=( (not A265)  and  A202 );
 a103907a <=( (not A268)  and  (not A266) );
 a103908a <=( a103907a  and  a103904a );
 a103911a <=( (not A299)  and  A298 );
 a103914a <=( A302  and  (not A301) );
 a103915a <=( a103914a  and  a103911a );
 a103916a <=( a103915a  and  a103908a );
 a103920a <=( (not A167)  and  A168 );
 a103921a <=( A170  and  a103920a );
 a103924a <=( (not A199)  and  A166 );
 a103927a <=( (not A201)  and  A200 );
 a103928a <=( a103927a  and  a103924a );
 a103929a <=( a103928a  and  a103921a );
 a103932a <=( (not A265)  and  A202 );
 a103935a <=( (not A268)  and  (not A266) );
 a103936a <=( a103935a  and  a103932a );
 a103939a <=( A299  and  (not A298) );
 a103942a <=( A302  and  (not A301) );
 a103943a <=( a103942a  and  a103939a );
 a103944a <=( a103943a  and  a103936a );
 a103948a <=( (not A167)  and  A168 );
 a103949a <=( A170  and  a103948a );
 a103952a <=( (not A199)  and  A166 );
 a103955a <=( (not A201)  and  A200 );
 a103956a <=( a103955a  and  a103952a );
 a103957a <=( a103956a  and  a103949a );
 a103960a <=( (not A265)  and  A202 );
 a103963a <=( (not A268)  and  (not A266) );
 a103964a <=( a103963a  and  a103960a );
 a103967a <=( (not A299)  and  (not A298) );
 a103970a <=( (not A302)  and  A301 );
 a103971a <=( a103970a  and  a103967a );
 a103972a <=( a103971a  and  a103964a );
 a103976a <=( (not A167)  and  A168 );
 a103977a <=( A170  and  a103976a );
 a103980a <=( (not A199)  and  A166 );
 a103983a <=( (not A201)  and  A200 );
 a103984a <=( a103983a  and  a103980a );
 a103985a <=( a103984a  and  a103977a );
 a103988a <=( (not A265)  and  A202 );
 a103991a <=( A269  and  (not A266) );
 a103992a <=( a103991a  and  a103988a );
 a103995a <=( A299  and  A298 );
 a103998a <=( (not A302)  and  A301 );
 a103999a <=( a103998a  and  a103995a );
 a104000a <=( a103999a  and  a103992a );
 a104004a <=( (not A167)  and  A168 );
 a104005a <=( A170  and  a104004a );
 a104008a <=( (not A199)  and  A166 );
 a104011a <=( (not A201)  and  A200 );
 a104012a <=( a104011a  and  a104008a );
 a104013a <=( a104012a  and  a104005a );
 a104016a <=( (not A265)  and  A202 );
 a104019a <=( A269  and  (not A266) );
 a104020a <=( a104019a  and  a104016a );
 a104023a <=( (not A299)  and  A298 );
 a104026a <=( A302  and  (not A301) );
 a104027a <=( a104026a  and  a104023a );
 a104028a <=( a104027a  and  a104020a );
 a104032a <=( (not A167)  and  A168 );
 a104033a <=( A170  and  a104032a );
 a104036a <=( (not A199)  and  A166 );
 a104039a <=( (not A201)  and  A200 );
 a104040a <=( a104039a  and  a104036a );
 a104041a <=( a104040a  and  a104033a );
 a104044a <=( (not A265)  and  A202 );
 a104047a <=( A269  and  (not A266) );
 a104048a <=( a104047a  and  a104044a );
 a104051a <=( A299  and  (not A298) );
 a104054a <=( A302  and  (not A301) );
 a104055a <=( a104054a  and  a104051a );
 a104056a <=( a104055a  and  a104048a );
 a104060a <=( (not A167)  and  A168 );
 a104061a <=( A170  and  a104060a );
 a104064a <=( (not A199)  and  A166 );
 a104067a <=( (not A201)  and  A200 );
 a104068a <=( a104067a  and  a104064a );
 a104069a <=( a104068a  and  a104061a );
 a104072a <=( (not A265)  and  A202 );
 a104075a <=( A269  and  (not A266) );
 a104076a <=( a104075a  and  a104072a );
 a104079a <=( (not A299)  and  (not A298) );
 a104082a <=( (not A302)  and  A301 );
 a104083a <=( a104082a  and  a104079a );
 a104084a <=( a104083a  and  a104076a );
 a104088a <=( (not A167)  and  A168 );
 a104089a <=( A170  and  a104088a );
 a104092a <=( (not A199)  and  A166 );
 a104095a <=( (not A201)  and  A200 );
 a104096a <=( a104095a  and  a104092a );
 a104097a <=( a104096a  and  a104089a );
 a104100a <=( (not A265)  and  (not A203) );
 a104103a <=( (not A268)  and  (not A266) );
 a104104a <=( a104103a  and  a104100a );
 a104107a <=( A299  and  A298 );
 a104110a <=( (not A302)  and  A301 );
 a104111a <=( a104110a  and  a104107a );
 a104112a <=( a104111a  and  a104104a );
 a104116a <=( (not A167)  and  A168 );
 a104117a <=( A170  and  a104116a );
 a104120a <=( (not A199)  and  A166 );
 a104123a <=( (not A201)  and  A200 );
 a104124a <=( a104123a  and  a104120a );
 a104125a <=( a104124a  and  a104117a );
 a104128a <=( (not A265)  and  (not A203) );
 a104131a <=( (not A268)  and  (not A266) );
 a104132a <=( a104131a  and  a104128a );
 a104135a <=( (not A299)  and  A298 );
 a104138a <=( A302  and  (not A301) );
 a104139a <=( a104138a  and  a104135a );
 a104140a <=( a104139a  and  a104132a );
 a104144a <=( (not A167)  and  A168 );
 a104145a <=( A170  and  a104144a );
 a104148a <=( (not A199)  and  A166 );
 a104151a <=( (not A201)  and  A200 );
 a104152a <=( a104151a  and  a104148a );
 a104153a <=( a104152a  and  a104145a );
 a104156a <=( (not A265)  and  (not A203) );
 a104159a <=( (not A268)  and  (not A266) );
 a104160a <=( a104159a  and  a104156a );
 a104163a <=( A299  and  (not A298) );
 a104166a <=( A302  and  (not A301) );
 a104167a <=( a104166a  and  a104163a );
 a104168a <=( a104167a  and  a104160a );
 a104172a <=( (not A167)  and  A168 );
 a104173a <=( A170  and  a104172a );
 a104176a <=( (not A199)  and  A166 );
 a104179a <=( (not A201)  and  A200 );
 a104180a <=( a104179a  and  a104176a );
 a104181a <=( a104180a  and  a104173a );
 a104184a <=( (not A265)  and  (not A203) );
 a104187a <=( (not A268)  and  (not A266) );
 a104188a <=( a104187a  and  a104184a );
 a104191a <=( (not A299)  and  (not A298) );
 a104194a <=( (not A302)  and  A301 );
 a104195a <=( a104194a  and  a104191a );
 a104196a <=( a104195a  and  a104188a );
 a104200a <=( (not A167)  and  A168 );
 a104201a <=( A170  and  a104200a );
 a104204a <=( (not A199)  and  A166 );
 a104207a <=( (not A201)  and  A200 );
 a104208a <=( a104207a  and  a104204a );
 a104209a <=( a104208a  and  a104201a );
 a104212a <=( (not A265)  and  (not A203) );
 a104215a <=( A269  and  (not A266) );
 a104216a <=( a104215a  and  a104212a );
 a104219a <=( A299  and  A298 );
 a104222a <=( (not A302)  and  A301 );
 a104223a <=( a104222a  and  a104219a );
 a104224a <=( a104223a  and  a104216a );
 a104228a <=( (not A167)  and  A168 );
 a104229a <=( A170  and  a104228a );
 a104232a <=( (not A199)  and  A166 );
 a104235a <=( (not A201)  and  A200 );
 a104236a <=( a104235a  and  a104232a );
 a104237a <=( a104236a  and  a104229a );
 a104240a <=( (not A265)  and  (not A203) );
 a104243a <=( A269  and  (not A266) );
 a104244a <=( a104243a  and  a104240a );
 a104247a <=( (not A299)  and  A298 );
 a104250a <=( A302  and  (not A301) );
 a104251a <=( a104250a  and  a104247a );
 a104252a <=( a104251a  and  a104244a );
 a104256a <=( (not A167)  and  A168 );
 a104257a <=( A170  and  a104256a );
 a104260a <=( (not A199)  and  A166 );
 a104263a <=( (not A201)  and  A200 );
 a104264a <=( a104263a  and  a104260a );
 a104265a <=( a104264a  and  a104257a );
 a104268a <=( (not A265)  and  (not A203) );
 a104271a <=( A269  and  (not A266) );
 a104272a <=( a104271a  and  a104268a );
 a104275a <=( A299  and  (not A298) );
 a104278a <=( A302  and  (not A301) );
 a104279a <=( a104278a  and  a104275a );
 a104280a <=( a104279a  and  a104272a );
 a104284a <=( (not A167)  and  A168 );
 a104285a <=( A170  and  a104284a );
 a104288a <=( (not A199)  and  A166 );
 a104291a <=( (not A201)  and  A200 );
 a104292a <=( a104291a  and  a104288a );
 a104293a <=( a104292a  and  a104285a );
 a104296a <=( (not A265)  and  (not A203) );
 a104299a <=( A269  and  (not A266) );
 a104300a <=( a104299a  and  a104296a );
 a104303a <=( (not A299)  and  (not A298) );
 a104306a <=( (not A302)  and  A301 );
 a104307a <=( a104306a  and  a104303a );
 a104308a <=( a104307a  and  a104300a );
 a104312a <=( (not A167)  and  A168 );
 a104313a <=( A170  and  a104312a );
 a104316a <=( A199  and  A166 );
 a104319a <=( (not A202)  and  (not A200) );
 a104320a <=( a104319a  and  a104316a );
 a104321a <=( a104320a  and  a104313a );
 a104324a <=( A265  and  A203 );
 a104327a <=( A268  and  A266 );
 a104328a <=( a104327a  and  a104324a );
 a104331a <=( (not A298)  and  (not A269) );
 a104334a <=( (not A301)  and  (not A299) );
 a104335a <=( a104334a  and  a104331a );
 a104336a <=( a104335a  and  a104328a );
 a104340a <=( (not A167)  and  A168 );
 a104341a <=( A170  and  a104340a );
 a104344a <=( A199  and  A166 );
 a104347a <=( (not A202)  and  (not A200) );
 a104348a <=( a104347a  and  a104344a );
 a104349a <=( a104348a  and  a104341a );
 a104352a <=( A265  and  A203 );
 a104355a <=( A268  and  A266 );
 a104356a <=( a104355a  and  a104352a );
 a104359a <=( (not A298)  and  (not A269) );
 a104362a <=( A302  and  (not A299) );
 a104363a <=( a104362a  and  a104359a );
 a104364a <=( a104363a  and  a104356a );
 a104368a <=( (not A167)  and  A168 );
 a104369a <=( A170  and  a104368a );
 a104372a <=( A199  and  A166 );
 a104375a <=( (not A202)  and  (not A200) );
 a104376a <=( a104375a  and  a104372a );
 a104377a <=( a104376a  and  a104369a );
 a104380a <=( (not A265)  and  A203 );
 a104383a <=( (not A268)  and  A266 );
 a104384a <=( a104383a  and  a104380a );
 a104387a <=( (not A298)  and  A269 );
 a104390a <=( (not A301)  and  (not A299) );
 a104391a <=( a104390a  and  a104387a );
 a104392a <=( a104391a  and  a104384a );
 a104396a <=( (not A167)  and  A168 );
 a104397a <=( A170  and  a104396a );
 a104400a <=( A199  and  A166 );
 a104403a <=( (not A202)  and  (not A200) );
 a104404a <=( a104403a  and  a104400a );
 a104405a <=( a104404a  and  a104397a );
 a104408a <=( (not A265)  and  A203 );
 a104411a <=( (not A268)  and  A266 );
 a104412a <=( a104411a  and  a104408a );
 a104415a <=( (not A298)  and  A269 );
 a104418a <=( A302  and  (not A299) );
 a104419a <=( a104418a  and  a104415a );
 a104420a <=( a104419a  and  a104412a );
 a104424a <=( (not A167)  and  A168 );
 a104425a <=( A170  and  a104424a );
 a104428a <=( A199  and  A166 );
 a104431a <=( (not A202)  and  (not A200) );
 a104432a <=( a104431a  and  a104428a );
 a104433a <=( a104432a  and  a104425a );
 a104436a <=( A265  and  A203 );
 a104439a <=( (not A268)  and  (not A266) );
 a104440a <=( a104439a  and  a104436a );
 a104443a <=( (not A298)  and  A269 );
 a104446a <=( (not A301)  and  (not A299) );
 a104447a <=( a104446a  and  a104443a );
 a104448a <=( a104447a  and  a104440a );
 a104452a <=( (not A167)  and  A168 );
 a104453a <=( A170  and  a104452a );
 a104456a <=( A199  and  A166 );
 a104459a <=( (not A202)  and  (not A200) );
 a104460a <=( a104459a  and  a104456a );
 a104461a <=( a104460a  and  a104453a );
 a104464a <=( A265  and  A203 );
 a104467a <=( (not A268)  and  (not A266) );
 a104468a <=( a104467a  and  a104464a );
 a104471a <=( (not A298)  and  A269 );
 a104474a <=( A302  and  (not A299) );
 a104475a <=( a104474a  and  a104471a );
 a104476a <=( a104475a  and  a104468a );
 a104480a <=( (not A167)  and  A168 );
 a104481a <=( A170  and  a104480a );
 a104484a <=( A199  and  A166 );
 a104487a <=( (not A202)  and  (not A200) );
 a104488a <=( a104487a  and  a104484a );
 a104489a <=( a104488a  and  a104481a );
 a104492a <=( (not A265)  and  A203 );
 a104495a <=( A268  and  (not A266) );
 a104496a <=( a104495a  and  a104492a );
 a104499a <=( (not A298)  and  (not A269) );
 a104502a <=( (not A301)  and  (not A299) );
 a104503a <=( a104502a  and  a104499a );
 a104504a <=( a104503a  and  a104496a );
 a104508a <=( (not A167)  and  A168 );
 a104509a <=( A170  and  a104508a );
 a104512a <=( A199  and  A166 );
 a104515a <=( (not A202)  and  (not A200) );
 a104516a <=( a104515a  and  a104512a );
 a104517a <=( a104516a  and  a104509a );
 a104520a <=( (not A265)  and  A203 );
 a104523a <=( A268  and  (not A266) );
 a104524a <=( a104523a  and  a104520a );
 a104527a <=( (not A298)  and  (not A269) );
 a104530a <=( A302  and  (not A299) );
 a104531a <=( a104530a  and  a104527a );
 a104532a <=( a104531a  and  a104524a );
 a104536a <=( (not A167)  and  A168 );
 a104537a <=( A170  and  a104536a );
 a104540a <=( A199  and  A166 );
 a104543a <=( (not A201)  and  (not A200) );
 a104544a <=( a104543a  and  a104540a );
 a104545a <=( a104544a  and  a104537a );
 a104548a <=( (not A265)  and  A202 );
 a104551a <=( (not A268)  and  (not A266) );
 a104552a <=( a104551a  and  a104548a );
 a104555a <=( A299  and  A298 );
 a104558a <=( (not A302)  and  A301 );
 a104559a <=( a104558a  and  a104555a );
 a104560a <=( a104559a  and  a104552a );
 a104564a <=( (not A167)  and  A168 );
 a104565a <=( A170  and  a104564a );
 a104568a <=( A199  and  A166 );
 a104571a <=( (not A201)  and  (not A200) );
 a104572a <=( a104571a  and  a104568a );
 a104573a <=( a104572a  and  a104565a );
 a104576a <=( (not A265)  and  A202 );
 a104579a <=( (not A268)  and  (not A266) );
 a104580a <=( a104579a  and  a104576a );
 a104583a <=( (not A299)  and  A298 );
 a104586a <=( A302  and  (not A301) );
 a104587a <=( a104586a  and  a104583a );
 a104588a <=( a104587a  and  a104580a );
 a104592a <=( (not A167)  and  A168 );
 a104593a <=( A170  and  a104592a );
 a104596a <=( A199  and  A166 );
 a104599a <=( (not A201)  and  (not A200) );
 a104600a <=( a104599a  and  a104596a );
 a104601a <=( a104600a  and  a104593a );
 a104604a <=( (not A265)  and  A202 );
 a104607a <=( (not A268)  and  (not A266) );
 a104608a <=( a104607a  and  a104604a );
 a104611a <=( A299  and  (not A298) );
 a104614a <=( A302  and  (not A301) );
 a104615a <=( a104614a  and  a104611a );
 a104616a <=( a104615a  and  a104608a );
 a104620a <=( (not A167)  and  A168 );
 a104621a <=( A170  and  a104620a );
 a104624a <=( A199  and  A166 );
 a104627a <=( (not A201)  and  (not A200) );
 a104628a <=( a104627a  and  a104624a );
 a104629a <=( a104628a  and  a104621a );
 a104632a <=( (not A265)  and  A202 );
 a104635a <=( (not A268)  and  (not A266) );
 a104636a <=( a104635a  and  a104632a );
 a104639a <=( (not A299)  and  (not A298) );
 a104642a <=( (not A302)  and  A301 );
 a104643a <=( a104642a  and  a104639a );
 a104644a <=( a104643a  and  a104636a );
 a104648a <=( (not A167)  and  A168 );
 a104649a <=( A170  and  a104648a );
 a104652a <=( A199  and  A166 );
 a104655a <=( (not A201)  and  (not A200) );
 a104656a <=( a104655a  and  a104652a );
 a104657a <=( a104656a  and  a104649a );
 a104660a <=( (not A265)  and  A202 );
 a104663a <=( A269  and  (not A266) );
 a104664a <=( a104663a  and  a104660a );
 a104667a <=( A299  and  A298 );
 a104670a <=( (not A302)  and  A301 );
 a104671a <=( a104670a  and  a104667a );
 a104672a <=( a104671a  and  a104664a );
 a104676a <=( (not A167)  and  A168 );
 a104677a <=( A170  and  a104676a );
 a104680a <=( A199  and  A166 );
 a104683a <=( (not A201)  and  (not A200) );
 a104684a <=( a104683a  and  a104680a );
 a104685a <=( a104684a  and  a104677a );
 a104688a <=( (not A265)  and  A202 );
 a104691a <=( A269  and  (not A266) );
 a104692a <=( a104691a  and  a104688a );
 a104695a <=( (not A299)  and  A298 );
 a104698a <=( A302  and  (not A301) );
 a104699a <=( a104698a  and  a104695a );
 a104700a <=( a104699a  and  a104692a );
 a104704a <=( (not A167)  and  A168 );
 a104705a <=( A170  and  a104704a );
 a104708a <=( A199  and  A166 );
 a104711a <=( (not A201)  and  (not A200) );
 a104712a <=( a104711a  and  a104708a );
 a104713a <=( a104712a  and  a104705a );
 a104716a <=( (not A265)  and  A202 );
 a104719a <=( A269  and  (not A266) );
 a104720a <=( a104719a  and  a104716a );
 a104723a <=( A299  and  (not A298) );
 a104726a <=( A302  and  (not A301) );
 a104727a <=( a104726a  and  a104723a );
 a104728a <=( a104727a  and  a104720a );
 a104732a <=( (not A167)  and  A168 );
 a104733a <=( A170  and  a104732a );
 a104736a <=( A199  and  A166 );
 a104739a <=( (not A201)  and  (not A200) );
 a104740a <=( a104739a  and  a104736a );
 a104741a <=( a104740a  and  a104733a );
 a104744a <=( (not A265)  and  A202 );
 a104747a <=( A269  and  (not A266) );
 a104748a <=( a104747a  and  a104744a );
 a104751a <=( (not A299)  and  (not A298) );
 a104754a <=( (not A302)  and  A301 );
 a104755a <=( a104754a  and  a104751a );
 a104756a <=( a104755a  and  a104748a );
 a104760a <=( (not A167)  and  A168 );
 a104761a <=( A170  and  a104760a );
 a104764a <=( A199  and  A166 );
 a104767a <=( (not A201)  and  (not A200) );
 a104768a <=( a104767a  and  a104764a );
 a104769a <=( a104768a  and  a104761a );
 a104772a <=( (not A265)  and  (not A203) );
 a104775a <=( (not A268)  and  (not A266) );
 a104776a <=( a104775a  and  a104772a );
 a104779a <=( A299  and  A298 );
 a104782a <=( (not A302)  and  A301 );
 a104783a <=( a104782a  and  a104779a );
 a104784a <=( a104783a  and  a104776a );
 a104788a <=( (not A167)  and  A168 );
 a104789a <=( A170  and  a104788a );
 a104792a <=( A199  and  A166 );
 a104795a <=( (not A201)  and  (not A200) );
 a104796a <=( a104795a  and  a104792a );
 a104797a <=( a104796a  and  a104789a );
 a104800a <=( (not A265)  and  (not A203) );
 a104803a <=( (not A268)  and  (not A266) );
 a104804a <=( a104803a  and  a104800a );
 a104807a <=( (not A299)  and  A298 );
 a104810a <=( A302  and  (not A301) );
 a104811a <=( a104810a  and  a104807a );
 a104812a <=( a104811a  and  a104804a );
 a104816a <=( (not A167)  and  A168 );
 a104817a <=( A170  and  a104816a );
 a104820a <=( A199  and  A166 );
 a104823a <=( (not A201)  and  (not A200) );
 a104824a <=( a104823a  and  a104820a );
 a104825a <=( a104824a  and  a104817a );
 a104828a <=( (not A265)  and  (not A203) );
 a104831a <=( (not A268)  and  (not A266) );
 a104832a <=( a104831a  and  a104828a );
 a104835a <=( A299  and  (not A298) );
 a104838a <=( A302  and  (not A301) );
 a104839a <=( a104838a  and  a104835a );
 a104840a <=( a104839a  and  a104832a );
 a104844a <=( (not A167)  and  A168 );
 a104845a <=( A170  and  a104844a );
 a104848a <=( A199  and  A166 );
 a104851a <=( (not A201)  and  (not A200) );
 a104852a <=( a104851a  and  a104848a );
 a104853a <=( a104852a  and  a104845a );
 a104856a <=( (not A265)  and  (not A203) );
 a104859a <=( (not A268)  and  (not A266) );
 a104860a <=( a104859a  and  a104856a );
 a104863a <=( (not A299)  and  (not A298) );
 a104866a <=( (not A302)  and  A301 );
 a104867a <=( a104866a  and  a104863a );
 a104868a <=( a104867a  and  a104860a );
 a104872a <=( (not A167)  and  A168 );
 a104873a <=( A170  and  a104872a );
 a104876a <=( A199  and  A166 );
 a104879a <=( (not A201)  and  (not A200) );
 a104880a <=( a104879a  and  a104876a );
 a104881a <=( a104880a  and  a104873a );
 a104884a <=( (not A265)  and  (not A203) );
 a104887a <=( A269  and  (not A266) );
 a104888a <=( a104887a  and  a104884a );
 a104891a <=( A299  and  A298 );
 a104894a <=( (not A302)  and  A301 );
 a104895a <=( a104894a  and  a104891a );
 a104896a <=( a104895a  and  a104888a );
 a104900a <=( (not A167)  and  A168 );
 a104901a <=( A170  and  a104900a );
 a104904a <=( A199  and  A166 );
 a104907a <=( (not A201)  and  (not A200) );
 a104908a <=( a104907a  and  a104904a );
 a104909a <=( a104908a  and  a104901a );
 a104912a <=( (not A265)  and  (not A203) );
 a104915a <=( A269  and  (not A266) );
 a104916a <=( a104915a  and  a104912a );
 a104919a <=( (not A299)  and  A298 );
 a104922a <=( A302  and  (not A301) );
 a104923a <=( a104922a  and  a104919a );
 a104924a <=( a104923a  and  a104916a );
 a104928a <=( (not A167)  and  A168 );
 a104929a <=( A170  and  a104928a );
 a104932a <=( A199  and  A166 );
 a104935a <=( (not A201)  and  (not A200) );
 a104936a <=( a104935a  and  a104932a );
 a104937a <=( a104936a  and  a104929a );
 a104940a <=( (not A265)  and  (not A203) );
 a104943a <=( A269  and  (not A266) );
 a104944a <=( a104943a  and  a104940a );
 a104947a <=( A299  and  (not A298) );
 a104950a <=( A302  and  (not A301) );
 a104951a <=( a104950a  and  a104947a );
 a104952a <=( a104951a  and  a104944a );
 a104956a <=( (not A167)  and  A168 );
 a104957a <=( A170  and  a104956a );
 a104960a <=( A199  and  A166 );
 a104963a <=( (not A201)  and  (not A200) );
 a104964a <=( a104963a  and  a104960a );
 a104965a <=( a104964a  and  a104957a );
 a104968a <=( (not A265)  and  (not A203) );
 a104971a <=( A269  and  (not A266) );
 a104972a <=( a104971a  and  a104968a );
 a104975a <=( (not A299)  and  (not A298) );
 a104978a <=( (not A302)  and  A301 );
 a104979a <=( a104978a  and  a104975a );
 a104980a <=( a104979a  and  a104972a );
 a104984a <=( (not A167)  and  A168 );
 a104985a <=( A170  and  a104984a );
 a104988a <=( (not A199)  and  A166 );
 a104991a <=( (not A202)  and  (not A200) );
 a104992a <=( a104991a  and  a104988a );
 a104993a <=( a104992a  and  a104985a );
 a104996a <=( A266  and  A265 );
 a104999a <=( (not A268)  and  (not A267) );
 a105000a <=( a104999a  and  a104996a );
 a105003a <=( A299  and  A298 );
 a105006a <=( (not A302)  and  A301 );
 a105007a <=( a105006a  and  a105003a );
 a105008a <=( a105007a  and  a105000a );
 a105012a <=( (not A167)  and  A168 );
 a105013a <=( A170  and  a105012a );
 a105016a <=( (not A199)  and  A166 );
 a105019a <=( (not A202)  and  (not A200) );
 a105020a <=( a105019a  and  a105016a );
 a105021a <=( a105020a  and  a105013a );
 a105024a <=( A266  and  A265 );
 a105027a <=( (not A268)  and  (not A267) );
 a105028a <=( a105027a  and  a105024a );
 a105031a <=( (not A299)  and  A298 );
 a105034a <=( A302  and  (not A301) );
 a105035a <=( a105034a  and  a105031a );
 a105036a <=( a105035a  and  a105028a );
 a105040a <=( (not A167)  and  A168 );
 a105041a <=( A170  and  a105040a );
 a105044a <=( (not A199)  and  A166 );
 a105047a <=( (not A202)  and  (not A200) );
 a105048a <=( a105047a  and  a105044a );
 a105049a <=( a105048a  and  a105041a );
 a105052a <=( A266  and  A265 );
 a105055a <=( (not A268)  and  (not A267) );
 a105056a <=( a105055a  and  a105052a );
 a105059a <=( A299  and  (not A298) );
 a105062a <=( A302  and  (not A301) );
 a105063a <=( a105062a  and  a105059a );
 a105064a <=( a105063a  and  a105056a );
 a105068a <=( (not A167)  and  A168 );
 a105069a <=( A170  and  a105068a );
 a105072a <=( (not A199)  and  A166 );
 a105075a <=( (not A202)  and  (not A200) );
 a105076a <=( a105075a  and  a105072a );
 a105077a <=( a105076a  and  a105069a );
 a105080a <=( A266  and  A265 );
 a105083a <=( (not A268)  and  (not A267) );
 a105084a <=( a105083a  and  a105080a );
 a105087a <=( (not A299)  and  (not A298) );
 a105090a <=( (not A302)  and  A301 );
 a105091a <=( a105090a  and  a105087a );
 a105092a <=( a105091a  and  a105084a );
 a105096a <=( (not A167)  and  A168 );
 a105097a <=( A170  and  a105096a );
 a105100a <=( (not A199)  and  A166 );
 a105103a <=( (not A202)  and  (not A200) );
 a105104a <=( a105103a  and  a105100a );
 a105105a <=( a105104a  and  a105097a );
 a105108a <=( A266  and  A265 );
 a105111a <=( A269  and  (not A267) );
 a105112a <=( a105111a  and  a105108a );
 a105115a <=( A299  and  A298 );
 a105118a <=( (not A302)  and  A301 );
 a105119a <=( a105118a  and  a105115a );
 a105120a <=( a105119a  and  a105112a );
 a105124a <=( (not A167)  and  A168 );
 a105125a <=( A170  and  a105124a );
 a105128a <=( (not A199)  and  A166 );
 a105131a <=( (not A202)  and  (not A200) );
 a105132a <=( a105131a  and  a105128a );
 a105133a <=( a105132a  and  a105125a );
 a105136a <=( A266  and  A265 );
 a105139a <=( A269  and  (not A267) );
 a105140a <=( a105139a  and  a105136a );
 a105143a <=( (not A299)  and  A298 );
 a105146a <=( A302  and  (not A301) );
 a105147a <=( a105146a  and  a105143a );
 a105148a <=( a105147a  and  a105140a );
 a105152a <=( (not A167)  and  A168 );
 a105153a <=( A170  and  a105152a );
 a105156a <=( (not A199)  and  A166 );
 a105159a <=( (not A202)  and  (not A200) );
 a105160a <=( a105159a  and  a105156a );
 a105161a <=( a105160a  and  a105153a );
 a105164a <=( A266  and  A265 );
 a105167a <=( A269  and  (not A267) );
 a105168a <=( a105167a  and  a105164a );
 a105171a <=( A299  and  (not A298) );
 a105174a <=( A302  and  (not A301) );
 a105175a <=( a105174a  and  a105171a );
 a105176a <=( a105175a  and  a105168a );
 a105180a <=( (not A167)  and  A168 );
 a105181a <=( A170  and  a105180a );
 a105184a <=( (not A199)  and  A166 );
 a105187a <=( (not A202)  and  (not A200) );
 a105188a <=( a105187a  and  a105184a );
 a105189a <=( a105188a  and  a105181a );
 a105192a <=( A266  and  A265 );
 a105195a <=( A269  and  (not A267) );
 a105196a <=( a105195a  and  a105192a );
 a105199a <=( (not A299)  and  (not A298) );
 a105202a <=( (not A302)  and  A301 );
 a105203a <=( a105202a  and  a105199a );
 a105204a <=( a105203a  and  a105196a );
 a105208a <=( (not A167)  and  A168 );
 a105209a <=( A170  and  a105208a );
 a105212a <=( (not A199)  and  A166 );
 a105215a <=( (not A202)  and  (not A200) );
 a105216a <=( a105215a  and  a105212a );
 a105217a <=( a105216a  and  a105209a );
 a105220a <=( A266  and  (not A265) );
 a105223a <=( A268  and  (not A267) );
 a105224a <=( a105223a  and  a105220a );
 a105227a <=( A299  and  A298 );
 a105230a <=( (not A302)  and  A301 );
 a105231a <=( a105230a  and  a105227a );
 a105232a <=( a105231a  and  a105224a );
 a105236a <=( (not A167)  and  A168 );
 a105237a <=( A170  and  a105236a );
 a105240a <=( (not A199)  and  A166 );
 a105243a <=( (not A202)  and  (not A200) );
 a105244a <=( a105243a  and  a105240a );
 a105245a <=( a105244a  and  a105237a );
 a105248a <=( A266  and  (not A265) );
 a105251a <=( A268  and  (not A267) );
 a105252a <=( a105251a  and  a105248a );
 a105255a <=( (not A299)  and  A298 );
 a105258a <=( A302  and  (not A301) );
 a105259a <=( a105258a  and  a105255a );
 a105260a <=( a105259a  and  a105252a );
 a105264a <=( (not A167)  and  A168 );
 a105265a <=( A170  and  a105264a );
 a105268a <=( (not A199)  and  A166 );
 a105271a <=( (not A202)  and  (not A200) );
 a105272a <=( a105271a  and  a105268a );
 a105273a <=( a105272a  and  a105265a );
 a105276a <=( A266  and  (not A265) );
 a105279a <=( A268  and  (not A267) );
 a105280a <=( a105279a  and  a105276a );
 a105283a <=( A299  and  (not A298) );
 a105286a <=( A302  and  (not A301) );
 a105287a <=( a105286a  and  a105283a );
 a105288a <=( a105287a  and  a105280a );
 a105292a <=( (not A167)  and  A168 );
 a105293a <=( A170  and  a105292a );
 a105296a <=( (not A199)  and  A166 );
 a105299a <=( (not A202)  and  (not A200) );
 a105300a <=( a105299a  and  a105296a );
 a105301a <=( a105300a  and  a105293a );
 a105304a <=( A266  and  (not A265) );
 a105307a <=( A268  and  (not A267) );
 a105308a <=( a105307a  and  a105304a );
 a105311a <=( (not A299)  and  (not A298) );
 a105314a <=( (not A302)  and  A301 );
 a105315a <=( a105314a  and  a105311a );
 a105316a <=( a105315a  and  a105308a );
 a105320a <=( (not A167)  and  A168 );
 a105321a <=( A170  and  a105320a );
 a105324a <=( (not A199)  and  A166 );
 a105327a <=( (not A202)  and  (not A200) );
 a105328a <=( a105327a  and  a105324a );
 a105329a <=( a105328a  and  a105321a );
 a105332a <=( A266  and  (not A265) );
 a105335a <=( (not A269)  and  (not A267) );
 a105336a <=( a105335a  and  a105332a );
 a105339a <=( A299  and  A298 );
 a105342a <=( (not A302)  and  A301 );
 a105343a <=( a105342a  and  a105339a );
 a105344a <=( a105343a  and  a105336a );
 a105348a <=( (not A167)  and  A168 );
 a105349a <=( A170  and  a105348a );
 a105352a <=( (not A199)  and  A166 );
 a105355a <=( (not A202)  and  (not A200) );
 a105356a <=( a105355a  and  a105352a );
 a105357a <=( a105356a  and  a105349a );
 a105360a <=( A266  and  (not A265) );
 a105363a <=( (not A269)  and  (not A267) );
 a105364a <=( a105363a  and  a105360a );
 a105367a <=( (not A299)  and  A298 );
 a105370a <=( A302  and  (not A301) );
 a105371a <=( a105370a  and  a105367a );
 a105372a <=( a105371a  and  a105364a );
 a105376a <=( (not A167)  and  A168 );
 a105377a <=( A170  and  a105376a );
 a105380a <=( (not A199)  and  A166 );
 a105383a <=( (not A202)  and  (not A200) );
 a105384a <=( a105383a  and  a105380a );
 a105385a <=( a105384a  and  a105377a );
 a105388a <=( A266  and  (not A265) );
 a105391a <=( (not A269)  and  (not A267) );
 a105392a <=( a105391a  and  a105388a );
 a105395a <=( A299  and  (not A298) );
 a105398a <=( A302  and  (not A301) );
 a105399a <=( a105398a  and  a105395a );
 a105400a <=( a105399a  and  a105392a );
 a105404a <=( (not A167)  and  A168 );
 a105405a <=( A170  and  a105404a );
 a105408a <=( (not A199)  and  A166 );
 a105411a <=( (not A202)  and  (not A200) );
 a105412a <=( a105411a  and  a105408a );
 a105413a <=( a105412a  and  a105405a );
 a105416a <=( A266  and  (not A265) );
 a105419a <=( (not A269)  and  (not A267) );
 a105420a <=( a105419a  and  a105416a );
 a105423a <=( (not A299)  and  (not A298) );
 a105426a <=( (not A302)  and  A301 );
 a105427a <=( a105426a  and  a105423a );
 a105428a <=( a105427a  and  a105420a );
 a105432a <=( (not A167)  and  A168 );
 a105433a <=( A170  and  a105432a );
 a105436a <=( (not A199)  and  A166 );
 a105439a <=( (not A202)  and  (not A200) );
 a105440a <=( a105439a  and  a105436a );
 a105441a <=( a105440a  and  a105433a );
 a105444a <=( (not A266)  and  A265 );
 a105447a <=( A268  and  (not A267) );
 a105448a <=( a105447a  and  a105444a );
 a105451a <=( A299  and  A298 );
 a105454a <=( (not A302)  and  A301 );
 a105455a <=( a105454a  and  a105451a );
 a105456a <=( a105455a  and  a105448a );
 a105460a <=( (not A167)  and  A168 );
 a105461a <=( A170  and  a105460a );
 a105464a <=( (not A199)  and  A166 );
 a105467a <=( (not A202)  and  (not A200) );
 a105468a <=( a105467a  and  a105464a );
 a105469a <=( a105468a  and  a105461a );
 a105472a <=( (not A266)  and  A265 );
 a105475a <=( A268  and  (not A267) );
 a105476a <=( a105475a  and  a105472a );
 a105479a <=( (not A299)  and  A298 );
 a105482a <=( A302  and  (not A301) );
 a105483a <=( a105482a  and  a105479a );
 a105484a <=( a105483a  and  a105476a );
 a105488a <=( (not A167)  and  A168 );
 a105489a <=( A170  and  a105488a );
 a105492a <=( (not A199)  and  A166 );
 a105495a <=( (not A202)  and  (not A200) );
 a105496a <=( a105495a  and  a105492a );
 a105497a <=( a105496a  and  a105489a );
 a105500a <=( (not A266)  and  A265 );
 a105503a <=( A268  and  (not A267) );
 a105504a <=( a105503a  and  a105500a );
 a105507a <=( A299  and  (not A298) );
 a105510a <=( A302  and  (not A301) );
 a105511a <=( a105510a  and  a105507a );
 a105512a <=( a105511a  and  a105504a );
 a105516a <=( (not A167)  and  A168 );
 a105517a <=( A170  and  a105516a );
 a105520a <=( (not A199)  and  A166 );
 a105523a <=( (not A202)  and  (not A200) );
 a105524a <=( a105523a  and  a105520a );
 a105525a <=( a105524a  and  a105517a );
 a105528a <=( (not A266)  and  A265 );
 a105531a <=( A268  and  (not A267) );
 a105532a <=( a105531a  and  a105528a );
 a105535a <=( (not A299)  and  (not A298) );
 a105538a <=( (not A302)  and  A301 );
 a105539a <=( a105538a  and  a105535a );
 a105540a <=( a105539a  and  a105532a );
 a105544a <=( (not A167)  and  A168 );
 a105545a <=( A170  and  a105544a );
 a105548a <=( (not A199)  and  A166 );
 a105551a <=( (not A202)  and  (not A200) );
 a105552a <=( a105551a  and  a105548a );
 a105553a <=( a105552a  and  a105545a );
 a105556a <=( (not A266)  and  A265 );
 a105559a <=( (not A269)  and  (not A267) );
 a105560a <=( a105559a  and  a105556a );
 a105563a <=( A299  and  A298 );
 a105566a <=( (not A302)  and  A301 );
 a105567a <=( a105566a  and  a105563a );
 a105568a <=( a105567a  and  a105560a );
 a105572a <=( (not A167)  and  A168 );
 a105573a <=( A170  and  a105572a );
 a105576a <=( (not A199)  and  A166 );
 a105579a <=( (not A202)  and  (not A200) );
 a105580a <=( a105579a  and  a105576a );
 a105581a <=( a105580a  and  a105573a );
 a105584a <=( (not A266)  and  A265 );
 a105587a <=( (not A269)  and  (not A267) );
 a105588a <=( a105587a  and  a105584a );
 a105591a <=( (not A299)  and  A298 );
 a105594a <=( A302  and  (not A301) );
 a105595a <=( a105594a  and  a105591a );
 a105596a <=( a105595a  and  a105588a );
 a105600a <=( (not A167)  and  A168 );
 a105601a <=( A170  and  a105600a );
 a105604a <=( (not A199)  and  A166 );
 a105607a <=( (not A202)  and  (not A200) );
 a105608a <=( a105607a  and  a105604a );
 a105609a <=( a105608a  and  a105601a );
 a105612a <=( (not A266)  and  A265 );
 a105615a <=( (not A269)  and  (not A267) );
 a105616a <=( a105615a  and  a105612a );
 a105619a <=( A299  and  (not A298) );
 a105622a <=( A302  and  (not A301) );
 a105623a <=( a105622a  and  a105619a );
 a105624a <=( a105623a  and  a105616a );
 a105628a <=( (not A167)  and  A168 );
 a105629a <=( A170  and  a105628a );
 a105632a <=( (not A199)  and  A166 );
 a105635a <=( (not A202)  and  (not A200) );
 a105636a <=( a105635a  and  a105632a );
 a105637a <=( a105636a  and  a105629a );
 a105640a <=( (not A266)  and  A265 );
 a105643a <=( (not A269)  and  (not A267) );
 a105644a <=( a105643a  and  a105640a );
 a105647a <=( (not A299)  and  (not A298) );
 a105650a <=( (not A302)  and  A301 );
 a105651a <=( a105650a  and  a105647a );
 a105652a <=( a105651a  and  a105644a );
 a105656a <=( (not A167)  and  A168 );
 a105657a <=( A170  and  a105656a );
 a105660a <=( (not A199)  and  A166 );
 a105663a <=( A203  and  (not A200) );
 a105664a <=( a105663a  and  a105660a );
 a105665a <=( a105664a  and  a105657a );
 a105668a <=( A266  and  A265 );
 a105671a <=( (not A268)  and  (not A267) );
 a105672a <=( a105671a  and  a105668a );
 a105675a <=( A299  and  A298 );
 a105678a <=( (not A302)  and  A301 );
 a105679a <=( a105678a  and  a105675a );
 a105680a <=( a105679a  and  a105672a );
 a105684a <=( (not A167)  and  A168 );
 a105685a <=( A170  and  a105684a );
 a105688a <=( (not A199)  and  A166 );
 a105691a <=( A203  and  (not A200) );
 a105692a <=( a105691a  and  a105688a );
 a105693a <=( a105692a  and  a105685a );
 a105696a <=( A266  and  A265 );
 a105699a <=( (not A268)  and  (not A267) );
 a105700a <=( a105699a  and  a105696a );
 a105703a <=( (not A299)  and  A298 );
 a105706a <=( A302  and  (not A301) );
 a105707a <=( a105706a  and  a105703a );
 a105708a <=( a105707a  and  a105700a );
 a105712a <=( (not A167)  and  A168 );
 a105713a <=( A170  and  a105712a );
 a105716a <=( (not A199)  and  A166 );
 a105719a <=( A203  and  (not A200) );
 a105720a <=( a105719a  and  a105716a );
 a105721a <=( a105720a  and  a105713a );
 a105724a <=( A266  and  A265 );
 a105727a <=( (not A268)  and  (not A267) );
 a105728a <=( a105727a  and  a105724a );
 a105731a <=( A299  and  (not A298) );
 a105734a <=( A302  and  (not A301) );
 a105735a <=( a105734a  and  a105731a );
 a105736a <=( a105735a  and  a105728a );
 a105740a <=( (not A167)  and  A168 );
 a105741a <=( A170  and  a105740a );
 a105744a <=( (not A199)  and  A166 );
 a105747a <=( A203  and  (not A200) );
 a105748a <=( a105747a  and  a105744a );
 a105749a <=( a105748a  and  a105741a );
 a105752a <=( A266  and  A265 );
 a105755a <=( (not A268)  and  (not A267) );
 a105756a <=( a105755a  and  a105752a );
 a105759a <=( (not A299)  and  (not A298) );
 a105762a <=( (not A302)  and  A301 );
 a105763a <=( a105762a  and  a105759a );
 a105764a <=( a105763a  and  a105756a );
 a105768a <=( (not A167)  and  A168 );
 a105769a <=( A170  and  a105768a );
 a105772a <=( (not A199)  and  A166 );
 a105775a <=( A203  and  (not A200) );
 a105776a <=( a105775a  and  a105772a );
 a105777a <=( a105776a  and  a105769a );
 a105780a <=( A266  and  A265 );
 a105783a <=( A269  and  (not A267) );
 a105784a <=( a105783a  and  a105780a );
 a105787a <=( A299  and  A298 );
 a105790a <=( (not A302)  and  A301 );
 a105791a <=( a105790a  and  a105787a );
 a105792a <=( a105791a  and  a105784a );
 a105796a <=( (not A167)  and  A168 );
 a105797a <=( A170  and  a105796a );
 a105800a <=( (not A199)  and  A166 );
 a105803a <=( A203  and  (not A200) );
 a105804a <=( a105803a  and  a105800a );
 a105805a <=( a105804a  and  a105797a );
 a105808a <=( A266  and  A265 );
 a105811a <=( A269  and  (not A267) );
 a105812a <=( a105811a  and  a105808a );
 a105815a <=( (not A299)  and  A298 );
 a105818a <=( A302  and  (not A301) );
 a105819a <=( a105818a  and  a105815a );
 a105820a <=( a105819a  and  a105812a );
 a105824a <=( (not A167)  and  A168 );
 a105825a <=( A170  and  a105824a );
 a105828a <=( (not A199)  and  A166 );
 a105831a <=( A203  and  (not A200) );
 a105832a <=( a105831a  and  a105828a );
 a105833a <=( a105832a  and  a105825a );
 a105836a <=( A266  and  A265 );
 a105839a <=( A269  and  (not A267) );
 a105840a <=( a105839a  and  a105836a );
 a105843a <=( A299  and  (not A298) );
 a105846a <=( A302  and  (not A301) );
 a105847a <=( a105846a  and  a105843a );
 a105848a <=( a105847a  and  a105840a );
 a105852a <=( (not A167)  and  A168 );
 a105853a <=( A170  and  a105852a );
 a105856a <=( (not A199)  and  A166 );
 a105859a <=( A203  and  (not A200) );
 a105860a <=( a105859a  and  a105856a );
 a105861a <=( a105860a  and  a105853a );
 a105864a <=( A266  and  A265 );
 a105867a <=( A269  and  (not A267) );
 a105868a <=( a105867a  and  a105864a );
 a105871a <=( (not A299)  and  (not A298) );
 a105874a <=( (not A302)  and  A301 );
 a105875a <=( a105874a  and  a105871a );
 a105876a <=( a105875a  and  a105868a );
 a105880a <=( (not A167)  and  A168 );
 a105881a <=( A170  and  a105880a );
 a105884a <=( (not A199)  and  A166 );
 a105887a <=( A203  and  (not A200) );
 a105888a <=( a105887a  and  a105884a );
 a105889a <=( a105888a  and  a105881a );
 a105892a <=( A266  and  (not A265) );
 a105895a <=( A268  and  (not A267) );
 a105896a <=( a105895a  and  a105892a );
 a105899a <=( A299  and  A298 );
 a105902a <=( (not A302)  and  A301 );
 a105903a <=( a105902a  and  a105899a );
 a105904a <=( a105903a  and  a105896a );
 a105908a <=( (not A167)  and  A168 );
 a105909a <=( A170  and  a105908a );
 a105912a <=( (not A199)  and  A166 );
 a105915a <=( A203  and  (not A200) );
 a105916a <=( a105915a  and  a105912a );
 a105917a <=( a105916a  and  a105909a );
 a105920a <=( A266  and  (not A265) );
 a105923a <=( A268  and  (not A267) );
 a105924a <=( a105923a  and  a105920a );
 a105927a <=( (not A299)  and  A298 );
 a105930a <=( A302  and  (not A301) );
 a105931a <=( a105930a  and  a105927a );
 a105932a <=( a105931a  and  a105924a );
 a105936a <=( (not A167)  and  A168 );
 a105937a <=( A170  and  a105936a );
 a105940a <=( (not A199)  and  A166 );
 a105943a <=( A203  and  (not A200) );
 a105944a <=( a105943a  and  a105940a );
 a105945a <=( a105944a  and  a105937a );
 a105948a <=( A266  and  (not A265) );
 a105951a <=( A268  and  (not A267) );
 a105952a <=( a105951a  and  a105948a );
 a105955a <=( A299  and  (not A298) );
 a105958a <=( A302  and  (not A301) );
 a105959a <=( a105958a  and  a105955a );
 a105960a <=( a105959a  and  a105952a );
 a105964a <=( (not A167)  and  A168 );
 a105965a <=( A170  and  a105964a );
 a105968a <=( (not A199)  and  A166 );
 a105971a <=( A203  and  (not A200) );
 a105972a <=( a105971a  and  a105968a );
 a105973a <=( a105972a  and  a105965a );
 a105976a <=( A266  and  (not A265) );
 a105979a <=( A268  and  (not A267) );
 a105980a <=( a105979a  and  a105976a );
 a105983a <=( (not A299)  and  (not A298) );
 a105986a <=( (not A302)  and  A301 );
 a105987a <=( a105986a  and  a105983a );
 a105988a <=( a105987a  and  a105980a );
 a105992a <=( (not A167)  and  A168 );
 a105993a <=( A170  and  a105992a );
 a105996a <=( (not A199)  and  A166 );
 a105999a <=( A203  and  (not A200) );
 a106000a <=( a105999a  and  a105996a );
 a106001a <=( a106000a  and  a105993a );
 a106004a <=( A266  and  (not A265) );
 a106007a <=( (not A269)  and  (not A267) );
 a106008a <=( a106007a  and  a106004a );
 a106011a <=( A299  and  A298 );
 a106014a <=( (not A302)  and  A301 );
 a106015a <=( a106014a  and  a106011a );
 a106016a <=( a106015a  and  a106008a );
 a106020a <=( (not A167)  and  A168 );
 a106021a <=( A170  and  a106020a );
 a106024a <=( (not A199)  and  A166 );
 a106027a <=( A203  and  (not A200) );
 a106028a <=( a106027a  and  a106024a );
 a106029a <=( a106028a  and  a106021a );
 a106032a <=( A266  and  (not A265) );
 a106035a <=( (not A269)  and  (not A267) );
 a106036a <=( a106035a  and  a106032a );
 a106039a <=( (not A299)  and  A298 );
 a106042a <=( A302  and  (not A301) );
 a106043a <=( a106042a  and  a106039a );
 a106044a <=( a106043a  and  a106036a );
 a106048a <=( (not A167)  and  A168 );
 a106049a <=( A170  and  a106048a );
 a106052a <=( (not A199)  and  A166 );
 a106055a <=( A203  and  (not A200) );
 a106056a <=( a106055a  and  a106052a );
 a106057a <=( a106056a  and  a106049a );
 a106060a <=( A266  and  (not A265) );
 a106063a <=( (not A269)  and  (not A267) );
 a106064a <=( a106063a  and  a106060a );
 a106067a <=( A299  and  (not A298) );
 a106070a <=( A302  and  (not A301) );
 a106071a <=( a106070a  and  a106067a );
 a106072a <=( a106071a  and  a106064a );
 a106076a <=( (not A167)  and  A168 );
 a106077a <=( A170  and  a106076a );
 a106080a <=( (not A199)  and  A166 );
 a106083a <=( A203  and  (not A200) );
 a106084a <=( a106083a  and  a106080a );
 a106085a <=( a106084a  and  a106077a );
 a106088a <=( A266  and  (not A265) );
 a106091a <=( (not A269)  and  (not A267) );
 a106092a <=( a106091a  and  a106088a );
 a106095a <=( (not A299)  and  (not A298) );
 a106098a <=( (not A302)  and  A301 );
 a106099a <=( a106098a  and  a106095a );
 a106100a <=( a106099a  and  a106092a );
 a106104a <=( (not A167)  and  A168 );
 a106105a <=( A170  and  a106104a );
 a106108a <=( (not A199)  and  A166 );
 a106111a <=( A203  and  (not A200) );
 a106112a <=( a106111a  and  a106108a );
 a106113a <=( a106112a  and  a106105a );
 a106116a <=( (not A266)  and  A265 );
 a106119a <=( A268  and  (not A267) );
 a106120a <=( a106119a  and  a106116a );
 a106123a <=( A299  and  A298 );
 a106126a <=( (not A302)  and  A301 );
 a106127a <=( a106126a  and  a106123a );
 a106128a <=( a106127a  and  a106120a );
 a106132a <=( (not A167)  and  A168 );
 a106133a <=( A170  and  a106132a );
 a106136a <=( (not A199)  and  A166 );
 a106139a <=( A203  and  (not A200) );
 a106140a <=( a106139a  and  a106136a );
 a106141a <=( a106140a  and  a106133a );
 a106144a <=( (not A266)  and  A265 );
 a106147a <=( A268  and  (not A267) );
 a106148a <=( a106147a  and  a106144a );
 a106151a <=( (not A299)  and  A298 );
 a106154a <=( A302  and  (not A301) );
 a106155a <=( a106154a  and  a106151a );
 a106156a <=( a106155a  and  a106148a );
 a106160a <=( (not A167)  and  A168 );
 a106161a <=( A170  and  a106160a );
 a106164a <=( (not A199)  and  A166 );
 a106167a <=( A203  and  (not A200) );
 a106168a <=( a106167a  and  a106164a );
 a106169a <=( a106168a  and  a106161a );
 a106172a <=( (not A266)  and  A265 );
 a106175a <=( A268  and  (not A267) );
 a106176a <=( a106175a  and  a106172a );
 a106179a <=( A299  and  (not A298) );
 a106182a <=( A302  and  (not A301) );
 a106183a <=( a106182a  and  a106179a );
 a106184a <=( a106183a  and  a106176a );
 a106188a <=( (not A167)  and  A168 );
 a106189a <=( A170  and  a106188a );
 a106192a <=( (not A199)  and  A166 );
 a106195a <=( A203  and  (not A200) );
 a106196a <=( a106195a  and  a106192a );
 a106197a <=( a106196a  and  a106189a );
 a106200a <=( (not A266)  and  A265 );
 a106203a <=( A268  and  (not A267) );
 a106204a <=( a106203a  and  a106200a );
 a106207a <=( (not A299)  and  (not A298) );
 a106210a <=( (not A302)  and  A301 );
 a106211a <=( a106210a  and  a106207a );
 a106212a <=( a106211a  and  a106204a );
 a106216a <=( (not A167)  and  A168 );
 a106217a <=( A170  and  a106216a );
 a106220a <=( (not A199)  and  A166 );
 a106223a <=( A203  and  (not A200) );
 a106224a <=( a106223a  and  a106220a );
 a106225a <=( a106224a  and  a106217a );
 a106228a <=( (not A266)  and  A265 );
 a106231a <=( (not A269)  and  (not A267) );
 a106232a <=( a106231a  and  a106228a );
 a106235a <=( A299  and  A298 );
 a106238a <=( (not A302)  and  A301 );
 a106239a <=( a106238a  and  a106235a );
 a106240a <=( a106239a  and  a106232a );
 a106244a <=( (not A167)  and  A168 );
 a106245a <=( A170  and  a106244a );
 a106248a <=( (not A199)  and  A166 );
 a106251a <=( A203  and  (not A200) );
 a106252a <=( a106251a  and  a106248a );
 a106253a <=( a106252a  and  a106245a );
 a106256a <=( (not A266)  and  A265 );
 a106259a <=( (not A269)  and  (not A267) );
 a106260a <=( a106259a  and  a106256a );
 a106263a <=( (not A299)  and  A298 );
 a106266a <=( A302  and  (not A301) );
 a106267a <=( a106266a  and  a106263a );
 a106268a <=( a106267a  and  a106260a );
 a106272a <=( (not A167)  and  A168 );
 a106273a <=( A170  and  a106272a );
 a106276a <=( (not A199)  and  A166 );
 a106279a <=( A203  and  (not A200) );
 a106280a <=( a106279a  and  a106276a );
 a106281a <=( a106280a  and  a106273a );
 a106284a <=( (not A266)  and  A265 );
 a106287a <=( (not A269)  and  (not A267) );
 a106288a <=( a106287a  and  a106284a );
 a106291a <=( A299  and  (not A298) );
 a106294a <=( A302  and  (not A301) );
 a106295a <=( a106294a  and  a106291a );
 a106296a <=( a106295a  and  a106288a );
 a106300a <=( (not A167)  and  A168 );
 a106301a <=( A170  and  a106300a );
 a106304a <=( (not A199)  and  A166 );
 a106307a <=( A203  and  (not A200) );
 a106308a <=( a106307a  and  a106304a );
 a106309a <=( a106308a  and  a106301a );
 a106312a <=( (not A266)  and  A265 );
 a106315a <=( (not A269)  and  (not A267) );
 a106316a <=( a106315a  and  a106312a );
 a106319a <=( (not A299)  and  (not A298) );
 a106322a <=( (not A302)  and  A301 );
 a106323a <=( a106322a  and  a106319a );
 a106324a <=( a106323a  and  a106316a );
 a106328a <=( (not A167)  and  A168 );
 a106329a <=( A170  and  a106328a );
 a106332a <=( (not A199)  and  A166 );
 a106335a <=( A202  and  (not A200) );
 a106336a <=( a106335a  and  a106332a );
 a106337a <=( a106336a  and  a106329a );
 a106340a <=( A265  and  (not A203) );
 a106343a <=( A268  and  A266 );
 a106344a <=( a106343a  and  a106340a );
 a106347a <=( (not A298)  and  (not A269) );
 a106350a <=( (not A301)  and  (not A299) );
 a106351a <=( a106350a  and  a106347a );
 a106352a <=( a106351a  and  a106344a );
 a106356a <=( (not A167)  and  A168 );
 a106357a <=( A170  and  a106356a );
 a106360a <=( (not A199)  and  A166 );
 a106363a <=( A202  and  (not A200) );
 a106364a <=( a106363a  and  a106360a );
 a106365a <=( a106364a  and  a106357a );
 a106368a <=( A265  and  (not A203) );
 a106371a <=( A268  and  A266 );
 a106372a <=( a106371a  and  a106368a );
 a106375a <=( (not A298)  and  (not A269) );
 a106378a <=( A302  and  (not A299) );
 a106379a <=( a106378a  and  a106375a );
 a106380a <=( a106379a  and  a106372a );
 a106384a <=( (not A167)  and  A168 );
 a106385a <=( A170  and  a106384a );
 a106388a <=( (not A199)  and  A166 );
 a106391a <=( A202  and  (not A200) );
 a106392a <=( a106391a  and  a106388a );
 a106393a <=( a106392a  and  a106385a );
 a106396a <=( (not A265)  and  (not A203) );
 a106399a <=( (not A268)  and  A266 );
 a106400a <=( a106399a  and  a106396a );
 a106403a <=( (not A298)  and  A269 );
 a106406a <=( (not A301)  and  (not A299) );
 a106407a <=( a106406a  and  a106403a );
 a106408a <=( a106407a  and  a106400a );
 a106412a <=( (not A167)  and  A168 );
 a106413a <=( A170  and  a106412a );
 a106416a <=( (not A199)  and  A166 );
 a106419a <=( A202  and  (not A200) );
 a106420a <=( a106419a  and  a106416a );
 a106421a <=( a106420a  and  a106413a );
 a106424a <=( (not A265)  and  (not A203) );
 a106427a <=( (not A268)  and  A266 );
 a106428a <=( a106427a  and  a106424a );
 a106431a <=( (not A298)  and  A269 );
 a106434a <=( A302  and  (not A299) );
 a106435a <=( a106434a  and  a106431a );
 a106436a <=( a106435a  and  a106428a );
 a106440a <=( (not A167)  and  A168 );
 a106441a <=( A170  and  a106440a );
 a106444a <=( (not A199)  and  A166 );
 a106447a <=( A202  and  (not A200) );
 a106448a <=( a106447a  and  a106444a );
 a106449a <=( a106448a  and  a106441a );
 a106452a <=( A265  and  (not A203) );
 a106455a <=( (not A268)  and  (not A266) );
 a106456a <=( a106455a  and  a106452a );
 a106459a <=( (not A298)  and  A269 );
 a106462a <=( (not A301)  and  (not A299) );
 a106463a <=( a106462a  and  a106459a );
 a106464a <=( a106463a  and  a106456a );
 a106468a <=( (not A167)  and  A168 );
 a106469a <=( A170  and  a106468a );
 a106472a <=( (not A199)  and  A166 );
 a106475a <=( A202  and  (not A200) );
 a106476a <=( a106475a  and  a106472a );
 a106477a <=( a106476a  and  a106469a );
 a106480a <=( A265  and  (not A203) );
 a106483a <=( (not A268)  and  (not A266) );
 a106484a <=( a106483a  and  a106480a );
 a106487a <=( (not A298)  and  A269 );
 a106490a <=( A302  and  (not A299) );
 a106491a <=( a106490a  and  a106487a );
 a106492a <=( a106491a  and  a106484a );
 a106496a <=( (not A167)  and  A168 );
 a106497a <=( A170  and  a106496a );
 a106500a <=( (not A199)  and  A166 );
 a106503a <=( A202  and  (not A200) );
 a106504a <=( a106503a  and  a106500a );
 a106505a <=( a106504a  and  a106497a );
 a106508a <=( (not A265)  and  (not A203) );
 a106511a <=( A268  and  (not A266) );
 a106512a <=( a106511a  and  a106508a );
 a106515a <=( (not A298)  and  (not A269) );
 a106518a <=( (not A301)  and  (not A299) );
 a106519a <=( a106518a  and  a106515a );
 a106520a <=( a106519a  and  a106512a );
 a106524a <=( (not A167)  and  A168 );
 a106525a <=( A170  and  a106524a );
 a106528a <=( (not A199)  and  A166 );
 a106531a <=( A202  and  (not A200) );
 a106532a <=( a106531a  and  a106528a );
 a106533a <=( a106532a  and  a106525a );
 a106536a <=( (not A265)  and  (not A203) );
 a106539a <=( A268  and  (not A266) );
 a106540a <=( a106539a  and  a106536a );
 a106543a <=( (not A298)  and  (not A269) );
 a106546a <=( A302  and  (not A299) );
 a106547a <=( a106546a  and  a106543a );
 a106548a <=( a106547a  and  a106540a );
 a106552a <=( (not A167)  and  A168 );
 a106553a <=( A169  and  a106552a );
 a106556a <=( A199  and  A166 );
 a106559a <=( A202  and  A200 );
 a106560a <=( a106559a  and  a106556a );
 a106561a <=( a106560a  and  a106553a );
 a106564a <=( A265  and  (not A203) );
 a106567a <=( A268  and  A266 );
 a106568a <=( a106567a  and  a106564a );
 a106571a <=( (not A298)  and  (not A269) );
 a106574a <=( (not A301)  and  (not A299) );
 a106575a <=( a106574a  and  a106571a );
 a106576a <=( a106575a  and  a106568a );
 a106580a <=( (not A167)  and  A168 );
 a106581a <=( A169  and  a106580a );
 a106584a <=( A199  and  A166 );
 a106587a <=( A202  and  A200 );
 a106588a <=( a106587a  and  a106584a );
 a106589a <=( a106588a  and  a106581a );
 a106592a <=( A265  and  (not A203) );
 a106595a <=( A268  and  A266 );
 a106596a <=( a106595a  and  a106592a );
 a106599a <=( (not A298)  and  (not A269) );
 a106602a <=( A302  and  (not A299) );
 a106603a <=( a106602a  and  a106599a );
 a106604a <=( a106603a  and  a106596a );
 a106608a <=( (not A167)  and  A168 );
 a106609a <=( A169  and  a106608a );
 a106612a <=( A199  and  A166 );
 a106615a <=( A202  and  A200 );
 a106616a <=( a106615a  and  a106612a );
 a106617a <=( a106616a  and  a106609a );
 a106620a <=( (not A265)  and  (not A203) );
 a106623a <=( (not A268)  and  A266 );
 a106624a <=( a106623a  and  a106620a );
 a106627a <=( (not A298)  and  A269 );
 a106630a <=( (not A301)  and  (not A299) );
 a106631a <=( a106630a  and  a106627a );
 a106632a <=( a106631a  and  a106624a );
 a106636a <=( (not A167)  and  A168 );
 a106637a <=( A169  and  a106636a );
 a106640a <=( A199  and  A166 );
 a106643a <=( A202  and  A200 );
 a106644a <=( a106643a  and  a106640a );
 a106645a <=( a106644a  and  a106637a );
 a106648a <=( (not A265)  and  (not A203) );
 a106651a <=( (not A268)  and  A266 );
 a106652a <=( a106651a  and  a106648a );
 a106655a <=( (not A298)  and  A269 );
 a106658a <=( A302  and  (not A299) );
 a106659a <=( a106658a  and  a106655a );
 a106660a <=( a106659a  and  a106652a );
 a106664a <=( (not A167)  and  A168 );
 a106665a <=( A169  and  a106664a );
 a106668a <=( A199  and  A166 );
 a106671a <=( A202  and  A200 );
 a106672a <=( a106671a  and  a106668a );
 a106673a <=( a106672a  and  a106665a );
 a106676a <=( A265  and  (not A203) );
 a106679a <=( (not A268)  and  (not A266) );
 a106680a <=( a106679a  and  a106676a );
 a106683a <=( (not A298)  and  A269 );
 a106686a <=( (not A301)  and  (not A299) );
 a106687a <=( a106686a  and  a106683a );
 a106688a <=( a106687a  and  a106680a );
 a106692a <=( (not A167)  and  A168 );
 a106693a <=( A169  and  a106692a );
 a106696a <=( A199  and  A166 );
 a106699a <=( A202  and  A200 );
 a106700a <=( a106699a  and  a106696a );
 a106701a <=( a106700a  and  a106693a );
 a106704a <=( A265  and  (not A203) );
 a106707a <=( (not A268)  and  (not A266) );
 a106708a <=( a106707a  and  a106704a );
 a106711a <=( (not A298)  and  A269 );
 a106714a <=( A302  and  (not A299) );
 a106715a <=( a106714a  and  a106711a );
 a106716a <=( a106715a  and  a106708a );
 a106720a <=( (not A167)  and  A168 );
 a106721a <=( A169  and  a106720a );
 a106724a <=( A199  and  A166 );
 a106727a <=( A202  and  A200 );
 a106728a <=( a106727a  and  a106724a );
 a106729a <=( a106728a  and  a106721a );
 a106732a <=( (not A265)  and  (not A203) );
 a106735a <=( A268  and  (not A266) );
 a106736a <=( a106735a  and  a106732a );
 a106739a <=( (not A298)  and  (not A269) );
 a106742a <=( (not A301)  and  (not A299) );
 a106743a <=( a106742a  and  a106739a );
 a106744a <=( a106743a  and  a106736a );
 a106748a <=( (not A167)  and  A168 );
 a106749a <=( A169  and  a106748a );
 a106752a <=( A199  and  A166 );
 a106755a <=( A202  and  A200 );
 a106756a <=( a106755a  and  a106752a );
 a106757a <=( a106756a  and  a106749a );
 a106760a <=( (not A265)  and  (not A203) );
 a106763a <=( A268  and  (not A266) );
 a106764a <=( a106763a  and  a106760a );
 a106767a <=( (not A298)  and  (not A269) );
 a106770a <=( A302  and  (not A299) );
 a106771a <=( a106770a  and  a106767a );
 a106772a <=( a106771a  and  a106764a );
 a106776a <=( (not A167)  and  A168 );
 a106777a <=( A169  and  a106776a );
 a106780a <=( A199  and  A166 );
 a106783a <=( (not A201)  and  A200 );
 a106784a <=( a106783a  and  a106780a );
 a106785a <=( a106784a  and  a106777a );
 a106788a <=( (not A265)  and  (not A202) );
 a106791a <=( (not A268)  and  (not A266) );
 a106792a <=( a106791a  and  a106788a );
 a106795a <=( A299  and  A298 );
 a106798a <=( (not A302)  and  A301 );
 a106799a <=( a106798a  and  a106795a );
 a106800a <=( a106799a  and  a106792a );
 a106804a <=( (not A167)  and  A168 );
 a106805a <=( A169  and  a106804a );
 a106808a <=( A199  and  A166 );
 a106811a <=( (not A201)  and  A200 );
 a106812a <=( a106811a  and  a106808a );
 a106813a <=( a106812a  and  a106805a );
 a106816a <=( (not A265)  and  (not A202) );
 a106819a <=( (not A268)  and  (not A266) );
 a106820a <=( a106819a  and  a106816a );
 a106823a <=( (not A299)  and  A298 );
 a106826a <=( A302  and  (not A301) );
 a106827a <=( a106826a  and  a106823a );
 a106828a <=( a106827a  and  a106820a );
 a106832a <=( (not A167)  and  A168 );
 a106833a <=( A169  and  a106832a );
 a106836a <=( A199  and  A166 );
 a106839a <=( (not A201)  and  A200 );
 a106840a <=( a106839a  and  a106836a );
 a106841a <=( a106840a  and  a106833a );
 a106844a <=( (not A265)  and  (not A202) );
 a106847a <=( (not A268)  and  (not A266) );
 a106848a <=( a106847a  and  a106844a );
 a106851a <=( A299  and  (not A298) );
 a106854a <=( A302  and  (not A301) );
 a106855a <=( a106854a  and  a106851a );
 a106856a <=( a106855a  and  a106848a );
 a106860a <=( (not A167)  and  A168 );
 a106861a <=( A169  and  a106860a );
 a106864a <=( A199  and  A166 );
 a106867a <=( (not A201)  and  A200 );
 a106868a <=( a106867a  and  a106864a );
 a106869a <=( a106868a  and  a106861a );
 a106872a <=( (not A265)  and  (not A202) );
 a106875a <=( (not A268)  and  (not A266) );
 a106876a <=( a106875a  and  a106872a );
 a106879a <=( (not A299)  and  (not A298) );
 a106882a <=( (not A302)  and  A301 );
 a106883a <=( a106882a  and  a106879a );
 a106884a <=( a106883a  and  a106876a );
 a106888a <=( (not A167)  and  A168 );
 a106889a <=( A169  and  a106888a );
 a106892a <=( A199  and  A166 );
 a106895a <=( (not A201)  and  A200 );
 a106896a <=( a106895a  and  a106892a );
 a106897a <=( a106896a  and  a106889a );
 a106900a <=( (not A265)  and  (not A202) );
 a106903a <=( A269  and  (not A266) );
 a106904a <=( a106903a  and  a106900a );
 a106907a <=( A299  and  A298 );
 a106910a <=( (not A302)  and  A301 );
 a106911a <=( a106910a  and  a106907a );
 a106912a <=( a106911a  and  a106904a );
 a106916a <=( (not A167)  and  A168 );
 a106917a <=( A169  and  a106916a );
 a106920a <=( A199  and  A166 );
 a106923a <=( (not A201)  and  A200 );
 a106924a <=( a106923a  and  a106920a );
 a106925a <=( a106924a  and  a106917a );
 a106928a <=( (not A265)  and  (not A202) );
 a106931a <=( A269  and  (not A266) );
 a106932a <=( a106931a  and  a106928a );
 a106935a <=( (not A299)  and  A298 );
 a106938a <=( A302  and  (not A301) );
 a106939a <=( a106938a  and  a106935a );
 a106940a <=( a106939a  and  a106932a );
 a106944a <=( (not A167)  and  A168 );
 a106945a <=( A169  and  a106944a );
 a106948a <=( A199  and  A166 );
 a106951a <=( (not A201)  and  A200 );
 a106952a <=( a106951a  and  a106948a );
 a106953a <=( a106952a  and  a106945a );
 a106956a <=( (not A265)  and  (not A202) );
 a106959a <=( A269  and  (not A266) );
 a106960a <=( a106959a  and  a106956a );
 a106963a <=( A299  and  (not A298) );
 a106966a <=( A302  and  (not A301) );
 a106967a <=( a106966a  and  a106963a );
 a106968a <=( a106967a  and  a106960a );
 a106972a <=( (not A167)  and  A168 );
 a106973a <=( A169  and  a106972a );
 a106976a <=( A199  and  A166 );
 a106979a <=( (not A201)  and  A200 );
 a106980a <=( a106979a  and  a106976a );
 a106981a <=( a106980a  and  a106973a );
 a106984a <=( (not A265)  and  (not A202) );
 a106987a <=( A269  and  (not A266) );
 a106988a <=( a106987a  and  a106984a );
 a106991a <=( (not A299)  and  (not A298) );
 a106994a <=( (not A302)  and  A301 );
 a106995a <=( a106994a  and  a106991a );
 a106996a <=( a106995a  and  a106988a );
 a107000a <=( (not A167)  and  A168 );
 a107001a <=( A169  and  a107000a );
 a107004a <=( A199  and  A166 );
 a107007a <=( (not A201)  and  A200 );
 a107008a <=( a107007a  and  a107004a );
 a107009a <=( a107008a  and  a107001a );
 a107012a <=( (not A265)  and  A203 );
 a107015a <=( (not A268)  and  (not A266) );
 a107016a <=( a107015a  and  a107012a );
 a107019a <=( A299  and  A298 );
 a107022a <=( (not A302)  and  A301 );
 a107023a <=( a107022a  and  a107019a );
 a107024a <=( a107023a  and  a107016a );
 a107028a <=( (not A167)  and  A168 );
 a107029a <=( A169  and  a107028a );
 a107032a <=( A199  and  A166 );
 a107035a <=( (not A201)  and  A200 );
 a107036a <=( a107035a  and  a107032a );
 a107037a <=( a107036a  and  a107029a );
 a107040a <=( (not A265)  and  A203 );
 a107043a <=( (not A268)  and  (not A266) );
 a107044a <=( a107043a  and  a107040a );
 a107047a <=( (not A299)  and  A298 );
 a107050a <=( A302  and  (not A301) );
 a107051a <=( a107050a  and  a107047a );
 a107052a <=( a107051a  and  a107044a );
 a107056a <=( (not A167)  and  A168 );
 a107057a <=( A169  and  a107056a );
 a107060a <=( A199  and  A166 );
 a107063a <=( (not A201)  and  A200 );
 a107064a <=( a107063a  and  a107060a );
 a107065a <=( a107064a  and  a107057a );
 a107068a <=( (not A265)  and  A203 );
 a107071a <=( (not A268)  and  (not A266) );
 a107072a <=( a107071a  and  a107068a );
 a107075a <=( A299  and  (not A298) );
 a107078a <=( A302  and  (not A301) );
 a107079a <=( a107078a  and  a107075a );
 a107080a <=( a107079a  and  a107072a );
 a107084a <=( (not A167)  and  A168 );
 a107085a <=( A169  and  a107084a );
 a107088a <=( A199  and  A166 );
 a107091a <=( (not A201)  and  A200 );
 a107092a <=( a107091a  and  a107088a );
 a107093a <=( a107092a  and  a107085a );
 a107096a <=( (not A265)  and  A203 );
 a107099a <=( (not A268)  and  (not A266) );
 a107100a <=( a107099a  and  a107096a );
 a107103a <=( (not A299)  and  (not A298) );
 a107106a <=( (not A302)  and  A301 );
 a107107a <=( a107106a  and  a107103a );
 a107108a <=( a107107a  and  a107100a );
 a107112a <=( (not A167)  and  A168 );
 a107113a <=( A169  and  a107112a );
 a107116a <=( A199  and  A166 );
 a107119a <=( (not A201)  and  A200 );
 a107120a <=( a107119a  and  a107116a );
 a107121a <=( a107120a  and  a107113a );
 a107124a <=( (not A265)  and  A203 );
 a107127a <=( A269  and  (not A266) );
 a107128a <=( a107127a  and  a107124a );
 a107131a <=( A299  and  A298 );
 a107134a <=( (not A302)  and  A301 );
 a107135a <=( a107134a  and  a107131a );
 a107136a <=( a107135a  and  a107128a );
 a107140a <=( (not A167)  and  A168 );
 a107141a <=( A169  and  a107140a );
 a107144a <=( A199  and  A166 );
 a107147a <=( (not A201)  and  A200 );
 a107148a <=( a107147a  and  a107144a );
 a107149a <=( a107148a  and  a107141a );
 a107152a <=( (not A265)  and  A203 );
 a107155a <=( A269  and  (not A266) );
 a107156a <=( a107155a  and  a107152a );
 a107159a <=( (not A299)  and  A298 );
 a107162a <=( A302  and  (not A301) );
 a107163a <=( a107162a  and  a107159a );
 a107164a <=( a107163a  and  a107156a );
 a107168a <=( (not A167)  and  A168 );
 a107169a <=( A169  and  a107168a );
 a107172a <=( A199  and  A166 );
 a107175a <=( (not A201)  and  A200 );
 a107176a <=( a107175a  and  a107172a );
 a107177a <=( a107176a  and  a107169a );
 a107180a <=( (not A265)  and  A203 );
 a107183a <=( A269  and  (not A266) );
 a107184a <=( a107183a  and  a107180a );
 a107187a <=( A299  and  (not A298) );
 a107190a <=( A302  and  (not A301) );
 a107191a <=( a107190a  and  a107187a );
 a107192a <=( a107191a  and  a107184a );
 a107196a <=( (not A167)  and  A168 );
 a107197a <=( A169  and  a107196a );
 a107200a <=( A199  and  A166 );
 a107203a <=( (not A201)  and  A200 );
 a107204a <=( a107203a  and  a107200a );
 a107205a <=( a107204a  and  a107197a );
 a107208a <=( (not A265)  and  A203 );
 a107211a <=( A269  and  (not A266) );
 a107212a <=( a107211a  and  a107208a );
 a107215a <=( (not A299)  and  (not A298) );
 a107218a <=( (not A302)  and  A301 );
 a107219a <=( a107218a  and  a107215a );
 a107220a <=( a107219a  and  a107212a );
 a107224a <=( (not A167)  and  A168 );
 a107225a <=( A169  and  a107224a );
 a107228a <=( (not A199)  and  A166 );
 a107231a <=( (not A202)  and  A200 );
 a107232a <=( a107231a  and  a107228a );
 a107233a <=( a107232a  and  a107225a );
 a107236a <=( A265  and  A203 );
 a107239a <=( A268  and  A266 );
 a107240a <=( a107239a  and  a107236a );
 a107243a <=( (not A298)  and  (not A269) );
 a107246a <=( (not A301)  and  (not A299) );
 a107247a <=( a107246a  and  a107243a );
 a107248a <=( a107247a  and  a107240a );
 a107252a <=( (not A167)  and  A168 );
 a107253a <=( A169  and  a107252a );
 a107256a <=( (not A199)  and  A166 );
 a107259a <=( (not A202)  and  A200 );
 a107260a <=( a107259a  and  a107256a );
 a107261a <=( a107260a  and  a107253a );
 a107264a <=( A265  and  A203 );
 a107267a <=( A268  and  A266 );
 a107268a <=( a107267a  and  a107264a );
 a107271a <=( (not A298)  and  (not A269) );
 a107274a <=( A302  and  (not A299) );
 a107275a <=( a107274a  and  a107271a );
 a107276a <=( a107275a  and  a107268a );
 a107280a <=( (not A167)  and  A168 );
 a107281a <=( A169  and  a107280a );
 a107284a <=( (not A199)  and  A166 );
 a107287a <=( (not A202)  and  A200 );
 a107288a <=( a107287a  and  a107284a );
 a107289a <=( a107288a  and  a107281a );
 a107292a <=( (not A265)  and  A203 );
 a107295a <=( (not A268)  and  A266 );
 a107296a <=( a107295a  and  a107292a );
 a107299a <=( (not A298)  and  A269 );
 a107302a <=( (not A301)  and  (not A299) );
 a107303a <=( a107302a  and  a107299a );
 a107304a <=( a107303a  and  a107296a );
 a107308a <=( (not A167)  and  A168 );
 a107309a <=( A169  and  a107308a );
 a107312a <=( (not A199)  and  A166 );
 a107315a <=( (not A202)  and  A200 );
 a107316a <=( a107315a  and  a107312a );
 a107317a <=( a107316a  and  a107309a );
 a107320a <=( (not A265)  and  A203 );
 a107323a <=( (not A268)  and  A266 );
 a107324a <=( a107323a  and  a107320a );
 a107327a <=( (not A298)  and  A269 );
 a107330a <=( A302  and  (not A299) );
 a107331a <=( a107330a  and  a107327a );
 a107332a <=( a107331a  and  a107324a );
 a107336a <=( (not A167)  and  A168 );
 a107337a <=( A169  and  a107336a );
 a107340a <=( (not A199)  and  A166 );
 a107343a <=( (not A202)  and  A200 );
 a107344a <=( a107343a  and  a107340a );
 a107345a <=( a107344a  and  a107337a );
 a107348a <=( A265  and  A203 );
 a107351a <=( (not A268)  and  (not A266) );
 a107352a <=( a107351a  and  a107348a );
 a107355a <=( (not A298)  and  A269 );
 a107358a <=( (not A301)  and  (not A299) );
 a107359a <=( a107358a  and  a107355a );
 a107360a <=( a107359a  and  a107352a );
 a107364a <=( (not A167)  and  A168 );
 a107365a <=( A169  and  a107364a );
 a107368a <=( (not A199)  and  A166 );
 a107371a <=( (not A202)  and  A200 );
 a107372a <=( a107371a  and  a107368a );
 a107373a <=( a107372a  and  a107365a );
 a107376a <=( A265  and  A203 );
 a107379a <=( (not A268)  and  (not A266) );
 a107380a <=( a107379a  and  a107376a );
 a107383a <=( (not A298)  and  A269 );
 a107386a <=( A302  and  (not A299) );
 a107387a <=( a107386a  and  a107383a );
 a107388a <=( a107387a  and  a107380a );
 a107392a <=( (not A167)  and  A168 );
 a107393a <=( A169  and  a107392a );
 a107396a <=( (not A199)  and  A166 );
 a107399a <=( (not A202)  and  A200 );
 a107400a <=( a107399a  and  a107396a );
 a107401a <=( a107400a  and  a107393a );
 a107404a <=( (not A265)  and  A203 );
 a107407a <=( A268  and  (not A266) );
 a107408a <=( a107407a  and  a107404a );
 a107411a <=( (not A298)  and  (not A269) );
 a107414a <=( (not A301)  and  (not A299) );
 a107415a <=( a107414a  and  a107411a );
 a107416a <=( a107415a  and  a107408a );
 a107420a <=( (not A167)  and  A168 );
 a107421a <=( A169  and  a107420a );
 a107424a <=( (not A199)  and  A166 );
 a107427a <=( (not A202)  and  A200 );
 a107428a <=( a107427a  and  a107424a );
 a107429a <=( a107428a  and  a107421a );
 a107432a <=( (not A265)  and  A203 );
 a107435a <=( A268  and  (not A266) );
 a107436a <=( a107435a  and  a107432a );
 a107439a <=( (not A298)  and  (not A269) );
 a107442a <=( A302  and  (not A299) );
 a107443a <=( a107442a  and  a107439a );
 a107444a <=( a107443a  and  a107436a );
 a107448a <=( (not A167)  and  A168 );
 a107449a <=( A169  and  a107448a );
 a107452a <=( (not A199)  and  A166 );
 a107455a <=( (not A201)  and  A200 );
 a107456a <=( a107455a  and  a107452a );
 a107457a <=( a107456a  and  a107449a );
 a107460a <=( (not A265)  and  A202 );
 a107463a <=( (not A268)  and  (not A266) );
 a107464a <=( a107463a  and  a107460a );
 a107467a <=( A299  and  A298 );
 a107470a <=( (not A302)  and  A301 );
 a107471a <=( a107470a  and  a107467a );
 a107472a <=( a107471a  and  a107464a );
 a107476a <=( (not A167)  and  A168 );
 a107477a <=( A169  and  a107476a );
 a107480a <=( (not A199)  and  A166 );
 a107483a <=( (not A201)  and  A200 );
 a107484a <=( a107483a  and  a107480a );
 a107485a <=( a107484a  and  a107477a );
 a107488a <=( (not A265)  and  A202 );
 a107491a <=( (not A268)  and  (not A266) );
 a107492a <=( a107491a  and  a107488a );
 a107495a <=( (not A299)  and  A298 );
 a107498a <=( A302  and  (not A301) );
 a107499a <=( a107498a  and  a107495a );
 a107500a <=( a107499a  and  a107492a );
 a107504a <=( (not A167)  and  A168 );
 a107505a <=( A169  and  a107504a );
 a107508a <=( (not A199)  and  A166 );
 a107511a <=( (not A201)  and  A200 );
 a107512a <=( a107511a  and  a107508a );
 a107513a <=( a107512a  and  a107505a );
 a107516a <=( (not A265)  and  A202 );
 a107519a <=( (not A268)  and  (not A266) );
 a107520a <=( a107519a  and  a107516a );
 a107523a <=( A299  and  (not A298) );
 a107526a <=( A302  and  (not A301) );
 a107527a <=( a107526a  and  a107523a );
 a107528a <=( a107527a  and  a107520a );
 a107532a <=( (not A167)  and  A168 );
 a107533a <=( A169  and  a107532a );
 a107536a <=( (not A199)  and  A166 );
 a107539a <=( (not A201)  and  A200 );
 a107540a <=( a107539a  and  a107536a );
 a107541a <=( a107540a  and  a107533a );
 a107544a <=( (not A265)  and  A202 );
 a107547a <=( (not A268)  and  (not A266) );
 a107548a <=( a107547a  and  a107544a );
 a107551a <=( (not A299)  and  (not A298) );
 a107554a <=( (not A302)  and  A301 );
 a107555a <=( a107554a  and  a107551a );
 a107556a <=( a107555a  and  a107548a );
 a107560a <=( (not A167)  and  A168 );
 a107561a <=( A169  and  a107560a );
 a107564a <=( (not A199)  and  A166 );
 a107567a <=( (not A201)  and  A200 );
 a107568a <=( a107567a  and  a107564a );
 a107569a <=( a107568a  and  a107561a );
 a107572a <=( (not A265)  and  A202 );
 a107575a <=( A269  and  (not A266) );
 a107576a <=( a107575a  and  a107572a );
 a107579a <=( A299  and  A298 );
 a107582a <=( (not A302)  and  A301 );
 a107583a <=( a107582a  and  a107579a );
 a107584a <=( a107583a  and  a107576a );
 a107588a <=( (not A167)  and  A168 );
 a107589a <=( A169  and  a107588a );
 a107592a <=( (not A199)  and  A166 );
 a107595a <=( (not A201)  and  A200 );
 a107596a <=( a107595a  and  a107592a );
 a107597a <=( a107596a  and  a107589a );
 a107600a <=( (not A265)  and  A202 );
 a107603a <=( A269  and  (not A266) );
 a107604a <=( a107603a  and  a107600a );
 a107607a <=( (not A299)  and  A298 );
 a107610a <=( A302  and  (not A301) );
 a107611a <=( a107610a  and  a107607a );
 a107612a <=( a107611a  and  a107604a );
 a107616a <=( (not A167)  and  A168 );
 a107617a <=( A169  and  a107616a );
 a107620a <=( (not A199)  and  A166 );
 a107623a <=( (not A201)  and  A200 );
 a107624a <=( a107623a  and  a107620a );
 a107625a <=( a107624a  and  a107617a );
 a107628a <=( (not A265)  and  A202 );
 a107631a <=( A269  and  (not A266) );
 a107632a <=( a107631a  and  a107628a );
 a107635a <=( A299  and  (not A298) );
 a107638a <=( A302  and  (not A301) );
 a107639a <=( a107638a  and  a107635a );
 a107640a <=( a107639a  and  a107632a );
 a107644a <=( (not A167)  and  A168 );
 a107645a <=( A169  and  a107644a );
 a107648a <=( (not A199)  and  A166 );
 a107651a <=( (not A201)  and  A200 );
 a107652a <=( a107651a  and  a107648a );
 a107653a <=( a107652a  and  a107645a );
 a107656a <=( (not A265)  and  A202 );
 a107659a <=( A269  and  (not A266) );
 a107660a <=( a107659a  and  a107656a );
 a107663a <=( (not A299)  and  (not A298) );
 a107666a <=( (not A302)  and  A301 );
 a107667a <=( a107666a  and  a107663a );
 a107668a <=( a107667a  and  a107660a );
 a107672a <=( (not A167)  and  A168 );
 a107673a <=( A169  and  a107672a );
 a107676a <=( (not A199)  and  A166 );
 a107679a <=( (not A201)  and  A200 );
 a107680a <=( a107679a  and  a107676a );
 a107681a <=( a107680a  and  a107673a );
 a107684a <=( (not A265)  and  (not A203) );
 a107687a <=( (not A268)  and  (not A266) );
 a107688a <=( a107687a  and  a107684a );
 a107691a <=( A299  and  A298 );
 a107694a <=( (not A302)  and  A301 );
 a107695a <=( a107694a  and  a107691a );
 a107696a <=( a107695a  and  a107688a );
 a107700a <=( (not A167)  and  A168 );
 a107701a <=( A169  and  a107700a );
 a107704a <=( (not A199)  and  A166 );
 a107707a <=( (not A201)  and  A200 );
 a107708a <=( a107707a  and  a107704a );
 a107709a <=( a107708a  and  a107701a );
 a107712a <=( (not A265)  and  (not A203) );
 a107715a <=( (not A268)  and  (not A266) );
 a107716a <=( a107715a  and  a107712a );
 a107719a <=( (not A299)  and  A298 );
 a107722a <=( A302  and  (not A301) );
 a107723a <=( a107722a  and  a107719a );
 a107724a <=( a107723a  and  a107716a );
 a107728a <=( (not A167)  and  A168 );
 a107729a <=( A169  and  a107728a );
 a107732a <=( (not A199)  and  A166 );
 a107735a <=( (not A201)  and  A200 );
 a107736a <=( a107735a  and  a107732a );
 a107737a <=( a107736a  and  a107729a );
 a107740a <=( (not A265)  and  (not A203) );
 a107743a <=( (not A268)  and  (not A266) );
 a107744a <=( a107743a  and  a107740a );
 a107747a <=( A299  and  (not A298) );
 a107750a <=( A302  and  (not A301) );
 a107751a <=( a107750a  and  a107747a );
 a107752a <=( a107751a  and  a107744a );
 a107756a <=( (not A167)  and  A168 );
 a107757a <=( A169  and  a107756a );
 a107760a <=( (not A199)  and  A166 );
 a107763a <=( (not A201)  and  A200 );
 a107764a <=( a107763a  and  a107760a );
 a107765a <=( a107764a  and  a107757a );
 a107768a <=( (not A265)  and  (not A203) );
 a107771a <=( (not A268)  and  (not A266) );
 a107772a <=( a107771a  and  a107768a );
 a107775a <=( (not A299)  and  (not A298) );
 a107778a <=( (not A302)  and  A301 );
 a107779a <=( a107778a  and  a107775a );
 a107780a <=( a107779a  and  a107772a );
 a107784a <=( (not A167)  and  A168 );
 a107785a <=( A169  and  a107784a );
 a107788a <=( (not A199)  and  A166 );
 a107791a <=( (not A201)  and  A200 );
 a107792a <=( a107791a  and  a107788a );
 a107793a <=( a107792a  and  a107785a );
 a107796a <=( (not A265)  and  (not A203) );
 a107799a <=( A269  and  (not A266) );
 a107800a <=( a107799a  and  a107796a );
 a107803a <=( A299  and  A298 );
 a107806a <=( (not A302)  and  A301 );
 a107807a <=( a107806a  and  a107803a );
 a107808a <=( a107807a  and  a107800a );
 a107812a <=( (not A167)  and  A168 );
 a107813a <=( A169  and  a107812a );
 a107816a <=( (not A199)  and  A166 );
 a107819a <=( (not A201)  and  A200 );
 a107820a <=( a107819a  and  a107816a );
 a107821a <=( a107820a  and  a107813a );
 a107824a <=( (not A265)  and  (not A203) );
 a107827a <=( A269  and  (not A266) );
 a107828a <=( a107827a  and  a107824a );
 a107831a <=( (not A299)  and  A298 );
 a107834a <=( A302  and  (not A301) );
 a107835a <=( a107834a  and  a107831a );
 a107836a <=( a107835a  and  a107828a );
 a107840a <=( (not A167)  and  A168 );
 a107841a <=( A169  and  a107840a );
 a107844a <=( (not A199)  and  A166 );
 a107847a <=( (not A201)  and  A200 );
 a107848a <=( a107847a  and  a107844a );
 a107849a <=( a107848a  and  a107841a );
 a107852a <=( (not A265)  and  (not A203) );
 a107855a <=( A269  and  (not A266) );
 a107856a <=( a107855a  and  a107852a );
 a107859a <=( A299  and  (not A298) );
 a107862a <=( A302  and  (not A301) );
 a107863a <=( a107862a  and  a107859a );
 a107864a <=( a107863a  and  a107856a );
 a107868a <=( (not A167)  and  A168 );
 a107869a <=( A169  and  a107868a );
 a107872a <=( (not A199)  and  A166 );
 a107875a <=( (not A201)  and  A200 );
 a107876a <=( a107875a  and  a107872a );
 a107877a <=( a107876a  and  a107869a );
 a107880a <=( (not A265)  and  (not A203) );
 a107883a <=( A269  and  (not A266) );
 a107884a <=( a107883a  and  a107880a );
 a107887a <=( (not A299)  and  (not A298) );
 a107890a <=( (not A302)  and  A301 );
 a107891a <=( a107890a  and  a107887a );
 a107892a <=( a107891a  and  a107884a );
 a107896a <=( (not A167)  and  A168 );
 a107897a <=( A169  and  a107896a );
 a107900a <=( A199  and  A166 );
 a107903a <=( (not A202)  and  (not A200) );
 a107904a <=( a107903a  and  a107900a );
 a107905a <=( a107904a  and  a107897a );
 a107908a <=( A265  and  A203 );
 a107911a <=( A268  and  A266 );
 a107912a <=( a107911a  and  a107908a );
 a107915a <=( (not A298)  and  (not A269) );
 a107918a <=( (not A301)  and  (not A299) );
 a107919a <=( a107918a  and  a107915a );
 a107920a <=( a107919a  and  a107912a );
 a107924a <=( (not A167)  and  A168 );
 a107925a <=( A169  and  a107924a );
 a107928a <=( A199  and  A166 );
 a107931a <=( (not A202)  and  (not A200) );
 a107932a <=( a107931a  and  a107928a );
 a107933a <=( a107932a  and  a107925a );
 a107936a <=( A265  and  A203 );
 a107939a <=( A268  and  A266 );
 a107940a <=( a107939a  and  a107936a );
 a107943a <=( (not A298)  and  (not A269) );
 a107946a <=( A302  and  (not A299) );
 a107947a <=( a107946a  and  a107943a );
 a107948a <=( a107947a  and  a107940a );
 a107952a <=( (not A167)  and  A168 );
 a107953a <=( A169  and  a107952a );
 a107956a <=( A199  and  A166 );
 a107959a <=( (not A202)  and  (not A200) );
 a107960a <=( a107959a  and  a107956a );
 a107961a <=( a107960a  and  a107953a );
 a107964a <=( (not A265)  and  A203 );
 a107967a <=( (not A268)  and  A266 );
 a107968a <=( a107967a  and  a107964a );
 a107971a <=( (not A298)  and  A269 );
 a107974a <=( (not A301)  and  (not A299) );
 a107975a <=( a107974a  and  a107971a );
 a107976a <=( a107975a  and  a107968a );
 a107980a <=( (not A167)  and  A168 );
 a107981a <=( A169  and  a107980a );
 a107984a <=( A199  and  A166 );
 a107987a <=( (not A202)  and  (not A200) );
 a107988a <=( a107987a  and  a107984a );
 a107989a <=( a107988a  and  a107981a );
 a107992a <=( (not A265)  and  A203 );
 a107995a <=( (not A268)  and  A266 );
 a107996a <=( a107995a  and  a107992a );
 a107999a <=( (not A298)  and  A269 );
 a108002a <=( A302  and  (not A299) );
 a108003a <=( a108002a  and  a107999a );
 a108004a <=( a108003a  and  a107996a );
 a108008a <=( (not A167)  and  A168 );
 a108009a <=( A169  and  a108008a );
 a108012a <=( A199  and  A166 );
 a108015a <=( (not A202)  and  (not A200) );
 a108016a <=( a108015a  and  a108012a );
 a108017a <=( a108016a  and  a108009a );
 a108020a <=( A265  and  A203 );
 a108023a <=( (not A268)  and  (not A266) );
 a108024a <=( a108023a  and  a108020a );
 a108027a <=( (not A298)  and  A269 );
 a108030a <=( (not A301)  and  (not A299) );
 a108031a <=( a108030a  and  a108027a );
 a108032a <=( a108031a  and  a108024a );
 a108036a <=( (not A167)  and  A168 );
 a108037a <=( A169  and  a108036a );
 a108040a <=( A199  and  A166 );
 a108043a <=( (not A202)  and  (not A200) );
 a108044a <=( a108043a  and  a108040a );
 a108045a <=( a108044a  and  a108037a );
 a108048a <=( A265  and  A203 );
 a108051a <=( (not A268)  and  (not A266) );
 a108052a <=( a108051a  and  a108048a );
 a108055a <=( (not A298)  and  A269 );
 a108058a <=( A302  and  (not A299) );
 a108059a <=( a108058a  and  a108055a );
 a108060a <=( a108059a  and  a108052a );
 a108064a <=( (not A167)  and  A168 );
 a108065a <=( A169  and  a108064a );
 a108068a <=( A199  and  A166 );
 a108071a <=( (not A202)  and  (not A200) );
 a108072a <=( a108071a  and  a108068a );
 a108073a <=( a108072a  and  a108065a );
 a108076a <=( (not A265)  and  A203 );
 a108079a <=( A268  and  (not A266) );
 a108080a <=( a108079a  and  a108076a );
 a108083a <=( (not A298)  and  (not A269) );
 a108086a <=( (not A301)  and  (not A299) );
 a108087a <=( a108086a  and  a108083a );
 a108088a <=( a108087a  and  a108080a );
 a108092a <=( (not A167)  and  A168 );
 a108093a <=( A169  and  a108092a );
 a108096a <=( A199  and  A166 );
 a108099a <=( (not A202)  and  (not A200) );
 a108100a <=( a108099a  and  a108096a );
 a108101a <=( a108100a  and  a108093a );
 a108104a <=( (not A265)  and  A203 );
 a108107a <=( A268  and  (not A266) );
 a108108a <=( a108107a  and  a108104a );
 a108111a <=( (not A298)  and  (not A269) );
 a108114a <=( A302  and  (not A299) );
 a108115a <=( a108114a  and  a108111a );
 a108116a <=( a108115a  and  a108108a );
 a108120a <=( (not A167)  and  A168 );
 a108121a <=( A169  and  a108120a );
 a108124a <=( A199  and  A166 );
 a108127a <=( (not A201)  and  (not A200) );
 a108128a <=( a108127a  and  a108124a );
 a108129a <=( a108128a  and  a108121a );
 a108132a <=( (not A265)  and  A202 );
 a108135a <=( (not A268)  and  (not A266) );
 a108136a <=( a108135a  and  a108132a );
 a108139a <=( A299  and  A298 );
 a108142a <=( (not A302)  and  A301 );
 a108143a <=( a108142a  and  a108139a );
 a108144a <=( a108143a  and  a108136a );
 a108148a <=( (not A167)  and  A168 );
 a108149a <=( A169  and  a108148a );
 a108152a <=( A199  and  A166 );
 a108155a <=( (not A201)  and  (not A200) );
 a108156a <=( a108155a  and  a108152a );
 a108157a <=( a108156a  and  a108149a );
 a108160a <=( (not A265)  and  A202 );
 a108163a <=( (not A268)  and  (not A266) );
 a108164a <=( a108163a  and  a108160a );
 a108167a <=( (not A299)  and  A298 );
 a108170a <=( A302  and  (not A301) );
 a108171a <=( a108170a  and  a108167a );
 a108172a <=( a108171a  and  a108164a );
 a108176a <=( (not A167)  and  A168 );
 a108177a <=( A169  and  a108176a );
 a108180a <=( A199  and  A166 );
 a108183a <=( (not A201)  and  (not A200) );
 a108184a <=( a108183a  and  a108180a );
 a108185a <=( a108184a  and  a108177a );
 a108188a <=( (not A265)  and  A202 );
 a108191a <=( (not A268)  and  (not A266) );
 a108192a <=( a108191a  and  a108188a );
 a108195a <=( A299  and  (not A298) );
 a108198a <=( A302  and  (not A301) );
 a108199a <=( a108198a  and  a108195a );
 a108200a <=( a108199a  and  a108192a );
 a108204a <=( (not A167)  and  A168 );
 a108205a <=( A169  and  a108204a );
 a108208a <=( A199  and  A166 );
 a108211a <=( (not A201)  and  (not A200) );
 a108212a <=( a108211a  and  a108208a );
 a108213a <=( a108212a  and  a108205a );
 a108216a <=( (not A265)  and  A202 );
 a108219a <=( (not A268)  and  (not A266) );
 a108220a <=( a108219a  and  a108216a );
 a108223a <=( (not A299)  and  (not A298) );
 a108226a <=( (not A302)  and  A301 );
 a108227a <=( a108226a  and  a108223a );
 a108228a <=( a108227a  and  a108220a );
 a108232a <=( (not A167)  and  A168 );
 a108233a <=( A169  and  a108232a );
 a108236a <=( A199  and  A166 );
 a108239a <=( (not A201)  and  (not A200) );
 a108240a <=( a108239a  and  a108236a );
 a108241a <=( a108240a  and  a108233a );
 a108244a <=( (not A265)  and  A202 );
 a108247a <=( A269  and  (not A266) );
 a108248a <=( a108247a  and  a108244a );
 a108251a <=( A299  and  A298 );
 a108254a <=( (not A302)  and  A301 );
 a108255a <=( a108254a  and  a108251a );
 a108256a <=( a108255a  and  a108248a );
 a108260a <=( (not A167)  and  A168 );
 a108261a <=( A169  and  a108260a );
 a108264a <=( A199  and  A166 );
 a108267a <=( (not A201)  and  (not A200) );
 a108268a <=( a108267a  and  a108264a );
 a108269a <=( a108268a  and  a108261a );
 a108272a <=( (not A265)  and  A202 );
 a108275a <=( A269  and  (not A266) );
 a108276a <=( a108275a  and  a108272a );
 a108279a <=( (not A299)  and  A298 );
 a108282a <=( A302  and  (not A301) );
 a108283a <=( a108282a  and  a108279a );
 a108284a <=( a108283a  and  a108276a );
 a108288a <=( (not A167)  and  A168 );
 a108289a <=( A169  and  a108288a );
 a108292a <=( A199  and  A166 );
 a108295a <=( (not A201)  and  (not A200) );
 a108296a <=( a108295a  and  a108292a );
 a108297a <=( a108296a  and  a108289a );
 a108300a <=( (not A265)  and  A202 );
 a108303a <=( A269  and  (not A266) );
 a108304a <=( a108303a  and  a108300a );
 a108307a <=( A299  and  (not A298) );
 a108310a <=( A302  and  (not A301) );
 a108311a <=( a108310a  and  a108307a );
 a108312a <=( a108311a  and  a108304a );
 a108316a <=( (not A167)  and  A168 );
 a108317a <=( A169  and  a108316a );
 a108320a <=( A199  and  A166 );
 a108323a <=( (not A201)  and  (not A200) );
 a108324a <=( a108323a  and  a108320a );
 a108325a <=( a108324a  and  a108317a );
 a108328a <=( (not A265)  and  A202 );
 a108331a <=( A269  and  (not A266) );
 a108332a <=( a108331a  and  a108328a );
 a108335a <=( (not A299)  and  (not A298) );
 a108338a <=( (not A302)  and  A301 );
 a108339a <=( a108338a  and  a108335a );
 a108340a <=( a108339a  and  a108332a );
 a108344a <=( (not A167)  and  A168 );
 a108345a <=( A169  and  a108344a );
 a108348a <=( A199  and  A166 );
 a108351a <=( (not A201)  and  (not A200) );
 a108352a <=( a108351a  and  a108348a );
 a108353a <=( a108352a  and  a108345a );
 a108356a <=( (not A265)  and  (not A203) );
 a108359a <=( (not A268)  and  (not A266) );
 a108360a <=( a108359a  and  a108356a );
 a108363a <=( A299  and  A298 );
 a108366a <=( (not A302)  and  A301 );
 a108367a <=( a108366a  and  a108363a );
 a108368a <=( a108367a  and  a108360a );
 a108372a <=( (not A167)  and  A168 );
 a108373a <=( A169  and  a108372a );
 a108376a <=( A199  and  A166 );
 a108379a <=( (not A201)  and  (not A200) );
 a108380a <=( a108379a  and  a108376a );
 a108381a <=( a108380a  and  a108373a );
 a108384a <=( (not A265)  and  (not A203) );
 a108387a <=( (not A268)  and  (not A266) );
 a108388a <=( a108387a  and  a108384a );
 a108391a <=( (not A299)  and  A298 );
 a108394a <=( A302  and  (not A301) );
 a108395a <=( a108394a  and  a108391a );
 a108396a <=( a108395a  and  a108388a );
 a108400a <=( (not A167)  and  A168 );
 a108401a <=( A169  and  a108400a );
 a108404a <=( A199  and  A166 );
 a108407a <=( (not A201)  and  (not A200) );
 a108408a <=( a108407a  and  a108404a );
 a108409a <=( a108408a  and  a108401a );
 a108412a <=( (not A265)  and  (not A203) );
 a108415a <=( (not A268)  and  (not A266) );
 a108416a <=( a108415a  and  a108412a );
 a108419a <=( A299  and  (not A298) );
 a108422a <=( A302  and  (not A301) );
 a108423a <=( a108422a  and  a108419a );
 a108424a <=( a108423a  and  a108416a );
 a108428a <=( (not A167)  and  A168 );
 a108429a <=( A169  and  a108428a );
 a108432a <=( A199  and  A166 );
 a108435a <=( (not A201)  and  (not A200) );
 a108436a <=( a108435a  and  a108432a );
 a108437a <=( a108436a  and  a108429a );
 a108440a <=( (not A265)  and  (not A203) );
 a108443a <=( (not A268)  and  (not A266) );
 a108444a <=( a108443a  and  a108440a );
 a108447a <=( (not A299)  and  (not A298) );
 a108450a <=( (not A302)  and  A301 );
 a108451a <=( a108450a  and  a108447a );
 a108452a <=( a108451a  and  a108444a );
 a108456a <=( (not A167)  and  A168 );
 a108457a <=( A169  and  a108456a );
 a108460a <=( A199  and  A166 );
 a108463a <=( (not A201)  and  (not A200) );
 a108464a <=( a108463a  and  a108460a );
 a108465a <=( a108464a  and  a108457a );
 a108468a <=( (not A265)  and  (not A203) );
 a108471a <=( A269  and  (not A266) );
 a108472a <=( a108471a  and  a108468a );
 a108475a <=( A299  and  A298 );
 a108478a <=( (not A302)  and  A301 );
 a108479a <=( a108478a  and  a108475a );
 a108480a <=( a108479a  and  a108472a );
 a108484a <=( (not A167)  and  A168 );
 a108485a <=( A169  and  a108484a );
 a108488a <=( A199  and  A166 );
 a108491a <=( (not A201)  and  (not A200) );
 a108492a <=( a108491a  and  a108488a );
 a108493a <=( a108492a  and  a108485a );
 a108496a <=( (not A265)  and  (not A203) );
 a108499a <=( A269  and  (not A266) );
 a108500a <=( a108499a  and  a108496a );
 a108503a <=( (not A299)  and  A298 );
 a108506a <=( A302  and  (not A301) );
 a108507a <=( a108506a  and  a108503a );
 a108508a <=( a108507a  and  a108500a );
 a108512a <=( (not A167)  and  A168 );
 a108513a <=( A169  and  a108512a );
 a108516a <=( A199  and  A166 );
 a108519a <=( (not A201)  and  (not A200) );
 a108520a <=( a108519a  and  a108516a );
 a108521a <=( a108520a  and  a108513a );
 a108524a <=( (not A265)  and  (not A203) );
 a108527a <=( A269  and  (not A266) );
 a108528a <=( a108527a  and  a108524a );
 a108531a <=( A299  and  (not A298) );
 a108534a <=( A302  and  (not A301) );
 a108535a <=( a108534a  and  a108531a );
 a108536a <=( a108535a  and  a108528a );
 a108540a <=( (not A167)  and  A168 );
 a108541a <=( A169  and  a108540a );
 a108544a <=( A199  and  A166 );
 a108547a <=( (not A201)  and  (not A200) );
 a108548a <=( a108547a  and  a108544a );
 a108549a <=( a108548a  and  a108541a );
 a108552a <=( (not A265)  and  (not A203) );
 a108555a <=( A269  and  (not A266) );
 a108556a <=( a108555a  and  a108552a );
 a108559a <=( (not A299)  and  (not A298) );
 a108562a <=( (not A302)  and  A301 );
 a108563a <=( a108562a  and  a108559a );
 a108564a <=( a108563a  and  a108556a );
 a108568a <=( (not A167)  and  A168 );
 a108569a <=( A169  and  a108568a );
 a108572a <=( (not A199)  and  A166 );
 a108575a <=( (not A202)  and  (not A200) );
 a108576a <=( a108575a  and  a108572a );
 a108577a <=( a108576a  and  a108569a );
 a108580a <=( A266  and  A265 );
 a108583a <=( (not A268)  and  (not A267) );
 a108584a <=( a108583a  and  a108580a );
 a108587a <=( A299  and  A298 );
 a108590a <=( (not A302)  and  A301 );
 a108591a <=( a108590a  and  a108587a );
 a108592a <=( a108591a  and  a108584a );
 a108596a <=( (not A167)  and  A168 );
 a108597a <=( A169  and  a108596a );
 a108600a <=( (not A199)  and  A166 );
 a108603a <=( (not A202)  and  (not A200) );
 a108604a <=( a108603a  and  a108600a );
 a108605a <=( a108604a  and  a108597a );
 a108608a <=( A266  and  A265 );
 a108611a <=( (not A268)  and  (not A267) );
 a108612a <=( a108611a  and  a108608a );
 a108615a <=( (not A299)  and  A298 );
 a108618a <=( A302  and  (not A301) );
 a108619a <=( a108618a  and  a108615a );
 a108620a <=( a108619a  and  a108612a );
 a108624a <=( (not A167)  and  A168 );
 a108625a <=( A169  and  a108624a );
 a108628a <=( (not A199)  and  A166 );
 a108631a <=( (not A202)  and  (not A200) );
 a108632a <=( a108631a  and  a108628a );
 a108633a <=( a108632a  and  a108625a );
 a108636a <=( A266  and  A265 );
 a108639a <=( (not A268)  and  (not A267) );
 a108640a <=( a108639a  and  a108636a );
 a108643a <=( A299  and  (not A298) );
 a108646a <=( A302  and  (not A301) );
 a108647a <=( a108646a  and  a108643a );
 a108648a <=( a108647a  and  a108640a );
 a108652a <=( (not A167)  and  A168 );
 a108653a <=( A169  and  a108652a );
 a108656a <=( (not A199)  and  A166 );
 a108659a <=( (not A202)  and  (not A200) );
 a108660a <=( a108659a  and  a108656a );
 a108661a <=( a108660a  and  a108653a );
 a108664a <=( A266  and  A265 );
 a108667a <=( (not A268)  and  (not A267) );
 a108668a <=( a108667a  and  a108664a );
 a108671a <=( (not A299)  and  (not A298) );
 a108674a <=( (not A302)  and  A301 );
 a108675a <=( a108674a  and  a108671a );
 a108676a <=( a108675a  and  a108668a );
 a108680a <=( (not A167)  and  A168 );
 a108681a <=( A169  and  a108680a );
 a108684a <=( (not A199)  and  A166 );
 a108687a <=( (not A202)  and  (not A200) );
 a108688a <=( a108687a  and  a108684a );
 a108689a <=( a108688a  and  a108681a );
 a108692a <=( A266  and  A265 );
 a108695a <=( A269  and  (not A267) );
 a108696a <=( a108695a  and  a108692a );
 a108699a <=( A299  and  A298 );
 a108702a <=( (not A302)  and  A301 );
 a108703a <=( a108702a  and  a108699a );
 a108704a <=( a108703a  and  a108696a );
 a108708a <=( (not A167)  and  A168 );
 a108709a <=( A169  and  a108708a );
 a108712a <=( (not A199)  and  A166 );
 a108715a <=( (not A202)  and  (not A200) );
 a108716a <=( a108715a  and  a108712a );
 a108717a <=( a108716a  and  a108709a );
 a108720a <=( A266  and  A265 );
 a108723a <=( A269  and  (not A267) );
 a108724a <=( a108723a  and  a108720a );
 a108727a <=( (not A299)  and  A298 );
 a108730a <=( A302  and  (not A301) );
 a108731a <=( a108730a  and  a108727a );
 a108732a <=( a108731a  and  a108724a );
 a108736a <=( (not A167)  and  A168 );
 a108737a <=( A169  and  a108736a );
 a108740a <=( (not A199)  and  A166 );
 a108743a <=( (not A202)  and  (not A200) );
 a108744a <=( a108743a  and  a108740a );
 a108745a <=( a108744a  and  a108737a );
 a108748a <=( A266  and  A265 );
 a108751a <=( A269  and  (not A267) );
 a108752a <=( a108751a  and  a108748a );
 a108755a <=( A299  and  (not A298) );
 a108758a <=( A302  and  (not A301) );
 a108759a <=( a108758a  and  a108755a );
 a108760a <=( a108759a  and  a108752a );
 a108764a <=( (not A167)  and  A168 );
 a108765a <=( A169  and  a108764a );
 a108768a <=( (not A199)  and  A166 );
 a108771a <=( (not A202)  and  (not A200) );
 a108772a <=( a108771a  and  a108768a );
 a108773a <=( a108772a  and  a108765a );
 a108776a <=( A266  and  A265 );
 a108779a <=( A269  and  (not A267) );
 a108780a <=( a108779a  and  a108776a );
 a108783a <=( (not A299)  and  (not A298) );
 a108786a <=( (not A302)  and  A301 );
 a108787a <=( a108786a  and  a108783a );
 a108788a <=( a108787a  and  a108780a );
 a108792a <=( (not A167)  and  A168 );
 a108793a <=( A169  and  a108792a );
 a108796a <=( (not A199)  and  A166 );
 a108799a <=( (not A202)  and  (not A200) );
 a108800a <=( a108799a  and  a108796a );
 a108801a <=( a108800a  and  a108793a );
 a108804a <=( A266  and  (not A265) );
 a108807a <=( A268  and  (not A267) );
 a108808a <=( a108807a  and  a108804a );
 a108811a <=( A299  and  A298 );
 a108814a <=( (not A302)  and  A301 );
 a108815a <=( a108814a  and  a108811a );
 a108816a <=( a108815a  and  a108808a );
 a108820a <=( (not A167)  and  A168 );
 a108821a <=( A169  and  a108820a );
 a108824a <=( (not A199)  and  A166 );
 a108827a <=( (not A202)  and  (not A200) );
 a108828a <=( a108827a  and  a108824a );
 a108829a <=( a108828a  and  a108821a );
 a108832a <=( A266  and  (not A265) );
 a108835a <=( A268  and  (not A267) );
 a108836a <=( a108835a  and  a108832a );
 a108839a <=( (not A299)  and  A298 );
 a108842a <=( A302  and  (not A301) );
 a108843a <=( a108842a  and  a108839a );
 a108844a <=( a108843a  and  a108836a );
 a108848a <=( (not A167)  and  A168 );
 a108849a <=( A169  and  a108848a );
 a108852a <=( (not A199)  and  A166 );
 a108855a <=( (not A202)  and  (not A200) );
 a108856a <=( a108855a  and  a108852a );
 a108857a <=( a108856a  and  a108849a );
 a108860a <=( A266  and  (not A265) );
 a108863a <=( A268  and  (not A267) );
 a108864a <=( a108863a  and  a108860a );
 a108867a <=( A299  and  (not A298) );
 a108870a <=( A302  and  (not A301) );
 a108871a <=( a108870a  and  a108867a );
 a108872a <=( a108871a  and  a108864a );
 a108876a <=( (not A167)  and  A168 );
 a108877a <=( A169  and  a108876a );
 a108880a <=( (not A199)  and  A166 );
 a108883a <=( (not A202)  and  (not A200) );
 a108884a <=( a108883a  and  a108880a );
 a108885a <=( a108884a  and  a108877a );
 a108888a <=( A266  and  (not A265) );
 a108891a <=( A268  and  (not A267) );
 a108892a <=( a108891a  and  a108888a );
 a108895a <=( (not A299)  and  (not A298) );
 a108898a <=( (not A302)  and  A301 );
 a108899a <=( a108898a  and  a108895a );
 a108900a <=( a108899a  and  a108892a );
 a108904a <=( (not A167)  and  A168 );
 a108905a <=( A169  and  a108904a );
 a108908a <=( (not A199)  and  A166 );
 a108911a <=( (not A202)  and  (not A200) );
 a108912a <=( a108911a  and  a108908a );
 a108913a <=( a108912a  and  a108905a );
 a108916a <=( A266  and  (not A265) );
 a108919a <=( (not A269)  and  (not A267) );
 a108920a <=( a108919a  and  a108916a );
 a108923a <=( A299  and  A298 );
 a108926a <=( (not A302)  and  A301 );
 a108927a <=( a108926a  and  a108923a );
 a108928a <=( a108927a  and  a108920a );
 a108932a <=( (not A167)  and  A168 );
 a108933a <=( A169  and  a108932a );
 a108936a <=( (not A199)  and  A166 );
 a108939a <=( (not A202)  and  (not A200) );
 a108940a <=( a108939a  and  a108936a );
 a108941a <=( a108940a  and  a108933a );
 a108944a <=( A266  and  (not A265) );
 a108947a <=( (not A269)  and  (not A267) );
 a108948a <=( a108947a  and  a108944a );
 a108951a <=( (not A299)  and  A298 );
 a108954a <=( A302  and  (not A301) );
 a108955a <=( a108954a  and  a108951a );
 a108956a <=( a108955a  and  a108948a );
 a108960a <=( (not A167)  and  A168 );
 a108961a <=( A169  and  a108960a );
 a108964a <=( (not A199)  and  A166 );
 a108967a <=( (not A202)  and  (not A200) );
 a108968a <=( a108967a  and  a108964a );
 a108969a <=( a108968a  and  a108961a );
 a108972a <=( A266  and  (not A265) );
 a108975a <=( (not A269)  and  (not A267) );
 a108976a <=( a108975a  and  a108972a );
 a108979a <=( A299  and  (not A298) );
 a108982a <=( A302  and  (not A301) );
 a108983a <=( a108982a  and  a108979a );
 a108984a <=( a108983a  and  a108976a );
 a108988a <=( (not A167)  and  A168 );
 a108989a <=( A169  and  a108988a );
 a108992a <=( (not A199)  and  A166 );
 a108995a <=( (not A202)  and  (not A200) );
 a108996a <=( a108995a  and  a108992a );
 a108997a <=( a108996a  and  a108989a );
 a109000a <=( A266  and  (not A265) );
 a109003a <=( (not A269)  and  (not A267) );
 a109004a <=( a109003a  and  a109000a );
 a109007a <=( (not A299)  and  (not A298) );
 a109010a <=( (not A302)  and  A301 );
 a109011a <=( a109010a  and  a109007a );
 a109012a <=( a109011a  and  a109004a );
 a109016a <=( (not A167)  and  A168 );
 a109017a <=( A169  and  a109016a );
 a109020a <=( (not A199)  and  A166 );
 a109023a <=( (not A202)  and  (not A200) );
 a109024a <=( a109023a  and  a109020a );
 a109025a <=( a109024a  and  a109017a );
 a109028a <=( (not A266)  and  A265 );
 a109031a <=( A268  and  (not A267) );
 a109032a <=( a109031a  and  a109028a );
 a109035a <=( A299  and  A298 );
 a109038a <=( (not A302)  and  A301 );
 a109039a <=( a109038a  and  a109035a );
 a109040a <=( a109039a  and  a109032a );
 a109044a <=( (not A167)  and  A168 );
 a109045a <=( A169  and  a109044a );
 a109048a <=( (not A199)  and  A166 );
 a109051a <=( (not A202)  and  (not A200) );
 a109052a <=( a109051a  and  a109048a );
 a109053a <=( a109052a  and  a109045a );
 a109056a <=( (not A266)  and  A265 );
 a109059a <=( A268  and  (not A267) );
 a109060a <=( a109059a  and  a109056a );
 a109063a <=( (not A299)  and  A298 );
 a109066a <=( A302  and  (not A301) );
 a109067a <=( a109066a  and  a109063a );
 a109068a <=( a109067a  and  a109060a );
 a109072a <=( (not A167)  and  A168 );
 a109073a <=( A169  and  a109072a );
 a109076a <=( (not A199)  and  A166 );
 a109079a <=( (not A202)  and  (not A200) );
 a109080a <=( a109079a  and  a109076a );
 a109081a <=( a109080a  and  a109073a );
 a109084a <=( (not A266)  and  A265 );
 a109087a <=( A268  and  (not A267) );
 a109088a <=( a109087a  and  a109084a );
 a109091a <=( A299  and  (not A298) );
 a109094a <=( A302  and  (not A301) );
 a109095a <=( a109094a  and  a109091a );
 a109096a <=( a109095a  and  a109088a );
 a109100a <=( (not A167)  and  A168 );
 a109101a <=( A169  and  a109100a );
 a109104a <=( (not A199)  and  A166 );
 a109107a <=( (not A202)  and  (not A200) );
 a109108a <=( a109107a  and  a109104a );
 a109109a <=( a109108a  and  a109101a );
 a109112a <=( (not A266)  and  A265 );
 a109115a <=( A268  and  (not A267) );
 a109116a <=( a109115a  and  a109112a );
 a109119a <=( (not A299)  and  (not A298) );
 a109122a <=( (not A302)  and  A301 );
 a109123a <=( a109122a  and  a109119a );
 a109124a <=( a109123a  and  a109116a );
 a109128a <=( (not A167)  and  A168 );
 a109129a <=( A169  and  a109128a );
 a109132a <=( (not A199)  and  A166 );
 a109135a <=( (not A202)  and  (not A200) );
 a109136a <=( a109135a  and  a109132a );
 a109137a <=( a109136a  and  a109129a );
 a109140a <=( (not A266)  and  A265 );
 a109143a <=( (not A269)  and  (not A267) );
 a109144a <=( a109143a  and  a109140a );
 a109147a <=( A299  and  A298 );
 a109150a <=( (not A302)  and  A301 );
 a109151a <=( a109150a  and  a109147a );
 a109152a <=( a109151a  and  a109144a );
 a109156a <=( (not A167)  and  A168 );
 a109157a <=( A169  and  a109156a );
 a109160a <=( (not A199)  and  A166 );
 a109163a <=( (not A202)  and  (not A200) );
 a109164a <=( a109163a  and  a109160a );
 a109165a <=( a109164a  and  a109157a );
 a109168a <=( (not A266)  and  A265 );
 a109171a <=( (not A269)  and  (not A267) );
 a109172a <=( a109171a  and  a109168a );
 a109175a <=( (not A299)  and  A298 );
 a109178a <=( A302  and  (not A301) );
 a109179a <=( a109178a  and  a109175a );
 a109180a <=( a109179a  and  a109172a );
 a109184a <=( (not A167)  and  A168 );
 a109185a <=( A169  and  a109184a );
 a109188a <=( (not A199)  and  A166 );
 a109191a <=( (not A202)  and  (not A200) );
 a109192a <=( a109191a  and  a109188a );
 a109193a <=( a109192a  and  a109185a );
 a109196a <=( (not A266)  and  A265 );
 a109199a <=( (not A269)  and  (not A267) );
 a109200a <=( a109199a  and  a109196a );
 a109203a <=( A299  and  (not A298) );
 a109206a <=( A302  and  (not A301) );
 a109207a <=( a109206a  and  a109203a );
 a109208a <=( a109207a  and  a109200a );
 a109212a <=( (not A167)  and  A168 );
 a109213a <=( A169  and  a109212a );
 a109216a <=( (not A199)  and  A166 );
 a109219a <=( (not A202)  and  (not A200) );
 a109220a <=( a109219a  and  a109216a );
 a109221a <=( a109220a  and  a109213a );
 a109224a <=( (not A266)  and  A265 );
 a109227a <=( (not A269)  and  (not A267) );
 a109228a <=( a109227a  and  a109224a );
 a109231a <=( (not A299)  and  (not A298) );
 a109234a <=( (not A302)  and  A301 );
 a109235a <=( a109234a  and  a109231a );
 a109236a <=( a109235a  and  a109228a );
 a109240a <=( (not A167)  and  A168 );
 a109241a <=( A169  and  a109240a );
 a109244a <=( (not A199)  and  A166 );
 a109247a <=( A203  and  (not A200) );
 a109248a <=( a109247a  and  a109244a );
 a109249a <=( a109248a  and  a109241a );
 a109252a <=( A266  and  A265 );
 a109255a <=( (not A268)  and  (not A267) );
 a109256a <=( a109255a  and  a109252a );
 a109259a <=( A299  and  A298 );
 a109262a <=( (not A302)  and  A301 );
 a109263a <=( a109262a  and  a109259a );
 a109264a <=( a109263a  and  a109256a );
 a109268a <=( (not A167)  and  A168 );
 a109269a <=( A169  and  a109268a );
 a109272a <=( (not A199)  and  A166 );
 a109275a <=( A203  and  (not A200) );
 a109276a <=( a109275a  and  a109272a );
 a109277a <=( a109276a  and  a109269a );
 a109280a <=( A266  and  A265 );
 a109283a <=( (not A268)  and  (not A267) );
 a109284a <=( a109283a  and  a109280a );
 a109287a <=( (not A299)  and  A298 );
 a109290a <=( A302  and  (not A301) );
 a109291a <=( a109290a  and  a109287a );
 a109292a <=( a109291a  and  a109284a );
 a109296a <=( (not A167)  and  A168 );
 a109297a <=( A169  and  a109296a );
 a109300a <=( (not A199)  and  A166 );
 a109303a <=( A203  and  (not A200) );
 a109304a <=( a109303a  and  a109300a );
 a109305a <=( a109304a  and  a109297a );
 a109308a <=( A266  and  A265 );
 a109311a <=( (not A268)  and  (not A267) );
 a109312a <=( a109311a  and  a109308a );
 a109315a <=( A299  and  (not A298) );
 a109318a <=( A302  and  (not A301) );
 a109319a <=( a109318a  and  a109315a );
 a109320a <=( a109319a  and  a109312a );
 a109324a <=( (not A167)  and  A168 );
 a109325a <=( A169  and  a109324a );
 a109328a <=( (not A199)  and  A166 );
 a109331a <=( A203  and  (not A200) );
 a109332a <=( a109331a  and  a109328a );
 a109333a <=( a109332a  and  a109325a );
 a109336a <=( A266  and  A265 );
 a109339a <=( (not A268)  and  (not A267) );
 a109340a <=( a109339a  and  a109336a );
 a109343a <=( (not A299)  and  (not A298) );
 a109346a <=( (not A302)  and  A301 );
 a109347a <=( a109346a  and  a109343a );
 a109348a <=( a109347a  and  a109340a );
 a109352a <=( (not A167)  and  A168 );
 a109353a <=( A169  and  a109352a );
 a109356a <=( (not A199)  and  A166 );
 a109359a <=( A203  and  (not A200) );
 a109360a <=( a109359a  and  a109356a );
 a109361a <=( a109360a  and  a109353a );
 a109364a <=( A266  and  A265 );
 a109367a <=( A269  and  (not A267) );
 a109368a <=( a109367a  and  a109364a );
 a109371a <=( A299  and  A298 );
 a109374a <=( (not A302)  and  A301 );
 a109375a <=( a109374a  and  a109371a );
 a109376a <=( a109375a  and  a109368a );
 a109380a <=( (not A167)  and  A168 );
 a109381a <=( A169  and  a109380a );
 a109384a <=( (not A199)  and  A166 );
 a109387a <=( A203  and  (not A200) );
 a109388a <=( a109387a  and  a109384a );
 a109389a <=( a109388a  and  a109381a );
 a109392a <=( A266  and  A265 );
 a109395a <=( A269  and  (not A267) );
 a109396a <=( a109395a  and  a109392a );
 a109399a <=( (not A299)  and  A298 );
 a109402a <=( A302  and  (not A301) );
 a109403a <=( a109402a  and  a109399a );
 a109404a <=( a109403a  and  a109396a );
 a109408a <=( (not A167)  and  A168 );
 a109409a <=( A169  and  a109408a );
 a109412a <=( (not A199)  and  A166 );
 a109415a <=( A203  and  (not A200) );
 a109416a <=( a109415a  and  a109412a );
 a109417a <=( a109416a  and  a109409a );
 a109420a <=( A266  and  A265 );
 a109423a <=( A269  and  (not A267) );
 a109424a <=( a109423a  and  a109420a );
 a109427a <=( A299  and  (not A298) );
 a109430a <=( A302  and  (not A301) );
 a109431a <=( a109430a  and  a109427a );
 a109432a <=( a109431a  and  a109424a );
 a109436a <=( (not A167)  and  A168 );
 a109437a <=( A169  and  a109436a );
 a109440a <=( (not A199)  and  A166 );
 a109443a <=( A203  and  (not A200) );
 a109444a <=( a109443a  and  a109440a );
 a109445a <=( a109444a  and  a109437a );
 a109448a <=( A266  and  A265 );
 a109451a <=( A269  and  (not A267) );
 a109452a <=( a109451a  and  a109448a );
 a109455a <=( (not A299)  and  (not A298) );
 a109458a <=( (not A302)  and  A301 );
 a109459a <=( a109458a  and  a109455a );
 a109460a <=( a109459a  and  a109452a );
 a109464a <=( (not A167)  and  A168 );
 a109465a <=( A169  and  a109464a );
 a109468a <=( (not A199)  and  A166 );
 a109471a <=( A203  and  (not A200) );
 a109472a <=( a109471a  and  a109468a );
 a109473a <=( a109472a  and  a109465a );
 a109476a <=( A266  and  (not A265) );
 a109479a <=( A268  and  (not A267) );
 a109480a <=( a109479a  and  a109476a );
 a109483a <=( A299  and  A298 );
 a109486a <=( (not A302)  and  A301 );
 a109487a <=( a109486a  and  a109483a );
 a109488a <=( a109487a  and  a109480a );
 a109492a <=( (not A167)  and  A168 );
 a109493a <=( A169  and  a109492a );
 a109496a <=( (not A199)  and  A166 );
 a109499a <=( A203  and  (not A200) );
 a109500a <=( a109499a  and  a109496a );
 a109501a <=( a109500a  and  a109493a );
 a109504a <=( A266  and  (not A265) );
 a109507a <=( A268  and  (not A267) );
 a109508a <=( a109507a  and  a109504a );
 a109511a <=( (not A299)  and  A298 );
 a109514a <=( A302  and  (not A301) );
 a109515a <=( a109514a  and  a109511a );
 a109516a <=( a109515a  and  a109508a );
 a109520a <=( (not A167)  and  A168 );
 a109521a <=( A169  and  a109520a );
 a109524a <=( (not A199)  and  A166 );
 a109527a <=( A203  and  (not A200) );
 a109528a <=( a109527a  and  a109524a );
 a109529a <=( a109528a  and  a109521a );
 a109532a <=( A266  and  (not A265) );
 a109535a <=( A268  and  (not A267) );
 a109536a <=( a109535a  and  a109532a );
 a109539a <=( A299  and  (not A298) );
 a109542a <=( A302  and  (not A301) );
 a109543a <=( a109542a  and  a109539a );
 a109544a <=( a109543a  and  a109536a );
 a109548a <=( (not A167)  and  A168 );
 a109549a <=( A169  and  a109548a );
 a109552a <=( (not A199)  and  A166 );
 a109555a <=( A203  and  (not A200) );
 a109556a <=( a109555a  and  a109552a );
 a109557a <=( a109556a  and  a109549a );
 a109560a <=( A266  and  (not A265) );
 a109563a <=( A268  and  (not A267) );
 a109564a <=( a109563a  and  a109560a );
 a109567a <=( (not A299)  and  (not A298) );
 a109570a <=( (not A302)  and  A301 );
 a109571a <=( a109570a  and  a109567a );
 a109572a <=( a109571a  and  a109564a );
 a109576a <=( (not A167)  and  A168 );
 a109577a <=( A169  and  a109576a );
 a109580a <=( (not A199)  and  A166 );
 a109583a <=( A203  and  (not A200) );
 a109584a <=( a109583a  and  a109580a );
 a109585a <=( a109584a  and  a109577a );
 a109588a <=( A266  and  (not A265) );
 a109591a <=( (not A269)  and  (not A267) );
 a109592a <=( a109591a  and  a109588a );
 a109595a <=( A299  and  A298 );
 a109598a <=( (not A302)  and  A301 );
 a109599a <=( a109598a  and  a109595a );
 a109600a <=( a109599a  and  a109592a );
 a109604a <=( (not A167)  and  A168 );
 a109605a <=( A169  and  a109604a );
 a109608a <=( (not A199)  and  A166 );
 a109611a <=( A203  and  (not A200) );
 a109612a <=( a109611a  and  a109608a );
 a109613a <=( a109612a  and  a109605a );
 a109616a <=( A266  and  (not A265) );
 a109619a <=( (not A269)  and  (not A267) );
 a109620a <=( a109619a  and  a109616a );
 a109623a <=( (not A299)  and  A298 );
 a109626a <=( A302  and  (not A301) );
 a109627a <=( a109626a  and  a109623a );
 a109628a <=( a109627a  and  a109620a );
 a109632a <=( (not A167)  and  A168 );
 a109633a <=( A169  and  a109632a );
 a109636a <=( (not A199)  and  A166 );
 a109639a <=( A203  and  (not A200) );
 a109640a <=( a109639a  and  a109636a );
 a109641a <=( a109640a  and  a109633a );
 a109644a <=( A266  and  (not A265) );
 a109647a <=( (not A269)  and  (not A267) );
 a109648a <=( a109647a  and  a109644a );
 a109651a <=( A299  and  (not A298) );
 a109654a <=( A302  and  (not A301) );
 a109655a <=( a109654a  and  a109651a );
 a109656a <=( a109655a  and  a109648a );
 a109660a <=( (not A167)  and  A168 );
 a109661a <=( A169  and  a109660a );
 a109664a <=( (not A199)  and  A166 );
 a109667a <=( A203  and  (not A200) );
 a109668a <=( a109667a  and  a109664a );
 a109669a <=( a109668a  and  a109661a );
 a109672a <=( A266  and  (not A265) );
 a109675a <=( (not A269)  and  (not A267) );
 a109676a <=( a109675a  and  a109672a );
 a109679a <=( (not A299)  and  (not A298) );
 a109682a <=( (not A302)  and  A301 );
 a109683a <=( a109682a  and  a109679a );
 a109684a <=( a109683a  and  a109676a );
 a109688a <=( (not A167)  and  A168 );
 a109689a <=( A169  and  a109688a );
 a109692a <=( (not A199)  and  A166 );
 a109695a <=( A203  and  (not A200) );
 a109696a <=( a109695a  and  a109692a );
 a109697a <=( a109696a  and  a109689a );
 a109700a <=( (not A266)  and  A265 );
 a109703a <=( A268  and  (not A267) );
 a109704a <=( a109703a  and  a109700a );
 a109707a <=( A299  and  A298 );
 a109710a <=( (not A302)  and  A301 );
 a109711a <=( a109710a  and  a109707a );
 a109712a <=( a109711a  and  a109704a );
 a109716a <=( (not A167)  and  A168 );
 a109717a <=( A169  and  a109716a );
 a109720a <=( (not A199)  and  A166 );
 a109723a <=( A203  and  (not A200) );
 a109724a <=( a109723a  and  a109720a );
 a109725a <=( a109724a  and  a109717a );
 a109728a <=( (not A266)  and  A265 );
 a109731a <=( A268  and  (not A267) );
 a109732a <=( a109731a  and  a109728a );
 a109735a <=( (not A299)  and  A298 );
 a109738a <=( A302  and  (not A301) );
 a109739a <=( a109738a  and  a109735a );
 a109740a <=( a109739a  and  a109732a );
 a109744a <=( (not A167)  and  A168 );
 a109745a <=( A169  and  a109744a );
 a109748a <=( (not A199)  and  A166 );
 a109751a <=( A203  and  (not A200) );
 a109752a <=( a109751a  and  a109748a );
 a109753a <=( a109752a  and  a109745a );
 a109756a <=( (not A266)  and  A265 );
 a109759a <=( A268  and  (not A267) );
 a109760a <=( a109759a  and  a109756a );
 a109763a <=( A299  and  (not A298) );
 a109766a <=( A302  and  (not A301) );
 a109767a <=( a109766a  and  a109763a );
 a109768a <=( a109767a  and  a109760a );
 a109772a <=( (not A167)  and  A168 );
 a109773a <=( A169  and  a109772a );
 a109776a <=( (not A199)  and  A166 );
 a109779a <=( A203  and  (not A200) );
 a109780a <=( a109779a  and  a109776a );
 a109781a <=( a109780a  and  a109773a );
 a109784a <=( (not A266)  and  A265 );
 a109787a <=( A268  and  (not A267) );
 a109788a <=( a109787a  and  a109784a );
 a109791a <=( (not A299)  and  (not A298) );
 a109794a <=( (not A302)  and  A301 );
 a109795a <=( a109794a  and  a109791a );
 a109796a <=( a109795a  and  a109788a );
 a109800a <=( (not A167)  and  A168 );
 a109801a <=( A169  and  a109800a );
 a109804a <=( (not A199)  and  A166 );
 a109807a <=( A203  and  (not A200) );
 a109808a <=( a109807a  and  a109804a );
 a109809a <=( a109808a  and  a109801a );
 a109812a <=( (not A266)  and  A265 );
 a109815a <=( (not A269)  and  (not A267) );
 a109816a <=( a109815a  and  a109812a );
 a109819a <=( A299  and  A298 );
 a109822a <=( (not A302)  and  A301 );
 a109823a <=( a109822a  and  a109819a );
 a109824a <=( a109823a  and  a109816a );
 a109828a <=( (not A167)  and  A168 );
 a109829a <=( A169  and  a109828a );
 a109832a <=( (not A199)  and  A166 );
 a109835a <=( A203  and  (not A200) );
 a109836a <=( a109835a  and  a109832a );
 a109837a <=( a109836a  and  a109829a );
 a109840a <=( (not A266)  and  A265 );
 a109843a <=( (not A269)  and  (not A267) );
 a109844a <=( a109843a  and  a109840a );
 a109847a <=( (not A299)  and  A298 );
 a109850a <=( A302  and  (not A301) );
 a109851a <=( a109850a  and  a109847a );
 a109852a <=( a109851a  and  a109844a );
 a109856a <=( (not A167)  and  A168 );
 a109857a <=( A169  and  a109856a );
 a109860a <=( (not A199)  and  A166 );
 a109863a <=( A203  and  (not A200) );
 a109864a <=( a109863a  and  a109860a );
 a109865a <=( a109864a  and  a109857a );
 a109868a <=( (not A266)  and  A265 );
 a109871a <=( (not A269)  and  (not A267) );
 a109872a <=( a109871a  and  a109868a );
 a109875a <=( A299  and  (not A298) );
 a109878a <=( A302  and  (not A301) );
 a109879a <=( a109878a  and  a109875a );
 a109880a <=( a109879a  and  a109872a );
 a109884a <=( (not A167)  and  A168 );
 a109885a <=( A169  and  a109884a );
 a109888a <=( (not A199)  and  A166 );
 a109891a <=( A203  and  (not A200) );
 a109892a <=( a109891a  and  a109888a );
 a109893a <=( a109892a  and  a109885a );
 a109896a <=( (not A266)  and  A265 );
 a109899a <=( (not A269)  and  (not A267) );
 a109900a <=( a109899a  and  a109896a );
 a109903a <=( (not A299)  and  (not A298) );
 a109906a <=( (not A302)  and  A301 );
 a109907a <=( a109906a  and  a109903a );
 a109908a <=( a109907a  and  a109900a );
 a109912a <=( (not A167)  and  A168 );
 a109913a <=( A169  and  a109912a );
 a109916a <=( (not A199)  and  A166 );
 a109919a <=( A202  and  (not A200) );
 a109920a <=( a109919a  and  a109916a );
 a109921a <=( a109920a  and  a109913a );
 a109924a <=( A265  and  (not A203) );
 a109927a <=( A268  and  A266 );
 a109928a <=( a109927a  and  a109924a );
 a109931a <=( (not A298)  and  (not A269) );
 a109934a <=( (not A301)  and  (not A299) );
 a109935a <=( a109934a  and  a109931a );
 a109936a <=( a109935a  and  a109928a );
 a109940a <=( (not A167)  and  A168 );
 a109941a <=( A169  and  a109940a );
 a109944a <=( (not A199)  and  A166 );
 a109947a <=( A202  and  (not A200) );
 a109948a <=( a109947a  and  a109944a );
 a109949a <=( a109948a  and  a109941a );
 a109952a <=( A265  and  (not A203) );
 a109955a <=( A268  and  A266 );
 a109956a <=( a109955a  and  a109952a );
 a109959a <=( (not A298)  and  (not A269) );
 a109962a <=( A302  and  (not A299) );
 a109963a <=( a109962a  and  a109959a );
 a109964a <=( a109963a  and  a109956a );
 a109968a <=( (not A167)  and  A168 );
 a109969a <=( A169  and  a109968a );
 a109972a <=( (not A199)  and  A166 );
 a109975a <=( A202  and  (not A200) );
 a109976a <=( a109975a  and  a109972a );
 a109977a <=( a109976a  and  a109969a );
 a109980a <=( (not A265)  and  (not A203) );
 a109983a <=( (not A268)  and  A266 );
 a109984a <=( a109983a  and  a109980a );
 a109987a <=( (not A298)  and  A269 );
 a109990a <=( (not A301)  and  (not A299) );
 a109991a <=( a109990a  and  a109987a );
 a109992a <=( a109991a  and  a109984a );
 a109996a <=( (not A167)  and  A168 );
 a109997a <=( A169  and  a109996a );
 a110000a <=( (not A199)  and  A166 );
 a110003a <=( A202  and  (not A200) );
 a110004a <=( a110003a  and  a110000a );
 a110005a <=( a110004a  and  a109997a );
 a110008a <=( (not A265)  and  (not A203) );
 a110011a <=( (not A268)  and  A266 );
 a110012a <=( a110011a  and  a110008a );
 a110015a <=( (not A298)  and  A269 );
 a110018a <=( A302  and  (not A299) );
 a110019a <=( a110018a  and  a110015a );
 a110020a <=( a110019a  and  a110012a );
 a110024a <=( (not A167)  and  A168 );
 a110025a <=( A169  and  a110024a );
 a110028a <=( (not A199)  and  A166 );
 a110031a <=( A202  and  (not A200) );
 a110032a <=( a110031a  and  a110028a );
 a110033a <=( a110032a  and  a110025a );
 a110036a <=( A265  and  (not A203) );
 a110039a <=( (not A268)  and  (not A266) );
 a110040a <=( a110039a  and  a110036a );
 a110043a <=( (not A298)  and  A269 );
 a110046a <=( (not A301)  and  (not A299) );
 a110047a <=( a110046a  and  a110043a );
 a110048a <=( a110047a  and  a110040a );
 a110052a <=( (not A167)  and  A168 );
 a110053a <=( A169  and  a110052a );
 a110056a <=( (not A199)  and  A166 );
 a110059a <=( A202  and  (not A200) );
 a110060a <=( a110059a  and  a110056a );
 a110061a <=( a110060a  and  a110053a );
 a110064a <=( A265  and  (not A203) );
 a110067a <=( (not A268)  and  (not A266) );
 a110068a <=( a110067a  and  a110064a );
 a110071a <=( (not A298)  and  A269 );
 a110074a <=( A302  and  (not A299) );
 a110075a <=( a110074a  and  a110071a );
 a110076a <=( a110075a  and  a110068a );
 a110080a <=( (not A167)  and  A168 );
 a110081a <=( A169  and  a110080a );
 a110084a <=( (not A199)  and  A166 );
 a110087a <=( A202  and  (not A200) );
 a110088a <=( a110087a  and  a110084a );
 a110089a <=( a110088a  and  a110081a );
 a110092a <=( (not A265)  and  (not A203) );
 a110095a <=( A268  and  (not A266) );
 a110096a <=( a110095a  and  a110092a );
 a110099a <=( (not A298)  and  (not A269) );
 a110102a <=( (not A301)  and  (not A299) );
 a110103a <=( a110102a  and  a110099a );
 a110104a <=( a110103a  and  a110096a );
 a110108a <=( (not A167)  and  A168 );
 a110109a <=( A169  and  a110108a );
 a110112a <=( (not A199)  and  A166 );
 a110115a <=( A202  and  (not A200) );
 a110116a <=( a110115a  and  a110112a );
 a110117a <=( a110116a  and  a110109a );
 a110120a <=( (not A265)  and  (not A203) );
 a110123a <=( A268  and  (not A266) );
 a110124a <=( a110123a  and  a110120a );
 a110127a <=( (not A298)  and  (not A269) );
 a110130a <=( A302  and  (not A299) );
 a110131a <=( a110130a  and  a110127a );
 a110132a <=( a110131a  and  a110124a );
 a110136a <=( (not A167)  and  (not A169) );
 a110137a <=( (not A170)  and  a110136a );
 a110140a <=( A200  and  A199 );
 a110143a <=( (not A203)  and  A202 );
 a110144a <=( a110143a  and  a110140a );
 a110145a <=( a110144a  and  a110137a );
 a110148a <=( A266  and  A265 );
 a110151a <=( (not A268)  and  (not A267) );
 a110152a <=( a110151a  and  a110148a );
 a110155a <=( A299  and  A298 );
 a110158a <=( (not A302)  and  A301 );
 a110159a <=( a110158a  and  a110155a );
 a110160a <=( a110159a  and  a110152a );
 a110164a <=( (not A167)  and  (not A169) );
 a110165a <=( (not A170)  and  a110164a );
 a110168a <=( A200  and  A199 );
 a110171a <=( (not A203)  and  A202 );
 a110172a <=( a110171a  and  a110168a );
 a110173a <=( a110172a  and  a110165a );
 a110176a <=( A266  and  A265 );
 a110179a <=( (not A268)  and  (not A267) );
 a110180a <=( a110179a  and  a110176a );
 a110183a <=( (not A299)  and  A298 );
 a110186a <=( A302  and  (not A301) );
 a110187a <=( a110186a  and  a110183a );
 a110188a <=( a110187a  and  a110180a );
 a110192a <=( (not A167)  and  (not A169) );
 a110193a <=( (not A170)  and  a110192a );
 a110196a <=( A200  and  A199 );
 a110199a <=( (not A203)  and  A202 );
 a110200a <=( a110199a  and  a110196a );
 a110201a <=( a110200a  and  a110193a );
 a110204a <=( A266  and  A265 );
 a110207a <=( (not A268)  and  (not A267) );
 a110208a <=( a110207a  and  a110204a );
 a110211a <=( A299  and  (not A298) );
 a110214a <=( A302  and  (not A301) );
 a110215a <=( a110214a  and  a110211a );
 a110216a <=( a110215a  and  a110208a );
 a110220a <=( (not A167)  and  (not A169) );
 a110221a <=( (not A170)  and  a110220a );
 a110224a <=( A200  and  A199 );
 a110227a <=( (not A203)  and  A202 );
 a110228a <=( a110227a  and  a110224a );
 a110229a <=( a110228a  and  a110221a );
 a110232a <=( A266  and  A265 );
 a110235a <=( (not A268)  and  (not A267) );
 a110236a <=( a110235a  and  a110232a );
 a110239a <=( (not A299)  and  (not A298) );
 a110242a <=( (not A302)  and  A301 );
 a110243a <=( a110242a  and  a110239a );
 a110244a <=( a110243a  and  a110236a );
 a110248a <=( (not A167)  and  (not A169) );
 a110249a <=( (not A170)  and  a110248a );
 a110252a <=( A200  and  A199 );
 a110255a <=( (not A203)  and  A202 );
 a110256a <=( a110255a  and  a110252a );
 a110257a <=( a110256a  and  a110249a );
 a110260a <=( A266  and  A265 );
 a110263a <=( A269  and  (not A267) );
 a110264a <=( a110263a  and  a110260a );
 a110267a <=( A299  and  A298 );
 a110270a <=( (not A302)  and  A301 );
 a110271a <=( a110270a  and  a110267a );
 a110272a <=( a110271a  and  a110264a );
 a110276a <=( (not A167)  and  (not A169) );
 a110277a <=( (not A170)  and  a110276a );
 a110280a <=( A200  and  A199 );
 a110283a <=( (not A203)  and  A202 );
 a110284a <=( a110283a  and  a110280a );
 a110285a <=( a110284a  and  a110277a );
 a110288a <=( A266  and  A265 );
 a110291a <=( A269  and  (not A267) );
 a110292a <=( a110291a  and  a110288a );
 a110295a <=( (not A299)  and  A298 );
 a110298a <=( A302  and  (not A301) );
 a110299a <=( a110298a  and  a110295a );
 a110300a <=( a110299a  and  a110292a );
 a110304a <=( (not A167)  and  (not A169) );
 a110305a <=( (not A170)  and  a110304a );
 a110308a <=( A200  and  A199 );
 a110311a <=( (not A203)  and  A202 );
 a110312a <=( a110311a  and  a110308a );
 a110313a <=( a110312a  and  a110305a );
 a110316a <=( A266  and  A265 );
 a110319a <=( A269  and  (not A267) );
 a110320a <=( a110319a  and  a110316a );
 a110323a <=( A299  and  (not A298) );
 a110326a <=( A302  and  (not A301) );
 a110327a <=( a110326a  and  a110323a );
 a110328a <=( a110327a  and  a110320a );
 a110332a <=( (not A167)  and  (not A169) );
 a110333a <=( (not A170)  and  a110332a );
 a110336a <=( A200  and  A199 );
 a110339a <=( (not A203)  and  A202 );
 a110340a <=( a110339a  and  a110336a );
 a110341a <=( a110340a  and  a110333a );
 a110344a <=( A266  and  A265 );
 a110347a <=( A269  and  (not A267) );
 a110348a <=( a110347a  and  a110344a );
 a110351a <=( (not A299)  and  (not A298) );
 a110354a <=( (not A302)  and  A301 );
 a110355a <=( a110354a  and  a110351a );
 a110356a <=( a110355a  and  a110348a );
 a110360a <=( (not A167)  and  (not A169) );
 a110361a <=( (not A170)  and  a110360a );
 a110364a <=( A200  and  A199 );
 a110367a <=( (not A203)  and  A202 );
 a110368a <=( a110367a  and  a110364a );
 a110369a <=( a110368a  and  a110361a );
 a110372a <=( A266  and  (not A265) );
 a110375a <=( A268  and  (not A267) );
 a110376a <=( a110375a  and  a110372a );
 a110379a <=( A299  and  A298 );
 a110382a <=( (not A302)  and  A301 );
 a110383a <=( a110382a  and  a110379a );
 a110384a <=( a110383a  and  a110376a );
 a110388a <=( (not A167)  and  (not A169) );
 a110389a <=( (not A170)  and  a110388a );
 a110392a <=( A200  and  A199 );
 a110395a <=( (not A203)  and  A202 );
 a110396a <=( a110395a  and  a110392a );
 a110397a <=( a110396a  and  a110389a );
 a110400a <=( A266  and  (not A265) );
 a110403a <=( A268  and  (not A267) );
 a110404a <=( a110403a  and  a110400a );
 a110407a <=( (not A299)  and  A298 );
 a110410a <=( A302  and  (not A301) );
 a110411a <=( a110410a  and  a110407a );
 a110412a <=( a110411a  and  a110404a );
 a110416a <=( (not A167)  and  (not A169) );
 a110417a <=( (not A170)  and  a110416a );
 a110420a <=( A200  and  A199 );
 a110423a <=( (not A203)  and  A202 );
 a110424a <=( a110423a  and  a110420a );
 a110425a <=( a110424a  and  a110417a );
 a110428a <=( A266  and  (not A265) );
 a110431a <=( A268  and  (not A267) );
 a110432a <=( a110431a  and  a110428a );
 a110435a <=( A299  and  (not A298) );
 a110438a <=( A302  and  (not A301) );
 a110439a <=( a110438a  and  a110435a );
 a110440a <=( a110439a  and  a110432a );
 a110444a <=( (not A167)  and  (not A169) );
 a110445a <=( (not A170)  and  a110444a );
 a110448a <=( A200  and  A199 );
 a110451a <=( (not A203)  and  A202 );
 a110452a <=( a110451a  and  a110448a );
 a110453a <=( a110452a  and  a110445a );
 a110456a <=( A266  and  (not A265) );
 a110459a <=( A268  and  (not A267) );
 a110460a <=( a110459a  and  a110456a );
 a110463a <=( (not A299)  and  (not A298) );
 a110466a <=( (not A302)  and  A301 );
 a110467a <=( a110466a  and  a110463a );
 a110468a <=( a110467a  and  a110460a );
 a110472a <=( (not A167)  and  (not A169) );
 a110473a <=( (not A170)  and  a110472a );
 a110476a <=( A200  and  A199 );
 a110479a <=( (not A203)  and  A202 );
 a110480a <=( a110479a  and  a110476a );
 a110481a <=( a110480a  and  a110473a );
 a110484a <=( A266  and  (not A265) );
 a110487a <=( (not A269)  and  (not A267) );
 a110488a <=( a110487a  and  a110484a );
 a110491a <=( A299  and  A298 );
 a110494a <=( (not A302)  and  A301 );
 a110495a <=( a110494a  and  a110491a );
 a110496a <=( a110495a  and  a110488a );
 a110500a <=( (not A167)  and  (not A169) );
 a110501a <=( (not A170)  and  a110500a );
 a110504a <=( A200  and  A199 );
 a110507a <=( (not A203)  and  A202 );
 a110508a <=( a110507a  and  a110504a );
 a110509a <=( a110508a  and  a110501a );
 a110512a <=( A266  and  (not A265) );
 a110515a <=( (not A269)  and  (not A267) );
 a110516a <=( a110515a  and  a110512a );
 a110519a <=( (not A299)  and  A298 );
 a110522a <=( A302  and  (not A301) );
 a110523a <=( a110522a  and  a110519a );
 a110524a <=( a110523a  and  a110516a );
 a110528a <=( (not A167)  and  (not A169) );
 a110529a <=( (not A170)  and  a110528a );
 a110532a <=( A200  and  A199 );
 a110535a <=( (not A203)  and  A202 );
 a110536a <=( a110535a  and  a110532a );
 a110537a <=( a110536a  and  a110529a );
 a110540a <=( A266  and  (not A265) );
 a110543a <=( (not A269)  and  (not A267) );
 a110544a <=( a110543a  and  a110540a );
 a110547a <=( A299  and  (not A298) );
 a110550a <=( A302  and  (not A301) );
 a110551a <=( a110550a  and  a110547a );
 a110552a <=( a110551a  and  a110544a );
 a110556a <=( (not A167)  and  (not A169) );
 a110557a <=( (not A170)  and  a110556a );
 a110560a <=( A200  and  A199 );
 a110563a <=( (not A203)  and  A202 );
 a110564a <=( a110563a  and  a110560a );
 a110565a <=( a110564a  and  a110557a );
 a110568a <=( A266  and  (not A265) );
 a110571a <=( (not A269)  and  (not A267) );
 a110572a <=( a110571a  and  a110568a );
 a110575a <=( (not A299)  and  (not A298) );
 a110578a <=( (not A302)  and  A301 );
 a110579a <=( a110578a  and  a110575a );
 a110580a <=( a110579a  and  a110572a );
 a110584a <=( (not A167)  and  (not A169) );
 a110585a <=( (not A170)  and  a110584a );
 a110588a <=( A200  and  A199 );
 a110591a <=( (not A203)  and  A202 );
 a110592a <=( a110591a  and  a110588a );
 a110593a <=( a110592a  and  a110585a );
 a110596a <=( (not A266)  and  A265 );
 a110599a <=( A268  and  (not A267) );
 a110600a <=( a110599a  and  a110596a );
 a110603a <=( A299  and  A298 );
 a110606a <=( (not A302)  and  A301 );
 a110607a <=( a110606a  and  a110603a );
 a110608a <=( a110607a  and  a110600a );
 a110612a <=( (not A167)  and  (not A169) );
 a110613a <=( (not A170)  and  a110612a );
 a110616a <=( A200  and  A199 );
 a110619a <=( (not A203)  and  A202 );
 a110620a <=( a110619a  and  a110616a );
 a110621a <=( a110620a  and  a110613a );
 a110624a <=( (not A266)  and  A265 );
 a110627a <=( A268  and  (not A267) );
 a110628a <=( a110627a  and  a110624a );
 a110631a <=( (not A299)  and  A298 );
 a110634a <=( A302  and  (not A301) );
 a110635a <=( a110634a  and  a110631a );
 a110636a <=( a110635a  and  a110628a );
 a110640a <=( (not A167)  and  (not A169) );
 a110641a <=( (not A170)  and  a110640a );
 a110644a <=( A200  and  A199 );
 a110647a <=( (not A203)  and  A202 );
 a110648a <=( a110647a  and  a110644a );
 a110649a <=( a110648a  and  a110641a );
 a110652a <=( (not A266)  and  A265 );
 a110655a <=( A268  and  (not A267) );
 a110656a <=( a110655a  and  a110652a );
 a110659a <=( A299  and  (not A298) );
 a110662a <=( A302  and  (not A301) );
 a110663a <=( a110662a  and  a110659a );
 a110664a <=( a110663a  and  a110656a );
 a110668a <=( (not A167)  and  (not A169) );
 a110669a <=( (not A170)  and  a110668a );
 a110672a <=( A200  and  A199 );
 a110675a <=( (not A203)  and  A202 );
 a110676a <=( a110675a  and  a110672a );
 a110677a <=( a110676a  and  a110669a );
 a110680a <=( (not A266)  and  A265 );
 a110683a <=( A268  and  (not A267) );
 a110684a <=( a110683a  and  a110680a );
 a110687a <=( (not A299)  and  (not A298) );
 a110690a <=( (not A302)  and  A301 );
 a110691a <=( a110690a  and  a110687a );
 a110692a <=( a110691a  and  a110684a );
 a110696a <=( (not A167)  and  (not A169) );
 a110697a <=( (not A170)  and  a110696a );
 a110700a <=( A200  and  A199 );
 a110703a <=( (not A203)  and  A202 );
 a110704a <=( a110703a  and  a110700a );
 a110705a <=( a110704a  and  a110697a );
 a110708a <=( (not A266)  and  A265 );
 a110711a <=( (not A269)  and  (not A267) );
 a110712a <=( a110711a  and  a110708a );
 a110715a <=( A299  and  A298 );
 a110718a <=( (not A302)  and  A301 );
 a110719a <=( a110718a  and  a110715a );
 a110720a <=( a110719a  and  a110712a );
 a110724a <=( (not A167)  and  (not A169) );
 a110725a <=( (not A170)  and  a110724a );
 a110728a <=( A200  and  A199 );
 a110731a <=( (not A203)  and  A202 );
 a110732a <=( a110731a  and  a110728a );
 a110733a <=( a110732a  and  a110725a );
 a110736a <=( (not A266)  and  A265 );
 a110739a <=( (not A269)  and  (not A267) );
 a110740a <=( a110739a  and  a110736a );
 a110743a <=( (not A299)  and  A298 );
 a110746a <=( A302  and  (not A301) );
 a110747a <=( a110746a  and  a110743a );
 a110748a <=( a110747a  and  a110740a );
 a110752a <=( (not A167)  and  (not A169) );
 a110753a <=( (not A170)  and  a110752a );
 a110756a <=( A200  and  A199 );
 a110759a <=( (not A203)  and  A202 );
 a110760a <=( a110759a  and  a110756a );
 a110761a <=( a110760a  and  a110753a );
 a110764a <=( (not A266)  and  A265 );
 a110767a <=( (not A269)  and  (not A267) );
 a110768a <=( a110767a  and  a110764a );
 a110771a <=( A299  and  (not A298) );
 a110774a <=( A302  and  (not A301) );
 a110775a <=( a110774a  and  a110771a );
 a110776a <=( a110775a  and  a110768a );
 a110780a <=( (not A167)  and  (not A169) );
 a110781a <=( (not A170)  and  a110780a );
 a110784a <=( A200  and  A199 );
 a110787a <=( (not A203)  and  A202 );
 a110788a <=( a110787a  and  a110784a );
 a110789a <=( a110788a  and  a110781a );
 a110792a <=( (not A266)  and  A265 );
 a110795a <=( (not A269)  and  (not A267) );
 a110796a <=( a110795a  and  a110792a );
 a110799a <=( (not A299)  and  (not A298) );
 a110802a <=( (not A302)  and  A301 );
 a110803a <=( a110802a  and  a110799a );
 a110804a <=( a110803a  and  a110796a );
 a110808a <=( (not A167)  and  (not A169) );
 a110809a <=( (not A170)  and  a110808a );
 a110812a <=( A200  and  A199 );
 a110815a <=( (not A202)  and  (not A201) );
 a110816a <=( a110815a  and  a110812a );
 a110817a <=( a110816a  and  a110809a );
 a110820a <=( A266  and  A265 );
 a110823a <=( (not A269)  and  A268 );
 a110824a <=( a110823a  and  a110820a );
 a110827a <=( A299  and  A298 );
 a110830a <=( (not A301)  and  (not A300) );
 a110831a <=( a110830a  and  a110827a );
 a110832a <=( a110831a  and  a110824a );
 a110836a <=( (not A167)  and  (not A169) );
 a110837a <=( (not A170)  and  a110836a );
 a110840a <=( A200  and  A199 );
 a110843a <=( (not A202)  and  (not A201) );
 a110844a <=( a110843a  and  a110840a );
 a110845a <=( a110844a  and  a110837a );
 a110848a <=( A266  and  A265 );
 a110851a <=( (not A269)  and  A268 );
 a110852a <=( a110851a  and  a110848a );
 a110855a <=( A299  and  A298 );
 a110858a <=( A302  and  (not A300) );
 a110859a <=( a110858a  and  a110855a );
 a110860a <=( a110859a  and  a110852a );
 a110864a <=( (not A167)  and  (not A169) );
 a110865a <=( (not A170)  and  a110864a );
 a110868a <=( A200  and  A199 );
 a110871a <=( (not A202)  and  (not A201) );
 a110872a <=( a110871a  and  a110868a );
 a110873a <=( a110872a  and  a110865a );
 a110876a <=( A266  and  A265 );
 a110879a <=( (not A269)  and  A268 );
 a110880a <=( a110879a  and  a110876a );
 a110883a <=( (not A299)  and  A298 );
 a110886a <=( A301  and  (not A300) );
 a110887a <=( a110886a  and  a110883a );
 a110888a <=( a110887a  and  a110880a );
 a110892a <=( (not A167)  and  (not A169) );
 a110893a <=( (not A170)  and  a110892a );
 a110896a <=( A200  and  A199 );
 a110899a <=( (not A202)  and  (not A201) );
 a110900a <=( a110899a  and  a110896a );
 a110901a <=( a110900a  and  a110893a );
 a110904a <=( A266  and  A265 );
 a110907a <=( (not A269)  and  A268 );
 a110908a <=( a110907a  and  a110904a );
 a110911a <=( (not A299)  and  A298 );
 a110914a <=( (not A302)  and  (not A300) );
 a110915a <=( a110914a  and  a110911a );
 a110916a <=( a110915a  and  a110908a );
 a110920a <=( (not A167)  and  (not A169) );
 a110921a <=( (not A170)  and  a110920a );
 a110924a <=( A200  and  A199 );
 a110927a <=( (not A202)  and  (not A201) );
 a110928a <=( a110927a  and  a110924a );
 a110929a <=( a110928a  and  a110921a );
 a110932a <=( A266  and  A265 );
 a110935a <=( (not A269)  and  A268 );
 a110936a <=( a110935a  and  a110932a );
 a110939a <=( A299  and  (not A298) );
 a110942a <=( A301  and  (not A300) );
 a110943a <=( a110942a  and  a110939a );
 a110944a <=( a110943a  and  a110936a );
 a110948a <=( (not A167)  and  (not A169) );
 a110949a <=( (not A170)  and  a110948a );
 a110952a <=( A200  and  A199 );
 a110955a <=( (not A202)  and  (not A201) );
 a110956a <=( a110955a  and  a110952a );
 a110957a <=( a110956a  and  a110949a );
 a110960a <=( A266  and  A265 );
 a110963a <=( (not A269)  and  A268 );
 a110964a <=( a110963a  and  a110960a );
 a110967a <=( A299  and  (not A298) );
 a110970a <=( (not A302)  and  (not A300) );
 a110971a <=( a110970a  and  a110967a );
 a110972a <=( a110971a  and  a110964a );
 a110976a <=( (not A167)  and  (not A169) );
 a110977a <=( (not A170)  and  a110976a );
 a110980a <=( A200  and  A199 );
 a110983a <=( (not A202)  and  (not A201) );
 a110984a <=( a110983a  and  a110980a );
 a110985a <=( a110984a  and  a110977a );
 a110988a <=( A266  and  (not A265) );
 a110991a <=( A269  and  (not A268) );
 a110992a <=( a110991a  and  a110988a );
 a110995a <=( A299  and  A298 );
 a110998a <=( (not A301)  and  (not A300) );
 a110999a <=( a110998a  and  a110995a );
 a111000a <=( a110999a  and  a110992a );
 a111004a <=( (not A167)  and  (not A169) );
 a111005a <=( (not A170)  and  a111004a );
 a111008a <=( A200  and  A199 );
 a111011a <=( (not A202)  and  (not A201) );
 a111012a <=( a111011a  and  a111008a );
 a111013a <=( a111012a  and  a111005a );
 a111016a <=( A266  and  (not A265) );
 a111019a <=( A269  and  (not A268) );
 a111020a <=( a111019a  and  a111016a );
 a111023a <=( A299  and  A298 );
 a111026a <=( A302  and  (not A300) );
 a111027a <=( a111026a  and  a111023a );
 a111028a <=( a111027a  and  a111020a );
 a111032a <=( (not A167)  and  (not A169) );
 a111033a <=( (not A170)  and  a111032a );
 a111036a <=( A200  and  A199 );
 a111039a <=( (not A202)  and  (not A201) );
 a111040a <=( a111039a  and  a111036a );
 a111041a <=( a111040a  and  a111033a );
 a111044a <=( A266  and  (not A265) );
 a111047a <=( A269  and  (not A268) );
 a111048a <=( a111047a  and  a111044a );
 a111051a <=( (not A299)  and  A298 );
 a111054a <=( A301  and  (not A300) );
 a111055a <=( a111054a  and  a111051a );
 a111056a <=( a111055a  and  a111048a );
 a111060a <=( (not A167)  and  (not A169) );
 a111061a <=( (not A170)  and  a111060a );
 a111064a <=( A200  and  A199 );
 a111067a <=( (not A202)  and  (not A201) );
 a111068a <=( a111067a  and  a111064a );
 a111069a <=( a111068a  and  a111061a );
 a111072a <=( A266  and  (not A265) );
 a111075a <=( A269  and  (not A268) );
 a111076a <=( a111075a  and  a111072a );
 a111079a <=( (not A299)  and  A298 );
 a111082a <=( (not A302)  and  (not A300) );
 a111083a <=( a111082a  and  a111079a );
 a111084a <=( a111083a  and  a111076a );
 a111088a <=( (not A167)  and  (not A169) );
 a111089a <=( (not A170)  and  a111088a );
 a111092a <=( A200  and  A199 );
 a111095a <=( (not A202)  and  (not A201) );
 a111096a <=( a111095a  and  a111092a );
 a111097a <=( a111096a  and  a111089a );
 a111100a <=( A266  and  (not A265) );
 a111103a <=( A269  and  (not A268) );
 a111104a <=( a111103a  and  a111100a );
 a111107a <=( A299  and  (not A298) );
 a111110a <=( A301  and  (not A300) );
 a111111a <=( a111110a  and  a111107a );
 a111112a <=( a111111a  and  a111104a );
 a111116a <=( (not A167)  and  (not A169) );
 a111117a <=( (not A170)  and  a111116a );
 a111120a <=( A200  and  A199 );
 a111123a <=( (not A202)  and  (not A201) );
 a111124a <=( a111123a  and  a111120a );
 a111125a <=( a111124a  and  a111117a );
 a111128a <=( A266  and  (not A265) );
 a111131a <=( A269  and  (not A268) );
 a111132a <=( a111131a  and  a111128a );
 a111135a <=( A299  and  (not A298) );
 a111138a <=( (not A302)  and  (not A300) );
 a111139a <=( a111138a  and  a111135a );
 a111140a <=( a111139a  and  a111132a );
 a111144a <=( (not A167)  and  (not A169) );
 a111145a <=( (not A170)  and  a111144a );
 a111148a <=( A200  and  A199 );
 a111151a <=( (not A202)  and  (not A201) );
 a111152a <=( a111151a  and  a111148a );
 a111153a <=( a111152a  and  a111145a );
 a111156a <=( (not A266)  and  A265 );
 a111159a <=( A269  and  (not A268) );
 a111160a <=( a111159a  and  a111156a );
 a111163a <=( A299  and  A298 );
 a111166a <=( (not A301)  and  (not A300) );
 a111167a <=( a111166a  and  a111163a );
 a111168a <=( a111167a  and  a111160a );
 a111172a <=( (not A167)  and  (not A169) );
 a111173a <=( (not A170)  and  a111172a );
 a111176a <=( A200  and  A199 );
 a111179a <=( (not A202)  and  (not A201) );
 a111180a <=( a111179a  and  a111176a );
 a111181a <=( a111180a  and  a111173a );
 a111184a <=( (not A266)  and  A265 );
 a111187a <=( A269  and  (not A268) );
 a111188a <=( a111187a  and  a111184a );
 a111191a <=( A299  and  A298 );
 a111194a <=( A302  and  (not A300) );
 a111195a <=( a111194a  and  a111191a );
 a111196a <=( a111195a  and  a111188a );
 a111200a <=( (not A167)  and  (not A169) );
 a111201a <=( (not A170)  and  a111200a );
 a111204a <=( A200  and  A199 );
 a111207a <=( (not A202)  and  (not A201) );
 a111208a <=( a111207a  and  a111204a );
 a111209a <=( a111208a  and  a111201a );
 a111212a <=( (not A266)  and  A265 );
 a111215a <=( A269  and  (not A268) );
 a111216a <=( a111215a  and  a111212a );
 a111219a <=( (not A299)  and  A298 );
 a111222a <=( A301  and  (not A300) );
 a111223a <=( a111222a  and  a111219a );
 a111224a <=( a111223a  and  a111216a );
 a111228a <=( (not A167)  and  (not A169) );
 a111229a <=( (not A170)  and  a111228a );
 a111232a <=( A200  and  A199 );
 a111235a <=( (not A202)  and  (not A201) );
 a111236a <=( a111235a  and  a111232a );
 a111237a <=( a111236a  and  a111229a );
 a111240a <=( (not A266)  and  A265 );
 a111243a <=( A269  and  (not A268) );
 a111244a <=( a111243a  and  a111240a );
 a111247a <=( (not A299)  and  A298 );
 a111250a <=( (not A302)  and  (not A300) );
 a111251a <=( a111250a  and  a111247a );
 a111252a <=( a111251a  and  a111244a );
 a111256a <=( (not A167)  and  (not A169) );
 a111257a <=( (not A170)  and  a111256a );
 a111260a <=( A200  and  A199 );
 a111263a <=( (not A202)  and  (not A201) );
 a111264a <=( a111263a  and  a111260a );
 a111265a <=( a111264a  and  a111257a );
 a111268a <=( (not A266)  and  A265 );
 a111271a <=( A269  and  (not A268) );
 a111272a <=( a111271a  and  a111268a );
 a111275a <=( A299  and  (not A298) );
 a111278a <=( A301  and  (not A300) );
 a111279a <=( a111278a  and  a111275a );
 a111280a <=( a111279a  and  a111272a );
 a111284a <=( (not A167)  and  (not A169) );
 a111285a <=( (not A170)  and  a111284a );
 a111288a <=( A200  and  A199 );
 a111291a <=( (not A202)  and  (not A201) );
 a111292a <=( a111291a  and  a111288a );
 a111293a <=( a111292a  and  a111285a );
 a111296a <=( (not A266)  and  A265 );
 a111299a <=( A269  and  (not A268) );
 a111300a <=( a111299a  and  a111296a );
 a111303a <=( A299  and  (not A298) );
 a111306a <=( (not A302)  and  (not A300) );
 a111307a <=( a111306a  and  a111303a );
 a111308a <=( a111307a  and  a111300a );
 a111312a <=( (not A167)  and  (not A169) );
 a111313a <=( (not A170)  and  a111312a );
 a111316a <=( A200  and  A199 );
 a111319a <=( (not A202)  and  (not A201) );
 a111320a <=( a111319a  and  a111316a );
 a111321a <=( a111320a  and  a111313a );
 a111324a <=( (not A266)  and  (not A265) );
 a111327a <=( (not A269)  and  A268 );
 a111328a <=( a111327a  and  a111324a );
 a111331a <=( A299  and  A298 );
 a111334a <=( (not A301)  and  (not A300) );
 a111335a <=( a111334a  and  a111331a );
 a111336a <=( a111335a  and  a111328a );
 a111340a <=( (not A167)  and  (not A169) );
 a111341a <=( (not A170)  and  a111340a );
 a111344a <=( A200  and  A199 );
 a111347a <=( (not A202)  and  (not A201) );
 a111348a <=( a111347a  and  a111344a );
 a111349a <=( a111348a  and  a111341a );
 a111352a <=( (not A266)  and  (not A265) );
 a111355a <=( (not A269)  and  A268 );
 a111356a <=( a111355a  and  a111352a );
 a111359a <=( A299  and  A298 );
 a111362a <=( A302  and  (not A300) );
 a111363a <=( a111362a  and  a111359a );
 a111364a <=( a111363a  and  a111356a );
 a111368a <=( (not A167)  and  (not A169) );
 a111369a <=( (not A170)  and  a111368a );
 a111372a <=( A200  and  A199 );
 a111375a <=( (not A202)  and  (not A201) );
 a111376a <=( a111375a  and  a111372a );
 a111377a <=( a111376a  and  a111369a );
 a111380a <=( (not A266)  and  (not A265) );
 a111383a <=( (not A269)  and  A268 );
 a111384a <=( a111383a  and  a111380a );
 a111387a <=( (not A299)  and  A298 );
 a111390a <=( A301  and  (not A300) );
 a111391a <=( a111390a  and  a111387a );
 a111392a <=( a111391a  and  a111384a );
 a111396a <=( (not A167)  and  (not A169) );
 a111397a <=( (not A170)  and  a111396a );
 a111400a <=( A200  and  A199 );
 a111403a <=( (not A202)  and  (not A201) );
 a111404a <=( a111403a  and  a111400a );
 a111405a <=( a111404a  and  a111397a );
 a111408a <=( (not A266)  and  (not A265) );
 a111411a <=( (not A269)  and  A268 );
 a111412a <=( a111411a  and  a111408a );
 a111415a <=( (not A299)  and  A298 );
 a111418a <=( (not A302)  and  (not A300) );
 a111419a <=( a111418a  and  a111415a );
 a111420a <=( a111419a  and  a111412a );
 a111424a <=( (not A167)  and  (not A169) );
 a111425a <=( (not A170)  and  a111424a );
 a111428a <=( A200  and  A199 );
 a111431a <=( (not A202)  and  (not A201) );
 a111432a <=( a111431a  and  a111428a );
 a111433a <=( a111432a  and  a111425a );
 a111436a <=( (not A266)  and  (not A265) );
 a111439a <=( (not A269)  and  A268 );
 a111440a <=( a111439a  and  a111436a );
 a111443a <=( A299  and  (not A298) );
 a111446a <=( A301  and  (not A300) );
 a111447a <=( a111446a  and  a111443a );
 a111448a <=( a111447a  and  a111440a );
 a111452a <=( (not A167)  and  (not A169) );
 a111453a <=( (not A170)  and  a111452a );
 a111456a <=( A200  and  A199 );
 a111459a <=( (not A202)  and  (not A201) );
 a111460a <=( a111459a  and  a111456a );
 a111461a <=( a111460a  and  a111453a );
 a111464a <=( (not A266)  and  (not A265) );
 a111467a <=( (not A269)  and  A268 );
 a111468a <=( a111467a  and  a111464a );
 a111471a <=( A299  and  (not A298) );
 a111474a <=( (not A302)  and  (not A300) );
 a111475a <=( a111474a  and  a111471a );
 a111476a <=( a111475a  and  a111468a );
 a111480a <=( (not A167)  and  (not A169) );
 a111481a <=( (not A170)  and  a111480a );
 a111484a <=( A200  and  A199 );
 a111487a <=( A203  and  (not A201) );
 a111488a <=( a111487a  and  a111484a );
 a111489a <=( a111488a  and  a111481a );
 a111492a <=( A266  and  A265 );
 a111495a <=( (not A269)  and  A268 );
 a111496a <=( a111495a  and  a111492a );
 a111499a <=( A299  and  A298 );
 a111502a <=( (not A301)  and  (not A300) );
 a111503a <=( a111502a  and  a111499a );
 a111504a <=( a111503a  and  a111496a );
 a111508a <=( (not A167)  and  (not A169) );
 a111509a <=( (not A170)  and  a111508a );
 a111512a <=( A200  and  A199 );
 a111515a <=( A203  and  (not A201) );
 a111516a <=( a111515a  and  a111512a );
 a111517a <=( a111516a  and  a111509a );
 a111520a <=( A266  and  A265 );
 a111523a <=( (not A269)  and  A268 );
 a111524a <=( a111523a  and  a111520a );
 a111527a <=( A299  and  A298 );
 a111530a <=( A302  and  (not A300) );
 a111531a <=( a111530a  and  a111527a );
 a111532a <=( a111531a  and  a111524a );
 a111536a <=( (not A167)  and  (not A169) );
 a111537a <=( (not A170)  and  a111536a );
 a111540a <=( A200  and  A199 );
 a111543a <=( A203  and  (not A201) );
 a111544a <=( a111543a  and  a111540a );
 a111545a <=( a111544a  and  a111537a );
 a111548a <=( A266  and  A265 );
 a111551a <=( (not A269)  and  A268 );
 a111552a <=( a111551a  and  a111548a );
 a111555a <=( (not A299)  and  A298 );
 a111558a <=( A301  and  (not A300) );
 a111559a <=( a111558a  and  a111555a );
 a111560a <=( a111559a  and  a111552a );
 a111564a <=( (not A167)  and  (not A169) );
 a111565a <=( (not A170)  and  a111564a );
 a111568a <=( A200  and  A199 );
 a111571a <=( A203  and  (not A201) );
 a111572a <=( a111571a  and  a111568a );
 a111573a <=( a111572a  and  a111565a );
 a111576a <=( A266  and  A265 );
 a111579a <=( (not A269)  and  A268 );
 a111580a <=( a111579a  and  a111576a );
 a111583a <=( (not A299)  and  A298 );
 a111586a <=( (not A302)  and  (not A300) );
 a111587a <=( a111586a  and  a111583a );
 a111588a <=( a111587a  and  a111580a );
 a111592a <=( (not A167)  and  (not A169) );
 a111593a <=( (not A170)  and  a111592a );
 a111596a <=( A200  and  A199 );
 a111599a <=( A203  and  (not A201) );
 a111600a <=( a111599a  and  a111596a );
 a111601a <=( a111600a  and  a111593a );
 a111604a <=( A266  and  A265 );
 a111607a <=( (not A269)  and  A268 );
 a111608a <=( a111607a  and  a111604a );
 a111611a <=( A299  and  (not A298) );
 a111614a <=( A301  and  (not A300) );
 a111615a <=( a111614a  and  a111611a );
 a111616a <=( a111615a  and  a111608a );
 a111620a <=( (not A167)  and  (not A169) );
 a111621a <=( (not A170)  and  a111620a );
 a111624a <=( A200  and  A199 );
 a111627a <=( A203  and  (not A201) );
 a111628a <=( a111627a  and  a111624a );
 a111629a <=( a111628a  and  a111621a );
 a111632a <=( A266  and  A265 );
 a111635a <=( (not A269)  and  A268 );
 a111636a <=( a111635a  and  a111632a );
 a111639a <=( A299  and  (not A298) );
 a111642a <=( (not A302)  and  (not A300) );
 a111643a <=( a111642a  and  a111639a );
 a111644a <=( a111643a  and  a111636a );
 a111648a <=( (not A167)  and  (not A169) );
 a111649a <=( (not A170)  and  a111648a );
 a111652a <=( A200  and  A199 );
 a111655a <=( A203  and  (not A201) );
 a111656a <=( a111655a  and  a111652a );
 a111657a <=( a111656a  and  a111649a );
 a111660a <=( A266  and  (not A265) );
 a111663a <=( A269  and  (not A268) );
 a111664a <=( a111663a  and  a111660a );
 a111667a <=( A299  and  A298 );
 a111670a <=( (not A301)  and  (not A300) );
 a111671a <=( a111670a  and  a111667a );
 a111672a <=( a111671a  and  a111664a );
 a111676a <=( (not A167)  and  (not A169) );
 a111677a <=( (not A170)  and  a111676a );
 a111680a <=( A200  and  A199 );
 a111683a <=( A203  and  (not A201) );
 a111684a <=( a111683a  and  a111680a );
 a111685a <=( a111684a  and  a111677a );
 a111688a <=( A266  and  (not A265) );
 a111691a <=( A269  and  (not A268) );
 a111692a <=( a111691a  and  a111688a );
 a111695a <=( A299  and  A298 );
 a111698a <=( A302  and  (not A300) );
 a111699a <=( a111698a  and  a111695a );
 a111700a <=( a111699a  and  a111692a );
 a111704a <=( (not A167)  and  (not A169) );
 a111705a <=( (not A170)  and  a111704a );
 a111708a <=( A200  and  A199 );
 a111711a <=( A203  and  (not A201) );
 a111712a <=( a111711a  and  a111708a );
 a111713a <=( a111712a  and  a111705a );
 a111716a <=( A266  and  (not A265) );
 a111719a <=( A269  and  (not A268) );
 a111720a <=( a111719a  and  a111716a );
 a111723a <=( (not A299)  and  A298 );
 a111726a <=( A301  and  (not A300) );
 a111727a <=( a111726a  and  a111723a );
 a111728a <=( a111727a  and  a111720a );
 a111732a <=( (not A167)  and  (not A169) );
 a111733a <=( (not A170)  and  a111732a );
 a111736a <=( A200  and  A199 );
 a111739a <=( A203  and  (not A201) );
 a111740a <=( a111739a  and  a111736a );
 a111741a <=( a111740a  and  a111733a );
 a111744a <=( A266  and  (not A265) );
 a111747a <=( A269  and  (not A268) );
 a111748a <=( a111747a  and  a111744a );
 a111751a <=( (not A299)  and  A298 );
 a111754a <=( (not A302)  and  (not A300) );
 a111755a <=( a111754a  and  a111751a );
 a111756a <=( a111755a  and  a111748a );
 a111760a <=( (not A167)  and  (not A169) );
 a111761a <=( (not A170)  and  a111760a );
 a111764a <=( A200  and  A199 );
 a111767a <=( A203  and  (not A201) );
 a111768a <=( a111767a  and  a111764a );
 a111769a <=( a111768a  and  a111761a );
 a111772a <=( A266  and  (not A265) );
 a111775a <=( A269  and  (not A268) );
 a111776a <=( a111775a  and  a111772a );
 a111779a <=( A299  and  (not A298) );
 a111782a <=( A301  and  (not A300) );
 a111783a <=( a111782a  and  a111779a );
 a111784a <=( a111783a  and  a111776a );
 a111788a <=( (not A167)  and  (not A169) );
 a111789a <=( (not A170)  and  a111788a );
 a111792a <=( A200  and  A199 );
 a111795a <=( A203  and  (not A201) );
 a111796a <=( a111795a  and  a111792a );
 a111797a <=( a111796a  and  a111789a );
 a111800a <=( A266  and  (not A265) );
 a111803a <=( A269  and  (not A268) );
 a111804a <=( a111803a  and  a111800a );
 a111807a <=( A299  and  (not A298) );
 a111810a <=( (not A302)  and  (not A300) );
 a111811a <=( a111810a  and  a111807a );
 a111812a <=( a111811a  and  a111804a );
 a111816a <=( (not A167)  and  (not A169) );
 a111817a <=( (not A170)  and  a111816a );
 a111820a <=( A200  and  A199 );
 a111823a <=( A203  and  (not A201) );
 a111824a <=( a111823a  and  a111820a );
 a111825a <=( a111824a  and  a111817a );
 a111828a <=( (not A266)  and  A265 );
 a111831a <=( A269  and  (not A268) );
 a111832a <=( a111831a  and  a111828a );
 a111835a <=( A299  and  A298 );
 a111838a <=( (not A301)  and  (not A300) );
 a111839a <=( a111838a  and  a111835a );
 a111840a <=( a111839a  and  a111832a );
 a111844a <=( (not A167)  and  (not A169) );
 a111845a <=( (not A170)  and  a111844a );
 a111848a <=( A200  and  A199 );
 a111851a <=( A203  and  (not A201) );
 a111852a <=( a111851a  and  a111848a );
 a111853a <=( a111852a  and  a111845a );
 a111856a <=( (not A266)  and  A265 );
 a111859a <=( A269  and  (not A268) );
 a111860a <=( a111859a  and  a111856a );
 a111863a <=( A299  and  A298 );
 a111866a <=( A302  and  (not A300) );
 a111867a <=( a111866a  and  a111863a );
 a111868a <=( a111867a  and  a111860a );
 a111872a <=( (not A167)  and  (not A169) );
 a111873a <=( (not A170)  and  a111872a );
 a111876a <=( A200  and  A199 );
 a111879a <=( A203  and  (not A201) );
 a111880a <=( a111879a  and  a111876a );
 a111881a <=( a111880a  and  a111873a );
 a111884a <=( (not A266)  and  A265 );
 a111887a <=( A269  and  (not A268) );
 a111888a <=( a111887a  and  a111884a );
 a111891a <=( (not A299)  and  A298 );
 a111894a <=( A301  and  (not A300) );
 a111895a <=( a111894a  and  a111891a );
 a111896a <=( a111895a  and  a111888a );
 a111900a <=( (not A167)  and  (not A169) );
 a111901a <=( (not A170)  and  a111900a );
 a111904a <=( A200  and  A199 );
 a111907a <=( A203  and  (not A201) );
 a111908a <=( a111907a  and  a111904a );
 a111909a <=( a111908a  and  a111901a );
 a111912a <=( (not A266)  and  A265 );
 a111915a <=( A269  and  (not A268) );
 a111916a <=( a111915a  and  a111912a );
 a111919a <=( (not A299)  and  A298 );
 a111922a <=( (not A302)  and  (not A300) );
 a111923a <=( a111922a  and  a111919a );
 a111924a <=( a111923a  and  a111916a );
 a111928a <=( (not A167)  and  (not A169) );
 a111929a <=( (not A170)  and  a111928a );
 a111932a <=( A200  and  A199 );
 a111935a <=( A203  and  (not A201) );
 a111936a <=( a111935a  and  a111932a );
 a111937a <=( a111936a  and  a111929a );
 a111940a <=( (not A266)  and  A265 );
 a111943a <=( A269  and  (not A268) );
 a111944a <=( a111943a  and  a111940a );
 a111947a <=( A299  and  (not A298) );
 a111950a <=( A301  and  (not A300) );
 a111951a <=( a111950a  and  a111947a );
 a111952a <=( a111951a  and  a111944a );
 a111956a <=( (not A167)  and  (not A169) );
 a111957a <=( (not A170)  and  a111956a );
 a111960a <=( A200  and  A199 );
 a111963a <=( A203  and  (not A201) );
 a111964a <=( a111963a  and  a111960a );
 a111965a <=( a111964a  and  a111957a );
 a111968a <=( (not A266)  and  A265 );
 a111971a <=( A269  and  (not A268) );
 a111972a <=( a111971a  and  a111968a );
 a111975a <=( A299  and  (not A298) );
 a111978a <=( (not A302)  and  (not A300) );
 a111979a <=( a111978a  and  a111975a );
 a111980a <=( a111979a  and  a111972a );
 a111984a <=( (not A167)  and  (not A169) );
 a111985a <=( (not A170)  and  a111984a );
 a111988a <=( A200  and  A199 );
 a111991a <=( A203  and  (not A201) );
 a111992a <=( a111991a  and  a111988a );
 a111993a <=( a111992a  and  a111985a );
 a111996a <=( (not A266)  and  (not A265) );
 a111999a <=( (not A269)  and  A268 );
 a112000a <=( a111999a  and  a111996a );
 a112003a <=( A299  and  A298 );
 a112006a <=( (not A301)  and  (not A300) );
 a112007a <=( a112006a  and  a112003a );
 a112008a <=( a112007a  and  a112000a );
 a112012a <=( (not A167)  and  (not A169) );
 a112013a <=( (not A170)  and  a112012a );
 a112016a <=( A200  and  A199 );
 a112019a <=( A203  and  (not A201) );
 a112020a <=( a112019a  and  a112016a );
 a112021a <=( a112020a  and  a112013a );
 a112024a <=( (not A266)  and  (not A265) );
 a112027a <=( (not A269)  and  A268 );
 a112028a <=( a112027a  and  a112024a );
 a112031a <=( A299  and  A298 );
 a112034a <=( A302  and  (not A300) );
 a112035a <=( a112034a  and  a112031a );
 a112036a <=( a112035a  and  a112028a );
 a112040a <=( (not A167)  and  (not A169) );
 a112041a <=( (not A170)  and  a112040a );
 a112044a <=( A200  and  A199 );
 a112047a <=( A203  and  (not A201) );
 a112048a <=( a112047a  and  a112044a );
 a112049a <=( a112048a  and  a112041a );
 a112052a <=( (not A266)  and  (not A265) );
 a112055a <=( (not A269)  and  A268 );
 a112056a <=( a112055a  and  a112052a );
 a112059a <=( (not A299)  and  A298 );
 a112062a <=( A301  and  (not A300) );
 a112063a <=( a112062a  and  a112059a );
 a112064a <=( a112063a  and  a112056a );
 a112068a <=( (not A167)  and  (not A169) );
 a112069a <=( (not A170)  and  a112068a );
 a112072a <=( A200  and  A199 );
 a112075a <=( A203  and  (not A201) );
 a112076a <=( a112075a  and  a112072a );
 a112077a <=( a112076a  and  a112069a );
 a112080a <=( (not A266)  and  (not A265) );
 a112083a <=( (not A269)  and  A268 );
 a112084a <=( a112083a  and  a112080a );
 a112087a <=( (not A299)  and  A298 );
 a112090a <=( (not A302)  and  (not A300) );
 a112091a <=( a112090a  and  a112087a );
 a112092a <=( a112091a  and  a112084a );
 a112096a <=( (not A167)  and  (not A169) );
 a112097a <=( (not A170)  and  a112096a );
 a112100a <=( A200  and  A199 );
 a112103a <=( A203  and  (not A201) );
 a112104a <=( a112103a  and  a112100a );
 a112105a <=( a112104a  and  a112097a );
 a112108a <=( (not A266)  and  (not A265) );
 a112111a <=( (not A269)  and  A268 );
 a112112a <=( a112111a  and  a112108a );
 a112115a <=( A299  and  (not A298) );
 a112118a <=( A301  and  (not A300) );
 a112119a <=( a112118a  and  a112115a );
 a112120a <=( a112119a  and  a112112a );
 a112124a <=( (not A167)  and  (not A169) );
 a112125a <=( (not A170)  and  a112124a );
 a112128a <=( A200  and  A199 );
 a112131a <=( A203  and  (not A201) );
 a112132a <=( a112131a  and  a112128a );
 a112133a <=( a112132a  and  a112125a );
 a112136a <=( (not A266)  and  (not A265) );
 a112139a <=( (not A269)  and  A268 );
 a112140a <=( a112139a  and  a112136a );
 a112143a <=( A299  and  (not A298) );
 a112146a <=( (not A302)  and  (not A300) );
 a112147a <=( a112146a  and  a112143a );
 a112148a <=( a112147a  and  a112140a );
 a112152a <=( (not A167)  and  (not A169) );
 a112153a <=( (not A170)  and  a112152a );
 a112156a <=( A200  and  (not A199) );
 a112159a <=( A203  and  (not A202) );
 a112160a <=( a112159a  and  a112156a );
 a112161a <=( a112160a  and  a112153a );
 a112164a <=( A266  and  A265 );
 a112167a <=( (not A268)  and  (not A267) );
 a112168a <=( a112167a  and  a112164a );
 a112171a <=( A299  and  A298 );
 a112174a <=( (not A302)  and  A301 );
 a112175a <=( a112174a  and  a112171a );
 a112176a <=( a112175a  and  a112168a );
 a112180a <=( (not A167)  and  (not A169) );
 a112181a <=( (not A170)  and  a112180a );
 a112184a <=( A200  and  (not A199) );
 a112187a <=( A203  and  (not A202) );
 a112188a <=( a112187a  and  a112184a );
 a112189a <=( a112188a  and  a112181a );
 a112192a <=( A266  and  A265 );
 a112195a <=( (not A268)  and  (not A267) );
 a112196a <=( a112195a  and  a112192a );
 a112199a <=( (not A299)  and  A298 );
 a112202a <=( A302  and  (not A301) );
 a112203a <=( a112202a  and  a112199a );
 a112204a <=( a112203a  and  a112196a );
 a112208a <=( (not A167)  and  (not A169) );
 a112209a <=( (not A170)  and  a112208a );
 a112212a <=( A200  and  (not A199) );
 a112215a <=( A203  and  (not A202) );
 a112216a <=( a112215a  and  a112212a );
 a112217a <=( a112216a  and  a112209a );
 a112220a <=( A266  and  A265 );
 a112223a <=( (not A268)  and  (not A267) );
 a112224a <=( a112223a  and  a112220a );
 a112227a <=( A299  and  (not A298) );
 a112230a <=( A302  and  (not A301) );
 a112231a <=( a112230a  and  a112227a );
 a112232a <=( a112231a  and  a112224a );
 a112236a <=( (not A167)  and  (not A169) );
 a112237a <=( (not A170)  and  a112236a );
 a112240a <=( A200  and  (not A199) );
 a112243a <=( A203  and  (not A202) );
 a112244a <=( a112243a  and  a112240a );
 a112245a <=( a112244a  and  a112237a );
 a112248a <=( A266  and  A265 );
 a112251a <=( (not A268)  and  (not A267) );
 a112252a <=( a112251a  and  a112248a );
 a112255a <=( (not A299)  and  (not A298) );
 a112258a <=( (not A302)  and  A301 );
 a112259a <=( a112258a  and  a112255a );
 a112260a <=( a112259a  and  a112252a );
 a112264a <=( (not A167)  and  (not A169) );
 a112265a <=( (not A170)  and  a112264a );
 a112268a <=( A200  and  (not A199) );
 a112271a <=( A203  and  (not A202) );
 a112272a <=( a112271a  and  a112268a );
 a112273a <=( a112272a  and  a112265a );
 a112276a <=( A266  and  A265 );
 a112279a <=( A269  and  (not A267) );
 a112280a <=( a112279a  and  a112276a );
 a112283a <=( A299  and  A298 );
 a112286a <=( (not A302)  and  A301 );
 a112287a <=( a112286a  and  a112283a );
 a112288a <=( a112287a  and  a112280a );
 a112292a <=( (not A167)  and  (not A169) );
 a112293a <=( (not A170)  and  a112292a );
 a112296a <=( A200  and  (not A199) );
 a112299a <=( A203  and  (not A202) );
 a112300a <=( a112299a  and  a112296a );
 a112301a <=( a112300a  and  a112293a );
 a112304a <=( A266  and  A265 );
 a112307a <=( A269  and  (not A267) );
 a112308a <=( a112307a  and  a112304a );
 a112311a <=( (not A299)  and  A298 );
 a112314a <=( A302  and  (not A301) );
 a112315a <=( a112314a  and  a112311a );
 a112316a <=( a112315a  and  a112308a );
 a112320a <=( (not A167)  and  (not A169) );
 a112321a <=( (not A170)  and  a112320a );
 a112324a <=( A200  and  (not A199) );
 a112327a <=( A203  and  (not A202) );
 a112328a <=( a112327a  and  a112324a );
 a112329a <=( a112328a  and  a112321a );
 a112332a <=( A266  and  A265 );
 a112335a <=( A269  and  (not A267) );
 a112336a <=( a112335a  and  a112332a );
 a112339a <=( A299  and  (not A298) );
 a112342a <=( A302  and  (not A301) );
 a112343a <=( a112342a  and  a112339a );
 a112344a <=( a112343a  and  a112336a );
 a112348a <=( (not A167)  and  (not A169) );
 a112349a <=( (not A170)  and  a112348a );
 a112352a <=( A200  and  (not A199) );
 a112355a <=( A203  and  (not A202) );
 a112356a <=( a112355a  and  a112352a );
 a112357a <=( a112356a  and  a112349a );
 a112360a <=( A266  and  A265 );
 a112363a <=( A269  and  (not A267) );
 a112364a <=( a112363a  and  a112360a );
 a112367a <=( (not A299)  and  (not A298) );
 a112370a <=( (not A302)  and  A301 );
 a112371a <=( a112370a  and  a112367a );
 a112372a <=( a112371a  and  a112364a );
 a112376a <=( (not A167)  and  (not A169) );
 a112377a <=( (not A170)  and  a112376a );
 a112380a <=( A200  and  (not A199) );
 a112383a <=( A203  and  (not A202) );
 a112384a <=( a112383a  and  a112380a );
 a112385a <=( a112384a  and  a112377a );
 a112388a <=( A266  and  (not A265) );
 a112391a <=( A268  and  (not A267) );
 a112392a <=( a112391a  and  a112388a );
 a112395a <=( A299  and  A298 );
 a112398a <=( (not A302)  and  A301 );
 a112399a <=( a112398a  and  a112395a );
 a112400a <=( a112399a  and  a112392a );
 a112404a <=( (not A167)  and  (not A169) );
 a112405a <=( (not A170)  and  a112404a );
 a112408a <=( A200  and  (not A199) );
 a112411a <=( A203  and  (not A202) );
 a112412a <=( a112411a  and  a112408a );
 a112413a <=( a112412a  and  a112405a );
 a112416a <=( A266  and  (not A265) );
 a112419a <=( A268  and  (not A267) );
 a112420a <=( a112419a  and  a112416a );
 a112423a <=( (not A299)  and  A298 );
 a112426a <=( A302  and  (not A301) );
 a112427a <=( a112426a  and  a112423a );
 a112428a <=( a112427a  and  a112420a );
 a112432a <=( (not A167)  and  (not A169) );
 a112433a <=( (not A170)  and  a112432a );
 a112436a <=( A200  and  (not A199) );
 a112439a <=( A203  and  (not A202) );
 a112440a <=( a112439a  and  a112436a );
 a112441a <=( a112440a  and  a112433a );
 a112444a <=( A266  and  (not A265) );
 a112447a <=( A268  and  (not A267) );
 a112448a <=( a112447a  and  a112444a );
 a112451a <=( A299  and  (not A298) );
 a112454a <=( A302  and  (not A301) );
 a112455a <=( a112454a  and  a112451a );
 a112456a <=( a112455a  and  a112448a );
 a112460a <=( (not A167)  and  (not A169) );
 a112461a <=( (not A170)  and  a112460a );
 a112464a <=( A200  and  (not A199) );
 a112467a <=( A203  and  (not A202) );
 a112468a <=( a112467a  and  a112464a );
 a112469a <=( a112468a  and  a112461a );
 a112472a <=( A266  and  (not A265) );
 a112475a <=( A268  and  (not A267) );
 a112476a <=( a112475a  and  a112472a );
 a112479a <=( (not A299)  and  (not A298) );
 a112482a <=( (not A302)  and  A301 );
 a112483a <=( a112482a  and  a112479a );
 a112484a <=( a112483a  and  a112476a );
 a112488a <=( (not A167)  and  (not A169) );
 a112489a <=( (not A170)  and  a112488a );
 a112492a <=( A200  and  (not A199) );
 a112495a <=( A203  and  (not A202) );
 a112496a <=( a112495a  and  a112492a );
 a112497a <=( a112496a  and  a112489a );
 a112500a <=( A266  and  (not A265) );
 a112503a <=( (not A269)  and  (not A267) );
 a112504a <=( a112503a  and  a112500a );
 a112507a <=( A299  and  A298 );
 a112510a <=( (not A302)  and  A301 );
 a112511a <=( a112510a  and  a112507a );
 a112512a <=( a112511a  and  a112504a );
 a112516a <=( (not A167)  and  (not A169) );
 a112517a <=( (not A170)  and  a112516a );
 a112520a <=( A200  and  (not A199) );
 a112523a <=( A203  and  (not A202) );
 a112524a <=( a112523a  and  a112520a );
 a112525a <=( a112524a  and  a112517a );
 a112528a <=( A266  and  (not A265) );
 a112531a <=( (not A269)  and  (not A267) );
 a112532a <=( a112531a  and  a112528a );
 a112535a <=( (not A299)  and  A298 );
 a112538a <=( A302  and  (not A301) );
 a112539a <=( a112538a  and  a112535a );
 a112540a <=( a112539a  and  a112532a );
 a112544a <=( (not A167)  and  (not A169) );
 a112545a <=( (not A170)  and  a112544a );
 a112548a <=( A200  and  (not A199) );
 a112551a <=( A203  and  (not A202) );
 a112552a <=( a112551a  and  a112548a );
 a112553a <=( a112552a  and  a112545a );
 a112556a <=( A266  and  (not A265) );
 a112559a <=( (not A269)  and  (not A267) );
 a112560a <=( a112559a  and  a112556a );
 a112563a <=( A299  and  (not A298) );
 a112566a <=( A302  and  (not A301) );
 a112567a <=( a112566a  and  a112563a );
 a112568a <=( a112567a  and  a112560a );
 a112572a <=( (not A167)  and  (not A169) );
 a112573a <=( (not A170)  and  a112572a );
 a112576a <=( A200  and  (not A199) );
 a112579a <=( A203  and  (not A202) );
 a112580a <=( a112579a  and  a112576a );
 a112581a <=( a112580a  and  a112573a );
 a112584a <=( A266  and  (not A265) );
 a112587a <=( (not A269)  and  (not A267) );
 a112588a <=( a112587a  and  a112584a );
 a112591a <=( (not A299)  and  (not A298) );
 a112594a <=( (not A302)  and  A301 );
 a112595a <=( a112594a  and  a112591a );
 a112596a <=( a112595a  and  a112588a );
 a112600a <=( (not A167)  and  (not A169) );
 a112601a <=( (not A170)  and  a112600a );
 a112604a <=( A200  and  (not A199) );
 a112607a <=( A203  and  (not A202) );
 a112608a <=( a112607a  and  a112604a );
 a112609a <=( a112608a  and  a112601a );
 a112612a <=( (not A266)  and  A265 );
 a112615a <=( A268  and  (not A267) );
 a112616a <=( a112615a  and  a112612a );
 a112619a <=( A299  and  A298 );
 a112622a <=( (not A302)  and  A301 );
 a112623a <=( a112622a  and  a112619a );
 a112624a <=( a112623a  and  a112616a );
 a112628a <=( (not A167)  and  (not A169) );
 a112629a <=( (not A170)  and  a112628a );
 a112632a <=( A200  and  (not A199) );
 a112635a <=( A203  and  (not A202) );
 a112636a <=( a112635a  and  a112632a );
 a112637a <=( a112636a  and  a112629a );
 a112640a <=( (not A266)  and  A265 );
 a112643a <=( A268  and  (not A267) );
 a112644a <=( a112643a  and  a112640a );
 a112647a <=( (not A299)  and  A298 );
 a112650a <=( A302  and  (not A301) );
 a112651a <=( a112650a  and  a112647a );
 a112652a <=( a112651a  and  a112644a );
 a112656a <=( (not A167)  and  (not A169) );
 a112657a <=( (not A170)  and  a112656a );
 a112660a <=( A200  and  (not A199) );
 a112663a <=( A203  and  (not A202) );
 a112664a <=( a112663a  and  a112660a );
 a112665a <=( a112664a  and  a112657a );
 a112668a <=( (not A266)  and  A265 );
 a112671a <=( A268  and  (not A267) );
 a112672a <=( a112671a  and  a112668a );
 a112675a <=( A299  and  (not A298) );
 a112678a <=( A302  and  (not A301) );
 a112679a <=( a112678a  and  a112675a );
 a112680a <=( a112679a  and  a112672a );
 a112684a <=( (not A167)  and  (not A169) );
 a112685a <=( (not A170)  and  a112684a );
 a112688a <=( A200  and  (not A199) );
 a112691a <=( A203  and  (not A202) );
 a112692a <=( a112691a  and  a112688a );
 a112693a <=( a112692a  and  a112685a );
 a112696a <=( (not A266)  and  A265 );
 a112699a <=( A268  and  (not A267) );
 a112700a <=( a112699a  and  a112696a );
 a112703a <=( (not A299)  and  (not A298) );
 a112706a <=( (not A302)  and  A301 );
 a112707a <=( a112706a  and  a112703a );
 a112708a <=( a112707a  and  a112700a );
 a112712a <=( (not A167)  and  (not A169) );
 a112713a <=( (not A170)  and  a112712a );
 a112716a <=( A200  and  (not A199) );
 a112719a <=( A203  and  (not A202) );
 a112720a <=( a112719a  and  a112716a );
 a112721a <=( a112720a  and  a112713a );
 a112724a <=( (not A266)  and  A265 );
 a112727a <=( (not A269)  and  (not A267) );
 a112728a <=( a112727a  and  a112724a );
 a112731a <=( A299  and  A298 );
 a112734a <=( (not A302)  and  A301 );
 a112735a <=( a112734a  and  a112731a );
 a112736a <=( a112735a  and  a112728a );
 a112740a <=( (not A167)  and  (not A169) );
 a112741a <=( (not A170)  and  a112740a );
 a112744a <=( A200  and  (not A199) );
 a112747a <=( A203  and  (not A202) );
 a112748a <=( a112747a  and  a112744a );
 a112749a <=( a112748a  and  a112741a );
 a112752a <=( (not A266)  and  A265 );
 a112755a <=( (not A269)  and  (not A267) );
 a112756a <=( a112755a  and  a112752a );
 a112759a <=( (not A299)  and  A298 );
 a112762a <=( A302  and  (not A301) );
 a112763a <=( a112762a  and  a112759a );
 a112764a <=( a112763a  and  a112756a );
 a112768a <=( (not A167)  and  (not A169) );
 a112769a <=( (not A170)  and  a112768a );
 a112772a <=( A200  and  (not A199) );
 a112775a <=( A203  and  (not A202) );
 a112776a <=( a112775a  and  a112772a );
 a112777a <=( a112776a  and  a112769a );
 a112780a <=( (not A266)  and  A265 );
 a112783a <=( (not A269)  and  (not A267) );
 a112784a <=( a112783a  and  a112780a );
 a112787a <=( A299  and  (not A298) );
 a112790a <=( A302  and  (not A301) );
 a112791a <=( a112790a  and  a112787a );
 a112792a <=( a112791a  and  a112784a );
 a112796a <=( (not A167)  and  (not A169) );
 a112797a <=( (not A170)  and  a112796a );
 a112800a <=( A200  and  (not A199) );
 a112803a <=( A203  and  (not A202) );
 a112804a <=( a112803a  and  a112800a );
 a112805a <=( a112804a  and  a112797a );
 a112808a <=( (not A266)  and  A265 );
 a112811a <=( (not A269)  and  (not A267) );
 a112812a <=( a112811a  and  a112808a );
 a112815a <=( (not A299)  and  (not A298) );
 a112818a <=( (not A302)  and  A301 );
 a112819a <=( a112818a  and  a112815a );
 a112820a <=( a112819a  and  a112812a );
 a112824a <=( (not A167)  and  (not A169) );
 a112825a <=( (not A170)  and  a112824a );
 a112828a <=( A200  and  (not A199) );
 a112831a <=( A202  and  (not A201) );
 a112832a <=( a112831a  and  a112828a );
 a112833a <=( a112832a  and  a112825a );
 a112836a <=( A266  and  A265 );
 a112839a <=( (not A269)  and  A268 );
 a112840a <=( a112839a  and  a112836a );
 a112843a <=( A299  and  A298 );
 a112846a <=( (not A301)  and  (not A300) );
 a112847a <=( a112846a  and  a112843a );
 a112848a <=( a112847a  and  a112840a );
 a112852a <=( (not A167)  and  (not A169) );
 a112853a <=( (not A170)  and  a112852a );
 a112856a <=( A200  and  (not A199) );
 a112859a <=( A202  and  (not A201) );
 a112860a <=( a112859a  and  a112856a );
 a112861a <=( a112860a  and  a112853a );
 a112864a <=( A266  and  A265 );
 a112867a <=( (not A269)  and  A268 );
 a112868a <=( a112867a  and  a112864a );
 a112871a <=( A299  and  A298 );
 a112874a <=( A302  and  (not A300) );
 a112875a <=( a112874a  and  a112871a );
 a112876a <=( a112875a  and  a112868a );
 a112880a <=( (not A167)  and  (not A169) );
 a112881a <=( (not A170)  and  a112880a );
 a112884a <=( A200  and  (not A199) );
 a112887a <=( A202  and  (not A201) );
 a112888a <=( a112887a  and  a112884a );
 a112889a <=( a112888a  and  a112881a );
 a112892a <=( A266  and  A265 );
 a112895a <=( (not A269)  and  A268 );
 a112896a <=( a112895a  and  a112892a );
 a112899a <=( (not A299)  and  A298 );
 a112902a <=( A301  and  (not A300) );
 a112903a <=( a112902a  and  a112899a );
 a112904a <=( a112903a  and  a112896a );
 a112908a <=( (not A167)  and  (not A169) );
 a112909a <=( (not A170)  and  a112908a );
 a112912a <=( A200  and  (not A199) );
 a112915a <=( A202  and  (not A201) );
 a112916a <=( a112915a  and  a112912a );
 a112917a <=( a112916a  and  a112909a );
 a112920a <=( A266  and  A265 );
 a112923a <=( (not A269)  and  A268 );
 a112924a <=( a112923a  and  a112920a );
 a112927a <=( (not A299)  and  A298 );
 a112930a <=( (not A302)  and  (not A300) );
 a112931a <=( a112930a  and  a112927a );
 a112932a <=( a112931a  and  a112924a );
 a112936a <=( (not A167)  and  (not A169) );
 a112937a <=( (not A170)  and  a112936a );
 a112940a <=( A200  and  (not A199) );
 a112943a <=( A202  and  (not A201) );
 a112944a <=( a112943a  and  a112940a );
 a112945a <=( a112944a  and  a112937a );
 a112948a <=( A266  and  A265 );
 a112951a <=( (not A269)  and  A268 );
 a112952a <=( a112951a  and  a112948a );
 a112955a <=( A299  and  (not A298) );
 a112958a <=( A301  and  (not A300) );
 a112959a <=( a112958a  and  a112955a );
 a112960a <=( a112959a  and  a112952a );
 a112964a <=( (not A167)  and  (not A169) );
 a112965a <=( (not A170)  and  a112964a );
 a112968a <=( A200  and  (not A199) );
 a112971a <=( A202  and  (not A201) );
 a112972a <=( a112971a  and  a112968a );
 a112973a <=( a112972a  and  a112965a );
 a112976a <=( A266  and  A265 );
 a112979a <=( (not A269)  and  A268 );
 a112980a <=( a112979a  and  a112976a );
 a112983a <=( A299  and  (not A298) );
 a112986a <=( (not A302)  and  (not A300) );
 a112987a <=( a112986a  and  a112983a );
 a112988a <=( a112987a  and  a112980a );
 a112992a <=( (not A167)  and  (not A169) );
 a112993a <=( (not A170)  and  a112992a );
 a112996a <=( A200  and  (not A199) );
 a112999a <=( A202  and  (not A201) );
 a113000a <=( a112999a  and  a112996a );
 a113001a <=( a113000a  and  a112993a );
 a113004a <=( A266  and  (not A265) );
 a113007a <=( A269  and  (not A268) );
 a113008a <=( a113007a  and  a113004a );
 a113011a <=( A299  and  A298 );
 a113014a <=( (not A301)  and  (not A300) );
 a113015a <=( a113014a  and  a113011a );
 a113016a <=( a113015a  and  a113008a );
 a113020a <=( (not A167)  and  (not A169) );
 a113021a <=( (not A170)  and  a113020a );
 a113024a <=( A200  and  (not A199) );
 a113027a <=( A202  and  (not A201) );
 a113028a <=( a113027a  and  a113024a );
 a113029a <=( a113028a  and  a113021a );
 a113032a <=( A266  and  (not A265) );
 a113035a <=( A269  and  (not A268) );
 a113036a <=( a113035a  and  a113032a );
 a113039a <=( A299  and  A298 );
 a113042a <=( A302  and  (not A300) );
 a113043a <=( a113042a  and  a113039a );
 a113044a <=( a113043a  and  a113036a );
 a113048a <=( (not A167)  and  (not A169) );
 a113049a <=( (not A170)  and  a113048a );
 a113052a <=( A200  and  (not A199) );
 a113055a <=( A202  and  (not A201) );
 a113056a <=( a113055a  and  a113052a );
 a113057a <=( a113056a  and  a113049a );
 a113060a <=( A266  and  (not A265) );
 a113063a <=( A269  and  (not A268) );
 a113064a <=( a113063a  and  a113060a );
 a113067a <=( (not A299)  and  A298 );
 a113070a <=( A301  and  (not A300) );
 a113071a <=( a113070a  and  a113067a );
 a113072a <=( a113071a  and  a113064a );
 a113076a <=( (not A167)  and  (not A169) );
 a113077a <=( (not A170)  and  a113076a );
 a113080a <=( A200  and  (not A199) );
 a113083a <=( A202  and  (not A201) );
 a113084a <=( a113083a  and  a113080a );
 a113085a <=( a113084a  and  a113077a );
 a113088a <=( A266  and  (not A265) );
 a113091a <=( A269  and  (not A268) );
 a113092a <=( a113091a  and  a113088a );
 a113095a <=( (not A299)  and  A298 );
 a113098a <=( (not A302)  and  (not A300) );
 a113099a <=( a113098a  and  a113095a );
 a113100a <=( a113099a  and  a113092a );
 a113104a <=( (not A167)  and  (not A169) );
 a113105a <=( (not A170)  and  a113104a );
 a113108a <=( A200  and  (not A199) );
 a113111a <=( A202  and  (not A201) );
 a113112a <=( a113111a  and  a113108a );
 a113113a <=( a113112a  and  a113105a );
 a113116a <=( A266  and  (not A265) );
 a113119a <=( A269  and  (not A268) );
 a113120a <=( a113119a  and  a113116a );
 a113123a <=( A299  and  (not A298) );
 a113126a <=( A301  and  (not A300) );
 a113127a <=( a113126a  and  a113123a );
 a113128a <=( a113127a  and  a113120a );
 a113132a <=( (not A167)  and  (not A169) );
 a113133a <=( (not A170)  and  a113132a );
 a113136a <=( A200  and  (not A199) );
 a113139a <=( A202  and  (not A201) );
 a113140a <=( a113139a  and  a113136a );
 a113141a <=( a113140a  and  a113133a );
 a113144a <=( A266  and  (not A265) );
 a113147a <=( A269  and  (not A268) );
 a113148a <=( a113147a  and  a113144a );
 a113151a <=( A299  and  (not A298) );
 a113154a <=( (not A302)  and  (not A300) );
 a113155a <=( a113154a  and  a113151a );
 a113156a <=( a113155a  and  a113148a );
 a113160a <=( (not A167)  and  (not A169) );
 a113161a <=( (not A170)  and  a113160a );
 a113164a <=( A200  and  (not A199) );
 a113167a <=( A202  and  (not A201) );
 a113168a <=( a113167a  and  a113164a );
 a113169a <=( a113168a  and  a113161a );
 a113172a <=( (not A266)  and  A265 );
 a113175a <=( A269  and  (not A268) );
 a113176a <=( a113175a  and  a113172a );
 a113179a <=( A299  and  A298 );
 a113182a <=( (not A301)  and  (not A300) );
 a113183a <=( a113182a  and  a113179a );
 a113184a <=( a113183a  and  a113176a );
 a113188a <=( (not A167)  and  (not A169) );
 a113189a <=( (not A170)  and  a113188a );
 a113192a <=( A200  and  (not A199) );
 a113195a <=( A202  and  (not A201) );
 a113196a <=( a113195a  and  a113192a );
 a113197a <=( a113196a  and  a113189a );
 a113200a <=( (not A266)  and  A265 );
 a113203a <=( A269  and  (not A268) );
 a113204a <=( a113203a  and  a113200a );
 a113207a <=( A299  and  A298 );
 a113210a <=( A302  and  (not A300) );
 a113211a <=( a113210a  and  a113207a );
 a113212a <=( a113211a  and  a113204a );
 a113216a <=( (not A167)  and  (not A169) );
 a113217a <=( (not A170)  and  a113216a );
 a113220a <=( A200  and  (not A199) );
 a113223a <=( A202  and  (not A201) );
 a113224a <=( a113223a  and  a113220a );
 a113225a <=( a113224a  and  a113217a );
 a113228a <=( (not A266)  and  A265 );
 a113231a <=( A269  and  (not A268) );
 a113232a <=( a113231a  and  a113228a );
 a113235a <=( (not A299)  and  A298 );
 a113238a <=( A301  and  (not A300) );
 a113239a <=( a113238a  and  a113235a );
 a113240a <=( a113239a  and  a113232a );
 a113244a <=( (not A167)  and  (not A169) );
 a113245a <=( (not A170)  and  a113244a );
 a113248a <=( A200  and  (not A199) );
 a113251a <=( A202  and  (not A201) );
 a113252a <=( a113251a  and  a113248a );
 a113253a <=( a113252a  and  a113245a );
 a113256a <=( (not A266)  and  A265 );
 a113259a <=( A269  and  (not A268) );
 a113260a <=( a113259a  and  a113256a );
 a113263a <=( (not A299)  and  A298 );
 a113266a <=( (not A302)  and  (not A300) );
 a113267a <=( a113266a  and  a113263a );
 a113268a <=( a113267a  and  a113260a );
 a113272a <=( (not A167)  and  (not A169) );
 a113273a <=( (not A170)  and  a113272a );
 a113276a <=( A200  and  (not A199) );
 a113279a <=( A202  and  (not A201) );
 a113280a <=( a113279a  and  a113276a );
 a113281a <=( a113280a  and  a113273a );
 a113284a <=( (not A266)  and  A265 );
 a113287a <=( A269  and  (not A268) );
 a113288a <=( a113287a  and  a113284a );
 a113291a <=( A299  and  (not A298) );
 a113294a <=( A301  and  (not A300) );
 a113295a <=( a113294a  and  a113291a );
 a113296a <=( a113295a  and  a113288a );
 a113300a <=( (not A167)  and  (not A169) );
 a113301a <=( (not A170)  and  a113300a );
 a113304a <=( A200  and  (not A199) );
 a113307a <=( A202  and  (not A201) );
 a113308a <=( a113307a  and  a113304a );
 a113309a <=( a113308a  and  a113301a );
 a113312a <=( (not A266)  and  A265 );
 a113315a <=( A269  and  (not A268) );
 a113316a <=( a113315a  and  a113312a );
 a113319a <=( A299  and  (not A298) );
 a113322a <=( (not A302)  and  (not A300) );
 a113323a <=( a113322a  and  a113319a );
 a113324a <=( a113323a  and  a113316a );
 a113328a <=( (not A167)  and  (not A169) );
 a113329a <=( (not A170)  and  a113328a );
 a113332a <=( A200  and  (not A199) );
 a113335a <=( A202  and  (not A201) );
 a113336a <=( a113335a  and  a113332a );
 a113337a <=( a113336a  and  a113329a );
 a113340a <=( (not A266)  and  (not A265) );
 a113343a <=( (not A269)  and  A268 );
 a113344a <=( a113343a  and  a113340a );
 a113347a <=( A299  and  A298 );
 a113350a <=( (not A301)  and  (not A300) );
 a113351a <=( a113350a  and  a113347a );
 a113352a <=( a113351a  and  a113344a );
 a113356a <=( (not A167)  and  (not A169) );
 a113357a <=( (not A170)  and  a113356a );
 a113360a <=( A200  and  (not A199) );
 a113363a <=( A202  and  (not A201) );
 a113364a <=( a113363a  and  a113360a );
 a113365a <=( a113364a  and  a113357a );
 a113368a <=( (not A266)  and  (not A265) );
 a113371a <=( (not A269)  and  A268 );
 a113372a <=( a113371a  and  a113368a );
 a113375a <=( A299  and  A298 );
 a113378a <=( A302  and  (not A300) );
 a113379a <=( a113378a  and  a113375a );
 a113380a <=( a113379a  and  a113372a );
 a113384a <=( (not A167)  and  (not A169) );
 a113385a <=( (not A170)  and  a113384a );
 a113388a <=( A200  and  (not A199) );
 a113391a <=( A202  and  (not A201) );
 a113392a <=( a113391a  and  a113388a );
 a113393a <=( a113392a  and  a113385a );
 a113396a <=( (not A266)  and  (not A265) );
 a113399a <=( (not A269)  and  A268 );
 a113400a <=( a113399a  and  a113396a );
 a113403a <=( (not A299)  and  A298 );
 a113406a <=( A301  and  (not A300) );
 a113407a <=( a113406a  and  a113403a );
 a113408a <=( a113407a  and  a113400a );
 a113412a <=( (not A167)  and  (not A169) );
 a113413a <=( (not A170)  and  a113412a );
 a113416a <=( A200  and  (not A199) );
 a113419a <=( A202  and  (not A201) );
 a113420a <=( a113419a  and  a113416a );
 a113421a <=( a113420a  and  a113413a );
 a113424a <=( (not A266)  and  (not A265) );
 a113427a <=( (not A269)  and  A268 );
 a113428a <=( a113427a  and  a113424a );
 a113431a <=( (not A299)  and  A298 );
 a113434a <=( (not A302)  and  (not A300) );
 a113435a <=( a113434a  and  a113431a );
 a113436a <=( a113435a  and  a113428a );
 a113440a <=( (not A167)  and  (not A169) );
 a113441a <=( (not A170)  and  a113440a );
 a113444a <=( A200  and  (not A199) );
 a113447a <=( A202  and  (not A201) );
 a113448a <=( a113447a  and  a113444a );
 a113449a <=( a113448a  and  a113441a );
 a113452a <=( (not A266)  and  (not A265) );
 a113455a <=( (not A269)  and  A268 );
 a113456a <=( a113455a  and  a113452a );
 a113459a <=( A299  and  (not A298) );
 a113462a <=( A301  and  (not A300) );
 a113463a <=( a113462a  and  a113459a );
 a113464a <=( a113463a  and  a113456a );
 a113468a <=( (not A167)  and  (not A169) );
 a113469a <=( (not A170)  and  a113468a );
 a113472a <=( A200  and  (not A199) );
 a113475a <=( A202  and  (not A201) );
 a113476a <=( a113475a  and  a113472a );
 a113477a <=( a113476a  and  a113469a );
 a113480a <=( (not A266)  and  (not A265) );
 a113483a <=( (not A269)  and  A268 );
 a113484a <=( a113483a  and  a113480a );
 a113487a <=( A299  and  (not A298) );
 a113490a <=( (not A302)  and  (not A300) );
 a113491a <=( a113490a  and  a113487a );
 a113492a <=( a113491a  and  a113484a );
 a113496a <=( (not A167)  and  (not A169) );
 a113497a <=( (not A170)  and  a113496a );
 a113500a <=( A200  and  (not A199) );
 a113503a <=( (not A203)  and  (not A201) );
 a113504a <=( a113503a  and  a113500a );
 a113505a <=( a113504a  and  a113497a );
 a113508a <=( A266  and  A265 );
 a113511a <=( (not A269)  and  A268 );
 a113512a <=( a113511a  and  a113508a );
 a113515a <=( A299  and  A298 );
 a113518a <=( (not A301)  and  (not A300) );
 a113519a <=( a113518a  and  a113515a );
 a113520a <=( a113519a  and  a113512a );
 a113524a <=( (not A167)  and  (not A169) );
 a113525a <=( (not A170)  and  a113524a );
 a113528a <=( A200  and  (not A199) );
 a113531a <=( (not A203)  and  (not A201) );
 a113532a <=( a113531a  and  a113528a );
 a113533a <=( a113532a  and  a113525a );
 a113536a <=( A266  and  A265 );
 a113539a <=( (not A269)  and  A268 );
 a113540a <=( a113539a  and  a113536a );
 a113543a <=( A299  and  A298 );
 a113546a <=( A302  and  (not A300) );
 a113547a <=( a113546a  and  a113543a );
 a113548a <=( a113547a  and  a113540a );
 a113552a <=( (not A167)  and  (not A169) );
 a113553a <=( (not A170)  and  a113552a );
 a113556a <=( A200  and  (not A199) );
 a113559a <=( (not A203)  and  (not A201) );
 a113560a <=( a113559a  and  a113556a );
 a113561a <=( a113560a  and  a113553a );
 a113564a <=( A266  and  A265 );
 a113567a <=( (not A269)  and  A268 );
 a113568a <=( a113567a  and  a113564a );
 a113571a <=( (not A299)  and  A298 );
 a113574a <=( A301  and  (not A300) );
 a113575a <=( a113574a  and  a113571a );
 a113576a <=( a113575a  and  a113568a );
 a113580a <=( (not A167)  and  (not A169) );
 a113581a <=( (not A170)  and  a113580a );
 a113584a <=( A200  and  (not A199) );
 a113587a <=( (not A203)  and  (not A201) );
 a113588a <=( a113587a  and  a113584a );
 a113589a <=( a113588a  and  a113581a );
 a113592a <=( A266  and  A265 );
 a113595a <=( (not A269)  and  A268 );
 a113596a <=( a113595a  and  a113592a );
 a113599a <=( (not A299)  and  A298 );
 a113602a <=( (not A302)  and  (not A300) );
 a113603a <=( a113602a  and  a113599a );
 a113604a <=( a113603a  and  a113596a );
 a113608a <=( (not A167)  and  (not A169) );
 a113609a <=( (not A170)  and  a113608a );
 a113612a <=( A200  and  (not A199) );
 a113615a <=( (not A203)  and  (not A201) );
 a113616a <=( a113615a  and  a113612a );
 a113617a <=( a113616a  and  a113609a );
 a113620a <=( A266  and  A265 );
 a113623a <=( (not A269)  and  A268 );
 a113624a <=( a113623a  and  a113620a );
 a113627a <=( A299  and  (not A298) );
 a113630a <=( A301  and  (not A300) );
 a113631a <=( a113630a  and  a113627a );
 a113632a <=( a113631a  and  a113624a );
 a113636a <=( (not A167)  and  (not A169) );
 a113637a <=( (not A170)  and  a113636a );
 a113640a <=( A200  and  (not A199) );
 a113643a <=( (not A203)  and  (not A201) );
 a113644a <=( a113643a  and  a113640a );
 a113645a <=( a113644a  and  a113637a );
 a113648a <=( A266  and  A265 );
 a113651a <=( (not A269)  and  A268 );
 a113652a <=( a113651a  and  a113648a );
 a113655a <=( A299  and  (not A298) );
 a113658a <=( (not A302)  and  (not A300) );
 a113659a <=( a113658a  and  a113655a );
 a113660a <=( a113659a  and  a113652a );
 a113664a <=( (not A167)  and  (not A169) );
 a113665a <=( (not A170)  and  a113664a );
 a113668a <=( A200  and  (not A199) );
 a113671a <=( (not A203)  and  (not A201) );
 a113672a <=( a113671a  and  a113668a );
 a113673a <=( a113672a  and  a113665a );
 a113676a <=( A266  and  (not A265) );
 a113679a <=( A269  and  (not A268) );
 a113680a <=( a113679a  and  a113676a );
 a113683a <=( A299  and  A298 );
 a113686a <=( (not A301)  and  (not A300) );
 a113687a <=( a113686a  and  a113683a );
 a113688a <=( a113687a  and  a113680a );
 a113692a <=( (not A167)  and  (not A169) );
 a113693a <=( (not A170)  and  a113692a );
 a113696a <=( A200  and  (not A199) );
 a113699a <=( (not A203)  and  (not A201) );
 a113700a <=( a113699a  and  a113696a );
 a113701a <=( a113700a  and  a113693a );
 a113704a <=( A266  and  (not A265) );
 a113707a <=( A269  and  (not A268) );
 a113708a <=( a113707a  and  a113704a );
 a113711a <=( A299  and  A298 );
 a113714a <=( A302  and  (not A300) );
 a113715a <=( a113714a  and  a113711a );
 a113716a <=( a113715a  and  a113708a );
 a113720a <=( (not A167)  and  (not A169) );
 a113721a <=( (not A170)  and  a113720a );
 a113724a <=( A200  and  (not A199) );
 a113727a <=( (not A203)  and  (not A201) );
 a113728a <=( a113727a  and  a113724a );
 a113729a <=( a113728a  and  a113721a );
 a113732a <=( A266  and  (not A265) );
 a113735a <=( A269  and  (not A268) );
 a113736a <=( a113735a  and  a113732a );
 a113739a <=( (not A299)  and  A298 );
 a113742a <=( A301  and  (not A300) );
 a113743a <=( a113742a  and  a113739a );
 a113744a <=( a113743a  and  a113736a );
 a113748a <=( (not A167)  and  (not A169) );
 a113749a <=( (not A170)  and  a113748a );
 a113752a <=( A200  and  (not A199) );
 a113755a <=( (not A203)  and  (not A201) );
 a113756a <=( a113755a  and  a113752a );
 a113757a <=( a113756a  and  a113749a );
 a113760a <=( A266  and  (not A265) );
 a113763a <=( A269  and  (not A268) );
 a113764a <=( a113763a  and  a113760a );
 a113767a <=( (not A299)  and  A298 );
 a113770a <=( (not A302)  and  (not A300) );
 a113771a <=( a113770a  and  a113767a );
 a113772a <=( a113771a  and  a113764a );
 a113776a <=( (not A167)  and  (not A169) );
 a113777a <=( (not A170)  and  a113776a );
 a113780a <=( A200  and  (not A199) );
 a113783a <=( (not A203)  and  (not A201) );
 a113784a <=( a113783a  and  a113780a );
 a113785a <=( a113784a  and  a113777a );
 a113788a <=( A266  and  (not A265) );
 a113791a <=( A269  and  (not A268) );
 a113792a <=( a113791a  and  a113788a );
 a113795a <=( A299  and  (not A298) );
 a113798a <=( A301  and  (not A300) );
 a113799a <=( a113798a  and  a113795a );
 a113800a <=( a113799a  and  a113792a );
 a113804a <=( (not A167)  and  (not A169) );
 a113805a <=( (not A170)  and  a113804a );
 a113808a <=( A200  and  (not A199) );
 a113811a <=( (not A203)  and  (not A201) );
 a113812a <=( a113811a  and  a113808a );
 a113813a <=( a113812a  and  a113805a );
 a113816a <=( A266  and  (not A265) );
 a113819a <=( A269  and  (not A268) );
 a113820a <=( a113819a  and  a113816a );
 a113823a <=( A299  and  (not A298) );
 a113826a <=( (not A302)  and  (not A300) );
 a113827a <=( a113826a  and  a113823a );
 a113828a <=( a113827a  and  a113820a );
 a113832a <=( (not A167)  and  (not A169) );
 a113833a <=( (not A170)  and  a113832a );
 a113836a <=( A200  and  (not A199) );
 a113839a <=( (not A203)  and  (not A201) );
 a113840a <=( a113839a  and  a113836a );
 a113841a <=( a113840a  and  a113833a );
 a113844a <=( (not A266)  and  A265 );
 a113847a <=( A269  and  (not A268) );
 a113848a <=( a113847a  and  a113844a );
 a113851a <=( A299  and  A298 );
 a113854a <=( (not A301)  and  (not A300) );
 a113855a <=( a113854a  and  a113851a );
 a113856a <=( a113855a  and  a113848a );
 a113860a <=( (not A167)  and  (not A169) );
 a113861a <=( (not A170)  and  a113860a );
 a113864a <=( A200  and  (not A199) );
 a113867a <=( (not A203)  and  (not A201) );
 a113868a <=( a113867a  and  a113864a );
 a113869a <=( a113868a  and  a113861a );
 a113872a <=( (not A266)  and  A265 );
 a113875a <=( A269  and  (not A268) );
 a113876a <=( a113875a  and  a113872a );
 a113879a <=( A299  and  A298 );
 a113882a <=( A302  and  (not A300) );
 a113883a <=( a113882a  and  a113879a );
 a113884a <=( a113883a  and  a113876a );
 a113888a <=( (not A167)  and  (not A169) );
 a113889a <=( (not A170)  and  a113888a );
 a113892a <=( A200  and  (not A199) );
 a113895a <=( (not A203)  and  (not A201) );
 a113896a <=( a113895a  and  a113892a );
 a113897a <=( a113896a  and  a113889a );
 a113900a <=( (not A266)  and  A265 );
 a113903a <=( A269  and  (not A268) );
 a113904a <=( a113903a  and  a113900a );
 a113907a <=( (not A299)  and  A298 );
 a113910a <=( A301  and  (not A300) );
 a113911a <=( a113910a  and  a113907a );
 a113912a <=( a113911a  and  a113904a );
 a113916a <=( (not A167)  and  (not A169) );
 a113917a <=( (not A170)  and  a113916a );
 a113920a <=( A200  and  (not A199) );
 a113923a <=( (not A203)  and  (not A201) );
 a113924a <=( a113923a  and  a113920a );
 a113925a <=( a113924a  and  a113917a );
 a113928a <=( (not A266)  and  A265 );
 a113931a <=( A269  and  (not A268) );
 a113932a <=( a113931a  and  a113928a );
 a113935a <=( (not A299)  and  A298 );
 a113938a <=( (not A302)  and  (not A300) );
 a113939a <=( a113938a  and  a113935a );
 a113940a <=( a113939a  and  a113932a );
 a113944a <=( (not A167)  and  (not A169) );
 a113945a <=( (not A170)  and  a113944a );
 a113948a <=( A200  and  (not A199) );
 a113951a <=( (not A203)  and  (not A201) );
 a113952a <=( a113951a  and  a113948a );
 a113953a <=( a113952a  and  a113945a );
 a113956a <=( (not A266)  and  A265 );
 a113959a <=( A269  and  (not A268) );
 a113960a <=( a113959a  and  a113956a );
 a113963a <=( A299  and  (not A298) );
 a113966a <=( A301  and  (not A300) );
 a113967a <=( a113966a  and  a113963a );
 a113968a <=( a113967a  and  a113960a );
 a113972a <=( (not A167)  and  (not A169) );
 a113973a <=( (not A170)  and  a113972a );
 a113976a <=( A200  and  (not A199) );
 a113979a <=( (not A203)  and  (not A201) );
 a113980a <=( a113979a  and  a113976a );
 a113981a <=( a113980a  and  a113973a );
 a113984a <=( (not A266)  and  A265 );
 a113987a <=( A269  and  (not A268) );
 a113988a <=( a113987a  and  a113984a );
 a113991a <=( A299  and  (not A298) );
 a113994a <=( (not A302)  and  (not A300) );
 a113995a <=( a113994a  and  a113991a );
 a113996a <=( a113995a  and  a113988a );
 a114000a <=( (not A167)  and  (not A169) );
 a114001a <=( (not A170)  and  a114000a );
 a114004a <=( A200  and  (not A199) );
 a114007a <=( (not A203)  and  (not A201) );
 a114008a <=( a114007a  and  a114004a );
 a114009a <=( a114008a  and  a114001a );
 a114012a <=( (not A266)  and  (not A265) );
 a114015a <=( (not A269)  and  A268 );
 a114016a <=( a114015a  and  a114012a );
 a114019a <=( A299  and  A298 );
 a114022a <=( (not A301)  and  (not A300) );
 a114023a <=( a114022a  and  a114019a );
 a114024a <=( a114023a  and  a114016a );
 a114028a <=( (not A167)  and  (not A169) );
 a114029a <=( (not A170)  and  a114028a );
 a114032a <=( A200  and  (not A199) );
 a114035a <=( (not A203)  and  (not A201) );
 a114036a <=( a114035a  and  a114032a );
 a114037a <=( a114036a  and  a114029a );
 a114040a <=( (not A266)  and  (not A265) );
 a114043a <=( (not A269)  and  A268 );
 a114044a <=( a114043a  and  a114040a );
 a114047a <=( A299  and  A298 );
 a114050a <=( A302  and  (not A300) );
 a114051a <=( a114050a  and  a114047a );
 a114052a <=( a114051a  and  a114044a );
 a114056a <=( (not A167)  and  (not A169) );
 a114057a <=( (not A170)  and  a114056a );
 a114060a <=( A200  and  (not A199) );
 a114063a <=( (not A203)  and  (not A201) );
 a114064a <=( a114063a  and  a114060a );
 a114065a <=( a114064a  and  a114057a );
 a114068a <=( (not A266)  and  (not A265) );
 a114071a <=( (not A269)  and  A268 );
 a114072a <=( a114071a  and  a114068a );
 a114075a <=( (not A299)  and  A298 );
 a114078a <=( A301  and  (not A300) );
 a114079a <=( a114078a  and  a114075a );
 a114080a <=( a114079a  and  a114072a );
 a114084a <=( (not A167)  and  (not A169) );
 a114085a <=( (not A170)  and  a114084a );
 a114088a <=( A200  and  (not A199) );
 a114091a <=( (not A203)  and  (not A201) );
 a114092a <=( a114091a  and  a114088a );
 a114093a <=( a114092a  and  a114085a );
 a114096a <=( (not A266)  and  (not A265) );
 a114099a <=( (not A269)  and  A268 );
 a114100a <=( a114099a  and  a114096a );
 a114103a <=( (not A299)  and  A298 );
 a114106a <=( (not A302)  and  (not A300) );
 a114107a <=( a114106a  and  a114103a );
 a114108a <=( a114107a  and  a114100a );
 a114112a <=( (not A167)  and  (not A169) );
 a114113a <=( (not A170)  and  a114112a );
 a114116a <=( A200  and  (not A199) );
 a114119a <=( (not A203)  and  (not A201) );
 a114120a <=( a114119a  and  a114116a );
 a114121a <=( a114120a  and  a114113a );
 a114124a <=( (not A266)  and  (not A265) );
 a114127a <=( (not A269)  and  A268 );
 a114128a <=( a114127a  and  a114124a );
 a114131a <=( A299  and  (not A298) );
 a114134a <=( A301  and  (not A300) );
 a114135a <=( a114134a  and  a114131a );
 a114136a <=( a114135a  and  a114128a );
 a114140a <=( (not A167)  and  (not A169) );
 a114141a <=( (not A170)  and  a114140a );
 a114144a <=( A200  and  (not A199) );
 a114147a <=( (not A203)  and  (not A201) );
 a114148a <=( a114147a  and  a114144a );
 a114149a <=( a114148a  and  a114141a );
 a114152a <=( (not A266)  and  (not A265) );
 a114155a <=( (not A269)  and  A268 );
 a114156a <=( a114155a  and  a114152a );
 a114159a <=( A299  and  (not A298) );
 a114162a <=( (not A302)  and  (not A300) );
 a114163a <=( a114162a  and  a114159a );
 a114164a <=( a114163a  and  a114156a );
 a114168a <=( (not A167)  and  (not A169) );
 a114169a <=( (not A170)  and  a114168a );
 a114172a <=( (not A200)  and  A199 );
 a114175a <=( A203  and  (not A202) );
 a114176a <=( a114175a  and  a114172a );
 a114177a <=( a114176a  and  a114169a );
 a114180a <=( A266  and  A265 );
 a114183a <=( (not A268)  and  (not A267) );
 a114184a <=( a114183a  and  a114180a );
 a114187a <=( A299  and  A298 );
 a114190a <=( (not A302)  and  A301 );
 a114191a <=( a114190a  and  a114187a );
 a114192a <=( a114191a  and  a114184a );
 a114196a <=( (not A167)  and  (not A169) );
 a114197a <=( (not A170)  and  a114196a );
 a114200a <=( (not A200)  and  A199 );
 a114203a <=( A203  and  (not A202) );
 a114204a <=( a114203a  and  a114200a );
 a114205a <=( a114204a  and  a114197a );
 a114208a <=( A266  and  A265 );
 a114211a <=( (not A268)  and  (not A267) );
 a114212a <=( a114211a  and  a114208a );
 a114215a <=( (not A299)  and  A298 );
 a114218a <=( A302  and  (not A301) );
 a114219a <=( a114218a  and  a114215a );
 a114220a <=( a114219a  and  a114212a );
 a114224a <=( (not A167)  and  (not A169) );
 a114225a <=( (not A170)  and  a114224a );
 a114228a <=( (not A200)  and  A199 );
 a114231a <=( A203  and  (not A202) );
 a114232a <=( a114231a  and  a114228a );
 a114233a <=( a114232a  and  a114225a );
 a114236a <=( A266  and  A265 );
 a114239a <=( (not A268)  and  (not A267) );
 a114240a <=( a114239a  and  a114236a );
 a114243a <=( A299  and  (not A298) );
 a114246a <=( A302  and  (not A301) );
 a114247a <=( a114246a  and  a114243a );
 a114248a <=( a114247a  and  a114240a );
 a114252a <=( (not A167)  and  (not A169) );
 a114253a <=( (not A170)  and  a114252a );
 a114256a <=( (not A200)  and  A199 );
 a114259a <=( A203  and  (not A202) );
 a114260a <=( a114259a  and  a114256a );
 a114261a <=( a114260a  and  a114253a );
 a114264a <=( A266  and  A265 );
 a114267a <=( (not A268)  and  (not A267) );
 a114268a <=( a114267a  and  a114264a );
 a114271a <=( (not A299)  and  (not A298) );
 a114274a <=( (not A302)  and  A301 );
 a114275a <=( a114274a  and  a114271a );
 a114276a <=( a114275a  and  a114268a );
 a114280a <=( (not A167)  and  (not A169) );
 a114281a <=( (not A170)  and  a114280a );
 a114284a <=( (not A200)  and  A199 );
 a114287a <=( A203  and  (not A202) );
 a114288a <=( a114287a  and  a114284a );
 a114289a <=( a114288a  and  a114281a );
 a114292a <=( A266  and  A265 );
 a114295a <=( A269  and  (not A267) );
 a114296a <=( a114295a  and  a114292a );
 a114299a <=( A299  and  A298 );
 a114302a <=( (not A302)  and  A301 );
 a114303a <=( a114302a  and  a114299a );
 a114304a <=( a114303a  and  a114296a );
 a114308a <=( (not A167)  and  (not A169) );
 a114309a <=( (not A170)  and  a114308a );
 a114312a <=( (not A200)  and  A199 );
 a114315a <=( A203  and  (not A202) );
 a114316a <=( a114315a  and  a114312a );
 a114317a <=( a114316a  and  a114309a );
 a114320a <=( A266  and  A265 );
 a114323a <=( A269  and  (not A267) );
 a114324a <=( a114323a  and  a114320a );
 a114327a <=( (not A299)  and  A298 );
 a114330a <=( A302  and  (not A301) );
 a114331a <=( a114330a  and  a114327a );
 a114332a <=( a114331a  and  a114324a );
 a114336a <=( (not A167)  and  (not A169) );
 a114337a <=( (not A170)  and  a114336a );
 a114340a <=( (not A200)  and  A199 );
 a114343a <=( A203  and  (not A202) );
 a114344a <=( a114343a  and  a114340a );
 a114345a <=( a114344a  and  a114337a );
 a114348a <=( A266  and  A265 );
 a114351a <=( A269  and  (not A267) );
 a114352a <=( a114351a  and  a114348a );
 a114355a <=( A299  and  (not A298) );
 a114358a <=( A302  and  (not A301) );
 a114359a <=( a114358a  and  a114355a );
 a114360a <=( a114359a  and  a114352a );
 a114364a <=( (not A167)  and  (not A169) );
 a114365a <=( (not A170)  and  a114364a );
 a114368a <=( (not A200)  and  A199 );
 a114371a <=( A203  and  (not A202) );
 a114372a <=( a114371a  and  a114368a );
 a114373a <=( a114372a  and  a114365a );
 a114376a <=( A266  and  A265 );
 a114379a <=( A269  and  (not A267) );
 a114380a <=( a114379a  and  a114376a );
 a114383a <=( (not A299)  and  (not A298) );
 a114386a <=( (not A302)  and  A301 );
 a114387a <=( a114386a  and  a114383a );
 a114388a <=( a114387a  and  a114380a );
 a114392a <=( (not A167)  and  (not A169) );
 a114393a <=( (not A170)  and  a114392a );
 a114396a <=( (not A200)  and  A199 );
 a114399a <=( A203  and  (not A202) );
 a114400a <=( a114399a  and  a114396a );
 a114401a <=( a114400a  and  a114393a );
 a114404a <=( A266  and  (not A265) );
 a114407a <=( A268  and  (not A267) );
 a114408a <=( a114407a  and  a114404a );
 a114411a <=( A299  and  A298 );
 a114414a <=( (not A302)  and  A301 );
 a114415a <=( a114414a  and  a114411a );
 a114416a <=( a114415a  and  a114408a );
 a114420a <=( (not A167)  and  (not A169) );
 a114421a <=( (not A170)  and  a114420a );
 a114424a <=( (not A200)  and  A199 );
 a114427a <=( A203  and  (not A202) );
 a114428a <=( a114427a  and  a114424a );
 a114429a <=( a114428a  and  a114421a );
 a114432a <=( A266  and  (not A265) );
 a114435a <=( A268  and  (not A267) );
 a114436a <=( a114435a  and  a114432a );
 a114439a <=( (not A299)  and  A298 );
 a114442a <=( A302  and  (not A301) );
 a114443a <=( a114442a  and  a114439a );
 a114444a <=( a114443a  and  a114436a );
 a114448a <=( (not A167)  and  (not A169) );
 a114449a <=( (not A170)  and  a114448a );
 a114452a <=( (not A200)  and  A199 );
 a114455a <=( A203  and  (not A202) );
 a114456a <=( a114455a  and  a114452a );
 a114457a <=( a114456a  and  a114449a );
 a114460a <=( A266  and  (not A265) );
 a114463a <=( A268  and  (not A267) );
 a114464a <=( a114463a  and  a114460a );
 a114467a <=( A299  and  (not A298) );
 a114470a <=( A302  and  (not A301) );
 a114471a <=( a114470a  and  a114467a );
 a114472a <=( a114471a  and  a114464a );
 a114476a <=( (not A167)  and  (not A169) );
 a114477a <=( (not A170)  and  a114476a );
 a114480a <=( (not A200)  and  A199 );
 a114483a <=( A203  and  (not A202) );
 a114484a <=( a114483a  and  a114480a );
 a114485a <=( a114484a  and  a114477a );
 a114488a <=( A266  and  (not A265) );
 a114491a <=( A268  and  (not A267) );
 a114492a <=( a114491a  and  a114488a );
 a114495a <=( (not A299)  and  (not A298) );
 a114498a <=( (not A302)  and  A301 );
 a114499a <=( a114498a  and  a114495a );
 a114500a <=( a114499a  and  a114492a );
 a114504a <=( (not A167)  and  (not A169) );
 a114505a <=( (not A170)  and  a114504a );
 a114508a <=( (not A200)  and  A199 );
 a114511a <=( A203  and  (not A202) );
 a114512a <=( a114511a  and  a114508a );
 a114513a <=( a114512a  and  a114505a );
 a114516a <=( A266  and  (not A265) );
 a114519a <=( (not A269)  and  (not A267) );
 a114520a <=( a114519a  and  a114516a );
 a114523a <=( A299  and  A298 );
 a114526a <=( (not A302)  and  A301 );
 a114527a <=( a114526a  and  a114523a );
 a114528a <=( a114527a  and  a114520a );
 a114532a <=( (not A167)  and  (not A169) );
 a114533a <=( (not A170)  and  a114532a );
 a114536a <=( (not A200)  and  A199 );
 a114539a <=( A203  and  (not A202) );
 a114540a <=( a114539a  and  a114536a );
 a114541a <=( a114540a  and  a114533a );
 a114544a <=( A266  and  (not A265) );
 a114547a <=( (not A269)  and  (not A267) );
 a114548a <=( a114547a  and  a114544a );
 a114551a <=( (not A299)  and  A298 );
 a114554a <=( A302  and  (not A301) );
 a114555a <=( a114554a  and  a114551a );
 a114556a <=( a114555a  and  a114548a );
 a114560a <=( (not A167)  and  (not A169) );
 a114561a <=( (not A170)  and  a114560a );
 a114564a <=( (not A200)  and  A199 );
 a114567a <=( A203  and  (not A202) );
 a114568a <=( a114567a  and  a114564a );
 a114569a <=( a114568a  and  a114561a );
 a114572a <=( A266  and  (not A265) );
 a114575a <=( (not A269)  and  (not A267) );
 a114576a <=( a114575a  and  a114572a );
 a114579a <=( A299  and  (not A298) );
 a114582a <=( A302  and  (not A301) );
 a114583a <=( a114582a  and  a114579a );
 a114584a <=( a114583a  and  a114576a );
 a114588a <=( (not A167)  and  (not A169) );
 a114589a <=( (not A170)  and  a114588a );
 a114592a <=( (not A200)  and  A199 );
 a114595a <=( A203  and  (not A202) );
 a114596a <=( a114595a  and  a114592a );
 a114597a <=( a114596a  and  a114589a );
 a114600a <=( A266  and  (not A265) );
 a114603a <=( (not A269)  and  (not A267) );
 a114604a <=( a114603a  and  a114600a );
 a114607a <=( (not A299)  and  (not A298) );
 a114610a <=( (not A302)  and  A301 );
 a114611a <=( a114610a  and  a114607a );
 a114612a <=( a114611a  and  a114604a );
 a114616a <=( (not A167)  and  (not A169) );
 a114617a <=( (not A170)  and  a114616a );
 a114620a <=( (not A200)  and  A199 );
 a114623a <=( A203  and  (not A202) );
 a114624a <=( a114623a  and  a114620a );
 a114625a <=( a114624a  and  a114617a );
 a114628a <=( (not A266)  and  A265 );
 a114631a <=( A268  and  (not A267) );
 a114632a <=( a114631a  and  a114628a );
 a114635a <=( A299  and  A298 );
 a114638a <=( (not A302)  and  A301 );
 a114639a <=( a114638a  and  a114635a );
 a114640a <=( a114639a  and  a114632a );
 a114644a <=( (not A167)  and  (not A169) );
 a114645a <=( (not A170)  and  a114644a );
 a114648a <=( (not A200)  and  A199 );
 a114651a <=( A203  and  (not A202) );
 a114652a <=( a114651a  and  a114648a );
 a114653a <=( a114652a  and  a114645a );
 a114656a <=( (not A266)  and  A265 );
 a114659a <=( A268  and  (not A267) );
 a114660a <=( a114659a  and  a114656a );
 a114663a <=( (not A299)  and  A298 );
 a114666a <=( A302  and  (not A301) );
 a114667a <=( a114666a  and  a114663a );
 a114668a <=( a114667a  and  a114660a );
 a114672a <=( (not A167)  and  (not A169) );
 a114673a <=( (not A170)  and  a114672a );
 a114676a <=( (not A200)  and  A199 );
 a114679a <=( A203  and  (not A202) );
 a114680a <=( a114679a  and  a114676a );
 a114681a <=( a114680a  and  a114673a );
 a114684a <=( (not A266)  and  A265 );
 a114687a <=( A268  and  (not A267) );
 a114688a <=( a114687a  and  a114684a );
 a114691a <=( A299  and  (not A298) );
 a114694a <=( A302  and  (not A301) );
 a114695a <=( a114694a  and  a114691a );
 a114696a <=( a114695a  and  a114688a );
 a114700a <=( (not A167)  and  (not A169) );
 a114701a <=( (not A170)  and  a114700a );
 a114704a <=( (not A200)  and  A199 );
 a114707a <=( A203  and  (not A202) );
 a114708a <=( a114707a  and  a114704a );
 a114709a <=( a114708a  and  a114701a );
 a114712a <=( (not A266)  and  A265 );
 a114715a <=( A268  and  (not A267) );
 a114716a <=( a114715a  and  a114712a );
 a114719a <=( (not A299)  and  (not A298) );
 a114722a <=( (not A302)  and  A301 );
 a114723a <=( a114722a  and  a114719a );
 a114724a <=( a114723a  and  a114716a );
 a114728a <=( (not A167)  and  (not A169) );
 a114729a <=( (not A170)  and  a114728a );
 a114732a <=( (not A200)  and  A199 );
 a114735a <=( A203  and  (not A202) );
 a114736a <=( a114735a  and  a114732a );
 a114737a <=( a114736a  and  a114729a );
 a114740a <=( (not A266)  and  A265 );
 a114743a <=( (not A269)  and  (not A267) );
 a114744a <=( a114743a  and  a114740a );
 a114747a <=( A299  and  A298 );
 a114750a <=( (not A302)  and  A301 );
 a114751a <=( a114750a  and  a114747a );
 a114752a <=( a114751a  and  a114744a );
 a114756a <=( (not A167)  and  (not A169) );
 a114757a <=( (not A170)  and  a114756a );
 a114760a <=( (not A200)  and  A199 );
 a114763a <=( A203  and  (not A202) );
 a114764a <=( a114763a  and  a114760a );
 a114765a <=( a114764a  and  a114757a );
 a114768a <=( (not A266)  and  A265 );
 a114771a <=( (not A269)  and  (not A267) );
 a114772a <=( a114771a  and  a114768a );
 a114775a <=( (not A299)  and  A298 );
 a114778a <=( A302  and  (not A301) );
 a114779a <=( a114778a  and  a114775a );
 a114780a <=( a114779a  and  a114772a );
 a114784a <=( (not A167)  and  (not A169) );
 a114785a <=( (not A170)  and  a114784a );
 a114788a <=( (not A200)  and  A199 );
 a114791a <=( A203  and  (not A202) );
 a114792a <=( a114791a  and  a114788a );
 a114793a <=( a114792a  and  a114785a );
 a114796a <=( (not A266)  and  A265 );
 a114799a <=( (not A269)  and  (not A267) );
 a114800a <=( a114799a  and  a114796a );
 a114803a <=( A299  and  (not A298) );
 a114806a <=( A302  and  (not A301) );
 a114807a <=( a114806a  and  a114803a );
 a114808a <=( a114807a  and  a114800a );
 a114812a <=( (not A167)  and  (not A169) );
 a114813a <=( (not A170)  and  a114812a );
 a114816a <=( (not A200)  and  A199 );
 a114819a <=( A203  and  (not A202) );
 a114820a <=( a114819a  and  a114816a );
 a114821a <=( a114820a  and  a114813a );
 a114824a <=( (not A266)  and  A265 );
 a114827a <=( (not A269)  and  (not A267) );
 a114828a <=( a114827a  and  a114824a );
 a114831a <=( (not A299)  and  (not A298) );
 a114834a <=( (not A302)  and  A301 );
 a114835a <=( a114834a  and  a114831a );
 a114836a <=( a114835a  and  a114828a );
 a114840a <=( (not A167)  and  (not A169) );
 a114841a <=( (not A170)  and  a114840a );
 a114844a <=( (not A200)  and  A199 );
 a114847a <=( A202  and  (not A201) );
 a114848a <=( a114847a  and  a114844a );
 a114849a <=( a114848a  and  a114841a );
 a114852a <=( A266  and  A265 );
 a114855a <=( (not A269)  and  A268 );
 a114856a <=( a114855a  and  a114852a );
 a114859a <=( A299  and  A298 );
 a114862a <=( (not A301)  and  (not A300) );
 a114863a <=( a114862a  and  a114859a );
 a114864a <=( a114863a  and  a114856a );
 a114868a <=( (not A167)  and  (not A169) );
 a114869a <=( (not A170)  and  a114868a );
 a114872a <=( (not A200)  and  A199 );
 a114875a <=( A202  and  (not A201) );
 a114876a <=( a114875a  and  a114872a );
 a114877a <=( a114876a  and  a114869a );
 a114880a <=( A266  and  A265 );
 a114883a <=( (not A269)  and  A268 );
 a114884a <=( a114883a  and  a114880a );
 a114887a <=( A299  and  A298 );
 a114890a <=( A302  and  (not A300) );
 a114891a <=( a114890a  and  a114887a );
 a114892a <=( a114891a  and  a114884a );
 a114896a <=( (not A167)  and  (not A169) );
 a114897a <=( (not A170)  and  a114896a );
 a114900a <=( (not A200)  and  A199 );
 a114903a <=( A202  and  (not A201) );
 a114904a <=( a114903a  and  a114900a );
 a114905a <=( a114904a  and  a114897a );
 a114908a <=( A266  and  A265 );
 a114911a <=( (not A269)  and  A268 );
 a114912a <=( a114911a  and  a114908a );
 a114915a <=( (not A299)  and  A298 );
 a114918a <=( A301  and  (not A300) );
 a114919a <=( a114918a  and  a114915a );
 a114920a <=( a114919a  and  a114912a );
 a114924a <=( (not A167)  and  (not A169) );
 a114925a <=( (not A170)  and  a114924a );
 a114928a <=( (not A200)  and  A199 );
 a114931a <=( A202  and  (not A201) );
 a114932a <=( a114931a  and  a114928a );
 a114933a <=( a114932a  and  a114925a );
 a114936a <=( A266  and  A265 );
 a114939a <=( (not A269)  and  A268 );
 a114940a <=( a114939a  and  a114936a );
 a114943a <=( (not A299)  and  A298 );
 a114946a <=( (not A302)  and  (not A300) );
 a114947a <=( a114946a  and  a114943a );
 a114948a <=( a114947a  and  a114940a );
 a114952a <=( (not A167)  and  (not A169) );
 a114953a <=( (not A170)  and  a114952a );
 a114956a <=( (not A200)  and  A199 );
 a114959a <=( A202  and  (not A201) );
 a114960a <=( a114959a  and  a114956a );
 a114961a <=( a114960a  and  a114953a );
 a114964a <=( A266  and  A265 );
 a114967a <=( (not A269)  and  A268 );
 a114968a <=( a114967a  and  a114964a );
 a114971a <=( A299  and  (not A298) );
 a114974a <=( A301  and  (not A300) );
 a114975a <=( a114974a  and  a114971a );
 a114976a <=( a114975a  and  a114968a );
 a114980a <=( (not A167)  and  (not A169) );
 a114981a <=( (not A170)  and  a114980a );
 a114984a <=( (not A200)  and  A199 );
 a114987a <=( A202  and  (not A201) );
 a114988a <=( a114987a  and  a114984a );
 a114989a <=( a114988a  and  a114981a );
 a114992a <=( A266  and  A265 );
 a114995a <=( (not A269)  and  A268 );
 a114996a <=( a114995a  and  a114992a );
 a114999a <=( A299  and  (not A298) );
 a115002a <=( (not A302)  and  (not A300) );
 a115003a <=( a115002a  and  a114999a );
 a115004a <=( a115003a  and  a114996a );
 a115008a <=( (not A167)  and  (not A169) );
 a115009a <=( (not A170)  and  a115008a );
 a115012a <=( (not A200)  and  A199 );
 a115015a <=( A202  and  (not A201) );
 a115016a <=( a115015a  and  a115012a );
 a115017a <=( a115016a  and  a115009a );
 a115020a <=( A266  and  (not A265) );
 a115023a <=( A269  and  (not A268) );
 a115024a <=( a115023a  and  a115020a );
 a115027a <=( A299  and  A298 );
 a115030a <=( (not A301)  and  (not A300) );
 a115031a <=( a115030a  and  a115027a );
 a115032a <=( a115031a  and  a115024a );
 a115036a <=( (not A167)  and  (not A169) );
 a115037a <=( (not A170)  and  a115036a );
 a115040a <=( (not A200)  and  A199 );
 a115043a <=( A202  and  (not A201) );
 a115044a <=( a115043a  and  a115040a );
 a115045a <=( a115044a  and  a115037a );
 a115048a <=( A266  and  (not A265) );
 a115051a <=( A269  and  (not A268) );
 a115052a <=( a115051a  and  a115048a );
 a115055a <=( A299  and  A298 );
 a115058a <=( A302  and  (not A300) );
 a115059a <=( a115058a  and  a115055a );
 a115060a <=( a115059a  and  a115052a );
 a115064a <=( (not A167)  and  (not A169) );
 a115065a <=( (not A170)  and  a115064a );
 a115068a <=( (not A200)  and  A199 );
 a115071a <=( A202  and  (not A201) );
 a115072a <=( a115071a  and  a115068a );
 a115073a <=( a115072a  and  a115065a );
 a115076a <=( A266  and  (not A265) );
 a115079a <=( A269  and  (not A268) );
 a115080a <=( a115079a  and  a115076a );
 a115083a <=( (not A299)  and  A298 );
 a115086a <=( A301  and  (not A300) );
 a115087a <=( a115086a  and  a115083a );
 a115088a <=( a115087a  and  a115080a );
 a115092a <=( (not A167)  and  (not A169) );
 a115093a <=( (not A170)  and  a115092a );
 a115096a <=( (not A200)  and  A199 );
 a115099a <=( A202  and  (not A201) );
 a115100a <=( a115099a  and  a115096a );
 a115101a <=( a115100a  and  a115093a );
 a115104a <=( A266  and  (not A265) );
 a115107a <=( A269  and  (not A268) );
 a115108a <=( a115107a  and  a115104a );
 a115111a <=( (not A299)  and  A298 );
 a115114a <=( (not A302)  and  (not A300) );
 a115115a <=( a115114a  and  a115111a );
 a115116a <=( a115115a  and  a115108a );
 a115120a <=( (not A167)  and  (not A169) );
 a115121a <=( (not A170)  and  a115120a );
 a115124a <=( (not A200)  and  A199 );
 a115127a <=( A202  and  (not A201) );
 a115128a <=( a115127a  and  a115124a );
 a115129a <=( a115128a  and  a115121a );
 a115132a <=( A266  and  (not A265) );
 a115135a <=( A269  and  (not A268) );
 a115136a <=( a115135a  and  a115132a );
 a115139a <=( A299  and  (not A298) );
 a115142a <=( A301  and  (not A300) );
 a115143a <=( a115142a  and  a115139a );
 a115144a <=( a115143a  and  a115136a );
 a115148a <=( (not A167)  and  (not A169) );
 a115149a <=( (not A170)  and  a115148a );
 a115152a <=( (not A200)  and  A199 );
 a115155a <=( A202  and  (not A201) );
 a115156a <=( a115155a  and  a115152a );
 a115157a <=( a115156a  and  a115149a );
 a115160a <=( A266  and  (not A265) );
 a115163a <=( A269  and  (not A268) );
 a115164a <=( a115163a  and  a115160a );
 a115167a <=( A299  and  (not A298) );
 a115170a <=( (not A302)  and  (not A300) );
 a115171a <=( a115170a  and  a115167a );
 a115172a <=( a115171a  and  a115164a );
 a115176a <=( (not A167)  and  (not A169) );
 a115177a <=( (not A170)  and  a115176a );
 a115180a <=( (not A200)  and  A199 );
 a115183a <=( A202  and  (not A201) );
 a115184a <=( a115183a  and  a115180a );
 a115185a <=( a115184a  and  a115177a );
 a115188a <=( (not A266)  and  A265 );
 a115191a <=( A269  and  (not A268) );
 a115192a <=( a115191a  and  a115188a );
 a115195a <=( A299  and  A298 );
 a115198a <=( (not A301)  and  (not A300) );
 a115199a <=( a115198a  and  a115195a );
 a115200a <=( a115199a  and  a115192a );
 a115204a <=( (not A167)  and  (not A169) );
 a115205a <=( (not A170)  and  a115204a );
 a115208a <=( (not A200)  and  A199 );
 a115211a <=( A202  and  (not A201) );
 a115212a <=( a115211a  and  a115208a );
 a115213a <=( a115212a  and  a115205a );
 a115216a <=( (not A266)  and  A265 );
 a115219a <=( A269  and  (not A268) );
 a115220a <=( a115219a  and  a115216a );
 a115223a <=( A299  and  A298 );
 a115226a <=( A302  and  (not A300) );
 a115227a <=( a115226a  and  a115223a );
 a115228a <=( a115227a  and  a115220a );
 a115232a <=( (not A167)  and  (not A169) );
 a115233a <=( (not A170)  and  a115232a );
 a115236a <=( (not A200)  and  A199 );
 a115239a <=( A202  and  (not A201) );
 a115240a <=( a115239a  and  a115236a );
 a115241a <=( a115240a  and  a115233a );
 a115244a <=( (not A266)  and  A265 );
 a115247a <=( A269  and  (not A268) );
 a115248a <=( a115247a  and  a115244a );
 a115251a <=( (not A299)  and  A298 );
 a115254a <=( A301  and  (not A300) );
 a115255a <=( a115254a  and  a115251a );
 a115256a <=( a115255a  and  a115248a );
 a115260a <=( (not A167)  and  (not A169) );
 a115261a <=( (not A170)  and  a115260a );
 a115264a <=( (not A200)  and  A199 );
 a115267a <=( A202  and  (not A201) );
 a115268a <=( a115267a  and  a115264a );
 a115269a <=( a115268a  and  a115261a );
 a115272a <=( (not A266)  and  A265 );
 a115275a <=( A269  and  (not A268) );
 a115276a <=( a115275a  and  a115272a );
 a115279a <=( (not A299)  and  A298 );
 a115282a <=( (not A302)  and  (not A300) );
 a115283a <=( a115282a  and  a115279a );
 a115284a <=( a115283a  and  a115276a );
 a115288a <=( (not A167)  and  (not A169) );
 a115289a <=( (not A170)  and  a115288a );
 a115292a <=( (not A200)  and  A199 );
 a115295a <=( A202  and  (not A201) );
 a115296a <=( a115295a  and  a115292a );
 a115297a <=( a115296a  and  a115289a );
 a115300a <=( (not A266)  and  A265 );
 a115303a <=( A269  and  (not A268) );
 a115304a <=( a115303a  and  a115300a );
 a115307a <=( A299  and  (not A298) );
 a115310a <=( A301  and  (not A300) );
 a115311a <=( a115310a  and  a115307a );
 a115312a <=( a115311a  and  a115304a );
 a115316a <=( (not A167)  and  (not A169) );
 a115317a <=( (not A170)  and  a115316a );
 a115320a <=( (not A200)  and  A199 );
 a115323a <=( A202  and  (not A201) );
 a115324a <=( a115323a  and  a115320a );
 a115325a <=( a115324a  and  a115317a );
 a115328a <=( (not A266)  and  A265 );
 a115331a <=( A269  and  (not A268) );
 a115332a <=( a115331a  and  a115328a );
 a115335a <=( A299  and  (not A298) );
 a115338a <=( (not A302)  and  (not A300) );
 a115339a <=( a115338a  and  a115335a );
 a115340a <=( a115339a  and  a115332a );
 a115344a <=( (not A167)  and  (not A169) );
 a115345a <=( (not A170)  and  a115344a );
 a115348a <=( (not A200)  and  A199 );
 a115351a <=( A202  and  (not A201) );
 a115352a <=( a115351a  and  a115348a );
 a115353a <=( a115352a  and  a115345a );
 a115356a <=( (not A266)  and  (not A265) );
 a115359a <=( (not A269)  and  A268 );
 a115360a <=( a115359a  and  a115356a );
 a115363a <=( A299  and  A298 );
 a115366a <=( (not A301)  and  (not A300) );
 a115367a <=( a115366a  and  a115363a );
 a115368a <=( a115367a  and  a115360a );
 a115372a <=( (not A167)  and  (not A169) );
 a115373a <=( (not A170)  and  a115372a );
 a115376a <=( (not A200)  and  A199 );
 a115379a <=( A202  and  (not A201) );
 a115380a <=( a115379a  and  a115376a );
 a115381a <=( a115380a  and  a115373a );
 a115384a <=( (not A266)  and  (not A265) );
 a115387a <=( (not A269)  and  A268 );
 a115388a <=( a115387a  and  a115384a );
 a115391a <=( A299  and  A298 );
 a115394a <=( A302  and  (not A300) );
 a115395a <=( a115394a  and  a115391a );
 a115396a <=( a115395a  and  a115388a );
 a115400a <=( (not A167)  and  (not A169) );
 a115401a <=( (not A170)  and  a115400a );
 a115404a <=( (not A200)  and  A199 );
 a115407a <=( A202  and  (not A201) );
 a115408a <=( a115407a  and  a115404a );
 a115409a <=( a115408a  and  a115401a );
 a115412a <=( (not A266)  and  (not A265) );
 a115415a <=( (not A269)  and  A268 );
 a115416a <=( a115415a  and  a115412a );
 a115419a <=( (not A299)  and  A298 );
 a115422a <=( A301  and  (not A300) );
 a115423a <=( a115422a  and  a115419a );
 a115424a <=( a115423a  and  a115416a );
 a115428a <=( (not A167)  and  (not A169) );
 a115429a <=( (not A170)  and  a115428a );
 a115432a <=( (not A200)  and  A199 );
 a115435a <=( A202  and  (not A201) );
 a115436a <=( a115435a  and  a115432a );
 a115437a <=( a115436a  and  a115429a );
 a115440a <=( (not A266)  and  (not A265) );
 a115443a <=( (not A269)  and  A268 );
 a115444a <=( a115443a  and  a115440a );
 a115447a <=( (not A299)  and  A298 );
 a115450a <=( (not A302)  and  (not A300) );
 a115451a <=( a115450a  and  a115447a );
 a115452a <=( a115451a  and  a115444a );
 a115456a <=( (not A167)  and  (not A169) );
 a115457a <=( (not A170)  and  a115456a );
 a115460a <=( (not A200)  and  A199 );
 a115463a <=( A202  and  (not A201) );
 a115464a <=( a115463a  and  a115460a );
 a115465a <=( a115464a  and  a115457a );
 a115468a <=( (not A266)  and  (not A265) );
 a115471a <=( (not A269)  and  A268 );
 a115472a <=( a115471a  and  a115468a );
 a115475a <=( A299  and  (not A298) );
 a115478a <=( A301  and  (not A300) );
 a115479a <=( a115478a  and  a115475a );
 a115480a <=( a115479a  and  a115472a );
 a115484a <=( (not A167)  and  (not A169) );
 a115485a <=( (not A170)  and  a115484a );
 a115488a <=( (not A200)  and  A199 );
 a115491a <=( A202  and  (not A201) );
 a115492a <=( a115491a  and  a115488a );
 a115493a <=( a115492a  and  a115485a );
 a115496a <=( (not A266)  and  (not A265) );
 a115499a <=( (not A269)  and  A268 );
 a115500a <=( a115499a  and  a115496a );
 a115503a <=( A299  and  (not A298) );
 a115506a <=( (not A302)  and  (not A300) );
 a115507a <=( a115506a  and  a115503a );
 a115508a <=( a115507a  and  a115500a );
 a115512a <=( (not A167)  and  (not A169) );
 a115513a <=( (not A170)  and  a115512a );
 a115516a <=( (not A200)  and  A199 );
 a115519a <=( (not A203)  and  (not A201) );
 a115520a <=( a115519a  and  a115516a );
 a115521a <=( a115520a  and  a115513a );
 a115524a <=( A266  and  A265 );
 a115527a <=( (not A269)  and  A268 );
 a115528a <=( a115527a  and  a115524a );
 a115531a <=( A299  and  A298 );
 a115534a <=( (not A301)  and  (not A300) );
 a115535a <=( a115534a  and  a115531a );
 a115536a <=( a115535a  and  a115528a );
 a115540a <=( (not A167)  and  (not A169) );
 a115541a <=( (not A170)  and  a115540a );
 a115544a <=( (not A200)  and  A199 );
 a115547a <=( (not A203)  and  (not A201) );
 a115548a <=( a115547a  and  a115544a );
 a115549a <=( a115548a  and  a115541a );
 a115552a <=( A266  and  A265 );
 a115555a <=( (not A269)  and  A268 );
 a115556a <=( a115555a  and  a115552a );
 a115559a <=( A299  and  A298 );
 a115562a <=( A302  and  (not A300) );
 a115563a <=( a115562a  and  a115559a );
 a115564a <=( a115563a  and  a115556a );
 a115568a <=( (not A167)  and  (not A169) );
 a115569a <=( (not A170)  and  a115568a );
 a115572a <=( (not A200)  and  A199 );
 a115575a <=( (not A203)  and  (not A201) );
 a115576a <=( a115575a  and  a115572a );
 a115577a <=( a115576a  and  a115569a );
 a115580a <=( A266  and  A265 );
 a115583a <=( (not A269)  and  A268 );
 a115584a <=( a115583a  and  a115580a );
 a115587a <=( (not A299)  and  A298 );
 a115590a <=( A301  and  (not A300) );
 a115591a <=( a115590a  and  a115587a );
 a115592a <=( a115591a  and  a115584a );
 a115596a <=( (not A167)  and  (not A169) );
 a115597a <=( (not A170)  and  a115596a );
 a115600a <=( (not A200)  and  A199 );
 a115603a <=( (not A203)  and  (not A201) );
 a115604a <=( a115603a  and  a115600a );
 a115605a <=( a115604a  and  a115597a );
 a115608a <=( A266  and  A265 );
 a115611a <=( (not A269)  and  A268 );
 a115612a <=( a115611a  and  a115608a );
 a115615a <=( (not A299)  and  A298 );
 a115618a <=( (not A302)  and  (not A300) );
 a115619a <=( a115618a  and  a115615a );
 a115620a <=( a115619a  and  a115612a );
 a115624a <=( (not A167)  and  (not A169) );
 a115625a <=( (not A170)  and  a115624a );
 a115628a <=( (not A200)  and  A199 );
 a115631a <=( (not A203)  and  (not A201) );
 a115632a <=( a115631a  and  a115628a );
 a115633a <=( a115632a  and  a115625a );
 a115636a <=( A266  and  A265 );
 a115639a <=( (not A269)  and  A268 );
 a115640a <=( a115639a  and  a115636a );
 a115643a <=( A299  and  (not A298) );
 a115646a <=( A301  and  (not A300) );
 a115647a <=( a115646a  and  a115643a );
 a115648a <=( a115647a  and  a115640a );
 a115652a <=( (not A167)  and  (not A169) );
 a115653a <=( (not A170)  and  a115652a );
 a115656a <=( (not A200)  and  A199 );
 a115659a <=( (not A203)  and  (not A201) );
 a115660a <=( a115659a  and  a115656a );
 a115661a <=( a115660a  and  a115653a );
 a115664a <=( A266  and  A265 );
 a115667a <=( (not A269)  and  A268 );
 a115668a <=( a115667a  and  a115664a );
 a115671a <=( A299  and  (not A298) );
 a115674a <=( (not A302)  and  (not A300) );
 a115675a <=( a115674a  and  a115671a );
 a115676a <=( a115675a  and  a115668a );
 a115680a <=( (not A167)  and  (not A169) );
 a115681a <=( (not A170)  and  a115680a );
 a115684a <=( (not A200)  and  A199 );
 a115687a <=( (not A203)  and  (not A201) );
 a115688a <=( a115687a  and  a115684a );
 a115689a <=( a115688a  and  a115681a );
 a115692a <=( A266  and  (not A265) );
 a115695a <=( A269  and  (not A268) );
 a115696a <=( a115695a  and  a115692a );
 a115699a <=( A299  and  A298 );
 a115702a <=( (not A301)  and  (not A300) );
 a115703a <=( a115702a  and  a115699a );
 a115704a <=( a115703a  and  a115696a );
 a115708a <=( (not A167)  and  (not A169) );
 a115709a <=( (not A170)  and  a115708a );
 a115712a <=( (not A200)  and  A199 );
 a115715a <=( (not A203)  and  (not A201) );
 a115716a <=( a115715a  and  a115712a );
 a115717a <=( a115716a  and  a115709a );
 a115720a <=( A266  and  (not A265) );
 a115723a <=( A269  and  (not A268) );
 a115724a <=( a115723a  and  a115720a );
 a115727a <=( A299  and  A298 );
 a115730a <=( A302  and  (not A300) );
 a115731a <=( a115730a  and  a115727a );
 a115732a <=( a115731a  and  a115724a );
 a115736a <=( (not A167)  and  (not A169) );
 a115737a <=( (not A170)  and  a115736a );
 a115740a <=( (not A200)  and  A199 );
 a115743a <=( (not A203)  and  (not A201) );
 a115744a <=( a115743a  and  a115740a );
 a115745a <=( a115744a  and  a115737a );
 a115748a <=( A266  and  (not A265) );
 a115751a <=( A269  and  (not A268) );
 a115752a <=( a115751a  and  a115748a );
 a115755a <=( (not A299)  and  A298 );
 a115758a <=( A301  and  (not A300) );
 a115759a <=( a115758a  and  a115755a );
 a115760a <=( a115759a  and  a115752a );
 a115764a <=( (not A167)  and  (not A169) );
 a115765a <=( (not A170)  and  a115764a );
 a115768a <=( (not A200)  and  A199 );
 a115771a <=( (not A203)  and  (not A201) );
 a115772a <=( a115771a  and  a115768a );
 a115773a <=( a115772a  and  a115765a );
 a115776a <=( A266  and  (not A265) );
 a115779a <=( A269  and  (not A268) );
 a115780a <=( a115779a  and  a115776a );
 a115783a <=( (not A299)  and  A298 );
 a115786a <=( (not A302)  and  (not A300) );
 a115787a <=( a115786a  and  a115783a );
 a115788a <=( a115787a  and  a115780a );
 a115792a <=( (not A167)  and  (not A169) );
 a115793a <=( (not A170)  and  a115792a );
 a115796a <=( (not A200)  and  A199 );
 a115799a <=( (not A203)  and  (not A201) );
 a115800a <=( a115799a  and  a115796a );
 a115801a <=( a115800a  and  a115793a );
 a115804a <=( A266  and  (not A265) );
 a115807a <=( A269  and  (not A268) );
 a115808a <=( a115807a  and  a115804a );
 a115811a <=( A299  and  (not A298) );
 a115814a <=( A301  and  (not A300) );
 a115815a <=( a115814a  and  a115811a );
 a115816a <=( a115815a  and  a115808a );
 a115820a <=( (not A167)  and  (not A169) );
 a115821a <=( (not A170)  and  a115820a );
 a115824a <=( (not A200)  and  A199 );
 a115827a <=( (not A203)  and  (not A201) );
 a115828a <=( a115827a  and  a115824a );
 a115829a <=( a115828a  and  a115821a );
 a115832a <=( A266  and  (not A265) );
 a115835a <=( A269  and  (not A268) );
 a115836a <=( a115835a  and  a115832a );
 a115839a <=( A299  and  (not A298) );
 a115842a <=( (not A302)  and  (not A300) );
 a115843a <=( a115842a  and  a115839a );
 a115844a <=( a115843a  and  a115836a );
 a115848a <=( (not A167)  and  (not A169) );
 a115849a <=( (not A170)  and  a115848a );
 a115852a <=( (not A200)  and  A199 );
 a115855a <=( (not A203)  and  (not A201) );
 a115856a <=( a115855a  and  a115852a );
 a115857a <=( a115856a  and  a115849a );
 a115860a <=( (not A266)  and  A265 );
 a115863a <=( A269  and  (not A268) );
 a115864a <=( a115863a  and  a115860a );
 a115867a <=( A299  and  A298 );
 a115870a <=( (not A301)  and  (not A300) );
 a115871a <=( a115870a  and  a115867a );
 a115872a <=( a115871a  and  a115864a );
 a115876a <=( (not A167)  and  (not A169) );
 a115877a <=( (not A170)  and  a115876a );
 a115880a <=( (not A200)  and  A199 );
 a115883a <=( (not A203)  and  (not A201) );
 a115884a <=( a115883a  and  a115880a );
 a115885a <=( a115884a  and  a115877a );
 a115888a <=( (not A266)  and  A265 );
 a115891a <=( A269  and  (not A268) );
 a115892a <=( a115891a  and  a115888a );
 a115895a <=( A299  and  A298 );
 a115898a <=( A302  and  (not A300) );
 a115899a <=( a115898a  and  a115895a );
 a115900a <=( a115899a  and  a115892a );
 a115904a <=( (not A167)  and  (not A169) );
 a115905a <=( (not A170)  and  a115904a );
 a115908a <=( (not A200)  and  A199 );
 a115911a <=( (not A203)  and  (not A201) );
 a115912a <=( a115911a  and  a115908a );
 a115913a <=( a115912a  and  a115905a );
 a115916a <=( (not A266)  and  A265 );
 a115919a <=( A269  and  (not A268) );
 a115920a <=( a115919a  and  a115916a );
 a115923a <=( (not A299)  and  A298 );
 a115926a <=( A301  and  (not A300) );
 a115927a <=( a115926a  and  a115923a );
 a115928a <=( a115927a  and  a115920a );
 a115932a <=( (not A167)  and  (not A169) );
 a115933a <=( (not A170)  and  a115932a );
 a115936a <=( (not A200)  and  A199 );
 a115939a <=( (not A203)  and  (not A201) );
 a115940a <=( a115939a  and  a115936a );
 a115941a <=( a115940a  and  a115933a );
 a115944a <=( (not A266)  and  A265 );
 a115947a <=( A269  and  (not A268) );
 a115948a <=( a115947a  and  a115944a );
 a115951a <=( (not A299)  and  A298 );
 a115954a <=( (not A302)  and  (not A300) );
 a115955a <=( a115954a  and  a115951a );
 a115956a <=( a115955a  and  a115948a );
 a115960a <=( (not A167)  and  (not A169) );
 a115961a <=( (not A170)  and  a115960a );
 a115964a <=( (not A200)  and  A199 );
 a115967a <=( (not A203)  and  (not A201) );
 a115968a <=( a115967a  and  a115964a );
 a115969a <=( a115968a  and  a115961a );
 a115972a <=( (not A266)  and  A265 );
 a115975a <=( A269  and  (not A268) );
 a115976a <=( a115975a  and  a115972a );
 a115979a <=( A299  and  (not A298) );
 a115982a <=( A301  and  (not A300) );
 a115983a <=( a115982a  and  a115979a );
 a115984a <=( a115983a  and  a115976a );
 a115988a <=( (not A167)  and  (not A169) );
 a115989a <=( (not A170)  and  a115988a );
 a115992a <=( (not A200)  and  A199 );
 a115995a <=( (not A203)  and  (not A201) );
 a115996a <=( a115995a  and  a115992a );
 a115997a <=( a115996a  and  a115989a );
 a116000a <=( (not A266)  and  A265 );
 a116003a <=( A269  and  (not A268) );
 a116004a <=( a116003a  and  a116000a );
 a116007a <=( A299  and  (not A298) );
 a116010a <=( (not A302)  and  (not A300) );
 a116011a <=( a116010a  and  a116007a );
 a116012a <=( a116011a  and  a116004a );
 a116016a <=( (not A167)  and  (not A169) );
 a116017a <=( (not A170)  and  a116016a );
 a116020a <=( (not A200)  and  A199 );
 a116023a <=( (not A203)  and  (not A201) );
 a116024a <=( a116023a  and  a116020a );
 a116025a <=( a116024a  and  a116017a );
 a116028a <=( (not A266)  and  (not A265) );
 a116031a <=( (not A269)  and  A268 );
 a116032a <=( a116031a  and  a116028a );
 a116035a <=( A299  and  A298 );
 a116038a <=( (not A301)  and  (not A300) );
 a116039a <=( a116038a  and  a116035a );
 a116040a <=( a116039a  and  a116032a );
 a116044a <=( (not A167)  and  (not A169) );
 a116045a <=( (not A170)  and  a116044a );
 a116048a <=( (not A200)  and  A199 );
 a116051a <=( (not A203)  and  (not A201) );
 a116052a <=( a116051a  and  a116048a );
 a116053a <=( a116052a  and  a116045a );
 a116056a <=( (not A266)  and  (not A265) );
 a116059a <=( (not A269)  and  A268 );
 a116060a <=( a116059a  and  a116056a );
 a116063a <=( A299  and  A298 );
 a116066a <=( A302  and  (not A300) );
 a116067a <=( a116066a  and  a116063a );
 a116068a <=( a116067a  and  a116060a );
 a116072a <=( (not A167)  and  (not A169) );
 a116073a <=( (not A170)  and  a116072a );
 a116076a <=( (not A200)  and  A199 );
 a116079a <=( (not A203)  and  (not A201) );
 a116080a <=( a116079a  and  a116076a );
 a116081a <=( a116080a  and  a116073a );
 a116084a <=( (not A266)  and  (not A265) );
 a116087a <=( (not A269)  and  A268 );
 a116088a <=( a116087a  and  a116084a );
 a116091a <=( (not A299)  and  A298 );
 a116094a <=( A301  and  (not A300) );
 a116095a <=( a116094a  and  a116091a );
 a116096a <=( a116095a  and  a116088a );
 a116100a <=( (not A167)  and  (not A169) );
 a116101a <=( (not A170)  and  a116100a );
 a116104a <=( (not A200)  and  A199 );
 a116107a <=( (not A203)  and  (not A201) );
 a116108a <=( a116107a  and  a116104a );
 a116109a <=( a116108a  and  a116101a );
 a116112a <=( (not A266)  and  (not A265) );
 a116115a <=( (not A269)  and  A268 );
 a116116a <=( a116115a  and  a116112a );
 a116119a <=( (not A299)  and  A298 );
 a116122a <=( (not A302)  and  (not A300) );
 a116123a <=( a116122a  and  a116119a );
 a116124a <=( a116123a  and  a116116a );
 a116128a <=( (not A167)  and  (not A169) );
 a116129a <=( (not A170)  and  a116128a );
 a116132a <=( (not A200)  and  A199 );
 a116135a <=( (not A203)  and  (not A201) );
 a116136a <=( a116135a  and  a116132a );
 a116137a <=( a116136a  and  a116129a );
 a116140a <=( (not A266)  and  (not A265) );
 a116143a <=( (not A269)  and  A268 );
 a116144a <=( a116143a  and  a116140a );
 a116147a <=( A299  and  (not A298) );
 a116150a <=( A301  and  (not A300) );
 a116151a <=( a116150a  and  a116147a );
 a116152a <=( a116151a  and  a116144a );
 a116156a <=( (not A167)  and  (not A169) );
 a116157a <=( (not A170)  and  a116156a );
 a116160a <=( (not A200)  and  A199 );
 a116163a <=( (not A203)  and  (not A201) );
 a116164a <=( a116163a  and  a116160a );
 a116165a <=( a116164a  and  a116157a );
 a116168a <=( (not A266)  and  (not A265) );
 a116171a <=( (not A269)  and  A268 );
 a116172a <=( a116171a  and  a116168a );
 a116175a <=( A299  and  (not A298) );
 a116178a <=( (not A302)  and  (not A300) );
 a116179a <=( a116178a  and  a116175a );
 a116180a <=( a116179a  and  a116172a );
 a116184a <=( (not A167)  and  (not A169) );
 a116185a <=( (not A170)  and  a116184a );
 a116188a <=( (not A200)  and  (not A199) );
 a116191a <=( (not A203)  and  A202 );
 a116192a <=( a116191a  and  a116188a );
 a116193a <=( a116192a  and  a116185a );
 a116196a <=( A266  and  A265 );
 a116199a <=( (not A268)  and  (not A267) );
 a116200a <=( a116199a  and  a116196a );
 a116203a <=( A299  and  A298 );
 a116206a <=( (not A302)  and  A301 );
 a116207a <=( a116206a  and  a116203a );
 a116208a <=( a116207a  and  a116200a );
 a116212a <=( (not A167)  and  (not A169) );
 a116213a <=( (not A170)  and  a116212a );
 a116216a <=( (not A200)  and  (not A199) );
 a116219a <=( (not A203)  and  A202 );
 a116220a <=( a116219a  and  a116216a );
 a116221a <=( a116220a  and  a116213a );
 a116224a <=( A266  and  A265 );
 a116227a <=( (not A268)  and  (not A267) );
 a116228a <=( a116227a  and  a116224a );
 a116231a <=( (not A299)  and  A298 );
 a116234a <=( A302  and  (not A301) );
 a116235a <=( a116234a  and  a116231a );
 a116236a <=( a116235a  and  a116228a );
 a116240a <=( (not A167)  and  (not A169) );
 a116241a <=( (not A170)  and  a116240a );
 a116244a <=( (not A200)  and  (not A199) );
 a116247a <=( (not A203)  and  A202 );
 a116248a <=( a116247a  and  a116244a );
 a116249a <=( a116248a  and  a116241a );
 a116252a <=( A266  and  A265 );
 a116255a <=( (not A268)  and  (not A267) );
 a116256a <=( a116255a  and  a116252a );
 a116259a <=( A299  and  (not A298) );
 a116262a <=( A302  and  (not A301) );
 a116263a <=( a116262a  and  a116259a );
 a116264a <=( a116263a  and  a116256a );
 a116268a <=( (not A167)  and  (not A169) );
 a116269a <=( (not A170)  and  a116268a );
 a116272a <=( (not A200)  and  (not A199) );
 a116275a <=( (not A203)  and  A202 );
 a116276a <=( a116275a  and  a116272a );
 a116277a <=( a116276a  and  a116269a );
 a116280a <=( A266  and  A265 );
 a116283a <=( (not A268)  and  (not A267) );
 a116284a <=( a116283a  and  a116280a );
 a116287a <=( (not A299)  and  (not A298) );
 a116290a <=( (not A302)  and  A301 );
 a116291a <=( a116290a  and  a116287a );
 a116292a <=( a116291a  and  a116284a );
 a116296a <=( (not A167)  and  (not A169) );
 a116297a <=( (not A170)  and  a116296a );
 a116300a <=( (not A200)  and  (not A199) );
 a116303a <=( (not A203)  and  A202 );
 a116304a <=( a116303a  and  a116300a );
 a116305a <=( a116304a  and  a116297a );
 a116308a <=( A266  and  A265 );
 a116311a <=( A269  and  (not A267) );
 a116312a <=( a116311a  and  a116308a );
 a116315a <=( A299  and  A298 );
 a116318a <=( (not A302)  and  A301 );
 a116319a <=( a116318a  and  a116315a );
 a116320a <=( a116319a  and  a116312a );
 a116324a <=( (not A167)  and  (not A169) );
 a116325a <=( (not A170)  and  a116324a );
 a116328a <=( (not A200)  and  (not A199) );
 a116331a <=( (not A203)  and  A202 );
 a116332a <=( a116331a  and  a116328a );
 a116333a <=( a116332a  and  a116325a );
 a116336a <=( A266  and  A265 );
 a116339a <=( A269  and  (not A267) );
 a116340a <=( a116339a  and  a116336a );
 a116343a <=( (not A299)  and  A298 );
 a116346a <=( A302  and  (not A301) );
 a116347a <=( a116346a  and  a116343a );
 a116348a <=( a116347a  and  a116340a );
 a116352a <=( (not A167)  and  (not A169) );
 a116353a <=( (not A170)  and  a116352a );
 a116356a <=( (not A200)  and  (not A199) );
 a116359a <=( (not A203)  and  A202 );
 a116360a <=( a116359a  and  a116356a );
 a116361a <=( a116360a  and  a116353a );
 a116364a <=( A266  and  A265 );
 a116367a <=( A269  and  (not A267) );
 a116368a <=( a116367a  and  a116364a );
 a116371a <=( A299  and  (not A298) );
 a116374a <=( A302  and  (not A301) );
 a116375a <=( a116374a  and  a116371a );
 a116376a <=( a116375a  and  a116368a );
 a116380a <=( (not A167)  and  (not A169) );
 a116381a <=( (not A170)  and  a116380a );
 a116384a <=( (not A200)  and  (not A199) );
 a116387a <=( (not A203)  and  A202 );
 a116388a <=( a116387a  and  a116384a );
 a116389a <=( a116388a  and  a116381a );
 a116392a <=( A266  and  A265 );
 a116395a <=( A269  and  (not A267) );
 a116396a <=( a116395a  and  a116392a );
 a116399a <=( (not A299)  and  (not A298) );
 a116402a <=( (not A302)  and  A301 );
 a116403a <=( a116402a  and  a116399a );
 a116404a <=( a116403a  and  a116396a );
 a116408a <=( (not A167)  and  (not A169) );
 a116409a <=( (not A170)  and  a116408a );
 a116412a <=( (not A200)  and  (not A199) );
 a116415a <=( (not A203)  and  A202 );
 a116416a <=( a116415a  and  a116412a );
 a116417a <=( a116416a  and  a116409a );
 a116420a <=( A266  and  (not A265) );
 a116423a <=( A268  and  (not A267) );
 a116424a <=( a116423a  and  a116420a );
 a116427a <=( A299  and  A298 );
 a116430a <=( (not A302)  and  A301 );
 a116431a <=( a116430a  and  a116427a );
 a116432a <=( a116431a  and  a116424a );
 a116436a <=( (not A167)  and  (not A169) );
 a116437a <=( (not A170)  and  a116436a );
 a116440a <=( (not A200)  and  (not A199) );
 a116443a <=( (not A203)  and  A202 );
 a116444a <=( a116443a  and  a116440a );
 a116445a <=( a116444a  and  a116437a );
 a116448a <=( A266  and  (not A265) );
 a116451a <=( A268  and  (not A267) );
 a116452a <=( a116451a  and  a116448a );
 a116455a <=( (not A299)  and  A298 );
 a116458a <=( A302  and  (not A301) );
 a116459a <=( a116458a  and  a116455a );
 a116460a <=( a116459a  and  a116452a );
 a116464a <=( (not A167)  and  (not A169) );
 a116465a <=( (not A170)  and  a116464a );
 a116468a <=( (not A200)  and  (not A199) );
 a116471a <=( (not A203)  and  A202 );
 a116472a <=( a116471a  and  a116468a );
 a116473a <=( a116472a  and  a116465a );
 a116476a <=( A266  and  (not A265) );
 a116479a <=( A268  and  (not A267) );
 a116480a <=( a116479a  and  a116476a );
 a116483a <=( A299  and  (not A298) );
 a116486a <=( A302  and  (not A301) );
 a116487a <=( a116486a  and  a116483a );
 a116488a <=( a116487a  and  a116480a );
 a116492a <=( (not A167)  and  (not A169) );
 a116493a <=( (not A170)  and  a116492a );
 a116496a <=( (not A200)  and  (not A199) );
 a116499a <=( (not A203)  and  A202 );
 a116500a <=( a116499a  and  a116496a );
 a116501a <=( a116500a  and  a116493a );
 a116504a <=( A266  and  (not A265) );
 a116507a <=( A268  and  (not A267) );
 a116508a <=( a116507a  and  a116504a );
 a116511a <=( (not A299)  and  (not A298) );
 a116514a <=( (not A302)  and  A301 );
 a116515a <=( a116514a  and  a116511a );
 a116516a <=( a116515a  and  a116508a );
 a116520a <=( (not A167)  and  (not A169) );
 a116521a <=( (not A170)  and  a116520a );
 a116524a <=( (not A200)  and  (not A199) );
 a116527a <=( (not A203)  and  A202 );
 a116528a <=( a116527a  and  a116524a );
 a116529a <=( a116528a  and  a116521a );
 a116532a <=( A266  and  (not A265) );
 a116535a <=( (not A269)  and  (not A267) );
 a116536a <=( a116535a  and  a116532a );
 a116539a <=( A299  and  A298 );
 a116542a <=( (not A302)  and  A301 );
 a116543a <=( a116542a  and  a116539a );
 a116544a <=( a116543a  and  a116536a );
 a116548a <=( (not A167)  and  (not A169) );
 a116549a <=( (not A170)  and  a116548a );
 a116552a <=( (not A200)  and  (not A199) );
 a116555a <=( (not A203)  and  A202 );
 a116556a <=( a116555a  and  a116552a );
 a116557a <=( a116556a  and  a116549a );
 a116560a <=( A266  and  (not A265) );
 a116563a <=( (not A269)  and  (not A267) );
 a116564a <=( a116563a  and  a116560a );
 a116567a <=( (not A299)  and  A298 );
 a116570a <=( A302  and  (not A301) );
 a116571a <=( a116570a  and  a116567a );
 a116572a <=( a116571a  and  a116564a );
 a116576a <=( (not A167)  and  (not A169) );
 a116577a <=( (not A170)  and  a116576a );
 a116580a <=( (not A200)  and  (not A199) );
 a116583a <=( (not A203)  and  A202 );
 a116584a <=( a116583a  and  a116580a );
 a116585a <=( a116584a  and  a116577a );
 a116588a <=( A266  and  (not A265) );
 a116591a <=( (not A269)  and  (not A267) );
 a116592a <=( a116591a  and  a116588a );
 a116595a <=( A299  and  (not A298) );
 a116598a <=( A302  and  (not A301) );
 a116599a <=( a116598a  and  a116595a );
 a116600a <=( a116599a  and  a116592a );
 a116604a <=( (not A167)  and  (not A169) );
 a116605a <=( (not A170)  and  a116604a );
 a116608a <=( (not A200)  and  (not A199) );
 a116611a <=( (not A203)  and  A202 );
 a116612a <=( a116611a  and  a116608a );
 a116613a <=( a116612a  and  a116605a );
 a116616a <=( A266  and  (not A265) );
 a116619a <=( (not A269)  and  (not A267) );
 a116620a <=( a116619a  and  a116616a );
 a116623a <=( (not A299)  and  (not A298) );
 a116626a <=( (not A302)  and  A301 );
 a116627a <=( a116626a  and  a116623a );
 a116628a <=( a116627a  and  a116620a );
 a116632a <=( (not A167)  and  (not A169) );
 a116633a <=( (not A170)  and  a116632a );
 a116636a <=( (not A200)  and  (not A199) );
 a116639a <=( (not A203)  and  A202 );
 a116640a <=( a116639a  and  a116636a );
 a116641a <=( a116640a  and  a116633a );
 a116644a <=( (not A266)  and  A265 );
 a116647a <=( A268  and  (not A267) );
 a116648a <=( a116647a  and  a116644a );
 a116651a <=( A299  and  A298 );
 a116654a <=( (not A302)  and  A301 );
 a116655a <=( a116654a  and  a116651a );
 a116656a <=( a116655a  and  a116648a );
 a116660a <=( (not A167)  and  (not A169) );
 a116661a <=( (not A170)  and  a116660a );
 a116664a <=( (not A200)  and  (not A199) );
 a116667a <=( (not A203)  and  A202 );
 a116668a <=( a116667a  and  a116664a );
 a116669a <=( a116668a  and  a116661a );
 a116672a <=( (not A266)  and  A265 );
 a116675a <=( A268  and  (not A267) );
 a116676a <=( a116675a  and  a116672a );
 a116679a <=( (not A299)  and  A298 );
 a116682a <=( A302  and  (not A301) );
 a116683a <=( a116682a  and  a116679a );
 a116684a <=( a116683a  and  a116676a );
 a116688a <=( (not A167)  and  (not A169) );
 a116689a <=( (not A170)  and  a116688a );
 a116692a <=( (not A200)  and  (not A199) );
 a116695a <=( (not A203)  and  A202 );
 a116696a <=( a116695a  and  a116692a );
 a116697a <=( a116696a  and  a116689a );
 a116700a <=( (not A266)  and  A265 );
 a116703a <=( A268  and  (not A267) );
 a116704a <=( a116703a  and  a116700a );
 a116707a <=( A299  and  (not A298) );
 a116710a <=( A302  and  (not A301) );
 a116711a <=( a116710a  and  a116707a );
 a116712a <=( a116711a  and  a116704a );
 a116716a <=( (not A167)  and  (not A169) );
 a116717a <=( (not A170)  and  a116716a );
 a116720a <=( (not A200)  and  (not A199) );
 a116723a <=( (not A203)  and  A202 );
 a116724a <=( a116723a  and  a116720a );
 a116725a <=( a116724a  and  a116717a );
 a116728a <=( (not A266)  and  A265 );
 a116731a <=( A268  and  (not A267) );
 a116732a <=( a116731a  and  a116728a );
 a116735a <=( (not A299)  and  (not A298) );
 a116738a <=( (not A302)  and  A301 );
 a116739a <=( a116738a  and  a116735a );
 a116740a <=( a116739a  and  a116732a );
 a116744a <=( (not A167)  and  (not A169) );
 a116745a <=( (not A170)  and  a116744a );
 a116748a <=( (not A200)  and  (not A199) );
 a116751a <=( (not A203)  and  A202 );
 a116752a <=( a116751a  and  a116748a );
 a116753a <=( a116752a  and  a116745a );
 a116756a <=( (not A266)  and  A265 );
 a116759a <=( (not A269)  and  (not A267) );
 a116760a <=( a116759a  and  a116756a );
 a116763a <=( A299  and  A298 );
 a116766a <=( (not A302)  and  A301 );
 a116767a <=( a116766a  and  a116763a );
 a116768a <=( a116767a  and  a116760a );
 a116772a <=( (not A167)  and  (not A169) );
 a116773a <=( (not A170)  and  a116772a );
 a116776a <=( (not A200)  and  (not A199) );
 a116779a <=( (not A203)  and  A202 );
 a116780a <=( a116779a  and  a116776a );
 a116781a <=( a116780a  and  a116773a );
 a116784a <=( (not A266)  and  A265 );
 a116787a <=( (not A269)  and  (not A267) );
 a116788a <=( a116787a  and  a116784a );
 a116791a <=( (not A299)  and  A298 );
 a116794a <=( A302  and  (not A301) );
 a116795a <=( a116794a  and  a116791a );
 a116796a <=( a116795a  and  a116788a );
 a116800a <=( (not A167)  and  (not A169) );
 a116801a <=( (not A170)  and  a116800a );
 a116804a <=( (not A200)  and  (not A199) );
 a116807a <=( (not A203)  and  A202 );
 a116808a <=( a116807a  and  a116804a );
 a116809a <=( a116808a  and  a116801a );
 a116812a <=( (not A266)  and  A265 );
 a116815a <=( (not A269)  and  (not A267) );
 a116816a <=( a116815a  and  a116812a );
 a116819a <=( A299  and  (not A298) );
 a116822a <=( A302  and  (not A301) );
 a116823a <=( a116822a  and  a116819a );
 a116824a <=( a116823a  and  a116816a );
 a116828a <=( (not A167)  and  (not A169) );
 a116829a <=( (not A170)  and  a116828a );
 a116832a <=( (not A200)  and  (not A199) );
 a116835a <=( (not A203)  and  A202 );
 a116836a <=( a116835a  and  a116832a );
 a116837a <=( a116836a  and  a116829a );
 a116840a <=( (not A266)  and  A265 );
 a116843a <=( (not A269)  and  (not A267) );
 a116844a <=( a116843a  and  a116840a );
 a116847a <=( (not A299)  and  (not A298) );
 a116850a <=( (not A302)  and  A301 );
 a116851a <=( a116850a  and  a116847a );
 a116852a <=( a116851a  and  a116844a );
 a116855a <=( A168  and  A170 );
 a116858a <=( A166  and  (not A167) );
 a116859a <=( a116858a  and  a116855a );
 a116862a <=( A200  and  A199 );
 a116865a <=( (not A203)  and  A202 );
 a116866a <=( a116865a  and  a116862a );
 a116867a <=( a116866a  and  a116859a );
 a116870a <=( A266  and  A265 );
 a116873a <=( (not A269)  and  A268 );
 a116874a <=( a116873a  and  a116870a );
 a116877a <=( A299  and  A298 );
 a116880a <=( (not A301)  and  (not A300) );
 a116881a <=( a116880a  and  a116877a );
 a116882a <=( a116881a  and  a116874a );
 a116885a <=( A168  and  A170 );
 a116888a <=( A166  and  (not A167) );
 a116889a <=( a116888a  and  a116885a );
 a116892a <=( A200  and  A199 );
 a116895a <=( (not A203)  and  A202 );
 a116896a <=( a116895a  and  a116892a );
 a116897a <=( a116896a  and  a116889a );
 a116900a <=( A266  and  A265 );
 a116903a <=( (not A269)  and  A268 );
 a116904a <=( a116903a  and  a116900a );
 a116907a <=( A299  and  A298 );
 a116910a <=( A302  and  (not A300) );
 a116911a <=( a116910a  and  a116907a );
 a116912a <=( a116911a  and  a116904a );
 a116915a <=( A168  and  A170 );
 a116918a <=( A166  and  (not A167) );
 a116919a <=( a116918a  and  a116915a );
 a116922a <=( A200  and  A199 );
 a116925a <=( (not A203)  and  A202 );
 a116926a <=( a116925a  and  a116922a );
 a116927a <=( a116926a  and  a116919a );
 a116930a <=( A266  and  A265 );
 a116933a <=( (not A269)  and  A268 );
 a116934a <=( a116933a  and  a116930a );
 a116937a <=( (not A299)  and  A298 );
 a116940a <=( A301  and  (not A300) );
 a116941a <=( a116940a  and  a116937a );
 a116942a <=( a116941a  and  a116934a );
 a116945a <=( A168  and  A170 );
 a116948a <=( A166  and  (not A167) );
 a116949a <=( a116948a  and  a116945a );
 a116952a <=( A200  and  A199 );
 a116955a <=( (not A203)  and  A202 );
 a116956a <=( a116955a  and  a116952a );
 a116957a <=( a116956a  and  a116949a );
 a116960a <=( A266  and  A265 );
 a116963a <=( (not A269)  and  A268 );
 a116964a <=( a116963a  and  a116960a );
 a116967a <=( (not A299)  and  A298 );
 a116970a <=( (not A302)  and  (not A300) );
 a116971a <=( a116970a  and  a116967a );
 a116972a <=( a116971a  and  a116964a );
 a116975a <=( A168  and  A170 );
 a116978a <=( A166  and  (not A167) );
 a116979a <=( a116978a  and  a116975a );
 a116982a <=( A200  and  A199 );
 a116985a <=( (not A203)  and  A202 );
 a116986a <=( a116985a  and  a116982a );
 a116987a <=( a116986a  and  a116979a );
 a116990a <=( A266  and  A265 );
 a116993a <=( (not A269)  and  A268 );
 a116994a <=( a116993a  and  a116990a );
 a116997a <=( A299  and  (not A298) );
 a117000a <=( A301  and  (not A300) );
 a117001a <=( a117000a  and  a116997a );
 a117002a <=( a117001a  and  a116994a );
 a117005a <=( A168  and  A170 );
 a117008a <=( A166  and  (not A167) );
 a117009a <=( a117008a  and  a117005a );
 a117012a <=( A200  and  A199 );
 a117015a <=( (not A203)  and  A202 );
 a117016a <=( a117015a  and  a117012a );
 a117017a <=( a117016a  and  a117009a );
 a117020a <=( A266  and  A265 );
 a117023a <=( (not A269)  and  A268 );
 a117024a <=( a117023a  and  a117020a );
 a117027a <=( A299  and  (not A298) );
 a117030a <=( (not A302)  and  (not A300) );
 a117031a <=( a117030a  and  a117027a );
 a117032a <=( a117031a  and  a117024a );
 a117035a <=( A168  and  A170 );
 a117038a <=( A166  and  (not A167) );
 a117039a <=( a117038a  and  a117035a );
 a117042a <=( A200  and  A199 );
 a117045a <=( (not A203)  and  A202 );
 a117046a <=( a117045a  and  a117042a );
 a117047a <=( a117046a  and  a117039a );
 a117050a <=( A266  and  (not A265) );
 a117053a <=( A269  and  (not A268) );
 a117054a <=( a117053a  and  a117050a );
 a117057a <=( A299  and  A298 );
 a117060a <=( (not A301)  and  (not A300) );
 a117061a <=( a117060a  and  a117057a );
 a117062a <=( a117061a  and  a117054a );
 a117065a <=( A168  and  A170 );
 a117068a <=( A166  and  (not A167) );
 a117069a <=( a117068a  and  a117065a );
 a117072a <=( A200  and  A199 );
 a117075a <=( (not A203)  and  A202 );
 a117076a <=( a117075a  and  a117072a );
 a117077a <=( a117076a  and  a117069a );
 a117080a <=( A266  and  (not A265) );
 a117083a <=( A269  and  (not A268) );
 a117084a <=( a117083a  and  a117080a );
 a117087a <=( A299  and  A298 );
 a117090a <=( A302  and  (not A300) );
 a117091a <=( a117090a  and  a117087a );
 a117092a <=( a117091a  and  a117084a );
 a117095a <=( A168  and  A170 );
 a117098a <=( A166  and  (not A167) );
 a117099a <=( a117098a  and  a117095a );
 a117102a <=( A200  and  A199 );
 a117105a <=( (not A203)  and  A202 );
 a117106a <=( a117105a  and  a117102a );
 a117107a <=( a117106a  and  a117099a );
 a117110a <=( A266  and  (not A265) );
 a117113a <=( A269  and  (not A268) );
 a117114a <=( a117113a  and  a117110a );
 a117117a <=( (not A299)  and  A298 );
 a117120a <=( A301  and  (not A300) );
 a117121a <=( a117120a  and  a117117a );
 a117122a <=( a117121a  and  a117114a );
 a117125a <=( A168  and  A170 );
 a117128a <=( A166  and  (not A167) );
 a117129a <=( a117128a  and  a117125a );
 a117132a <=( A200  and  A199 );
 a117135a <=( (not A203)  and  A202 );
 a117136a <=( a117135a  and  a117132a );
 a117137a <=( a117136a  and  a117129a );
 a117140a <=( A266  and  (not A265) );
 a117143a <=( A269  and  (not A268) );
 a117144a <=( a117143a  and  a117140a );
 a117147a <=( (not A299)  and  A298 );
 a117150a <=( (not A302)  and  (not A300) );
 a117151a <=( a117150a  and  a117147a );
 a117152a <=( a117151a  and  a117144a );
 a117155a <=( A168  and  A170 );
 a117158a <=( A166  and  (not A167) );
 a117159a <=( a117158a  and  a117155a );
 a117162a <=( A200  and  A199 );
 a117165a <=( (not A203)  and  A202 );
 a117166a <=( a117165a  and  a117162a );
 a117167a <=( a117166a  and  a117159a );
 a117170a <=( A266  and  (not A265) );
 a117173a <=( A269  and  (not A268) );
 a117174a <=( a117173a  and  a117170a );
 a117177a <=( A299  and  (not A298) );
 a117180a <=( A301  and  (not A300) );
 a117181a <=( a117180a  and  a117177a );
 a117182a <=( a117181a  and  a117174a );
 a117185a <=( A168  and  A170 );
 a117188a <=( A166  and  (not A167) );
 a117189a <=( a117188a  and  a117185a );
 a117192a <=( A200  and  A199 );
 a117195a <=( (not A203)  and  A202 );
 a117196a <=( a117195a  and  a117192a );
 a117197a <=( a117196a  and  a117189a );
 a117200a <=( A266  and  (not A265) );
 a117203a <=( A269  and  (not A268) );
 a117204a <=( a117203a  and  a117200a );
 a117207a <=( A299  and  (not A298) );
 a117210a <=( (not A302)  and  (not A300) );
 a117211a <=( a117210a  and  a117207a );
 a117212a <=( a117211a  and  a117204a );
 a117215a <=( A168  and  A170 );
 a117218a <=( A166  and  (not A167) );
 a117219a <=( a117218a  and  a117215a );
 a117222a <=( A200  and  A199 );
 a117225a <=( (not A203)  and  A202 );
 a117226a <=( a117225a  and  a117222a );
 a117227a <=( a117226a  and  a117219a );
 a117230a <=( (not A266)  and  A265 );
 a117233a <=( A269  and  (not A268) );
 a117234a <=( a117233a  and  a117230a );
 a117237a <=( A299  and  A298 );
 a117240a <=( (not A301)  and  (not A300) );
 a117241a <=( a117240a  and  a117237a );
 a117242a <=( a117241a  and  a117234a );
 a117245a <=( A168  and  A170 );
 a117248a <=( A166  and  (not A167) );
 a117249a <=( a117248a  and  a117245a );
 a117252a <=( A200  and  A199 );
 a117255a <=( (not A203)  and  A202 );
 a117256a <=( a117255a  and  a117252a );
 a117257a <=( a117256a  and  a117249a );
 a117260a <=( (not A266)  and  A265 );
 a117263a <=( A269  and  (not A268) );
 a117264a <=( a117263a  and  a117260a );
 a117267a <=( A299  and  A298 );
 a117270a <=( A302  and  (not A300) );
 a117271a <=( a117270a  and  a117267a );
 a117272a <=( a117271a  and  a117264a );
 a117275a <=( A168  and  A170 );
 a117278a <=( A166  and  (not A167) );
 a117279a <=( a117278a  and  a117275a );
 a117282a <=( A200  and  A199 );
 a117285a <=( (not A203)  and  A202 );
 a117286a <=( a117285a  and  a117282a );
 a117287a <=( a117286a  and  a117279a );
 a117290a <=( (not A266)  and  A265 );
 a117293a <=( A269  and  (not A268) );
 a117294a <=( a117293a  and  a117290a );
 a117297a <=( (not A299)  and  A298 );
 a117300a <=( A301  and  (not A300) );
 a117301a <=( a117300a  and  a117297a );
 a117302a <=( a117301a  and  a117294a );
 a117305a <=( A168  and  A170 );
 a117308a <=( A166  and  (not A167) );
 a117309a <=( a117308a  and  a117305a );
 a117312a <=( A200  and  A199 );
 a117315a <=( (not A203)  and  A202 );
 a117316a <=( a117315a  and  a117312a );
 a117317a <=( a117316a  and  a117309a );
 a117320a <=( (not A266)  and  A265 );
 a117323a <=( A269  and  (not A268) );
 a117324a <=( a117323a  and  a117320a );
 a117327a <=( (not A299)  and  A298 );
 a117330a <=( (not A302)  and  (not A300) );
 a117331a <=( a117330a  and  a117327a );
 a117332a <=( a117331a  and  a117324a );
 a117335a <=( A168  and  A170 );
 a117338a <=( A166  and  (not A167) );
 a117339a <=( a117338a  and  a117335a );
 a117342a <=( A200  and  A199 );
 a117345a <=( (not A203)  and  A202 );
 a117346a <=( a117345a  and  a117342a );
 a117347a <=( a117346a  and  a117339a );
 a117350a <=( (not A266)  and  A265 );
 a117353a <=( A269  and  (not A268) );
 a117354a <=( a117353a  and  a117350a );
 a117357a <=( A299  and  (not A298) );
 a117360a <=( A301  and  (not A300) );
 a117361a <=( a117360a  and  a117357a );
 a117362a <=( a117361a  and  a117354a );
 a117365a <=( A168  and  A170 );
 a117368a <=( A166  and  (not A167) );
 a117369a <=( a117368a  and  a117365a );
 a117372a <=( A200  and  A199 );
 a117375a <=( (not A203)  and  A202 );
 a117376a <=( a117375a  and  a117372a );
 a117377a <=( a117376a  and  a117369a );
 a117380a <=( (not A266)  and  A265 );
 a117383a <=( A269  and  (not A268) );
 a117384a <=( a117383a  and  a117380a );
 a117387a <=( A299  and  (not A298) );
 a117390a <=( (not A302)  and  (not A300) );
 a117391a <=( a117390a  and  a117387a );
 a117392a <=( a117391a  and  a117384a );
 a117395a <=( A168  and  A170 );
 a117398a <=( A166  and  (not A167) );
 a117399a <=( a117398a  and  a117395a );
 a117402a <=( A200  and  A199 );
 a117405a <=( (not A203)  and  A202 );
 a117406a <=( a117405a  and  a117402a );
 a117407a <=( a117406a  and  a117399a );
 a117410a <=( (not A266)  and  (not A265) );
 a117413a <=( (not A269)  and  A268 );
 a117414a <=( a117413a  and  a117410a );
 a117417a <=( A299  and  A298 );
 a117420a <=( (not A301)  and  (not A300) );
 a117421a <=( a117420a  and  a117417a );
 a117422a <=( a117421a  and  a117414a );
 a117425a <=( A168  and  A170 );
 a117428a <=( A166  and  (not A167) );
 a117429a <=( a117428a  and  a117425a );
 a117432a <=( A200  and  A199 );
 a117435a <=( (not A203)  and  A202 );
 a117436a <=( a117435a  and  a117432a );
 a117437a <=( a117436a  and  a117429a );
 a117440a <=( (not A266)  and  (not A265) );
 a117443a <=( (not A269)  and  A268 );
 a117444a <=( a117443a  and  a117440a );
 a117447a <=( A299  and  A298 );
 a117450a <=( A302  and  (not A300) );
 a117451a <=( a117450a  and  a117447a );
 a117452a <=( a117451a  and  a117444a );
 a117455a <=( A168  and  A170 );
 a117458a <=( A166  and  (not A167) );
 a117459a <=( a117458a  and  a117455a );
 a117462a <=( A200  and  A199 );
 a117465a <=( (not A203)  and  A202 );
 a117466a <=( a117465a  and  a117462a );
 a117467a <=( a117466a  and  a117459a );
 a117470a <=( (not A266)  and  (not A265) );
 a117473a <=( (not A269)  and  A268 );
 a117474a <=( a117473a  and  a117470a );
 a117477a <=( (not A299)  and  A298 );
 a117480a <=( A301  and  (not A300) );
 a117481a <=( a117480a  and  a117477a );
 a117482a <=( a117481a  and  a117474a );
 a117485a <=( A168  and  A170 );
 a117488a <=( A166  and  (not A167) );
 a117489a <=( a117488a  and  a117485a );
 a117492a <=( A200  and  A199 );
 a117495a <=( (not A203)  and  A202 );
 a117496a <=( a117495a  and  a117492a );
 a117497a <=( a117496a  and  a117489a );
 a117500a <=( (not A266)  and  (not A265) );
 a117503a <=( (not A269)  and  A268 );
 a117504a <=( a117503a  and  a117500a );
 a117507a <=( (not A299)  and  A298 );
 a117510a <=( (not A302)  and  (not A300) );
 a117511a <=( a117510a  and  a117507a );
 a117512a <=( a117511a  and  a117504a );
 a117515a <=( A168  and  A170 );
 a117518a <=( A166  and  (not A167) );
 a117519a <=( a117518a  and  a117515a );
 a117522a <=( A200  and  A199 );
 a117525a <=( (not A203)  and  A202 );
 a117526a <=( a117525a  and  a117522a );
 a117527a <=( a117526a  and  a117519a );
 a117530a <=( (not A266)  and  (not A265) );
 a117533a <=( (not A269)  and  A268 );
 a117534a <=( a117533a  and  a117530a );
 a117537a <=( A299  and  (not A298) );
 a117540a <=( A301  and  (not A300) );
 a117541a <=( a117540a  and  a117537a );
 a117542a <=( a117541a  and  a117534a );
 a117545a <=( A168  and  A170 );
 a117548a <=( A166  and  (not A167) );
 a117549a <=( a117548a  and  a117545a );
 a117552a <=( A200  and  A199 );
 a117555a <=( (not A203)  and  A202 );
 a117556a <=( a117555a  and  a117552a );
 a117557a <=( a117556a  and  a117549a );
 a117560a <=( (not A266)  and  (not A265) );
 a117563a <=( (not A269)  and  A268 );
 a117564a <=( a117563a  and  a117560a );
 a117567a <=( A299  and  (not A298) );
 a117570a <=( (not A302)  and  (not A300) );
 a117571a <=( a117570a  and  a117567a );
 a117572a <=( a117571a  and  a117564a );
 a117575a <=( A168  and  A170 );
 a117578a <=( A166  and  (not A167) );
 a117579a <=( a117578a  and  a117575a );
 a117582a <=( A200  and  A199 );
 a117585a <=( (not A202)  and  (not A201) );
 a117586a <=( a117585a  and  a117582a );
 a117587a <=( a117586a  and  a117579a );
 a117590a <=( A266  and  A265 );
 a117593a <=( (not A268)  and  (not A267) );
 a117594a <=( a117593a  and  a117590a );
 a117597a <=( A299  and  A298 );
 a117600a <=( (not A302)  and  A301 );
 a117601a <=( a117600a  and  a117597a );
 a117602a <=( a117601a  and  a117594a );
 a117605a <=( A168  and  A170 );
 a117608a <=( A166  and  (not A167) );
 a117609a <=( a117608a  and  a117605a );
 a117612a <=( A200  and  A199 );
 a117615a <=( (not A202)  and  (not A201) );
 a117616a <=( a117615a  and  a117612a );
 a117617a <=( a117616a  and  a117609a );
 a117620a <=( A266  and  A265 );
 a117623a <=( (not A268)  and  (not A267) );
 a117624a <=( a117623a  and  a117620a );
 a117627a <=( (not A299)  and  A298 );
 a117630a <=( A302  and  (not A301) );
 a117631a <=( a117630a  and  a117627a );
 a117632a <=( a117631a  and  a117624a );
 a117635a <=( A168  and  A170 );
 a117638a <=( A166  and  (not A167) );
 a117639a <=( a117638a  and  a117635a );
 a117642a <=( A200  and  A199 );
 a117645a <=( (not A202)  and  (not A201) );
 a117646a <=( a117645a  and  a117642a );
 a117647a <=( a117646a  and  a117639a );
 a117650a <=( A266  and  A265 );
 a117653a <=( (not A268)  and  (not A267) );
 a117654a <=( a117653a  and  a117650a );
 a117657a <=( A299  and  (not A298) );
 a117660a <=( A302  and  (not A301) );
 a117661a <=( a117660a  and  a117657a );
 a117662a <=( a117661a  and  a117654a );
 a117665a <=( A168  and  A170 );
 a117668a <=( A166  and  (not A167) );
 a117669a <=( a117668a  and  a117665a );
 a117672a <=( A200  and  A199 );
 a117675a <=( (not A202)  and  (not A201) );
 a117676a <=( a117675a  and  a117672a );
 a117677a <=( a117676a  and  a117669a );
 a117680a <=( A266  and  A265 );
 a117683a <=( (not A268)  and  (not A267) );
 a117684a <=( a117683a  and  a117680a );
 a117687a <=( (not A299)  and  (not A298) );
 a117690a <=( (not A302)  and  A301 );
 a117691a <=( a117690a  and  a117687a );
 a117692a <=( a117691a  and  a117684a );
 a117695a <=( A168  and  A170 );
 a117698a <=( A166  and  (not A167) );
 a117699a <=( a117698a  and  a117695a );
 a117702a <=( A200  and  A199 );
 a117705a <=( (not A202)  and  (not A201) );
 a117706a <=( a117705a  and  a117702a );
 a117707a <=( a117706a  and  a117699a );
 a117710a <=( A266  and  A265 );
 a117713a <=( A269  and  (not A267) );
 a117714a <=( a117713a  and  a117710a );
 a117717a <=( A299  and  A298 );
 a117720a <=( (not A302)  and  A301 );
 a117721a <=( a117720a  and  a117717a );
 a117722a <=( a117721a  and  a117714a );
 a117725a <=( A168  and  A170 );
 a117728a <=( A166  and  (not A167) );
 a117729a <=( a117728a  and  a117725a );
 a117732a <=( A200  and  A199 );
 a117735a <=( (not A202)  and  (not A201) );
 a117736a <=( a117735a  and  a117732a );
 a117737a <=( a117736a  and  a117729a );
 a117740a <=( A266  and  A265 );
 a117743a <=( A269  and  (not A267) );
 a117744a <=( a117743a  and  a117740a );
 a117747a <=( (not A299)  and  A298 );
 a117750a <=( A302  and  (not A301) );
 a117751a <=( a117750a  and  a117747a );
 a117752a <=( a117751a  and  a117744a );
 a117755a <=( A168  and  A170 );
 a117758a <=( A166  and  (not A167) );
 a117759a <=( a117758a  and  a117755a );
 a117762a <=( A200  and  A199 );
 a117765a <=( (not A202)  and  (not A201) );
 a117766a <=( a117765a  and  a117762a );
 a117767a <=( a117766a  and  a117759a );
 a117770a <=( A266  and  A265 );
 a117773a <=( A269  and  (not A267) );
 a117774a <=( a117773a  and  a117770a );
 a117777a <=( A299  and  (not A298) );
 a117780a <=( A302  and  (not A301) );
 a117781a <=( a117780a  and  a117777a );
 a117782a <=( a117781a  and  a117774a );
 a117785a <=( A168  and  A170 );
 a117788a <=( A166  and  (not A167) );
 a117789a <=( a117788a  and  a117785a );
 a117792a <=( A200  and  A199 );
 a117795a <=( (not A202)  and  (not A201) );
 a117796a <=( a117795a  and  a117792a );
 a117797a <=( a117796a  and  a117789a );
 a117800a <=( A266  and  A265 );
 a117803a <=( A269  and  (not A267) );
 a117804a <=( a117803a  and  a117800a );
 a117807a <=( (not A299)  and  (not A298) );
 a117810a <=( (not A302)  and  A301 );
 a117811a <=( a117810a  and  a117807a );
 a117812a <=( a117811a  and  a117804a );
 a117815a <=( A168  and  A170 );
 a117818a <=( A166  and  (not A167) );
 a117819a <=( a117818a  and  a117815a );
 a117822a <=( A200  and  A199 );
 a117825a <=( (not A202)  and  (not A201) );
 a117826a <=( a117825a  and  a117822a );
 a117827a <=( a117826a  and  a117819a );
 a117830a <=( A266  and  (not A265) );
 a117833a <=( A268  and  (not A267) );
 a117834a <=( a117833a  and  a117830a );
 a117837a <=( A299  and  A298 );
 a117840a <=( (not A302)  and  A301 );
 a117841a <=( a117840a  and  a117837a );
 a117842a <=( a117841a  and  a117834a );
 a117845a <=( A168  and  A170 );
 a117848a <=( A166  and  (not A167) );
 a117849a <=( a117848a  and  a117845a );
 a117852a <=( A200  and  A199 );
 a117855a <=( (not A202)  and  (not A201) );
 a117856a <=( a117855a  and  a117852a );
 a117857a <=( a117856a  and  a117849a );
 a117860a <=( A266  and  (not A265) );
 a117863a <=( A268  and  (not A267) );
 a117864a <=( a117863a  and  a117860a );
 a117867a <=( (not A299)  and  A298 );
 a117870a <=( A302  and  (not A301) );
 a117871a <=( a117870a  and  a117867a );
 a117872a <=( a117871a  and  a117864a );
 a117875a <=( A168  and  A170 );
 a117878a <=( A166  and  (not A167) );
 a117879a <=( a117878a  and  a117875a );
 a117882a <=( A200  and  A199 );
 a117885a <=( (not A202)  and  (not A201) );
 a117886a <=( a117885a  and  a117882a );
 a117887a <=( a117886a  and  a117879a );
 a117890a <=( A266  and  (not A265) );
 a117893a <=( A268  and  (not A267) );
 a117894a <=( a117893a  and  a117890a );
 a117897a <=( A299  and  (not A298) );
 a117900a <=( A302  and  (not A301) );
 a117901a <=( a117900a  and  a117897a );
 a117902a <=( a117901a  and  a117894a );
 a117905a <=( A168  and  A170 );
 a117908a <=( A166  and  (not A167) );
 a117909a <=( a117908a  and  a117905a );
 a117912a <=( A200  and  A199 );
 a117915a <=( (not A202)  and  (not A201) );
 a117916a <=( a117915a  and  a117912a );
 a117917a <=( a117916a  and  a117909a );
 a117920a <=( A266  and  (not A265) );
 a117923a <=( A268  and  (not A267) );
 a117924a <=( a117923a  and  a117920a );
 a117927a <=( (not A299)  and  (not A298) );
 a117930a <=( (not A302)  and  A301 );
 a117931a <=( a117930a  and  a117927a );
 a117932a <=( a117931a  and  a117924a );
 a117935a <=( A168  and  A170 );
 a117938a <=( A166  and  (not A167) );
 a117939a <=( a117938a  and  a117935a );
 a117942a <=( A200  and  A199 );
 a117945a <=( (not A202)  and  (not A201) );
 a117946a <=( a117945a  and  a117942a );
 a117947a <=( a117946a  and  a117939a );
 a117950a <=( A266  and  (not A265) );
 a117953a <=( (not A269)  and  (not A267) );
 a117954a <=( a117953a  and  a117950a );
 a117957a <=( A299  and  A298 );
 a117960a <=( (not A302)  and  A301 );
 a117961a <=( a117960a  and  a117957a );
 a117962a <=( a117961a  and  a117954a );
 a117965a <=( A168  and  A170 );
 a117968a <=( A166  and  (not A167) );
 a117969a <=( a117968a  and  a117965a );
 a117972a <=( A200  and  A199 );
 a117975a <=( (not A202)  and  (not A201) );
 a117976a <=( a117975a  and  a117972a );
 a117977a <=( a117976a  and  a117969a );
 a117980a <=( A266  and  (not A265) );
 a117983a <=( (not A269)  and  (not A267) );
 a117984a <=( a117983a  and  a117980a );
 a117987a <=( (not A299)  and  A298 );
 a117990a <=( A302  and  (not A301) );
 a117991a <=( a117990a  and  a117987a );
 a117992a <=( a117991a  and  a117984a );
 a117995a <=( A168  and  A170 );
 a117998a <=( A166  and  (not A167) );
 a117999a <=( a117998a  and  a117995a );
 a118002a <=( A200  and  A199 );
 a118005a <=( (not A202)  and  (not A201) );
 a118006a <=( a118005a  and  a118002a );
 a118007a <=( a118006a  and  a117999a );
 a118010a <=( A266  and  (not A265) );
 a118013a <=( (not A269)  and  (not A267) );
 a118014a <=( a118013a  and  a118010a );
 a118017a <=( A299  and  (not A298) );
 a118020a <=( A302  and  (not A301) );
 a118021a <=( a118020a  and  a118017a );
 a118022a <=( a118021a  and  a118014a );
 a118025a <=( A168  and  A170 );
 a118028a <=( A166  and  (not A167) );
 a118029a <=( a118028a  and  a118025a );
 a118032a <=( A200  and  A199 );
 a118035a <=( (not A202)  and  (not A201) );
 a118036a <=( a118035a  and  a118032a );
 a118037a <=( a118036a  and  a118029a );
 a118040a <=( A266  and  (not A265) );
 a118043a <=( (not A269)  and  (not A267) );
 a118044a <=( a118043a  and  a118040a );
 a118047a <=( (not A299)  and  (not A298) );
 a118050a <=( (not A302)  and  A301 );
 a118051a <=( a118050a  and  a118047a );
 a118052a <=( a118051a  and  a118044a );
 a118055a <=( A168  and  A170 );
 a118058a <=( A166  and  (not A167) );
 a118059a <=( a118058a  and  a118055a );
 a118062a <=( A200  and  A199 );
 a118065a <=( (not A202)  and  (not A201) );
 a118066a <=( a118065a  and  a118062a );
 a118067a <=( a118066a  and  a118059a );
 a118070a <=( (not A266)  and  A265 );
 a118073a <=( A268  and  (not A267) );
 a118074a <=( a118073a  and  a118070a );
 a118077a <=( A299  and  A298 );
 a118080a <=( (not A302)  and  A301 );
 a118081a <=( a118080a  and  a118077a );
 a118082a <=( a118081a  and  a118074a );
 a118085a <=( A168  and  A170 );
 a118088a <=( A166  and  (not A167) );
 a118089a <=( a118088a  and  a118085a );
 a118092a <=( A200  and  A199 );
 a118095a <=( (not A202)  and  (not A201) );
 a118096a <=( a118095a  and  a118092a );
 a118097a <=( a118096a  and  a118089a );
 a118100a <=( (not A266)  and  A265 );
 a118103a <=( A268  and  (not A267) );
 a118104a <=( a118103a  and  a118100a );
 a118107a <=( (not A299)  and  A298 );
 a118110a <=( A302  and  (not A301) );
 a118111a <=( a118110a  and  a118107a );
 a118112a <=( a118111a  and  a118104a );
 a118115a <=( A168  and  A170 );
 a118118a <=( A166  and  (not A167) );
 a118119a <=( a118118a  and  a118115a );
 a118122a <=( A200  and  A199 );
 a118125a <=( (not A202)  and  (not A201) );
 a118126a <=( a118125a  and  a118122a );
 a118127a <=( a118126a  and  a118119a );
 a118130a <=( (not A266)  and  A265 );
 a118133a <=( A268  and  (not A267) );
 a118134a <=( a118133a  and  a118130a );
 a118137a <=( A299  and  (not A298) );
 a118140a <=( A302  and  (not A301) );
 a118141a <=( a118140a  and  a118137a );
 a118142a <=( a118141a  and  a118134a );
 a118145a <=( A168  and  A170 );
 a118148a <=( A166  and  (not A167) );
 a118149a <=( a118148a  and  a118145a );
 a118152a <=( A200  and  A199 );
 a118155a <=( (not A202)  and  (not A201) );
 a118156a <=( a118155a  and  a118152a );
 a118157a <=( a118156a  and  a118149a );
 a118160a <=( (not A266)  and  A265 );
 a118163a <=( A268  and  (not A267) );
 a118164a <=( a118163a  and  a118160a );
 a118167a <=( (not A299)  and  (not A298) );
 a118170a <=( (not A302)  and  A301 );
 a118171a <=( a118170a  and  a118167a );
 a118172a <=( a118171a  and  a118164a );
 a118175a <=( A168  and  A170 );
 a118178a <=( A166  and  (not A167) );
 a118179a <=( a118178a  and  a118175a );
 a118182a <=( A200  and  A199 );
 a118185a <=( (not A202)  and  (not A201) );
 a118186a <=( a118185a  and  a118182a );
 a118187a <=( a118186a  and  a118179a );
 a118190a <=( (not A266)  and  A265 );
 a118193a <=( (not A269)  and  (not A267) );
 a118194a <=( a118193a  and  a118190a );
 a118197a <=( A299  and  A298 );
 a118200a <=( (not A302)  and  A301 );
 a118201a <=( a118200a  and  a118197a );
 a118202a <=( a118201a  and  a118194a );
 a118205a <=( A168  and  A170 );
 a118208a <=( A166  and  (not A167) );
 a118209a <=( a118208a  and  a118205a );
 a118212a <=( A200  and  A199 );
 a118215a <=( (not A202)  and  (not A201) );
 a118216a <=( a118215a  and  a118212a );
 a118217a <=( a118216a  and  a118209a );
 a118220a <=( (not A266)  and  A265 );
 a118223a <=( (not A269)  and  (not A267) );
 a118224a <=( a118223a  and  a118220a );
 a118227a <=( (not A299)  and  A298 );
 a118230a <=( A302  and  (not A301) );
 a118231a <=( a118230a  and  a118227a );
 a118232a <=( a118231a  and  a118224a );
 a118235a <=( A168  and  A170 );
 a118238a <=( A166  and  (not A167) );
 a118239a <=( a118238a  and  a118235a );
 a118242a <=( A200  and  A199 );
 a118245a <=( (not A202)  and  (not A201) );
 a118246a <=( a118245a  and  a118242a );
 a118247a <=( a118246a  and  a118239a );
 a118250a <=( (not A266)  and  A265 );
 a118253a <=( (not A269)  and  (not A267) );
 a118254a <=( a118253a  and  a118250a );
 a118257a <=( A299  and  (not A298) );
 a118260a <=( A302  and  (not A301) );
 a118261a <=( a118260a  and  a118257a );
 a118262a <=( a118261a  and  a118254a );
 a118265a <=( A168  and  A170 );
 a118268a <=( A166  and  (not A167) );
 a118269a <=( a118268a  and  a118265a );
 a118272a <=( A200  and  A199 );
 a118275a <=( (not A202)  and  (not A201) );
 a118276a <=( a118275a  and  a118272a );
 a118277a <=( a118276a  and  a118269a );
 a118280a <=( (not A266)  and  A265 );
 a118283a <=( (not A269)  and  (not A267) );
 a118284a <=( a118283a  and  a118280a );
 a118287a <=( (not A299)  and  (not A298) );
 a118290a <=( (not A302)  and  A301 );
 a118291a <=( a118290a  and  a118287a );
 a118292a <=( a118291a  and  a118284a );
 a118295a <=( A168  and  A170 );
 a118298a <=( A166  and  (not A167) );
 a118299a <=( a118298a  and  a118295a );
 a118302a <=( A200  and  A199 );
 a118305a <=( A203  and  (not A201) );
 a118306a <=( a118305a  and  a118302a );
 a118307a <=( a118306a  and  a118299a );
 a118310a <=( A266  and  A265 );
 a118313a <=( (not A268)  and  (not A267) );
 a118314a <=( a118313a  and  a118310a );
 a118317a <=( A299  and  A298 );
 a118320a <=( (not A302)  and  A301 );
 a118321a <=( a118320a  and  a118317a );
 a118322a <=( a118321a  and  a118314a );
 a118325a <=( A168  and  A170 );
 a118328a <=( A166  and  (not A167) );
 a118329a <=( a118328a  and  a118325a );
 a118332a <=( A200  and  A199 );
 a118335a <=( A203  and  (not A201) );
 a118336a <=( a118335a  and  a118332a );
 a118337a <=( a118336a  and  a118329a );
 a118340a <=( A266  and  A265 );
 a118343a <=( (not A268)  and  (not A267) );
 a118344a <=( a118343a  and  a118340a );
 a118347a <=( (not A299)  and  A298 );
 a118350a <=( A302  and  (not A301) );
 a118351a <=( a118350a  and  a118347a );
 a118352a <=( a118351a  and  a118344a );
 a118355a <=( A168  and  A170 );
 a118358a <=( A166  and  (not A167) );
 a118359a <=( a118358a  and  a118355a );
 a118362a <=( A200  and  A199 );
 a118365a <=( A203  and  (not A201) );
 a118366a <=( a118365a  and  a118362a );
 a118367a <=( a118366a  and  a118359a );
 a118370a <=( A266  and  A265 );
 a118373a <=( (not A268)  and  (not A267) );
 a118374a <=( a118373a  and  a118370a );
 a118377a <=( A299  and  (not A298) );
 a118380a <=( A302  and  (not A301) );
 a118381a <=( a118380a  and  a118377a );
 a118382a <=( a118381a  and  a118374a );
 a118385a <=( A168  and  A170 );
 a118388a <=( A166  and  (not A167) );
 a118389a <=( a118388a  and  a118385a );
 a118392a <=( A200  and  A199 );
 a118395a <=( A203  and  (not A201) );
 a118396a <=( a118395a  and  a118392a );
 a118397a <=( a118396a  and  a118389a );
 a118400a <=( A266  and  A265 );
 a118403a <=( (not A268)  and  (not A267) );
 a118404a <=( a118403a  and  a118400a );
 a118407a <=( (not A299)  and  (not A298) );
 a118410a <=( (not A302)  and  A301 );
 a118411a <=( a118410a  and  a118407a );
 a118412a <=( a118411a  and  a118404a );
 a118415a <=( A168  and  A170 );
 a118418a <=( A166  and  (not A167) );
 a118419a <=( a118418a  and  a118415a );
 a118422a <=( A200  and  A199 );
 a118425a <=( A203  and  (not A201) );
 a118426a <=( a118425a  and  a118422a );
 a118427a <=( a118426a  and  a118419a );
 a118430a <=( A266  and  A265 );
 a118433a <=( A269  and  (not A267) );
 a118434a <=( a118433a  and  a118430a );
 a118437a <=( A299  and  A298 );
 a118440a <=( (not A302)  and  A301 );
 a118441a <=( a118440a  and  a118437a );
 a118442a <=( a118441a  and  a118434a );
 a118445a <=( A168  and  A170 );
 a118448a <=( A166  and  (not A167) );
 a118449a <=( a118448a  and  a118445a );
 a118452a <=( A200  and  A199 );
 a118455a <=( A203  and  (not A201) );
 a118456a <=( a118455a  and  a118452a );
 a118457a <=( a118456a  and  a118449a );
 a118460a <=( A266  and  A265 );
 a118463a <=( A269  and  (not A267) );
 a118464a <=( a118463a  and  a118460a );
 a118467a <=( (not A299)  and  A298 );
 a118470a <=( A302  and  (not A301) );
 a118471a <=( a118470a  and  a118467a );
 a118472a <=( a118471a  and  a118464a );
 a118475a <=( A168  and  A170 );
 a118478a <=( A166  and  (not A167) );
 a118479a <=( a118478a  and  a118475a );
 a118482a <=( A200  and  A199 );
 a118485a <=( A203  and  (not A201) );
 a118486a <=( a118485a  and  a118482a );
 a118487a <=( a118486a  and  a118479a );
 a118490a <=( A266  and  A265 );
 a118493a <=( A269  and  (not A267) );
 a118494a <=( a118493a  and  a118490a );
 a118497a <=( A299  and  (not A298) );
 a118500a <=( A302  and  (not A301) );
 a118501a <=( a118500a  and  a118497a );
 a118502a <=( a118501a  and  a118494a );
 a118505a <=( A168  and  A170 );
 a118508a <=( A166  and  (not A167) );
 a118509a <=( a118508a  and  a118505a );
 a118512a <=( A200  and  A199 );
 a118515a <=( A203  and  (not A201) );
 a118516a <=( a118515a  and  a118512a );
 a118517a <=( a118516a  and  a118509a );
 a118520a <=( A266  and  A265 );
 a118523a <=( A269  and  (not A267) );
 a118524a <=( a118523a  and  a118520a );
 a118527a <=( (not A299)  and  (not A298) );
 a118530a <=( (not A302)  and  A301 );
 a118531a <=( a118530a  and  a118527a );
 a118532a <=( a118531a  and  a118524a );
 a118535a <=( A168  and  A170 );
 a118538a <=( A166  and  (not A167) );
 a118539a <=( a118538a  and  a118535a );
 a118542a <=( A200  and  A199 );
 a118545a <=( A203  and  (not A201) );
 a118546a <=( a118545a  and  a118542a );
 a118547a <=( a118546a  and  a118539a );
 a118550a <=( A266  and  (not A265) );
 a118553a <=( A268  and  (not A267) );
 a118554a <=( a118553a  and  a118550a );
 a118557a <=( A299  and  A298 );
 a118560a <=( (not A302)  and  A301 );
 a118561a <=( a118560a  and  a118557a );
 a118562a <=( a118561a  and  a118554a );
 a118565a <=( A168  and  A170 );
 a118568a <=( A166  and  (not A167) );
 a118569a <=( a118568a  and  a118565a );
 a118572a <=( A200  and  A199 );
 a118575a <=( A203  and  (not A201) );
 a118576a <=( a118575a  and  a118572a );
 a118577a <=( a118576a  and  a118569a );
 a118580a <=( A266  and  (not A265) );
 a118583a <=( A268  and  (not A267) );
 a118584a <=( a118583a  and  a118580a );
 a118587a <=( (not A299)  and  A298 );
 a118590a <=( A302  and  (not A301) );
 a118591a <=( a118590a  and  a118587a );
 a118592a <=( a118591a  and  a118584a );
 a118595a <=( A168  and  A170 );
 a118598a <=( A166  and  (not A167) );
 a118599a <=( a118598a  and  a118595a );
 a118602a <=( A200  and  A199 );
 a118605a <=( A203  and  (not A201) );
 a118606a <=( a118605a  and  a118602a );
 a118607a <=( a118606a  and  a118599a );
 a118610a <=( A266  and  (not A265) );
 a118613a <=( A268  and  (not A267) );
 a118614a <=( a118613a  and  a118610a );
 a118617a <=( A299  and  (not A298) );
 a118620a <=( A302  and  (not A301) );
 a118621a <=( a118620a  and  a118617a );
 a118622a <=( a118621a  and  a118614a );
 a118625a <=( A168  and  A170 );
 a118628a <=( A166  and  (not A167) );
 a118629a <=( a118628a  and  a118625a );
 a118632a <=( A200  and  A199 );
 a118635a <=( A203  and  (not A201) );
 a118636a <=( a118635a  and  a118632a );
 a118637a <=( a118636a  and  a118629a );
 a118640a <=( A266  and  (not A265) );
 a118643a <=( A268  and  (not A267) );
 a118644a <=( a118643a  and  a118640a );
 a118647a <=( (not A299)  and  (not A298) );
 a118650a <=( (not A302)  and  A301 );
 a118651a <=( a118650a  and  a118647a );
 a118652a <=( a118651a  and  a118644a );
 a118655a <=( A168  and  A170 );
 a118658a <=( A166  and  (not A167) );
 a118659a <=( a118658a  and  a118655a );
 a118662a <=( A200  and  A199 );
 a118665a <=( A203  and  (not A201) );
 a118666a <=( a118665a  and  a118662a );
 a118667a <=( a118666a  and  a118659a );
 a118670a <=( A266  and  (not A265) );
 a118673a <=( (not A269)  and  (not A267) );
 a118674a <=( a118673a  and  a118670a );
 a118677a <=( A299  and  A298 );
 a118680a <=( (not A302)  and  A301 );
 a118681a <=( a118680a  and  a118677a );
 a118682a <=( a118681a  and  a118674a );
 a118685a <=( A168  and  A170 );
 a118688a <=( A166  and  (not A167) );
 a118689a <=( a118688a  and  a118685a );
 a118692a <=( A200  and  A199 );
 a118695a <=( A203  and  (not A201) );
 a118696a <=( a118695a  and  a118692a );
 a118697a <=( a118696a  and  a118689a );
 a118700a <=( A266  and  (not A265) );
 a118703a <=( (not A269)  and  (not A267) );
 a118704a <=( a118703a  and  a118700a );
 a118707a <=( (not A299)  and  A298 );
 a118710a <=( A302  and  (not A301) );
 a118711a <=( a118710a  and  a118707a );
 a118712a <=( a118711a  and  a118704a );
 a118715a <=( A168  and  A170 );
 a118718a <=( A166  and  (not A167) );
 a118719a <=( a118718a  and  a118715a );
 a118722a <=( A200  and  A199 );
 a118725a <=( A203  and  (not A201) );
 a118726a <=( a118725a  and  a118722a );
 a118727a <=( a118726a  and  a118719a );
 a118730a <=( A266  and  (not A265) );
 a118733a <=( (not A269)  and  (not A267) );
 a118734a <=( a118733a  and  a118730a );
 a118737a <=( A299  and  (not A298) );
 a118740a <=( A302  and  (not A301) );
 a118741a <=( a118740a  and  a118737a );
 a118742a <=( a118741a  and  a118734a );
 a118745a <=( A168  and  A170 );
 a118748a <=( A166  and  (not A167) );
 a118749a <=( a118748a  and  a118745a );
 a118752a <=( A200  and  A199 );
 a118755a <=( A203  and  (not A201) );
 a118756a <=( a118755a  and  a118752a );
 a118757a <=( a118756a  and  a118749a );
 a118760a <=( A266  and  (not A265) );
 a118763a <=( (not A269)  and  (not A267) );
 a118764a <=( a118763a  and  a118760a );
 a118767a <=( (not A299)  and  (not A298) );
 a118770a <=( (not A302)  and  A301 );
 a118771a <=( a118770a  and  a118767a );
 a118772a <=( a118771a  and  a118764a );
 a118775a <=( A168  and  A170 );
 a118778a <=( A166  and  (not A167) );
 a118779a <=( a118778a  and  a118775a );
 a118782a <=( A200  and  A199 );
 a118785a <=( A203  and  (not A201) );
 a118786a <=( a118785a  and  a118782a );
 a118787a <=( a118786a  and  a118779a );
 a118790a <=( (not A266)  and  A265 );
 a118793a <=( A268  and  (not A267) );
 a118794a <=( a118793a  and  a118790a );
 a118797a <=( A299  and  A298 );
 a118800a <=( (not A302)  and  A301 );
 a118801a <=( a118800a  and  a118797a );
 a118802a <=( a118801a  and  a118794a );
 a118805a <=( A168  and  A170 );
 a118808a <=( A166  and  (not A167) );
 a118809a <=( a118808a  and  a118805a );
 a118812a <=( A200  and  A199 );
 a118815a <=( A203  and  (not A201) );
 a118816a <=( a118815a  and  a118812a );
 a118817a <=( a118816a  and  a118809a );
 a118820a <=( (not A266)  and  A265 );
 a118823a <=( A268  and  (not A267) );
 a118824a <=( a118823a  and  a118820a );
 a118827a <=( (not A299)  and  A298 );
 a118830a <=( A302  and  (not A301) );
 a118831a <=( a118830a  and  a118827a );
 a118832a <=( a118831a  and  a118824a );
 a118835a <=( A168  and  A170 );
 a118838a <=( A166  and  (not A167) );
 a118839a <=( a118838a  and  a118835a );
 a118842a <=( A200  and  A199 );
 a118845a <=( A203  and  (not A201) );
 a118846a <=( a118845a  and  a118842a );
 a118847a <=( a118846a  and  a118839a );
 a118850a <=( (not A266)  and  A265 );
 a118853a <=( A268  and  (not A267) );
 a118854a <=( a118853a  and  a118850a );
 a118857a <=( A299  and  (not A298) );
 a118860a <=( A302  and  (not A301) );
 a118861a <=( a118860a  and  a118857a );
 a118862a <=( a118861a  and  a118854a );
 a118865a <=( A168  and  A170 );
 a118868a <=( A166  and  (not A167) );
 a118869a <=( a118868a  and  a118865a );
 a118872a <=( A200  and  A199 );
 a118875a <=( A203  and  (not A201) );
 a118876a <=( a118875a  and  a118872a );
 a118877a <=( a118876a  and  a118869a );
 a118880a <=( (not A266)  and  A265 );
 a118883a <=( A268  and  (not A267) );
 a118884a <=( a118883a  and  a118880a );
 a118887a <=( (not A299)  and  (not A298) );
 a118890a <=( (not A302)  and  A301 );
 a118891a <=( a118890a  and  a118887a );
 a118892a <=( a118891a  and  a118884a );
 a118895a <=( A168  and  A170 );
 a118898a <=( A166  and  (not A167) );
 a118899a <=( a118898a  and  a118895a );
 a118902a <=( A200  and  A199 );
 a118905a <=( A203  and  (not A201) );
 a118906a <=( a118905a  and  a118902a );
 a118907a <=( a118906a  and  a118899a );
 a118910a <=( (not A266)  and  A265 );
 a118913a <=( (not A269)  and  (not A267) );
 a118914a <=( a118913a  and  a118910a );
 a118917a <=( A299  and  A298 );
 a118920a <=( (not A302)  and  A301 );
 a118921a <=( a118920a  and  a118917a );
 a118922a <=( a118921a  and  a118914a );
 a118925a <=( A168  and  A170 );
 a118928a <=( A166  and  (not A167) );
 a118929a <=( a118928a  and  a118925a );
 a118932a <=( A200  and  A199 );
 a118935a <=( A203  and  (not A201) );
 a118936a <=( a118935a  and  a118932a );
 a118937a <=( a118936a  and  a118929a );
 a118940a <=( (not A266)  and  A265 );
 a118943a <=( (not A269)  and  (not A267) );
 a118944a <=( a118943a  and  a118940a );
 a118947a <=( (not A299)  and  A298 );
 a118950a <=( A302  and  (not A301) );
 a118951a <=( a118950a  and  a118947a );
 a118952a <=( a118951a  and  a118944a );
 a118955a <=( A168  and  A170 );
 a118958a <=( A166  and  (not A167) );
 a118959a <=( a118958a  and  a118955a );
 a118962a <=( A200  and  A199 );
 a118965a <=( A203  and  (not A201) );
 a118966a <=( a118965a  and  a118962a );
 a118967a <=( a118966a  and  a118959a );
 a118970a <=( (not A266)  and  A265 );
 a118973a <=( (not A269)  and  (not A267) );
 a118974a <=( a118973a  and  a118970a );
 a118977a <=( A299  and  (not A298) );
 a118980a <=( A302  and  (not A301) );
 a118981a <=( a118980a  and  a118977a );
 a118982a <=( a118981a  and  a118974a );
 a118985a <=( A168  and  A170 );
 a118988a <=( A166  and  (not A167) );
 a118989a <=( a118988a  and  a118985a );
 a118992a <=( A200  and  A199 );
 a118995a <=( A203  and  (not A201) );
 a118996a <=( a118995a  and  a118992a );
 a118997a <=( a118996a  and  a118989a );
 a119000a <=( (not A266)  and  A265 );
 a119003a <=( (not A269)  and  (not A267) );
 a119004a <=( a119003a  and  a119000a );
 a119007a <=( (not A299)  and  (not A298) );
 a119010a <=( (not A302)  and  A301 );
 a119011a <=( a119010a  and  a119007a );
 a119012a <=( a119011a  and  a119004a );
 a119015a <=( A168  and  A170 );
 a119018a <=( A166  and  (not A167) );
 a119019a <=( a119018a  and  a119015a );
 a119022a <=( A200  and  (not A199) );
 a119025a <=( A203  and  (not A202) );
 a119026a <=( a119025a  and  a119022a );
 a119027a <=( a119026a  and  a119019a );
 a119030a <=( A266  and  A265 );
 a119033a <=( (not A269)  and  A268 );
 a119034a <=( a119033a  and  a119030a );
 a119037a <=( A299  and  A298 );
 a119040a <=( (not A301)  and  (not A300) );
 a119041a <=( a119040a  and  a119037a );
 a119042a <=( a119041a  and  a119034a );
 a119045a <=( A168  and  A170 );
 a119048a <=( A166  and  (not A167) );
 a119049a <=( a119048a  and  a119045a );
 a119052a <=( A200  and  (not A199) );
 a119055a <=( A203  and  (not A202) );
 a119056a <=( a119055a  and  a119052a );
 a119057a <=( a119056a  and  a119049a );
 a119060a <=( A266  and  A265 );
 a119063a <=( (not A269)  and  A268 );
 a119064a <=( a119063a  and  a119060a );
 a119067a <=( A299  and  A298 );
 a119070a <=( A302  and  (not A300) );
 a119071a <=( a119070a  and  a119067a );
 a119072a <=( a119071a  and  a119064a );
 a119075a <=( A168  and  A170 );
 a119078a <=( A166  and  (not A167) );
 a119079a <=( a119078a  and  a119075a );
 a119082a <=( A200  and  (not A199) );
 a119085a <=( A203  and  (not A202) );
 a119086a <=( a119085a  and  a119082a );
 a119087a <=( a119086a  and  a119079a );
 a119090a <=( A266  and  A265 );
 a119093a <=( (not A269)  and  A268 );
 a119094a <=( a119093a  and  a119090a );
 a119097a <=( (not A299)  and  A298 );
 a119100a <=( A301  and  (not A300) );
 a119101a <=( a119100a  and  a119097a );
 a119102a <=( a119101a  and  a119094a );
 a119105a <=( A168  and  A170 );
 a119108a <=( A166  and  (not A167) );
 a119109a <=( a119108a  and  a119105a );
 a119112a <=( A200  and  (not A199) );
 a119115a <=( A203  and  (not A202) );
 a119116a <=( a119115a  and  a119112a );
 a119117a <=( a119116a  and  a119109a );
 a119120a <=( A266  and  A265 );
 a119123a <=( (not A269)  and  A268 );
 a119124a <=( a119123a  and  a119120a );
 a119127a <=( (not A299)  and  A298 );
 a119130a <=( (not A302)  and  (not A300) );
 a119131a <=( a119130a  and  a119127a );
 a119132a <=( a119131a  and  a119124a );
 a119135a <=( A168  and  A170 );
 a119138a <=( A166  and  (not A167) );
 a119139a <=( a119138a  and  a119135a );
 a119142a <=( A200  and  (not A199) );
 a119145a <=( A203  and  (not A202) );
 a119146a <=( a119145a  and  a119142a );
 a119147a <=( a119146a  and  a119139a );
 a119150a <=( A266  and  A265 );
 a119153a <=( (not A269)  and  A268 );
 a119154a <=( a119153a  and  a119150a );
 a119157a <=( A299  and  (not A298) );
 a119160a <=( A301  and  (not A300) );
 a119161a <=( a119160a  and  a119157a );
 a119162a <=( a119161a  and  a119154a );
 a119165a <=( A168  and  A170 );
 a119168a <=( A166  and  (not A167) );
 a119169a <=( a119168a  and  a119165a );
 a119172a <=( A200  and  (not A199) );
 a119175a <=( A203  and  (not A202) );
 a119176a <=( a119175a  and  a119172a );
 a119177a <=( a119176a  and  a119169a );
 a119180a <=( A266  and  A265 );
 a119183a <=( (not A269)  and  A268 );
 a119184a <=( a119183a  and  a119180a );
 a119187a <=( A299  and  (not A298) );
 a119190a <=( (not A302)  and  (not A300) );
 a119191a <=( a119190a  and  a119187a );
 a119192a <=( a119191a  and  a119184a );
 a119195a <=( A168  and  A170 );
 a119198a <=( A166  and  (not A167) );
 a119199a <=( a119198a  and  a119195a );
 a119202a <=( A200  and  (not A199) );
 a119205a <=( A203  and  (not A202) );
 a119206a <=( a119205a  and  a119202a );
 a119207a <=( a119206a  and  a119199a );
 a119210a <=( A266  and  (not A265) );
 a119213a <=( A269  and  (not A268) );
 a119214a <=( a119213a  and  a119210a );
 a119217a <=( A299  and  A298 );
 a119220a <=( (not A301)  and  (not A300) );
 a119221a <=( a119220a  and  a119217a );
 a119222a <=( a119221a  and  a119214a );
 a119225a <=( A168  and  A170 );
 a119228a <=( A166  and  (not A167) );
 a119229a <=( a119228a  and  a119225a );
 a119232a <=( A200  and  (not A199) );
 a119235a <=( A203  and  (not A202) );
 a119236a <=( a119235a  and  a119232a );
 a119237a <=( a119236a  and  a119229a );
 a119240a <=( A266  and  (not A265) );
 a119243a <=( A269  and  (not A268) );
 a119244a <=( a119243a  and  a119240a );
 a119247a <=( A299  and  A298 );
 a119250a <=( A302  and  (not A300) );
 a119251a <=( a119250a  and  a119247a );
 a119252a <=( a119251a  and  a119244a );
 a119255a <=( A168  and  A170 );
 a119258a <=( A166  and  (not A167) );
 a119259a <=( a119258a  and  a119255a );
 a119262a <=( A200  and  (not A199) );
 a119265a <=( A203  and  (not A202) );
 a119266a <=( a119265a  and  a119262a );
 a119267a <=( a119266a  and  a119259a );
 a119270a <=( A266  and  (not A265) );
 a119273a <=( A269  and  (not A268) );
 a119274a <=( a119273a  and  a119270a );
 a119277a <=( (not A299)  and  A298 );
 a119280a <=( A301  and  (not A300) );
 a119281a <=( a119280a  and  a119277a );
 a119282a <=( a119281a  and  a119274a );
 a119285a <=( A168  and  A170 );
 a119288a <=( A166  and  (not A167) );
 a119289a <=( a119288a  and  a119285a );
 a119292a <=( A200  and  (not A199) );
 a119295a <=( A203  and  (not A202) );
 a119296a <=( a119295a  and  a119292a );
 a119297a <=( a119296a  and  a119289a );
 a119300a <=( A266  and  (not A265) );
 a119303a <=( A269  and  (not A268) );
 a119304a <=( a119303a  and  a119300a );
 a119307a <=( (not A299)  and  A298 );
 a119310a <=( (not A302)  and  (not A300) );
 a119311a <=( a119310a  and  a119307a );
 a119312a <=( a119311a  and  a119304a );
 a119315a <=( A168  and  A170 );
 a119318a <=( A166  and  (not A167) );
 a119319a <=( a119318a  and  a119315a );
 a119322a <=( A200  and  (not A199) );
 a119325a <=( A203  and  (not A202) );
 a119326a <=( a119325a  and  a119322a );
 a119327a <=( a119326a  and  a119319a );
 a119330a <=( A266  and  (not A265) );
 a119333a <=( A269  and  (not A268) );
 a119334a <=( a119333a  and  a119330a );
 a119337a <=( A299  and  (not A298) );
 a119340a <=( A301  and  (not A300) );
 a119341a <=( a119340a  and  a119337a );
 a119342a <=( a119341a  and  a119334a );
 a119345a <=( A168  and  A170 );
 a119348a <=( A166  and  (not A167) );
 a119349a <=( a119348a  and  a119345a );
 a119352a <=( A200  and  (not A199) );
 a119355a <=( A203  and  (not A202) );
 a119356a <=( a119355a  and  a119352a );
 a119357a <=( a119356a  and  a119349a );
 a119360a <=( A266  and  (not A265) );
 a119363a <=( A269  and  (not A268) );
 a119364a <=( a119363a  and  a119360a );
 a119367a <=( A299  and  (not A298) );
 a119370a <=( (not A302)  and  (not A300) );
 a119371a <=( a119370a  and  a119367a );
 a119372a <=( a119371a  and  a119364a );
 a119375a <=( A168  and  A170 );
 a119378a <=( A166  and  (not A167) );
 a119379a <=( a119378a  and  a119375a );
 a119382a <=( A200  and  (not A199) );
 a119385a <=( A203  and  (not A202) );
 a119386a <=( a119385a  and  a119382a );
 a119387a <=( a119386a  and  a119379a );
 a119390a <=( (not A266)  and  A265 );
 a119393a <=( A269  and  (not A268) );
 a119394a <=( a119393a  and  a119390a );
 a119397a <=( A299  and  A298 );
 a119400a <=( (not A301)  and  (not A300) );
 a119401a <=( a119400a  and  a119397a );
 a119402a <=( a119401a  and  a119394a );
 a119405a <=( A168  and  A170 );
 a119408a <=( A166  and  (not A167) );
 a119409a <=( a119408a  and  a119405a );
 a119412a <=( A200  and  (not A199) );
 a119415a <=( A203  and  (not A202) );
 a119416a <=( a119415a  and  a119412a );
 a119417a <=( a119416a  and  a119409a );
 a119420a <=( (not A266)  and  A265 );
 a119423a <=( A269  and  (not A268) );
 a119424a <=( a119423a  and  a119420a );
 a119427a <=( A299  and  A298 );
 a119430a <=( A302  and  (not A300) );
 a119431a <=( a119430a  and  a119427a );
 a119432a <=( a119431a  and  a119424a );
 a119435a <=( A168  and  A170 );
 a119438a <=( A166  and  (not A167) );
 a119439a <=( a119438a  and  a119435a );
 a119442a <=( A200  and  (not A199) );
 a119445a <=( A203  and  (not A202) );
 a119446a <=( a119445a  and  a119442a );
 a119447a <=( a119446a  and  a119439a );
 a119450a <=( (not A266)  and  A265 );
 a119453a <=( A269  and  (not A268) );
 a119454a <=( a119453a  and  a119450a );
 a119457a <=( (not A299)  and  A298 );
 a119460a <=( A301  and  (not A300) );
 a119461a <=( a119460a  and  a119457a );
 a119462a <=( a119461a  and  a119454a );
 a119465a <=( A168  and  A170 );
 a119468a <=( A166  and  (not A167) );
 a119469a <=( a119468a  and  a119465a );
 a119472a <=( A200  and  (not A199) );
 a119475a <=( A203  and  (not A202) );
 a119476a <=( a119475a  and  a119472a );
 a119477a <=( a119476a  and  a119469a );
 a119480a <=( (not A266)  and  A265 );
 a119483a <=( A269  and  (not A268) );
 a119484a <=( a119483a  and  a119480a );
 a119487a <=( (not A299)  and  A298 );
 a119490a <=( (not A302)  and  (not A300) );
 a119491a <=( a119490a  and  a119487a );
 a119492a <=( a119491a  and  a119484a );
 a119495a <=( A168  and  A170 );
 a119498a <=( A166  and  (not A167) );
 a119499a <=( a119498a  and  a119495a );
 a119502a <=( A200  and  (not A199) );
 a119505a <=( A203  and  (not A202) );
 a119506a <=( a119505a  and  a119502a );
 a119507a <=( a119506a  and  a119499a );
 a119510a <=( (not A266)  and  A265 );
 a119513a <=( A269  and  (not A268) );
 a119514a <=( a119513a  and  a119510a );
 a119517a <=( A299  and  (not A298) );
 a119520a <=( A301  and  (not A300) );
 a119521a <=( a119520a  and  a119517a );
 a119522a <=( a119521a  and  a119514a );
 a119525a <=( A168  and  A170 );
 a119528a <=( A166  and  (not A167) );
 a119529a <=( a119528a  and  a119525a );
 a119532a <=( A200  and  (not A199) );
 a119535a <=( A203  and  (not A202) );
 a119536a <=( a119535a  and  a119532a );
 a119537a <=( a119536a  and  a119529a );
 a119540a <=( (not A266)  and  A265 );
 a119543a <=( A269  and  (not A268) );
 a119544a <=( a119543a  and  a119540a );
 a119547a <=( A299  and  (not A298) );
 a119550a <=( (not A302)  and  (not A300) );
 a119551a <=( a119550a  and  a119547a );
 a119552a <=( a119551a  and  a119544a );
 a119555a <=( A168  and  A170 );
 a119558a <=( A166  and  (not A167) );
 a119559a <=( a119558a  and  a119555a );
 a119562a <=( A200  and  (not A199) );
 a119565a <=( A203  and  (not A202) );
 a119566a <=( a119565a  and  a119562a );
 a119567a <=( a119566a  and  a119559a );
 a119570a <=( (not A266)  and  (not A265) );
 a119573a <=( (not A269)  and  A268 );
 a119574a <=( a119573a  and  a119570a );
 a119577a <=( A299  and  A298 );
 a119580a <=( (not A301)  and  (not A300) );
 a119581a <=( a119580a  and  a119577a );
 a119582a <=( a119581a  and  a119574a );
 a119585a <=( A168  and  A170 );
 a119588a <=( A166  and  (not A167) );
 a119589a <=( a119588a  and  a119585a );
 a119592a <=( A200  and  (not A199) );
 a119595a <=( A203  and  (not A202) );
 a119596a <=( a119595a  and  a119592a );
 a119597a <=( a119596a  and  a119589a );
 a119600a <=( (not A266)  and  (not A265) );
 a119603a <=( (not A269)  and  A268 );
 a119604a <=( a119603a  and  a119600a );
 a119607a <=( A299  and  A298 );
 a119610a <=( A302  and  (not A300) );
 a119611a <=( a119610a  and  a119607a );
 a119612a <=( a119611a  and  a119604a );
 a119615a <=( A168  and  A170 );
 a119618a <=( A166  and  (not A167) );
 a119619a <=( a119618a  and  a119615a );
 a119622a <=( A200  and  (not A199) );
 a119625a <=( A203  and  (not A202) );
 a119626a <=( a119625a  and  a119622a );
 a119627a <=( a119626a  and  a119619a );
 a119630a <=( (not A266)  and  (not A265) );
 a119633a <=( (not A269)  and  A268 );
 a119634a <=( a119633a  and  a119630a );
 a119637a <=( (not A299)  and  A298 );
 a119640a <=( A301  and  (not A300) );
 a119641a <=( a119640a  and  a119637a );
 a119642a <=( a119641a  and  a119634a );
 a119645a <=( A168  and  A170 );
 a119648a <=( A166  and  (not A167) );
 a119649a <=( a119648a  and  a119645a );
 a119652a <=( A200  and  (not A199) );
 a119655a <=( A203  and  (not A202) );
 a119656a <=( a119655a  and  a119652a );
 a119657a <=( a119656a  and  a119649a );
 a119660a <=( (not A266)  and  (not A265) );
 a119663a <=( (not A269)  and  A268 );
 a119664a <=( a119663a  and  a119660a );
 a119667a <=( (not A299)  and  A298 );
 a119670a <=( (not A302)  and  (not A300) );
 a119671a <=( a119670a  and  a119667a );
 a119672a <=( a119671a  and  a119664a );
 a119675a <=( A168  and  A170 );
 a119678a <=( A166  and  (not A167) );
 a119679a <=( a119678a  and  a119675a );
 a119682a <=( A200  and  (not A199) );
 a119685a <=( A203  and  (not A202) );
 a119686a <=( a119685a  and  a119682a );
 a119687a <=( a119686a  and  a119679a );
 a119690a <=( (not A266)  and  (not A265) );
 a119693a <=( (not A269)  and  A268 );
 a119694a <=( a119693a  and  a119690a );
 a119697a <=( A299  and  (not A298) );
 a119700a <=( A301  and  (not A300) );
 a119701a <=( a119700a  and  a119697a );
 a119702a <=( a119701a  and  a119694a );
 a119705a <=( A168  and  A170 );
 a119708a <=( A166  and  (not A167) );
 a119709a <=( a119708a  and  a119705a );
 a119712a <=( A200  and  (not A199) );
 a119715a <=( A203  and  (not A202) );
 a119716a <=( a119715a  and  a119712a );
 a119717a <=( a119716a  and  a119709a );
 a119720a <=( (not A266)  and  (not A265) );
 a119723a <=( (not A269)  and  A268 );
 a119724a <=( a119723a  and  a119720a );
 a119727a <=( A299  and  (not A298) );
 a119730a <=( (not A302)  and  (not A300) );
 a119731a <=( a119730a  and  a119727a );
 a119732a <=( a119731a  and  a119724a );
 a119735a <=( A168  and  A170 );
 a119738a <=( A166  and  (not A167) );
 a119739a <=( a119738a  and  a119735a );
 a119742a <=( A200  and  (not A199) );
 a119745a <=( A202  and  (not A201) );
 a119746a <=( a119745a  and  a119742a );
 a119747a <=( a119746a  and  a119739a );
 a119750a <=( A266  and  A265 );
 a119753a <=( (not A268)  and  (not A267) );
 a119754a <=( a119753a  and  a119750a );
 a119757a <=( A299  and  A298 );
 a119760a <=( (not A302)  and  A301 );
 a119761a <=( a119760a  and  a119757a );
 a119762a <=( a119761a  and  a119754a );
 a119765a <=( A168  and  A170 );
 a119768a <=( A166  and  (not A167) );
 a119769a <=( a119768a  and  a119765a );
 a119772a <=( A200  and  (not A199) );
 a119775a <=( A202  and  (not A201) );
 a119776a <=( a119775a  and  a119772a );
 a119777a <=( a119776a  and  a119769a );
 a119780a <=( A266  and  A265 );
 a119783a <=( (not A268)  and  (not A267) );
 a119784a <=( a119783a  and  a119780a );
 a119787a <=( (not A299)  and  A298 );
 a119790a <=( A302  and  (not A301) );
 a119791a <=( a119790a  and  a119787a );
 a119792a <=( a119791a  and  a119784a );
 a119795a <=( A168  and  A170 );
 a119798a <=( A166  and  (not A167) );
 a119799a <=( a119798a  and  a119795a );
 a119802a <=( A200  and  (not A199) );
 a119805a <=( A202  and  (not A201) );
 a119806a <=( a119805a  and  a119802a );
 a119807a <=( a119806a  and  a119799a );
 a119810a <=( A266  and  A265 );
 a119813a <=( (not A268)  and  (not A267) );
 a119814a <=( a119813a  and  a119810a );
 a119817a <=( A299  and  (not A298) );
 a119820a <=( A302  and  (not A301) );
 a119821a <=( a119820a  and  a119817a );
 a119822a <=( a119821a  and  a119814a );
 a119825a <=( A168  and  A170 );
 a119828a <=( A166  and  (not A167) );
 a119829a <=( a119828a  and  a119825a );
 a119832a <=( A200  and  (not A199) );
 a119835a <=( A202  and  (not A201) );
 a119836a <=( a119835a  and  a119832a );
 a119837a <=( a119836a  and  a119829a );
 a119840a <=( A266  and  A265 );
 a119843a <=( (not A268)  and  (not A267) );
 a119844a <=( a119843a  and  a119840a );
 a119847a <=( (not A299)  and  (not A298) );
 a119850a <=( (not A302)  and  A301 );
 a119851a <=( a119850a  and  a119847a );
 a119852a <=( a119851a  and  a119844a );
 a119855a <=( A168  and  A170 );
 a119858a <=( A166  and  (not A167) );
 a119859a <=( a119858a  and  a119855a );
 a119862a <=( A200  and  (not A199) );
 a119865a <=( A202  and  (not A201) );
 a119866a <=( a119865a  and  a119862a );
 a119867a <=( a119866a  and  a119859a );
 a119870a <=( A266  and  A265 );
 a119873a <=( A269  and  (not A267) );
 a119874a <=( a119873a  and  a119870a );
 a119877a <=( A299  and  A298 );
 a119880a <=( (not A302)  and  A301 );
 a119881a <=( a119880a  and  a119877a );
 a119882a <=( a119881a  and  a119874a );
 a119885a <=( A168  and  A170 );
 a119888a <=( A166  and  (not A167) );
 a119889a <=( a119888a  and  a119885a );
 a119892a <=( A200  and  (not A199) );
 a119895a <=( A202  and  (not A201) );
 a119896a <=( a119895a  and  a119892a );
 a119897a <=( a119896a  and  a119889a );
 a119900a <=( A266  and  A265 );
 a119903a <=( A269  and  (not A267) );
 a119904a <=( a119903a  and  a119900a );
 a119907a <=( (not A299)  and  A298 );
 a119910a <=( A302  and  (not A301) );
 a119911a <=( a119910a  and  a119907a );
 a119912a <=( a119911a  and  a119904a );
 a119915a <=( A168  and  A170 );
 a119918a <=( A166  and  (not A167) );
 a119919a <=( a119918a  and  a119915a );
 a119922a <=( A200  and  (not A199) );
 a119925a <=( A202  and  (not A201) );
 a119926a <=( a119925a  and  a119922a );
 a119927a <=( a119926a  and  a119919a );
 a119930a <=( A266  and  A265 );
 a119933a <=( A269  and  (not A267) );
 a119934a <=( a119933a  and  a119930a );
 a119937a <=( A299  and  (not A298) );
 a119940a <=( A302  and  (not A301) );
 a119941a <=( a119940a  and  a119937a );
 a119942a <=( a119941a  and  a119934a );
 a119945a <=( A168  and  A170 );
 a119948a <=( A166  and  (not A167) );
 a119949a <=( a119948a  and  a119945a );
 a119952a <=( A200  and  (not A199) );
 a119955a <=( A202  and  (not A201) );
 a119956a <=( a119955a  and  a119952a );
 a119957a <=( a119956a  and  a119949a );
 a119960a <=( A266  and  A265 );
 a119963a <=( A269  and  (not A267) );
 a119964a <=( a119963a  and  a119960a );
 a119967a <=( (not A299)  and  (not A298) );
 a119970a <=( (not A302)  and  A301 );
 a119971a <=( a119970a  and  a119967a );
 a119972a <=( a119971a  and  a119964a );
 a119975a <=( A168  and  A170 );
 a119978a <=( A166  and  (not A167) );
 a119979a <=( a119978a  and  a119975a );
 a119982a <=( A200  and  (not A199) );
 a119985a <=( A202  and  (not A201) );
 a119986a <=( a119985a  and  a119982a );
 a119987a <=( a119986a  and  a119979a );
 a119990a <=( A266  and  (not A265) );
 a119993a <=( A268  and  (not A267) );
 a119994a <=( a119993a  and  a119990a );
 a119997a <=( A299  and  A298 );
 a120000a <=( (not A302)  and  A301 );
 a120001a <=( a120000a  and  a119997a );
 a120002a <=( a120001a  and  a119994a );
 a120005a <=( A168  and  A170 );
 a120008a <=( A166  and  (not A167) );
 a120009a <=( a120008a  and  a120005a );
 a120012a <=( A200  and  (not A199) );
 a120015a <=( A202  and  (not A201) );
 a120016a <=( a120015a  and  a120012a );
 a120017a <=( a120016a  and  a120009a );
 a120020a <=( A266  and  (not A265) );
 a120023a <=( A268  and  (not A267) );
 a120024a <=( a120023a  and  a120020a );
 a120027a <=( (not A299)  and  A298 );
 a120030a <=( A302  and  (not A301) );
 a120031a <=( a120030a  and  a120027a );
 a120032a <=( a120031a  and  a120024a );
 a120035a <=( A168  and  A170 );
 a120038a <=( A166  and  (not A167) );
 a120039a <=( a120038a  and  a120035a );
 a120042a <=( A200  and  (not A199) );
 a120045a <=( A202  and  (not A201) );
 a120046a <=( a120045a  and  a120042a );
 a120047a <=( a120046a  and  a120039a );
 a120050a <=( A266  and  (not A265) );
 a120053a <=( A268  and  (not A267) );
 a120054a <=( a120053a  and  a120050a );
 a120057a <=( A299  and  (not A298) );
 a120060a <=( A302  and  (not A301) );
 a120061a <=( a120060a  and  a120057a );
 a120062a <=( a120061a  and  a120054a );
 a120065a <=( A168  and  A170 );
 a120068a <=( A166  and  (not A167) );
 a120069a <=( a120068a  and  a120065a );
 a120072a <=( A200  and  (not A199) );
 a120075a <=( A202  and  (not A201) );
 a120076a <=( a120075a  and  a120072a );
 a120077a <=( a120076a  and  a120069a );
 a120080a <=( A266  and  (not A265) );
 a120083a <=( A268  and  (not A267) );
 a120084a <=( a120083a  and  a120080a );
 a120087a <=( (not A299)  and  (not A298) );
 a120090a <=( (not A302)  and  A301 );
 a120091a <=( a120090a  and  a120087a );
 a120092a <=( a120091a  and  a120084a );
 a120095a <=( A168  and  A170 );
 a120098a <=( A166  and  (not A167) );
 a120099a <=( a120098a  and  a120095a );
 a120102a <=( A200  and  (not A199) );
 a120105a <=( A202  and  (not A201) );
 a120106a <=( a120105a  and  a120102a );
 a120107a <=( a120106a  and  a120099a );
 a120110a <=( A266  and  (not A265) );
 a120113a <=( (not A269)  and  (not A267) );
 a120114a <=( a120113a  and  a120110a );
 a120117a <=( A299  and  A298 );
 a120120a <=( (not A302)  and  A301 );
 a120121a <=( a120120a  and  a120117a );
 a120122a <=( a120121a  and  a120114a );
 a120125a <=( A168  and  A170 );
 a120128a <=( A166  and  (not A167) );
 a120129a <=( a120128a  and  a120125a );
 a120132a <=( A200  and  (not A199) );
 a120135a <=( A202  and  (not A201) );
 a120136a <=( a120135a  and  a120132a );
 a120137a <=( a120136a  and  a120129a );
 a120140a <=( A266  and  (not A265) );
 a120143a <=( (not A269)  and  (not A267) );
 a120144a <=( a120143a  and  a120140a );
 a120147a <=( (not A299)  and  A298 );
 a120150a <=( A302  and  (not A301) );
 a120151a <=( a120150a  and  a120147a );
 a120152a <=( a120151a  and  a120144a );
 a120155a <=( A168  and  A170 );
 a120158a <=( A166  and  (not A167) );
 a120159a <=( a120158a  and  a120155a );
 a120162a <=( A200  and  (not A199) );
 a120165a <=( A202  and  (not A201) );
 a120166a <=( a120165a  and  a120162a );
 a120167a <=( a120166a  and  a120159a );
 a120170a <=( A266  and  (not A265) );
 a120173a <=( (not A269)  and  (not A267) );
 a120174a <=( a120173a  and  a120170a );
 a120177a <=( A299  and  (not A298) );
 a120180a <=( A302  and  (not A301) );
 a120181a <=( a120180a  and  a120177a );
 a120182a <=( a120181a  and  a120174a );
 a120185a <=( A168  and  A170 );
 a120188a <=( A166  and  (not A167) );
 a120189a <=( a120188a  and  a120185a );
 a120192a <=( A200  and  (not A199) );
 a120195a <=( A202  and  (not A201) );
 a120196a <=( a120195a  and  a120192a );
 a120197a <=( a120196a  and  a120189a );
 a120200a <=( A266  and  (not A265) );
 a120203a <=( (not A269)  and  (not A267) );
 a120204a <=( a120203a  and  a120200a );
 a120207a <=( (not A299)  and  (not A298) );
 a120210a <=( (not A302)  and  A301 );
 a120211a <=( a120210a  and  a120207a );
 a120212a <=( a120211a  and  a120204a );
 a120215a <=( A168  and  A170 );
 a120218a <=( A166  and  (not A167) );
 a120219a <=( a120218a  and  a120215a );
 a120222a <=( A200  and  (not A199) );
 a120225a <=( A202  and  (not A201) );
 a120226a <=( a120225a  and  a120222a );
 a120227a <=( a120226a  and  a120219a );
 a120230a <=( (not A266)  and  A265 );
 a120233a <=( A268  and  (not A267) );
 a120234a <=( a120233a  and  a120230a );
 a120237a <=( A299  and  A298 );
 a120240a <=( (not A302)  and  A301 );
 a120241a <=( a120240a  and  a120237a );
 a120242a <=( a120241a  and  a120234a );
 a120245a <=( A168  and  A170 );
 a120248a <=( A166  and  (not A167) );
 a120249a <=( a120248a  and  a120245a );
 a120252a <=( A200  and  (not A199) );
 a120255a <=( A202  and  (not A201) );
 a120256a <=( a120255a  and  a120252a );
 a120257a <=( a120256a  and  a120249a );
 a120260a <=( (not A266)  and  A265 );
 a120263a <=( A268  and  (not A267) );
 a120264a <=( a120263a  and  a120260a );
 a120267a <=( (not A299)  and  A298 );
 a120270a <=( A302  and  (not A301) );
 a120271a <=( a120270a  and  a120267a );
 a120272a <=( a120271a  and  a120264a );
 a120275a <=( A168  and  A170 );
 a120278a <=( A166  and  (not A167) );
 a120279a <=( a120278a  and  a120275a );
 a120282a <=( A200  and  (not A199) );
 a120285a <=( A202  and  (not A201) );
 a120286a <=( a120285a  and  a120282a );
 a120287a <=( a120286a  and  a120279a );
 a120290a <=( (not A266)  and  A265 );
 a120293a <=( A268  and  (not A267) );
 a120294a <=( a120293a  and  a120290a );
 a120297a <=( A299  and  (not A298) );
 a120300a <=( A302  and  (not A301) );
 a120301a <=( a120300a  and  a120297a );
 a120302a <=( a120301a  and  a120294a );
 a120305a <=( A168  and  A170 );
 a120308a <=( A166  and  (not A167) );
 a120309a <=( a120308a  and  a120305a );
 a120312a <=( A200  and  (not A199) );
 a120315a <=( A202  and  (not A201) );
 a120316a <=( a120315a  and  a120312a );
 a120317a <=( a120316a  and  a120309a );
 a120320a <=( (not A266)  and  A265 );
 a120323a <=( A268  and  (not A267) );
 a120324a <=( a120323a  and  a120320a );
 a120327a <=( (not A299)  and  (not A298) );
 a120330a <=( (not A302)  and  A301 );
 a120331a <=( a120330a  and  a120327a );
 a120332a <=( a120331a  and  a120324a );
 a120335a <=( A168  and  A170 );
 a120338a <=( A166  and  (not A167) );
 a120339a <=( a120338a  and  a120335a );
 a120342a <=( A200  and  (not A199) );
 a120345a <=( A202  and  (not A201) );
 a120346a <=( a120345a  and  a120342a );
 a120347a <=( a120346a  and  a120339a );
 a120350a <=( (not A266)  and  A265 );
 a120353a <=( (not A269)  and  (not A267) );
 a120354a <=( a120353a  and  a120350a );
 a120357a <=( A299  and  A298 );
 a120360a <=( (not A302)  and  A301 );
 a120361a <=( a120360a  and  a120357a );
 a120362a <=( a120361a  and  a120354a );
 a120365a <=( A168  and  A170 );
 a120368a <=( A166  and  (not A167) );
 a120369a <=( a120368a  and  a120365a );
 a120372a <=( A200  and  (not A199) );
 a120375a <=( A202  and  (not A201) );
 a120376a <=( a120375a  and  a120372a );
 a120377a <=( a120376a  and  a120369a );
 a120380a <=( (not A266)  and  A265 );
 a120383a <=( (not A269)  and  (not A267) );
 a120384a <=( a120383a  and  a120380a );
 a120387a <=( (not A299)  and  A298 );
 a120390a <=( A302  and  (not A301) );
 a120391a <=( a120390a  and  a120387a );
 a120392a <=( a120391a  and  a120384a );
 a120395a <=( A168  and  A170 );
 a120398a <=( A166  and  (not A167) );
 a120399a <=( a120398a  and  a120395a );
 a120402a <=( A200  and  (not A199) );
 a120405a <=( A202  and  (not A201) );
 a120406a <=( a120405a  and  a120402a );
 a120407a <=( a120406a  and  a120399a );
 a120410a <=( (not A266)  and  A265 );
 a120413a <=( (not A269)  and  (not A267) );
 a120414a <=( a120413a  and  a120410a );
 a120417a <=( A299  and  (not A298) );
 a120420a <=( A302  and  (not A301) );
 a120421a <=( a120420a  and  a120417a );
 a120422a <=( a120421a  and  a120414a );
 a120425a <=( A168  and  A170 );
 a120428a <=( A166  and  (not A167) );
 a120429a <=( a120428a  and  a120425a );
 a120432a <=( A200  and  (not A199) );
 a120435a <=( A202  and  (not A201) );
 a120436a <=( a120435a  and  a120432a );
 a120437a <=( a120436a  and  a120429a );
 a120440a <=( (not A266)  and  A265 );
 a120443a <=( (not A269)  and  (not A267) );
 a120444a <=( a120443a  and  a120440a );
 a120447a <=( (not A299)  and  (not A298) );
 a120450a <=( (not A302)  and  A301 );
 a120451a <=( a120450a  and  a120447a );
 a120452a <=( a120451a  and  a120444a );
 a120455a <=( A168  and  A170 );
 a120458a <=( A166  and  (not A167) );
 a120459a <=( a120458a  and  a120455a );
 a120462a <=( A200  and  (not A199) );
 a120465a <=( (not A203)  and  (not A201) );
 a120466a <=( a120465a  and  a120462a );
 a120467a <=( a120466a  and  a120459a );
 a120470a <=( A266  and  A265 );
 a120473a <=( (not A268)  and  (not A267) );
 a120474a <=( a120473a  and  a120470a );
 a120477a <=( A299  and  A298 );
 a120480a <=( (not A302)  and  A301 );
 a120481a <=( a120480a  and  a120477a );
 a120482a <=( a120481a  and  a120474a );
 a120485a <=( A168  and  A170 );
 a120488a <=( A166  and  (not A167) );
 a120489a <=( a120488a  and  a120485a );
 a120492a <=( A200  and  (not A199) );
 a120495a <=( (not A203)  and  (not A201) );
 a120496a <=( a120495a  and  a120492a );
 a120497a <=( a120496a  and  a120489a );
 a120500a <=( A266  and  A265 );
 a120503a <=( (not A268)  and  (not A267) );
 a120504a <=( a120503a  and  a120500a );
 a120507a <=( (not A299)  and  A298 );
 a120510a <=( A302  and  (not A301) );
 a120511a <=( a120510a  and  a120507a );
 a120512a <=( a120511a  and  a120504a );
 a120515a <=( A168  and  A170 );
 a120518a <=( A166  and  (not A167) );
 a120519a <=( a120518a  and  a120515a );
 a120522a <=( A200  and  (not A199) );
 a120525a <=( (not A203)  and  (not A201) );
 a120526a <=( a120525a  and  a120522a );
 a120527a <=( a120526a  and  a120519a );
 a120530a <=( A266  and  A265 );
 a120533a <=( (not A268)  and  (not A267) );
 a120534a <=( a120533a  and  a120530a );
 a120537a <=( A299  and  (not A298) );
 a120540a <=( A302  and  (not A301) );
 a120541a <=( a120540a  and  a120537a );
 a120542a <=( a120541a  and  a120534a );
 a120545a <=( A168  and  A170 );
 a120548a <=( A166  and  (not A167) );
 a120549a <=( a120548a  and  a120545a );
 a120552a <=( A200  and  (not A199) );
 a120555a <=( (not A203)  and  (not A201) );
 a120556a <=( a120555a  and  a120552a );
 a120557a <=( a120556a  and  a120549a );
 a120560a <=( A266  and  A265 );
 a120563a <=( (not A268)  and  (not A267) );
 a120564a <=( a120563a  and  a120560a );
 a120567a <=( (not A299)  and  (not A298) );
 a120570a <=( (not A302)  and  A301 );
 a120571a <=( a120570a  and  a120567a );
 a120572a <=( a120571a  and  a120564a );
 a120575a <=( A168  and  A170 );
 a120578a <=( A166  and  (not A167) );
 a120579a <=( a120578a  and  a120575a );
 a120582a <=( A200  and  (not A199) );
 a120585a <=( (not A203)  and  (not A201) );
 a120586a <=( a120585a  and  a120582a );
 a120587a <=( a120586a  and  a120579a );
 a120590a <=( A266  and  A265 );
 a120593a <=( A269  and  (not A267) );
 a120594a <=( a120593a  and  a120590a );
 a120597a <=( A299  and  A298 );
 a120600a <=( (not A302)  and  A301 );
 a120601a <=( a120600a  and  a120597a );
 a120602a <=( a120601a  and  a120594a );
 a120605a <=( A168  and  A170 );
 a120608a <=( A166  and  (not A167) );
 a120609a <=( a120608a  and  a120605a );
 a120612a <=( A200  and  (not A199) );
 a120615a <=( (not A203)  and  (not A201) );
 a120616a <=( a120615a  and  a120612a );
 a120617a <=( a120616a  and  a120609a );
 a120620a <=( A266  and  A265 );
 a120623a <=( A269  and  (not A267) );
 a120624a <=( a120623a  and  a120620a );
 a120627a <=( (not A299)  and  A298 );
 a120630a <=( A302  and  (not A301) );
 a120631a <=( a120630a  and  a120627a );
 a120632a <=( a120631a  and  a120624a );
 a120635a <=( A168  and  A170 );
 a120638a <=( A166  and  (not A167) );
 a120639a <=( a120638a  and  a120635a );
 a120642a <=( A200  and  (not A199) );
 a120645a <=( (not A203)  and  (not A201) );
 a120646a <=( a120645a  and  a120642a );
 a120647a <=( a120646a  and  a120639a );
 a120650a <=( A266  and  A265 );
 a120653a <=( A269  and  (not A267) );
 a120654a <=( a120653a  and  a120650a );
 a120657a <=( A299  and  (not A298) );
 a120660a <=( A302  and  (not A301) );
 a120661a <=( a120660a  and  a120657a );
 a120662a <=( a120661a  and  a120654a );
 a120665a <=( A168  and  A170 );
 a120668a <=( A166  and  (not A167) );
 a120669a <=( a120668a  and  a120665a );
 a120672a <=( A200  and  (not A199) );
 a120675a <=( (not A203)  and  (not A201) );
 a120676a <=( a120675a  and  a120672a );
 a120677a <=( a120676a  and  a120669a );
 a120680a <=( A266  and  A265 );
 a120683a <=( A269  and  (not A267) );
 a120684a <=( a120683a  and  a120680a );
 a120687a <=( (not A299)  and  (not A298) );
 a120690a <=( (not A302)  and  A301 );
 a120691a <=( a120690a  and  a120687a );
 a120692a <=( a120691a  and  a120684a );
 a120695a <=( A168  and  A170 );
 a120698a <=( A166  and  (not A167) );
 a120699a <=( a120698a  and  a120695a );
 a120702a <=( A200  and  (not A199) );
 a120705a <=( (not A203)  and  (not A201) );
 a120706a <=( a120705a  and  a120702a );
 a120707a <=( a120706a  and  a120699a );
 a120710a <=( A266  and  (not A265) );
 a120713a <=( A268  and  (not A267) );
 a120714a <=( a120713a  and  a120710a );
 a120717a <=( A299  and  A298 );
 a120720a <=( (not A302)  and  A301 );
 a120721a <=( a120720a  and  a120717a );
 a120722a <=( a120721a  and  a120714a );
 a120725a <=( A168  and  A170 );
 a120728a <=( A166  and  (not A167) );
 a120729a <=( a120728a  and  a120725a );
 a120732a <=( A200  and  (not A199) );
 a120735a <=( (not A203)  and  (not A201) );
 a120736a <=( a120735a  and  a120732a );
 a120737a <=( a120736a  and  a120729a );
 a120740a <=( A266  and  (not A265) );
 a120743a <=( A268  and  (not A267) );
 a120744a <=( a120743a  and  a120740a );
 a120747a <=( (not A299)  and  A298 );
 a120750a <=( A302  and  (not A301) );
 a120751a <=( a120750a  and  a120747a );
 a120752a <=( a120751a  and  a120744a );
 a120755a <=( A168  and  A170 );
 a120758a <=( A166  and  (not A167) );
 a120759a <=( a120758a  and  a120755a );
 a120762a <=( A200  and  (not A199) );
 a120765a <=( (not A203)  and  (not A201) );
 a120766a <=( a120765a  and  a120762a );
 a120767a <=( a120766a  and  a120759a );
 a120770a <=( A266  and  (not A265) );
 a120773a <=( A268  and  (not A267) );
 a120774a <=( a120773a  and  a120770a );
 a120777a <=( A299  and  (not A298) );
 a120780a <=( A302  and  (not A301) );
 a120781a <=( a120780a  and  a120777a );
 a120782a <=( a120781a  and  a120774a );
 a120785a <=( A168  and  A170 );
 a120788a <=( A166  and  (not A167) );
 a120789a <=( a120788a  and  a120785a );
 a120792a <=( A200  and  (not A199) );
 a120795a <=( (not A203)  and  (not A201) );
 a120796a <=( a120795a  and  a120792a );
 a120797a <=( a120796a  and  a120789a );
 a120800a <=( A266  and  (not A265) );
 a120803a <=( A268  and  (not A267) );
 a120804a <=( a120803a  and  a120800a );
 a120807a <=( (not A299)  and  (not A298) );
 a120810a <=( (not A302)  and  A301 );
 a120811a <=( a120810a  and  a120807a );
 a120812a <=( a120811a  and  a120804a );
 a120815a <=( A168  and  A170 );
 a120818a <=( A166  and  (not A167) );
 a120819a <=( a120818a  and  a120815a );
 a120822a <=( A200  and  (not A199) );
 a120825a <=( (not A203)  and  (not A201) );
 a120826a <=( a120825a  and  a120822a );
 a120827a <=( a120826a  and  a120819a );
 a120830a <=( A266  and  (not A265) );
 a120833a <=( (not A269)  and  (not A267) );
 a120834a <=( a120833a  and  a120830a );
 a120837a <=( A299  and  A298 );
 a120840a <=( (not A302)  and  A301 );
 a120841a <=( a120840a  and  a120837a );
 a120842a <=( a120841a  and  a120834a );
 a120845a <=( A168  and  A170 );
 a120848a <=( A166  and  (not A167) );
 a120849a <=( a120848a  and  a120845a );
 a120852a <=( A200  and  (not A199) );
 a120855a <=( (not A203)  and  (not A201) );
 a120856a <=( a120855a  and  a120852a );
 a120857a <=( a120856a  and  a120849a );
 a120860a <=( A266  and  (not A265) );
 a120863a <=( (not A269)  and  (not A267) );
 a120864a <=( a120863a  and  a120860a );
 a120867a <=( (not A299)  and  A298 );
 a120870a <=( A302  and  (not A301) );
 a120871a <=( a120870a  and  a120867a );
 a120872a <=( a120871a  and  a120864a );
 a120875a <=( A168  and  A170 );
 a120878a <=( A166  and  (not A167) );
 a120879a <=( a120878a  and  a120875a );
 a120882a <=( A200  and  (not A199) );
 a120885a <=( (not A203)  and  (not A201) );
 a120886a <=( a120885a  and  a120882a );
 a120887a <=( a120886a  and  a120879a );
 a120890a <=( A266  and  (not A265) );
 a120893a <=( (not A269)  and  (not A267) );
 a120894a <=( a120893a  and  a120890a );
 a120897a <=( A299  and  (not A298) );
 a120900a <=( A302  and  (not A301) );
 a120901a <=( a120900a  and  a120897a );
 a120902a <=( a120901a  and  a120894a );
 a120905a <=( A168  and  A170 );
 a120908a <=( A166  and  (not A167) );
 a120909a <=( a120908a  and  a120905a );
 a120912a <=( A200  and  (not A199) );
 a120915a <=( (not A203)  and  (not A201) );
 a120916a <=( a120915a  and  a120912a );
 a120917a <=( a120916a  and  a120909a );
 a120920a <=( A266  and  (not A265) );
 a120923a <=( (not A269)  and  (not A267) );
 a120924a <=( a120923a  and  a120920a );
 a120927a <=( (not A299)  and  (not A298) );
 a120930a <=( (not A302)  and  A301 );
 a120931a <=( a120930a  and  a120927a );
 a120932a <=( a120931a  and  a120924a );
 a120935a <=( A168  and  A170 );
 a120938a <=( A166  and  (not A167) );
 a120939a <=( a120938a  and  a120935a );
 a120942a <=( A200  and  (not A199) );
 a120945a <=( (not A203)  and  (not A201) );
 a120946a <=( a120945a  and  a120942a );
 a120947a <=( a120946a  and  a120939a );
 a120950a <=( (not A266)  and  A265 );
 a120953a <=( A268  and  (not A267) );
 a120954a <=( a120953a  and  a120950a );
 a120957a <=( A299  and  A298 );
 a120960a <=( (not A302)  and  A301 );
 a120961a <=( a120960a  and  a120957a );
 a120962a <=( a120961a  and  a120954a );
 a120965a <=( A168  and  A170 );
 a120968a <=( A166  and  (not A167) );
 a120969a <=( a120968a  and  a120965a );
 a120972a <=( A200  and  (not A199) );
 a120975a <=( (not A203)  and  (not A201) );
 a120976a <=( a120975a  and  a120972a );
 a120977a <=( a120976a  and  a120969a );
 a120980a <=( (not A266)  and  A265 );
 a120983a <=( A268  and  (not A267) );
 a120984a <=( a120983a  and  a120980a );
 a120987a <=( (not A299)  and  A298 );
 a120990a <=( A302  and  (not A301) );
 a120991a <=( a120990a  and  a120987a );
 a120992a <=( a120991a  and  a120984a );
 a120995a <=( A168  and  A170 );
 a120998a <=( A166  and  (not A167) );
 a120999a <=( a120998a  and  a120995a );
 a121002a <=( A200  and  (not A199) );
 a121005a <=( (not A203)  and  (not A201) );
 a121006a <=( a121005a  and  a121002a );
 a121007a <=( a121006a  and  a120999a );
 a121010a <=( (not A266)  and  A265 );
 a121013a <=( A268  and  (not A267) );
 a121014a <=( a121013a  and  a121010a );
 a121017a <=( A299  and  (not A298) );
 a121020a <=( A302  and  (not A301) );
 a121021a <=( a121020a  and  a121017a );
 a121022a <=( a121021a  and  a121014a );
 a121025a <=( A168  and  A170 );
 a121028a <=( A166  and  (not A167) );
 a121029a <=( a121028a  and  a121025a );
 a121032a <=( A200  and  (not A199) );
 a121035a <=( (not A203)  and  (not A201) );
 a121036a <=( a121035a  and  a121032a );
 a121037a <=( a121036a  and  a121029a );
 a121040a <=( (not A266)  and  A265 );
 a121043a <=( A268  and  (not A267) );
 a121044a <=( a121043a  and  a121040a );
 a121047a <=( (not A299)  and  (not A298) );
 a121050a <=( (not A302)  and  A301 );
 a121051a <=( a121050a  and  a121047a );
 a121052a <=( a121051a  and  a121044a );
 a121055a <=( A168  and  A170 );
 a121058a <=( A166  and  (not A167) );
 a121059a <=( a121058a  and  a121055a );
 a121062a <=( A200  and  (not A199) );
 a121065a <=( (not A203)  and  (not A201) );
 a121066a <=( a121065a  and  a121062a );
 a121067a <=( a121066a  and  a121059a );
 a121070a <=( (not A266)  and  A265 );
 a121073a <=( (not A269)  and  (not A267) );
 a121074a <=( a121073a  and  a121070a );
 a121077a <=( A299  and  A298 );
 a121080a <=( (not A302)  and  A301 );
 a121081a <=( a121080a  and  a121077a );
 a121082a <=( a121081a  and  a121074a );
 a121085a <=( A168  and  A170 );
 a121088a <=( A166  and  (not A167) );
 a121089a <=( a121088a  and  a121085a );
 a121092a <=( A200  and  (not A199) );
 a121095a <=( (not A203)  and  (not A201) );
 a121096a <=( a121095a  and  a121092a );
 a121097a <=( a121096a  and  a121089a );
 a121100a <=( (not A266)  and  A265 );
 a121103a <=( (not A269)  and  (not A267) );
 a121104a <=( a121103a  and  a121100a );
 a121107a <=( (not A299)  and  A298 );
 a121110a <=( A302  and  (not A301) );
 a121111a <=( a121110a  and  a121107a );
 a121112a <=( a121111a  and  a121104a );
 a121115a <=( A168  and  A170 );
 a121118a <=( A166  and  (not A167) );
 a121119a <=( a121118a  and  a121115a );
 a121122a <=( A200  and  (not A199) );
 a121125a <=( (not A203)  and  (not A201) );
 a121126a <=( a121125a  and  a121122a );
 a121127a <=( a121126a  and  a121119a );
 a121130a <=( (not A266)  and  A265 );
 a121133a <=( (not A269)  and  (not A267) );
 a121134a <=( a121133a  and  a121130a );
 a121137a <=( A299  and  (not A298) );
 a121140a <=( A302  and  (not A301) );
 a121141a <=( a121140a  and  a121137a );
 a121142a <=( a121141a  and  a121134a );
 a121145a <=( A168  and  A170 );
 a121148a <=( A166  and  (not A167) );
 a121149a <=( a121148a  and  a121145a );
 a121152a <=( A200  and  (not A199) );
 a121155a <=( (not A203)  and  (not A201) );
 a121156a <=( a121155a  and  a121152a );
 a121157a <=( a121156a  and  a121149a );
 a121160a <=( (not A266)  and  A265 );
 a121163a <=( (not A269)  and  (not A267) );
 a121164a <=( a121163a  and  a121160a );
 a121167a <=( (not A299)  and  (not A298) );
 a121170a <=( (not A302)  and  A301 );
 a121171a <=( a121170a  and  a121167a );
 a121172a <=( a121171a  and  a121164a );
 a121175a <=( A168  and  A170 );
 a121178a <=( A166  and  (not A167) );
 a121179a <=( a121178a  and  a121175a );
 a121182a <=( (not A200)  and  A199 );
 a121185a <=( A203  and  (not A202) );
 a121186a <=( a121185a  and  a121182a );
 a121187a <=( a121186a  and  a121179a );
 a121190a <=( A266  and  A265 );
 a121193a <=( (not A269)  and  A268 );
 a121194a <=( a121193a  and  a121190a );
 a121197a <=( A299  and  A298 );
 a121200a <=( (not A301)  and  (not A300) );
 a121201a <=( a121200a  and  a121197a );
 a121202a <=( a121201a  and  a121194a );
 a121205a <=( A168  and  A170 );
 a121208a <=( A166  and  (not A167) );
 a121209a <=( a121208a  and  a121205a );
 a121212a <=( (not A200)  and  A199 );
 a121215a <=( A203  and  (not A202) );
 a121216a <=( a121215a  and  a121212a );
 a121217a <=( a121216a  and  a121209a );
 a121220a <=( A266  and  A265 );
 a121223a <=( (not A269)  and  A268 );
 a121224a <=( a121223a  and  a121220a );
 a121227a <=( A299  and  A298 );
 a121230a <=( A302  and  (not A300) );
 a121231a <=( a121230a  and  a121227a );
 a121232a <=( a121231a  and  a121224a );
 a121235a <=( A168  and  A170 );
 a121238a <=( A166  and  (not A167) );
 a121239a <=( a121238a  and  a121235a );
 a121242a <=( (not A200)  and  A199 );
 a121245a <=( A203  and  (not A202) );
 a121246a <=( a121245a  and  a121242a );
 a121247a <=( a121246a  and  a121239a );
 a121250a <=( A266  and  A265 );
 a121253a <=( (not A269)  and  A268 );
 a121254a <=( a121253a  and  a121250a );
 a121257a <=( (not A299)  and  A298 );
 a121260a <=( A301  and  (not A300) );
 a121261a <=( a121260a  and  a121257a );
 a121262a <=( a121261a  and  a121254a );
 a121265a <=( A168  and  A170 );
 a121268a <=( A166  and  (not A167) );
 a121269a <=( a121268a  and  a121265a );
 a121272a <=( (not A200)  and  A199 );
 a121275a <=( A203  and  (not A202) );
 a121276a <=( a121275a  and  a121272a );
 a121277a <=( a121276a  and  a121269a );
 a121280a <=( A266  and  A265 );
 a121283a <=( (not A269)  and  A268 );
 a121284a <=( a121283a  and  a121280a );
 a121287a <=( (not A299)  and  A298 );
 a121290a <=( (not A302)  and  (not A300) );
 a121291a <=( a121290a  and  a121287a );
 a121292a <=( a121291a  and  a121284a );
 a121295a <=( A168  and  A170 );
 a121298a <=( A166  and  (not A167) );
 a121299a <=( a121298a  and  a121295a );
 a121302a <=( (not A200)  and  A199 );
 a121305a <=( A203  and  (not A202) );
 a121306a <=( a121305a  and  a121302a );
 a121307a <=( a121306a  and  a121299a );
 a121310a <=( A266  and  A265 );
 a121313a <=( (not A269)  and  A268 );
 a121314a <=( a121313a  and  a121310a );
 a121317a <=( A299  and  (not A298) );
 a121320a <=( A301  and  (not A300) );
 a121321a <=( a121320a  and  a121317a );
 a121322a <=( a121321a  and  a121314a );
 a121325a <=( A168  and  A170 );
 a121328a <=( A166  and  (not A167) );
 a121329a <=( a121328a  and  a121325a );
 a121332a <=( (not A200)  and  A199 );
 a121335a <=( A203  and  (not A202) );
 a121336a <=( a121335a  and  a121332a );
 a121337a <=( a121336a  and  a121329a );
 a121340a <=( A266  and  A265 );
 a121343a <=( (not A269)  and  A268 );
 a121344a <=( a121343a  and  a121340a );
 a121347a <=( A299  and  (not A298) );
 a121350a <=( (not A302)  and  (not A300) );
 a121351a <=( a121350a  and  a121347a );
 a121352a <=( a121351a  and  a121344a );
 a121355a <=( A168  and  A170 );
 a121358a <=( A166  and  (not A167) );
 a121359a <=( a121358a  and  a121355a );
 a121362a <=( (not A200)  and  A199 );
 a121365a <=( A203  and  (not A202) );
 a121366a <=( a121365a  and  a121362a );
 a121367a <=( a121366a  and  a121359a );
 a121370a <=( A266  and  (not A265) );
 a121373a <=( A269  and  (not A268) );
 a121374a <=( a121373a  and  a121370a );
 a121377a <=( A299  and  A298 );
 a121380a <=( (not A301)  and  (not A300) );
 a121381a <=( a121380a  and  a121377a );
 a121382a <=( a121381a  and  a121374a );
 a121385a <=( A168  and  A170 );
 a121388a <=( A166  and  (not A167) );
 a121389a <=( a121388a  and  a121385a );
 a121392a <=( (not A200)  and  A199 );
 a121395a <=( A203  and  (not A202) );
 a121396a <=( a121395a  and  a121392a );
 a121397a <=( a121396a  and  a121389a );
 a121400a <=( A266  and  (not A265) );
 a121403a <=( A269  and  (not A268) );
 a121404a <=( a121403a  and  a121400a );
 a121407a <=( A299  and  A298 );
 a121410a <=( A302  and  (not A300) );
 a121411a <=( a121410a  and  a121407a );
 a121412a <=( a121411a  and  a121404a );
 a121415a <=( A168  and  A170 );
 a121418a <=( A166  and  (not A167) );
 a121419a <=( a121418a  and  a121415a );
 a121422a <=( (not A200)  and  A199 );
 a121425a <=( A203  and  (not A202) );
 a121426a <=( a121425a  and  a121422a );
 a121427a <=( a121426a  and  a121419a );
 a121430a <=( A266  and  (not A265) );
 a121433a <=( A269  and  (not A268) );
 a121434a <=( a121433a  and  a121430a );
 a121437a <=( (not A299)  and  A298 );
 a121440a <=( A301  and  (not A300) );
 a121441a <=( a121440a  and  a121437a );
 a121442a <=( a121441a  and  a121434a );
 a121445a <=( A168  and  A170 );
 a121448a <=( A166  and  (not A167) );
 a121449a <=( a121448a  and  a121445a );
 a121452a <=( (not A200)  and  A199 );
 a121455a <=( A203  and  (not A202) );
 a121456a <=( a121455a  and  a121452a );
 a121457a <=( a121456a  and  a121449a );
 a121460a <=( A266  and  (not A265) );
 a121463a <=( A269  and  (not A268) );
 a121464a <=( a121463a  and  a121460a );
 a121467a <=( (not A299)  and  A298 );
 a121470a <=( (not A302)  and  (not A300) );
 a121471a <=( a121470a  and  a121467a );
 a121472a <=( a121471a  and  a121464a );
 a121475a <=( A168  and  A170 );
 a121478a <=( A166  and  (not A167) );
 a121479a <=( a121478a  and  a121475a );
 a121482a <=( (not A200)  and  A199 );
 a121485a <=( A203  and  (not A202) );
 a121486a <=( a121485a  and  a121482a );
 a121487a <=( a121486a  and  a121479a );
 a121490a <=( A266  and  (not A265) );
 a121493a <=( A269  and  (not A268) );
 a121494a <=( a121493a  and  a121490a );
 a121497a <=( A299  and  (not A298) );
 a121500a <=( A301  and  (not A300) );
 a121501a <=( a121500a  and  a121497a );
 a121502a <=( a121501a  and  a121494a );
 a121505a <=( A168  and  A170 );
 a121508a <=( A166  and  (not A167) );
 a121509a <=( a121508a  and  a121505a );
 a121512a <=( (not A200)  and  A199 );
 a121515a <=( A203  and  (not A202) );
 a121516a <=( a121515a  and  a121512a );
 a121517a <=( a121516a  and  a121509a );
 a121520a <=( A266  and  (not A265) );
 a121523a <=( A269  and  (not A268) );
 a121524a <=( a121523a  and  a121520a );
 a121527a <=( A299  and  (not A298) );
 a121530a <=( (not A302)  and  (not A300) );
 a121531a <=( a121530a  and  a121527a );
 a121532a <=( a121531a  and  a121524a );
 a121535a <=( A168  and  A170 );
 a121538a <=( A166  and  (not A167) );
 a121539a <=( a121538a  and  a121535a );
 a121542a <=( (not A200)  and  A199 );
 a121545a <=( A203  and  (not A202) );
 a121546a <=( a121545a  and  a121542a );
 a121547a <=( a121546a  and  a121539a );
 a121550a <=( (not A266)  and  A265 );
 a121553a <=( A269  and  (not A268) );
 a121554a <=( a121553a  and  a121550a );
 a121557a <=( A299  and  A298 );
 a121560a <=( (not A301)  and  (not A300) );
 a121561a <=( a121560a  and  a121557a );
 a121562a <=( a121561a  and  a121554a );
 a121565a <=( A168  and  A170 );
 a121568a <=( A166  and  (not A167) );
 a121569a <=( a121568a  and  a121565a );
 a121572a <=( (not A200)  and  A199 );
 a121575a <=( A203  and  (not A202) );
 a121576a <=( a121575a  and  a121572a );
 a121577a <=( a121576a  and  a121569a );
 a121580a <=( (not A266)  and  A265 );
 a121583a <=( A269  and  (not A268) );
 a121584a <=( a121583a  and  a121580a );
 a121587a <=( A299  and  A298 );
 a121590a <=( A302  and  (not A300) );
 a121591a <=( a121590a  and  a121587a );
 a121592a <=( a121591a  and  a121584a );
 a121595a <=( A168  and  A170 );
 a121598a <=( A166  and  (not A167) );
 a121599a <=( a121598a  and  a121595a );
 a121602a <=( (not A200)  and  A199 );
 a121605a <=( A203  and  (not A202) );
 a121606a <=( a121605a  and  a121602a );
 a121607a <=( a121606a  and  a121599a );
 a121610a <=( (not A266)  and  A265 );
 a121613a <=( A269  and  (not A268) );
 a121614a <=( a121613a  and  a121610a );
 a121617a <=( (not A299)  and  A298 );
 a121620a <=( A301  and  (not A300) );
 a121621a <=( a121620a  and  a121617a );
 a121622a <=( a121621a  and  a121614a );
 a121625a <=( A168  and  A170 );
 a121628a <=( A166  and  (not A167) );
 a121629a <=( a121628a  and  a121625a );
 a121632a <=( (not A200)  and  A199 );
 a121635a <=( A203  and  (not A202) );
 a121636a <=( a121635a  and  a121632a );
 a121637a <=( a121636a  and  a121629a );
 a121640a <=( (not A266)  and  A265 );
 a121643a <=( A269  and  (not A268) );
 a121644a <=( a121643a  and  a121640a );
 a121647a <=( (not A299)  and  A298 );
 a121650a <=( (not A302)  and  (not A300) );
 a121651a <=( a121650a  and  a121647a );
 a121652a <=( a121651a  and  a121644a );
 a121655a <=( A168  and  A170 );
 a121658a <=( A166  and  (not A167) );
 a121659a <=( a121658a  and  a121655a );
 a121662a <=( (not A200)  and  A199 );
 a121665a <=( A203  and  (not A202) );
 a121666a <=( a121665a  and  a121662a );
 a121667a <=( a121666a  and  a121659a );
 a121670a <=( (not A266)  and  A265 );
 a121673a <=( A269  and  (not A268) );
 a121674a <=( a121673a  and  a121670a );
 a121677a <=( A299  and  (not A298) );
 a121680a <=( A301  and  (not A300) );
 a121681a <=( a121680a  and  a121677a );
 a121682a <=( a121681a  and  a121674a );
 a121685a <=( A168  and  A170 );
 a121688a <=( A166  and  (not A167) );
 a121689a <=( a121688a  and  a121685a );
 a121692a <=( (not A200)  and  A199 );
 a121695a <=( A203  and  (not A202) );
 a121696a <=( a121695a  and  a121692a );
 a121697a <=( a121696a  and  a121689a );
 a121700a <=( (not A266)  and  A265 );
 a121703a <=( A269  and  (not A268) );
 a121704a <=( a121703a  and  a121700a );
 a121707a <=( A299  and  (not A298) );
 a121710a <=( (not A302)  and  (not A300) );
 a121711a <=( a121710a  and  a121707a );
 a121712a <=( a121711a  and  a121704a );
 a121715a <=( A168  and  A170 );
 a121718a <=( A166  and  (not A167) );
 a121719a <=( a121718a  and  a121715a );
 a121722a <=( (not A200)  and  A199 );
 a121725a <=( A203  and  (not A202) );
 a121726a <=( a121725a  and  a121722a );
 a121727a <=( a121726a  and  a121719a );
 a121730a <=( (not A266)  and  (not A265) );
 a121733a <=( (not A269)  and  A268 );
 a121734a <=( a121733a  and  a121730a );
 a121737a <=( A299  and  A298 );
 a121740a <=( (not A301)  and  (not A300) );
 a121741a <=( a121740a  and  a121737a );
 a121742a <=( a121741a  and  a121734a );
 a121745a <=( A168  and  A170 );
 a121748a <=( A166  and  (not A167) );
 a121749a <=( a121748a  and  a121745a );
 a121752a <=( (not A200)  and  A199 );
 a121755a <=( A203  and  (not A202) );
 a121756a <=( a121755a  and  a121752a );
 a121757a <=( a121756a  and  a121749a );
 a121760a <=( (not A266)  and  (not A265) );
 a121763a <=( (not A269)  and  A268 );
 a121764a <=( a121763a  and  a121760a );
 a121767a <=( A299  and  A298 );
 a121770a <=( A302  and  (not A300) );
 a121771a <=( a121770a  and  a121767a );
 a121772a <=( a121771a  and  a121764a );
 a121775a <=( A168  and  A170 );
 a121778a <=( A166  and  (not A167) );
 a121779a <=( a121778a  and  a121775a );
 a121782a <=( (not A200)  and  A199 );
 a121785a <=( A203  and  (not A202) );
 a121786a <=( a121785a  and  a121782a );
 a121787a <=( a121786a  and  a121779a );
 a121790a <=( (not A266)  and  (not A265) );
 a121793a <=( (not A269)  and  A268 );
 a121794a <=( a121793a  and  a121790a );
 a121797a <=( (not A299)  and  A298 );
 a121800a <=( A301  and  (not A300) );
 a121801a <=( a121800a  and  a121797a );
 a121802a <=( a121801a  and  a121794a );
 a121805a <=( A168  and  A170 );
 a121808a <=( A166  and  (not A167) );
 a121809a <=( a121808a  and  a121805a );
 a121812a <=( (not A200)  and  A199 );
 a121815a <=( A203  and  (not A202) );
 a121816a <=( a121815a  and  a121812a );
 a121817a <=( a121816a  and  a121809a );
 a121820a <=( (not A266)  and  (not A265) );
 a121823a <=( (not A269)  and  A268 );
 a121824a <=( a121823a  and  a121820a );
 a121827a <=( (not A299)  and  A298 );
 a121830a <=( (not A302)  and  (not A300) );
 a121831a <=( a121830a  and  a121827a );
 a121832a <=( a121831a  and  a121824a );
 a121835a <=( A168  and  A170 );
 a121838a <=( A166  and  (not A167) );
 a121839a <=( a121838a  and  a121835a );
 a121842a <=( (not A200)  and  A199 );
 a121845a <=( A203  and  (not A202) );
 a121846a <=( a121845a  and  a121842a );
 a121847a <=( a121846a  and  a121839a );
 a121850a <=( (not A266)  and  (not A265) );
 a121853a <=( (not A269)  and  A268 );
 a121854a <=( a121853a  and  a121850a );
 a121857a <=( A299  and  (not A298) );
 a121860a <=( A301  and  (not A300) );
 a121861a <=( a121860a  and  a121857a );
 a121862a <=( a121861a  and  a121854a );
 a121865a <=( A168  and  A170 );
 a121868a <=( A166  and  (not A167) );
 a121869a <=( a121868a  and  a121865a );
 a121872a <=( (not A200)  and  A199 );
 a121875a <=( A203  and  (not A202) );
 a121876a <=( a121875a  and  a121872a );
 a121877a <=( a121876a  and  a121869a );
 a121880a <=( (not A266)  and  (not A265) );
 a121883a <=( (not A269)  and  A268 );
 a121884a <=( a121883a  and  a121880a );
 a121887a <=( A299  and  (not A298) );
 a121890a <=( (not A302)  and  (not A300) );
 a121891a <=( a121890a  and  a121887a );
 a121892a <=( a121891a  and  a121884a );
 a121895a <=( A168  and  A170 );
 a121898a <=( A166  and  (not A167) );
 a121899a <=( a121898a  and  a121895a );
 a121902a <=( (not A200)  and  A199 );
 a121905a <=( A202  and  (not A201) );
 a121906a <=( a121905a  and  a121902a );
 a121907a <=( a121906a  and  a121899a );
 a121910a <=( A266  and  A265 );
 a121913a <=( (not A268)  and  (not A267) );
 a121914a <=( a121913a  and  a121910a );
 a121917a <=( A299  and  A298 );
 a121920a <=( (not A302)  and  A301 );
 a121921a <=( a121920a  and  a121917a );
 a121922a <=( a121921a  and  a121914a );
 a121925a <=( A168  and  A170 );
 a121928a <=( A166  and  (not A167) );
 a121929a <=( a121928a  and  a121925a );
 a121932a <=( (not A200)  and  A199 );
 a121935a <=( A202  and  (not A201) );
 a121936a <=( a121935a  and  a121932a );
 a121937a <=( a121936a  and  a121929a );
 a121940a <=( A266  and  A265 );
 a121943a <=( (not A268)  and  (not A267) );
 a121944a <=( a121943a  and  a121940a );
 a121947a <=( (not A299)  and  A298 );
 a121950a <=( A302  and  (not A301) );
 a121951a <=( a121950a  and  a121947a );
 a121952a <=( a121951a  and  a121944a );
 a121955a <=( A168  and  A170 );
 a121958a <=( A166  and  (not A167) );
 a121959a <=( a121958a  and  a121955a );
 a121962a <=( (not A200)  and  A199 );
 a121965a <=( A202  and  (not A201) );
 a121966a <=( a121965a  and  a121962a );
 a121967a <=( a121966a  and  a121959a );
 a121970a <=( A266  and  A265 );
 a121973a <=( (not A268)  and  (not A267) );
 a121974a <=( a121973a  and  a121970a );
 a121977a <=( A299  and  (not A298) );
 a121980a <=( A302  and  (not A301) );
 a121981a <=( a121980a  and  a121977a );
 a121982a <=( a121981a  and  a121974a );
 a121985a <=( A168  and  A170 );
 a121988a <=( A166  and  (not A167) );
 a121989a <=( a121988a  and  a121985a );
 a121992a <=( (not A200)  and  A199 );
 a121995a <=( A202  and  (not A201) );
 a121996a <=( a121995a  and  a121992a );
 a121997a <=( a121996a  and  a121989a );
 a122000a <=( A266  and  A265 );
 a122003a <=( (not A268)  and  (not A267) );
 a122004a <=( a122003a  and  a122000a );
 a122007a <=( (not A299)  and  (not A298) );
 a122010a <=( (not A302)  and  A301 );
 a122011a <=( a122010a  and  a122007a );
 a122012a <=( a122011a  and  a122004a );
 a122015a <=( A168  and  A170 );
 a122018a <=( A166  and  (not A167) );
 a122019a <=( a122018a  and  a122015a );
 a122022a <=( (not A200)  and  A199 );
 a122025a <=( A202  and  (not A201) );
 a122026a <=( a122025a  and  a122022a );
 a122027a <=( a122026a  and  a122019a );
 a122030a <=( A266  and  A265 );
 a122033a <=( A269  and  (not A267) );
 a122034a <=( a122033a  and  a122030a );
 a122037a <=( A299  and  A298 );
 a122040a <=( (not A302)  and  A301 );
 a122041a <=( a122040a  and  a122037a );
 a122042a <=( a122041a  and  a122034a );
 a122045a <=( A168  and  A170 );
 a122048a <=( A166  and  (not A167) );
 a122049a <=( a122048a  and  a122045a );
 a122052a <=( (not A200)  and  A199 );
 a122055a <=( A202  and  (not A201) );
 a122056a <=( a122055a  and  a122052a );
 a122057a <=( a122056a  and  a122049a );
 a122060a <=( A266  and  A265 );
 a122063a <=( A269  and  (not A267) );
 a122064a <=( a122063a  and  a122060a );
 a122067a <=( (not A299)  and  A298 );
 a122070a <=( A302  and  (not A301) );
 a122071a <=( a122070a  and  a122067a );
 a122072a <=( a122071a  and  a122064a );
 a122075a <=( A168  and  A170 );
 a122078a <=( A166  and  (not A167) );
 a122079a <=( a122078a  and  a122075a );
 a122082a <=( (not A200)  and  A199 );
 a122085a <=( A202  and  (not A201) );
 a122086a <=( a122085a  and  a122082a );
 a122087a <=( a122086a  and  a122079a );
 a122090a <=( A266  and  A265 );
 a122093a <=( A269  and  (not A267) );
 a122094a <=( a122093a  and  a122090a );
 a122097a <=( A299  and  (not A298) );
 a122100a <=( A302  and  (not A301) );
 a122101a <=( a122100a  and  a122097a );
 a122102a <=( a122101a  and  a122094a );
 a122105a <=( A168  and  A170 );
 a122108a <=( A166  and  (not A167) );
 a122109a <=( a122108a  and  a122105a );
 a122112a <=( (not A200)  and  A199 );
 a122115a <=( A202  and  (not A201) );
 a122116a <=( a122115a  and  a122112a );
 a122117a <=( a122116a  and  a122109a );
 a122120a <=( A266  and  A265 );
 a122123a <=( A269  and  (not A267) );
 a122124a <=( a122123a  and  a122120a );
 a122127a <=( (not A299)  and  (not A298) );
 a122130a <=( (not A302)  and  A301 );
 a122131a <=( a122130a  and  a122127a );
 a122132a <=( a122131a  and  a122124a );
 a122135a <=( A168  and  A170 );
 a122138a <=( A166  and  (not A167) );
 a122139a <=( a122138a  and  a122135a );
 a122142a <=( (not A200)  and  A199 );
 a122145a <=( A202  and  (not A201) );
 a122146a <=( a122145a  and  a122142a );
 a122147a <=( a122146a  and  a122139a );
 a122150a <=( A266  and  (not A265) );
 a122153a <=( A268  and  (not A267) );
 a122154a <=( a122153a  and  a122150a );
 a122157a <=( A299  and  A298 );
 a122160a <=( (not A302)  and  A301 );
 a122161a <=( a122160a  and  a122157a );
 a122162a <=( a122161a  and  a122154a );
 a122165a <=( A168  and  A170 );
 a122168a <=( A166  and  (not A167) );
 a122169a <=( a122168a  and  a122165a );
 a122172a <=( (not A200)  and  A199 );
 a122175a <=( A202  and  (not A201) );
 a122176a <=( a122175a  and  a122172a );
 a122177a <=( a122176a  and  a122169a );
 a122180a <=( A266  and  (not A265) );
 a122183a <=( A268  and  (not A267) );
 a122184a <=( a122183a  and  a122180a );
 a122187a <=( (not A299)  and  A298 );
 a122190a <=( A302  and  (not A301) );
 a122191a <=( a122190a  and  a122187a );
 a122192a <=( a122191a  and  a122184a );
 a122195a <=( A168  and  A170 );
 a122198a <=( A166  and  (not A167) );
 a122199a <=( a122198a  and  a122195a );
 a122202a <=( (not A200)  and  A199 );
 a122205a <=( A202  and  (not A201) );
 a122206a <=( a122205a  and  a122202a );
 a122207a <=( a122206a  and  a122199a );
 a122210a <=( A266  and  (not A265) );
 a122213a <=( A268  and  (not A267) );
 a122214a <=( a122213a  and  a122210a );
 a122217a <=( A299  and  (not A298) );
 a122220a <=( A302  and  (not A301) );
 a122221a <=( a122220a  and  a122217a );
 a122222a <=( a122221a  and  a122214a );
 a122225a <=( A168  and  A170 );
 a122228a <=( A166  and  (not A167) );
 a122229a <=( a122228a  and  a122225a );
 a122232a <=( (not A200)  and  A199 );
 a122235a <=( A202  and  (not A201) );
 a122236a <=( a122235a  and  a122232a );
 a122237a <=( a122236a  and  a122229a );
 a122240a <=( A266  and  (not A265) );
 a122243a <=( A268  and  (not A267) );
 a122244a <=( a122243a  and  a122240a );
 a122247a <=( (not A299)  and  (not A298) );
 a122250a <=( (not A302)  and  A301 );
 a122251a <=( a122250a  and  a122247a );
 a122252a <=( a122251a  and  a122244a );
 a122255a <=( A168  and  A170 );
 a122258a <=( A166  and  (not A167) );
 a122259a <=( a122258a  and  a122255a );
 a122262a <=( (not A200)  and  A199 );
 a122265a <=( A202  and  (not A201) );
 a122266a <=( a122265a  and  a122262a );
 a122267a <=( a122266a  and  a122259a );
 a122270a <=( A266  and  (not A265) );
 a122273a <=( (not A269)  and  (not A267) );
 a122274a <=( a122273a  and  a122270a );
 a122277a <=( A299  and  A298 );
 a122280a <=( (not A302)  and  A301 );
 a122281a <=( a122280a  and  a122277a );
 a122282a <=( a122281a  and  a122274a );
 a122285a <=( A168  and  A170 );
 a122288a <=( A166  and  (not A167) );
 a122289a <=( a122288a  and  a122285a );
 a122292a <=( (not A200)  and  A199 );
 a122295a <=( A202  and  (not A201) );
 a122296a <=( a122295a  and  a122292a );
 a122297a <=( a122296a  and  a122289a );
 a122300a <=( A266  and  (not A265) );
 a122303a <=( (not A269)  and  (not A267) );
 a122304a <=( a122303a  and  a122300a );
 a122307a <=( (not A299)  and  A298 );
 a122310a <=( A302  and  (not A301) );
 a122311a <=( a122310a  and  a122307a );
 a122312a <=( a122311a  and  a122304a );
 a122315a <=( A168  and  A170 );
 a122318a <=( A166  and  (not A167) );
 a122319a <=( a122318a  and  a122315a );
 a122322a <=( (not A200)  and  A199 );
 a122325a <=( A202  and  (not A201) );
 a122326a <=( a122325a  and  a122322a );
 a122327a <=( a122326a  and  a122319a );
 a122330a <=( A266  and  (not A265) );
 a122333a <=( (not A269)  and  (not A267) );
 a122334a <=( a122333a  and  a122330a );
 a122337a <=( A299  and  (not A298) );
 a122340a <=( A302  and  (not A301) );
 a122341a <=( a122340a  and  a122337a );
 a122342a <=( a122341a  and  a122334a );
 a122345a <=( A168  and  A170 );
 a122348a <=( A166  and  (not A167) );
 a122349a <=( a122348a  and  a122345a );
 a122352a <=( (not A200)  and  A199 );
 a122355a <=( A202  and  (not A201) );
 a122356a <=( a122355a  and  a122352a );
 a122357a <=( a122356a  and  a122349a );
 a122360a <=( A266  and  (not A265) );
 a122363a <=( (not A269)  and  (not A267) );
 a122364a <=( a122363a  and  a122360a );
 a122367a <=( (not A299)  and  (not A298) );
 a122370a <=( (not A302)  and  A301 );
 a122371a <=( a122370a  and  a122367a );
 a122372a <=( a122371a  and  a122364a );
 a122375a <=( A168  and  A170 );
 a122378a <=( A166  and  (not A167) );
 a122379a <=( a122378a  and  a122375a );
 a122382a <=( (not A200)  and  A199 );
 a122385a <=( A202  and  (not A201) );
 a122386a <=( a122385a  and  a122382a );
 a122387a <=( a122386a  and  a122379a );
 a122390a <=( (not A266)  and  A265 );
 a122393a <=( A268  and  (not A267) );
 a122394a <=( a122393a  and  a122390a );
 a122397a <=( A299  and  A298 );
 a122400a <=( (not A302)  and  A301 );
 a122401a <=( a122400a  and  a122397a );
 a122402a <=( a122401a  and  a122394a );
 a122405a <=( A168  and  A170 );
 a122408a <=( A166  and  (not A167) );
 a122409a <=( a122408a  and  a122405a );
 a122412a <=( (not A200)  and  A199 );
 a122415a <=( A202  and  (not A201) );
 a122416a <=( a122415a  and  a122412a );
 a122417a <=( a122416a  and  a122409a );
 a122420a <=( (not A266)  and  A265 );
 a122423a <=( A268  and  (not A267) );
 a122424a <=( a122423a  and  a122420a );
 a122427a <=( (not A299)  and  A298 );
 a122430a <=( A302  and  (not A301) );
 a122431a <=( a122430a  and  a122427a );
 a122432a <=( a122431a  and  a122424a );
 a122435a <=( A168  and  A170 );
 a122438a <=( A166  and  (not A167) );
 a122439a <=( a122438a  and  a122435a );
 a122442a <=( (not A200)  and  A199 );
 a122445a <=( A202  and  (not A201) );
 a122446a <=( a122445a  and  a122442a );
 a122447a <=( a122446a  and  a122439a );
 a122450a <=( (not A266)  and  A265 );
 a122453a <=( A268  and  (not A267) );
 a122454a <=( a122453a  and  a122450a );
 a122457a <=( A299  and  (not A298) );
 a122460a <=( A302  and  (not A301) );
 a122461a <=( a122460a  and  a122457a );
 a122462a <=( a122461a  and  a122454a );
 a122465a <=( A168  and  A170 );
 a122468a <=( A166  and  (not A167) );
 a122469a <=( a122468a  and  a122465a );
 a122472a <=( (not A200)  and  A199 );
 a122475a <=( A202  and  (not A201) );
 a122476a <=( a122475a  and  a122472a );
 a122477a <=( a122476a  and  a122469a );
 a122480a <=( (not A266)  and  A265 );
 a122483a <=( A268  and  (not A267) );
 a122484a <=( a122483a  and  a122480a );
 a122487a <=( (not A299)  and  (not A298) );
 a122490a <=( (not A302)  and  A301 );
 a122491a <=( a122490a  and  a122487a );
 a122492a <=( a122491a  and  a122484a );
 a122495a <=( A168  and  A170 );
 a122498a <=( A166  and  (not A167) );
 a122499a <=( a122498a  and  a122495a );
 a122502a <=( (not A200)  and  A199 );
 a122505a <=( A202  and  (not A201) );
 a122506a <=( a122505a  and  a122502a );
 a122507a <=( a122506a  and  a122499a );
 a122510a <=( (not A266)  and  A265 );
 a122513a <=( (not A269)  and  (not A267) );
 a122514a <=( a122513a  and  a122510a );
 a122517a <=( A299  and  A298 );
 a122520a <=( (not A302)  and  A301 );
 a122521a <=( a122520a  and  a122517a );
 a122522a <=( a122521a  and  a122514a );
 a122525a <=( A168  and  A170 );
 a122528a <=( A166  and  (not A167) );
 a122529a <=( a122528a  and  a122525a );
 a122532a <=( (not A200)  and  A199 );
 a122535a <=( A202  and  (not A201) );
 a122536a <=( a122535a  and  a122532a );
 a122537a <=( a122536a  and  a122529a );
 a122540a <=( (not A266)  and  A265 );
 a122543a <=( (not A269)  and  (not A267) );
 a122544a <=( a122543a  and  a122540a );
 a122547a <=( (not A299)  and  A298 );
 a122550a <=( A302  and  (not A301) );
 a122551a <=( a122550a  and  a122547a );
 a122552a <=( a122551a  and  a122544a );
 a122555a <=( A168  and  A170 );
 a122558a <=( A166  and  (not A167) );
 a122559a <=( a122558a  and  a122555a );
 a122562a <=( (not A200)  and  A199 );
 a122565a <=( A202  and  (not A201) );
 a122566a <=( a122565a  and  a122562a );
 a122567a <=( a122566a  and  a122559a );
 a122570a <=( (not A266)  and  A265 );
 a122573a <=( (not A269)  and  (not A267) );
 a122574a <=( a122573a  and  a122570a );
 a122577a <=( A299  and  (not A298) );
 a122580a <=( A302  and  (not A301) );
 a122581a <=( a122580a  and  a122577a );
 a122582a <=( a122581a  and  a122574a );
 a122585a <=( A168  and  A170 );
 a122588a <=( A166  and  (not A167) );
 a122589a <=( a122588a  and  a122585a );
 a122592a <=( (not A200)  and  A199 );
 a122595a <=( A202  and  (not A201) );
 a122596a <=( a122595a  and  a122592a );
 a122597a <=( a122596a  and  a122589a );
 a122600a <=( (not A266)  and  A265 );
 a122603a <=( (not A269)  and  (not A267) );
 a122604a <=( a122603a  and  a122600a );
 a122607a <=( (not A299)  and  (not A298) );
 a122610a <=( (not A302)  and  A301 );
 a122611a <=( a122610a  and  a122607a );
 a122612a <=( a122611a  and  a122604a );
 a122615a <=( A168  and  A170 );
 a122618a <=( A166  and  (not A167) );
 a122619a <=( a122618a  and  a122615a );
 a122622a <=( (not A200)  and  A199 );
 a122625a <=( (not A203)  and  (not A201) );
 a122626a <=( a122625a  and  a122622a );
 a122627a <=( a122626a  and  a122619a );
 a122630a <=( A266  and  A265 );
 a122633a <=( (not A268)  and  (not A267) );
 a122634a <=( a122633a  and  a122630a );
 a122637a <=( A299  and  A298 );
 a122640a <=( (not A302)  and  A301 );
 a122641a <=( a122640a  and  a122637a );
 a122642a <=( a122641a  and  a122634a );
 a122645a <=( A168  and  A170 );
 a122648a <=( A166  and  (not A167) );
 a122649a <=( a122648a  and  a122645a );
 a122652a <=( (not A200)  and  A199 );
 a122655a <=( (not A203)  and  (not A201) );
 a122656a <=( a122655a  and  a122652a );
 a122657a <=( a122656a  and  a122649a );
 a122660a <=( A266  and  A265 );
 a122663a <=( (not A268)  and  (not A267) );
 a122664a <=( a122663a  and  a122660a );
 a122667a <=( (not A299)  and  A298 );
 a122670a <=( A302  and  (not A301) );
 a122671a <=( a122670a  and  a122667a );
 a122672a <=( a122671a  and  a122664a );
 a122675a <=( A168  and  A170 );
 a122678a <=( A166  and  (not A167) );
 a122679a <=( a122678a  and  a122675a );
 a122682a <=( (not A200)  and  A199 );
 a122685a <=( (not A203)  and  (not A201) );
 a122686a <=( a122685a  and  a122682a );
 a122687a <=( a122686a  and  a122679a );
 a122690a <=( A266  and  A265 );
 a122693a <=( (not A268)  and  (not A267) );
 a122694a <=( a122693a  and  a122690a );
 a122697a <=( A299  and  (not A298) );
 a122700a <=( A302  and  (not A301) );
 a122701a <=( a122700a  and  a122697a );
 a122702a <=( a122701a  and  a122694a );
 a122705a <=( A168  and  A170 );
 a122708a <=( A166  and  (not A167) );
 a122709a <=( a122708a  and  a122705a );
 a122712a <=( (not A200)  and  A199 );
 a122715a <=( (not A203)  and  (not A201) );
 a122716a <=( a122715a  and  a122712a );
 a122717a <=( a122716a  and  a122709a );
 a122720a <=( A266  and  A265 );
 a122723a <=( (not A268)  and  (not A267) );
 a122724a <=( a122723a  and  a122720a );
 a122727a <=( (not A299)  and  (not A298) );
 a122730a <=( (not A302)  and  A301 );
 a122731a <=( a122730a  and  a122727a );
 a122732a <=( a122731a  and  a122724a );
 a122735a <=( A168  and  A170 );
 a122738a <=( A166  and  (not A167) );
 a122739a <=( a122738a  and  a122735a );
 a122742a <=( (not A200)  and  A199 );
 a122745a <=( (not A203)  and  (not A201) );
 a122746a <=( a122745a  and  a122742a );
 a122747a <=( a122746a  and  a122739a );
 a122750a <=( A266  and  A265 );
 a122753a <=( A269  and  (not A267) );
 a122754a <=( a122753a  and  a122750a );
 a122757a <=( A299  and  A298 );
 a122760a <=( (not A302)  and  A301 );
 a122761a <=( a122760a  and  a122757a );
 a122762a <=( a122761a  and  a122754a );
 a122765a <=( A168  and  A170 );
 a122768a <=( A166  and  (not A167) );
 a122769a <=( a122768a  and  a122765a );
 a122772a <=( (not A200)  and  A199 );
 a122775a <=( (not A203)  and  (not A201) );
 a122776a <=( a122775a  and  a122772a );
 a122777a <=( a122776a  and  a122769a );
 a122780a <=( A266  and  A265 );
 a122783a <=( A269  and  (not A267) );
 a122784a <=( a122783a  and  a122780a );
 a122787a <=( (not A299)  and  A298 );
 a122790a <=( A302  and  (not A301) );
 a122791a <=( a122790a  and  a122787a );
 a122792a <=( a122791a  and  a122784a );
 a122795a <=( A168  and  A170 );
 a122798a <=( A166  and  (not A167) );
 a122799a <=( a122798a  and  a122795a );
 a122802a <=( (not A200)  and  A199 );
 a122805a <=( (not A203)  and  (not A201) );
 a122806a <=( a122805a  and  a122802a );
 a122807a <=( a122806a  and  a122799a );
 a122810a <=( A266  and  A265 );
 a122813a <=( A269  and  (not A267) );
 a122814a <=( a122813a  and  a122810a );
 a122817a <=( A299  and  (not A298) );
 a122820a <=( A302  and  (not A301) );
 a122821a <=( a122820a  and  a122817a );
 a122822a <=( a122821a  and  a122814a );
 a122825a <=( A168  and  A170 );
 a122828a <=( A166  and  (not A167) );
 a122829a <=( a122828a  and  a122825a );
 a122832a <=( (not A200)  and  A199 );
 a122835a <=( (not A203)  and  (not A201) );
 a122836a <=( a122835a  and  a122832a );
 a122837a <=( a122836a  and  a122829a );
 a122840a <=( A266  and  A265 );
 a122843a <=( A269  and  (not A267) );
 a122844a <=( a122843a  and  a122840a );
 a122847a <=( (not A299)  and  (not A298) );
 a122850a <=( (not A302)  and  A301 );
 a122851a <=( a122850a  and  a122847a );
 a122852a <=( a122851a  and  a122844a );
 a122855a <=( A168  and  A170 );
 a122858a <=( A166  and  (not A167) );
 a122859a <=( a122858a  and  a122855a );
 a122862a <=( (not A200)  and  A199 );
 a122865a <=( (not A203)  and  (not A201) );
 a122866a <=( a122865a  and  a122862a );
 a122867a <=( a122866a  and  a122859a );
 a122870a <=( A266  and  (not A265) );
 a122873a <=( A268  and  (not A267) );
 a122874a <=( a122873a  and  a122870a );
 a122877a <=( A299  and  A298 );
 a122880a <=( (not A302)  and  A301 );
 a122881a <=( a122880a  and  a122877a );
 a122882a <=( a122881a  and  a122874a );
 a122885a <=( A168  and  A170 );
 a122888a <=( A166  and  (not A167) );
 a122889a <=( a122888a  and  a122885a );
 a122892a <=( (not A200)  and  A199 );
 a122895a <=( (not A203)  and  (not A201) );
 a122896a <=( a122895a  and  a122892a );
 a122897a <=( a122896a  and  a122889a );
 a122900a <=( A266  and  (not A265) );
 a122903a <=( A268  and  (not A267) );
 a122904a <=( a122903a  and  a122900a );
 a122907a <=( (not A299)  and  A298 );
 a122910a <=( A302  and  (not A301) );
 a122911a <=( a122910a  and  a122907a );
 a122912a <=( a122911a  and  a122904a );
 a122915a <=( A168  and  A170 );
 a122918a <=( A166  and  (not A167) );
 a122919a <=( a122918a  and  a122915a );
 a122922a <=( (not A200)  and  A199 );
 a122925a <=( (not A203)  and  (not A201) );
 a122926a <=( a122925a  and  a122922a );
 a122927a <=( a122926a  and  a122919a );
 a122930a <=( A266  and  (not A265) );
 a122933a <=( A268  and  (not A267) );
 a122934a <=( a122933a  and  a122930a );
 a122937a <=( A299  and  (not A298) );
 a122940a <=( A302  and  (not A301) );
 a122941a <=( a122940a  and  a122937a );
 a122942a <=( a122941a  and  a122934a );
 a122945a <=( A168  and  A170 );
 a122948a <=( A166  and  (not A167) );
 a122949a <=( a122948a  and  a122945a );
 a122952a <=( (not A200)  and  A199 );
 a122955a <=( (not A203)  and  (not A201) );
 a122956a <=( a122955a  and  a122952a );
 a122957a <=( a122956a  and  a122949a );
 a122960a <=( A266  and  (not A265) );
 a122963a <=( A268  and  (not A267) );
 a122964a <=( a122963a  and  a122960a );
 a122967a <=( (not A299)  and  (not A298) );
 a122970a <=( (not A302)  and  A301 );
 a122971a <=( a122970a  and  a122967a );
 a122972a <=( a122971a  and  a122964a );
 a122975a <=( A168  and  A170 );
 a122978a <=( A166  and  (not A167) );
 a122979a <=( a122978a  and  a122975a );
 a122982a <=( (not A200)  and  A199 );
 a122985a <=( (not A203)  and  (not A201) );
 a122986a <=( a122985a  and  a122982a );
 a122987a <=( a122986a  and  a122979a );
 a122990a <=( A266  and  (not A265) );
 a122993a <=( (not A269)  and  (not A267) );
 a122994a <=( a122993a  and  a122990a );
 a122997a <=( A299  and  A298 );
 a123000a <=( (not A302)  and  A301 );
 a123001a <=( a123000a  and  a122997a );
 a123002a <=( a123001a  and  a122994a );
 a123005a <=( A168  and  A170 );
 a123008a <=( A166  and  (not A167) );
 a123009a <=( a123008a  and  a123005a );
 a123012a <=( (not A200)  and  A199 );
 a123015a <=( (not A203)  and  (not A201) );
 a123016a <=( a123015a  and  a123012a );
 a123017a <=( a123016a  and  a123009a );
 a123020a <=( A266  and  (not A265) );
 a123023a <=( (not A269)  and  (not A267) );
 a123024a <=( a123023a  and  a123020a );
 a123027a <=( (not A299)  and  A298 );
 a123030a <=( A302  and  (not A301) );
 a123031a <=( a123030a  and  a123027a );
 a123032a <=( a123031a  and  a123024a );
 a123035a <=( A168  and  A170 );
 a123038a <=( A166  and  (not A167) );
 a123039a <=( a123038a  and  a123035a );
 a123042a <=( (not A200)  and  A199 );
 a123045a <=( (not A203)  and  (not A201) );
 a123046a <=( a123045a  and  a123042a );
 a123047a <=( a123046a  and  a123039a );
 a123050a <=( A266  and  (not A265) );
 a123053a <=( (not A269)  and  (not A267) );
 a123054a <=( a123053a  and  a123050a );
 a123057a <=( A299  and  (not A298) );
 a123060a <=( A302  and  (not A301) );
 a123061a <=( a123060a  and  a123057a );
 a123062a <=( a123061a  and  a123054a );
 a123065a <=( A168  and  A170 );
 a123068a <=( A166  and  (not A167) );
 a123069a <=( a123068a  and  a123065a );
 a123072a <=( (not A200)  and  A199 );
 a123075a <=( (not A203)  and  (not A201) );
 a123076a <=( a123075a  and  a123072a );
 a123077a <=( a123076a  and  a123069a );
 a123080a <=( A266  and  (not A265) );
 a123083a <=( (not A269)  and  (not A267) );
 a123084a <=( a123083a  and  a123080a );
 a123087a <=( (not A299)  and  (not A298) );
 a123090a <=( (not A302)  and  A301 );
 a123091a <=( a123090a  and  a123087a );
 a123092a <=( a123091a  and  a123084a );
 a123095a <=( A168  and  A170 );
 a123098a <=( A166  and  (not A167) );
 a123099a <=( a123098a  and  a123095a );
 a123102a <=( (not A200)  and  A199 );
 a123105a <=( (not A203)  and  (not A201) );
 a123106a <=( a123105a  and  a123102a );
 a123107a <=( a123106a  and  a123099a );
 a123110a <=( (not A266)  and  A265 );
 a123113a <=( A268  and  (not A267) );
 a123114a <=( a123113a  and  a123110a );
 a123117a <=( A299  and  A298 );
 a123120a <=( (not A302)  and  A301 );
 a123121a <=( a123120a  and  a123117a );
 a123122a <=( a123121a  and  a123114a );
 a123125a <=( A168  and  A170 );
 a123128a <=( A166  and  (not A167) );
 a123129a <=( a123128a  and  a123125a );
 a123132a <=( (not A200)  and  A199 );
 a123135a <=( (not A203)  and  (not A201) );
 a123136a <=( a123135a  and  a123132a );
 a123137a <=( a123136a  and  a123129a );
 a123140a <=( (not A266)  and  A265 );
 a123143a <=( A268  and  (not A267) );
 a123144a <=( a123143a  and  a123140a );
 a123147a <=( (not A299)  and  A298 );
 a123150a <=( A302  and  (not A301) );
 a123151a <=( a123150a  and  a123147a );
 a123152a <=( a123151a  and  a123144a );
 a123155a <=( A168  and  A170 );
 a123158a <=( A166  and  (not A167) );
 a123159a <=( a123158a  and  a123155a );
 a123162a <=( (not A200)  and  A199 );
 a123165a <=( (not A203)  and  (not A201) );
 a123166a <=( a123165a  and  a123162a );
 a123167a <=( a123166a  and  a123159a );
 a123170a <=( (not A266)  and  A265 );
 a123173a <=( A268  and  (not A267) );
 a123174a <=( a123173a  and  a123170a );
 a123177a <=( A299  and  (not A298) );
 a123180a <=( A302  and  (not A301) );
 a123181a <=( a123180a  and  a123177a );
 a123182a <=( a123181a  and  a123174a );
 a123185a <=( A168  and  A170 );
 a123188a <=( A166  and  (not A167) );
 a123189a <=( a123188a  and  a123185a );
 a123192a <=( (not A200)  and  A199 );
 a123195a <=( (not A203)  and  (not A201) );
 a123196a <=( a123195a  and  a123192a );
 a123197a <=( a123196a  and  a123189a );
 a123200a <=( (not A266)  and  A265 );
 a123203a <=( A268  and  (not A267) );
 a123204a <=( a123203a  and  a123200a );
 a123207a <=( (not A299)  and  (not A298) );
 a123210a <=( (not A302)  and  A301 );
 a123211a <=( a123210a  and  a123207a );
 a123212a <=( a123211a  and  a123204a );
 a123215a <=( A168  and  A170 );
 a123218a <=( A166  and  (not A167) );
 a123219a <=( a123218a  and  a123215a );
 a123222a <=( (not A200)  and  A199 );
 a123225a <=( (not A203)  and  (not A201) );
 a123226a <=( a123225a  and  a123222a );
 a123227a <=( a123226a  and  a123219a );
 a123230a <=( (not A266)  and  A265 );
 a123233a <=( (not A269)  and  (not A267) );
 a123234a <=( a123233a  and  a123230a );
 a123237a <=( A299  and  A298 );
 a123240a <=( (not A302)  and  A301 );
 a123241a <=( a123240a  and  a123237a );
 a123242a <=( a123241a  and  a123234a );
 a123245a <=( A168  and  A170 );
 a123248a <=( A166  and  (not A167) );
 a123249a <=( a123248a  and  a123245a );
 a123252a <=( (not A200)  and  A199 );
 a123255a <=( (not A203)  and  (not A201) );
 a123256a <=( a123255a  and  a123252a );
 a123257a <=( a123256a  and  a123249a );
 a123260a <=( (not A266)  and  A265 );
 a123263a <=( (not A269)  and  (not A267) );
 a123264a <=( a123263a  and  a123260a );
 a123267a <=( (not A299)  and  A298 );
 a123270a <=( A302  and  (not A301) );
 a123271a <=( a123270a  and  a123267a );
 a123272a <=( a123271a  and  a123264a );
 a123275a <=( A168  and  A170 );
 a123278a <=( A166  and  (not A167) );
 a123279a <=( a123278a  and  a123275a );
 a123282a <=( (not A200)  and  A199 );
 a123285a <=( (not A203)  and  (not A201) );
 a123286a <=( a123285a  and  a123282a );
 a123287a <=( a123286a  and  a123279a );
 a123290a <=( (not A266)  and  A265 );
 a123293a <=( (not A269)  and  (not A267) );
 a123294a <=( a123293a  and  a123290a );
 a123297a <=( A299  and  (not A298) );
 a123300a <=( A302  and  (not A301) );
 a123301a <=( a123300a  and  a123297a );
 a123302a <=( a123301a  and  a123294a );
 a123305a <=( A168  and  A170 );
 a123308a <=( A166  and  (not A167) );
 a123309a <=( a123308a  and  a123305a );
 a123312a <=( (not A200)  and  A199 );
 a123315a <=( (not A203)  and  (not A201) );
 a123316a <=( a123315a  and  a123312a );
 a123317a <=( a123316a  and  a123309a );
 a123320a <=( (not A266)  and  A265 );
 a123323a <=( (not A269)  and  (not A267) );
 a123324a <=( a123323a  and  a123320a );
 a123327a <=( (not A299)  and  (not A298) );
 a123330a <=( (not A302)  and  A301 );
 a123331a <=( a123330a  and  a123327a );
 a123332a <=( a123331a  and  a123324a );
 a123335a <=( A168  and  A170 );
 a123338a <=( A166  and  (not A167) );
 a123339a <=( a123338a  and  a123335a );
 a123342a <=( (not A200)  and  (not A199) );
 a123345a <=( (not A203)  and  A202 );
 a123346a <=( a123345a  and  a123342a );
 a123347a <=( a123346a  and  a123339a );
 a123350a <=( A266  and  A265 );
 a123353a <=( (not A269)  and  A268 );
 a123354a <=( a123353a  and  a123350a );
 a123357a <=( A299  and  A298 );
 a123360a <=( (not A301)  and  (not A300) );
 a123361a <=( a123360a  and  a123357a );
 a123362a <=( a123361a  and  a123354a );
 a123365a <=( A168  and  A170 );
 a123368a <=( A166  and  (not A167) );
 a123369a <=( a123368a  and  a123365a );
 a123372a <=( (not A200)  and  (not A199) );
 a123375a <=( (not A203)  and  A202 );
 a123376a <=( a123375a  and  a123372a );
 a123377a <=( a123376a  and  a123369a );
 a123380a <=( A266  and  A265 );
 a123383a <=( (not A269)  and  A268 );
 a123384a <=( a123383a  and  a123380a );
 a123387a <=( A299  and  A298 );
 a123390a <=( A302  and  (not A300) );
 a123391a <=( a123390a  and  a123387a );
 a123392a <=( a123391a  and  a123384a );
 a123395a <=( A168  and  A170 );
 a123398a <=( A166  and  (not A167) );
 a123399a <=( a123398a  and  a123395a );
 a123402a <=( (not A200)  and  (not A199) );
 a123405a <=( (not A203)  and  A202 );
 a123406a <=( a123405a  and  a123402a );
 a123407a <=( a123406a  and  a123399a );
 a123410a <=( A266  and  A265 );
 a123413a <=( (not A269)  and  A268 );
 a123414a <=( a123413a  and  a123410a );
 a123417a <=( (not A299)  and  A298 );
 a123420a <=( A301  and  (not A300) );
 a123421a <=( a123420a  and  a123417a );
 a123422a <=( a123421a  and  a123414a );
 a123425a <=( A168  and  A170 );
 a123428a <=( A166  and  (not A167) );
 a123429a <=( a123428a  and  a123425a );
 a123432a <=( (not A200)  and  (not A199) );
 a123435a <=( (not A203)  and  A202 );
 a123436a <=( a123435a  and  a123432a );
 a123437a <=( a123436a  and  a123429a );
 a123440a <=( A266  and  A265 );
 a123443a <=( (not A269)  and  A268 );
 a123444a <=( a123443a  and  a123440a );
 a123447a <=( (not A299)  and  A298 );
 a123450a <=( (not A302)  and  (not A300) );
 a123451a <=( a123450a  and  a123447a );
 a123452a <=( a123451a  and  a123444a );
 a123455a <=( A168  and  A170 );
 a123458a <=( A166  and  (not A167) );
 a123459a <=( a123458a  and  a123455a );
 a123462a <=( (not A200)  and  (not A199) );
 a123465a <=( (not A203)  and  A202 );
 a123466a <=( a123465a  and  a123462a );
 a123467a <=( a123466a  and  a123459a );
 a123470a <=( A266  and  A265 );
 a123473a <=( (not A269)  and  A268 );
 a123474a <=( a123473a  and  a123470a );
 a123477a <=( A299  and  (not A298) );
 a123480a <=( A301  and  (not A300) );
 a123481a <=( a123480a  and  a123477a );
 a123482a <=( a123481a  and  a123474a );
 a123485a <=( A168  and  A170 );
 a123488a <=( A166  and  (not A167) );
 a123489a <=( a123488a  and  a123485a );
 a123492a <=( (not A200)  and  (not A199) );
 a123495a <=( (not A203)  and  A202 );
 a123496a <=( a123495a  and  a123492a );
 a123497a <=( a123496a  and  a123489a );
 a123500a <=( A266  and  A265 );
 a123503a <=( (not A269)  and  A268 );
 a123504a <=( a123503a  and  a123500a );
 a123507a <=( A299  and  (not A298) );
 a123510a <=( (not A302)  and  (not A300) );
 a123511a <=( a123510a  and  a123507a );
 a123512a <=( a123511a  and  a123504a );
 a123515a <=( A168  and  A170 );
 a123518a <=( A166  and  (not A167) );
 a123519a <=( a123518a  and  a123515a );
 a123522a <=( (not A200)  and  (not A199) );
 a123525a <=( (not A203)  and  A202 );
 a123526a <=( a123525a  and  a123522a );
 a123527a <=( a123526a  and  a123519a );
 a123530a <=( A266  and  (not A265) );
 a123533a <=( A269  and  (not A268) );
 a123534a <=( a123533a  and  a123530a );
 a123537a <=( A299  and  A298 );
 a123540a <=( (not A301)  and  (not A300) );
 a123541a <=( a123540a  and  a123537a );
 a123542a <=( a123541a  and  a123534a );
 a123545a <=( A168  and  A170 );
 a123548a <=( A166  and  (not A167) );
 a123549a <=( a123548a  and  a123545a );
 a123552a <=( (not A200)  and  (not A199) );
 a123555a <=( (not A203)  and  A202 );
 a123556a <=( a123555a  and  a123552a );
 a123557a <=( a123556a  and  a123549a );
 a123560a <=( A266  and  (not A265) );
 a123563a <=( A269  and  (not A268) );
 a123564a <=( a123563a  and  a123560a );
 a123567a <=( A299  and  A298 );
 a123570a <=( A302  and  (not A300) );
 a123571a <=( a123570a  and  a123567a );
 a123572a <=( a123571a  and  a123564a );
 a123575a <=( A168  and  A170 );
 a123578a <=( A166  and  (not A167) );
 a123579a <=( a123578a  and  a123575a );
 a123582a <=( (not A200)  and  (not A199) );
 a123585a <=( (not A203)  and  A202 );
 a123586a <=( a123585a  and  a123582a );
 a123587a <=( a123586a  and  a123579a );
 a123590a <=( A266  and  (not A265) );
 a123593a <=( A269  and  (not A268) );
 a123594a <=( a123593a  and  a123590a );
 a123597a <=( (not A299)  and  A298 );
 a123600a <=( A301  and  (not A300) );
 a123601a <=( a123600a  and  a123597a );
 a123602a <=( a123601a  and  a123594a );
 a123605a <=( A168  and  A170 );
 a123608a <=( A166  and  (not A167) );
 a123609a <=( a123608a  and  a123605a );
 a123612a <=( (not A200)  and  (not A199) );
 a123615a <=( (not A203)  and  A202 );
 a123616a <=( a123615a  and  a123612a );
 a123617a <=( a123616a  and  a123609a );
 a123620a <=( A266  and  (not A265) );
 a123623a <=( A269  and  (not A268) );
 a123624a <=( a123623a  and  a123620a );
 a123627a <=( (not A299)  and  A298 );
 a123630a <=( (not A302)  and  (not A300) );
 a123631a <=( a123630a  and  a123627a );
 a123632a <=( a123631a  and  a123624a );
 a123635a <=( A168  and  A170 );
 a123638a <=( A166  and  (not A167) );
 a123639a <=( a123638a  and  a123635a );
 a123642a <=( (not A200)  and  (not A199) );
 a123645a <=( (not A203)  and  A202 );
 a123646a <=( a123645a  and  a123642a );
 a123647a <=( a123646a  and  a123639a );
 a123650a <=( A266  and  (not A265) );
 a123653a <=( A269  and  (not A268) );
 a123654a <=( a123653a  and  a123650a );
 a123657a <=( A299  and  (not A298) );
 a123660a <=( A301  and  (not A300) );
 a123661a <=( a123660a  and  a123657a );
 a123662a <=( a123661a  and  a123654a );
 a123665a <=( A168  and  A170 );
 a123668a <=( A166  and  (not A167) );
 a123669a <=( a123668a  and  a123665a );
 a123672a <=( (not A200)  and  (not A199) );
 a123675a <=( (not A203)  and  A202 );
 a123676a <=( a123675a  and  a123672a );
 a123677a <=( a123676a  and  a123669a );
 a123680a <=( A266  and  (not A265) );
 a123683a <=( A269  and  (not A268) );
 a123684a <=( a123683a  and  a123680a );
 a123687a <=( A299  and  (not A298) );
 a123690a <=( (not A302)  and  (not A300) );
 a123691a <=( a123690a  and  a123687a );
 a123692a <=( a123691a  and  a123684a );
 a123695a <=( A168  and  A170 );
 a123698a <=( A166  and  (not A167) );
 a123699a <=( a123698a  and  a123695a );
 a123702a <=( (not A200)  and  (not A199) );
 a123705a <=( (not A203)  and  A202 );
 a123706a <=( a123705a  and  a123702a );
 a123707a <=( a123706a  and  a123699a );
 a123710a <=( (not A266)  and  A265 );
 a123713a <=( A269  and  (not A268) );
 a123714a <=( a123713a  and  a123710a );
 a123717a <=( A299  and  A298 );
 a123720a <=( (not A301)  and  (not A300) );
 a123721a <=( a123720a  and  a123717a );
 a123722a <=( a123721a  and  a123714a );
 a123725a <=( A168  and  A170 );
 a123728a <=( A166  and  (not A167) );
 a123729a <=( a123728a  and  a123725a );
 a123732a <=( (not A200)  and  (not A199) );
 a123735a <=( (not A203)  and  A202 );
 a123736a <=( a123735a  and  a123732a );
 a123737a <=( a123736a  and  a123729a );
 a123740a <=( (not A266)  and  A265 );
 a123743a <=( A269  and  (not A268) );
 a123744a <=( a123743a  and  a123740a );
 a123747a <=( A299  and  A298 );
 a123750a <=( A302  and  (not A300) );
 a123751a <=( a123750a  and  a123747a );
 a123752a <=( a123751a  and  a123744a );
 a123755a <=( A168  and  A170 );
 a123758a <=( A166  and  (not A167) );
 a123759a <=( a123758a  and  a123755a );
 a123762a <=( (not A200)  and  (not A199) );
 a123765a <=( (not A203)  and  A202 );
 a123766a <=( a123765a  and  a123762a );
 a123767a <=( a123766a  and  a123759a );
 a123770a <=( (not A266)  and  A265 );
 a123773a <=( A269  and  (not A268) );
 a123774a <=( a123773a  and  a123770a );
 a123777a <=( (not A299)  and  A298 );
 a123780a <=( A301  and  (not A300) );
 a123781a <=( a123780a  and  a123777a );
 a123782a <=( a123781a  and  a123774a );
 a123785a <=( A168  and  A170 );
 a123788a <=( A166  and  (not A167) );
 a123789a <=( a123788a  and  a123785a );
 a123792a <=( (not A200)  and  (not A199) );
 a123795a <=( (not A203)  and  A202 );
 a123796a <=( a123795a  and  a123792a );
 a123797a <=( a123796a  and  a123789a );
 a123800a <=( (not A266)  and  A265 );
 a123803a <=( A269  and  (not A268) );
 a123804a <=( a123803a  and  a123800a );
 a123807a <=( (not A299)  and  A298 );
 a123810a <=( (not A302)  and  (not A300) );
 a123811a <=( a123810a  and  a123807a );
 a123812a <=( a123811a  and  a123804a );
 a123815a <=( A168  and  A170 );
 a123818a <=( A166  and  (not A167) );
 a123819a <=( a123818a  and  a123815a );
 a123822a <=( (not A200)  and  (not A199) );
 a123825a <=( (not A203)  and  A202 );
 a123826a <=( a123825a  and  a123822a );
 a123827a <=( a123826a  and  a123819a );
 a123830a <=( (not A266)  and  A265 );
 a123833a <=( A269  and  (not A268) );
 a123834a <=( a123833a  and  a123830a );
 a123837a <=( A299  and  (not A298) );
 a123840a <=( A301  and  (not A300) );
 a123841a <=( a123840a  and  a123837a );
 a123842a <=( a123841a  and  a123834a );
 a123845a <=( A168  and  A170 );
 a123848a <=( A166  and  (not A167) );
 a123849a <=( a123848a  and  a123845a );
 a123852a <=( (not A200)  and  (not A199) );
 a123855a <=( (not A203)  and  A202 );
 a123856a <=( a123855a  and  a123852a );
 a123857a <=( a123856a  and  a123849a );
 a123860a <=( (not A266)  and  A265 );
 a123863a <=( A269  and  (not A268) );
 a123864a <=( a123863a  and  a123860a );
 a123867a <=( A299  and  (not A298) );
 a123870a <=( (not A302)  and  (not A300) );
 a123871a <=( a123870a  and  a123867a );
 a123872a <=( a123871a  and  a123864a );
 a123875a <=( A168  and  A170 );
 a123878a <=( A166  and  (not A167) );
 a123879a <=( a123878a  and  a123875a );
 a123882a <=( (not A200)  and  (not A199) );
 a123885a <=( (not A203)  and  A202 );
 a123886a <=( a123885a  and  a123882a );
 a123887a <=( a123886a  and  a123879a );
 a123890a <=( (not A266)  and  (not A265) );
 a123893a <=( (not A269)  and  A268 );
 a123894a <=( a123893a  and  a123890a );
 a123897a <=( A299  and  A298 );
 a123900a <=( (not A301)  and  (not A300) );
 a123901a <=( a123900a  and  a123897a );
 a123902a <=( a123901a  and  a123894a );
 a123905a <=( A168  and  A170 );
 a123908a <=( A166  and  (not A167) );
 a123909a <=( a123908a  and  a123905a );
 a123912a <=( (not A200)  and  (not A199) );
 a123915a <=( (not A203)  and  A202 );
 a123916a <=( a123915a  and  a123912a );
 a123917a <=( a123916a  and  a123909a );
 a123920a <=( (not A266)  and  (not A265) );
 a123923a <=( (not A269)  and  A268 );
 a123924a <=( a123923a  and  a123920a );
 a123927a <=( A299  and  A298 );
 a123930a <=( A302  and  (not A300) );
 a123931a <=( a123930a  and  a123927a );
 a123932a <=( a123931a  and  a123924a );
 a123935a <=( A168  and  A170 );
 a123938a <=( A166  and  (not A167) );
 a123939a <=( a123938a  and  a123935a );
 a123942a <=( (not A200)  and  (not A199) );
 a123945a <=( (not A203)  and  A202 );
 a123946a <=( a123945a  and  a123942a );
 a123947a <=( a123946a  and  a123939a );
 a123950a <=( (not A266)  and  (not A265) );
 a123953a <=( (not A269)  and  A268 );
 a123954a <=( a123953a  and  a123950a );
 a123957a <=( (not A299)  and  A298 );
 a123960a <=( A301  and  (not A300) );
 a123961a <=( a123960a  and  a123957a );
 a123962a <=( a123961a  and  a123954a );
 a123965a <=( A168  and  A170 );
 a123968a <=( A166  and  (not A167) );
 a123969a <=( a123968a  and  a123965a );
 a123972a <=( (not A200)  and  (not A199) );
 a123975a <=( (not A203)  and  A202 );
 a123976a <=( a123975a  and  a123972a );
 a123977a <=( a123976a  and  a123969a );
 a123980a <=( (not A266)  and  (not A265) );
 a123983a <=( (not A269)  and  A268 );
 a123984a <=( a123983a  and  a123980a );
 a123987a <=( (not A299)  and  A298 );
 a123990a <=( (not A302)  and  (not A300) );
 a123991a <=( a123990a  and  a123987a );
 a123992a <=( a123991a  and  a123984a );
 a123995a <=( A168  and  A170 );
 a123998a <=( A166  and  (not A167) );
 a123999a <=( a123998a  and  a123995a );
 a124002a <=( (not A200)  and  (not A199) );
 a124005a <=( (not A203)  and  A202 );
 a124006a <=( a124005a  and  a124002a );
 a124007a <=( a124006a  and  a123999a );
 a124010a <=( (not A266)  and  (not A265) );
 a124013a <=( (not A269)  and  A268 );
 a124014a <=( a124013a  and  a124010a );
 a124017a <=( A299  and  (not A298) );
 a124020a <=( A301  and  (not A300) );
 a124021a <=( a124020a  and  a124017a );
 a124022a <=( a124021a  and  a124014a );
 a124025a <=( A168  and  A170 );
 a124028a <=( A166  and  (not A167) );
 a124029a <=( a124028a  and  a124025a );
 a124032a <=( (not A200)  and  (not A199) );
 a124035a <=( (not A203)  and  A202 );
 a124036a <=( a124035a  and  a124032a );
 a124037a <=( a124036a  and  a124029a );
 a124040a <=( (not A266)  and  (not A265) );
 a124043a <=( (not A269)  and  A268 );
 a124044a <=( a124043a  and  a124040a );
 a124047a <=( A299  and  (not A298) );
 a124050a <=( (not A302)  and  (not A300) );
 a124051a <=( a124050a  and  a124047a );
 a124052a <=( a124051a  and  a124044a );
 a124055a <=( A168  and  A169 );
 a124058a <=( A166  and  (not A167) );
 a124059a <=( a124058a  and  a124055a );
 a124062a <=( A200  and  A199 );
 a124065a <=( (not A203)  and  A202 );
 a124066a <=( a124065a  and  a124062a );
 a124067a <=( a124066a  and  a124059a );
 a124070a <=( A266  and  A265 );
 a124073a <=( (not A269)  and  A268 );
 a124074a <=( a124073a  and  a124070a );
 a124077a <=( A299  and  A298 );
 a124080a <=( (not A301)  and  (not A300) );
 a124081a <=( a124080a  and  a124077a );
 a124082a <=( a124081a  and  a124074a );
 a124085a <=( A168  and  A169 );
 a124088a <=( A166  and  (not A167) );
 a124089a <=( a124088a  and  a124085a );
 a124092a <=( A200  and  A199 );
 a124095a <=( (not A203)  and  A202 );
 a124096a <=( a124095a  and  a124092a );
 a124097a <=( a124096a  and  a124089a );
 a124100a <=( A266  and  A265 );
 a124103a <=( (not A269)  and  A268 );
 a124104a <=( a124103a  and  a124100a );
 a124107a <=( A299  and  A298 );
 a124110a <=( A302  and  (not A300) );
 a124111a <=( a124110a  and  a124107a );
 a124112a <=( a124111a  and  a124104a );
 a124115a <=( A168  and  A169 );
 a124118a <=( A166  and  (not A167) );
 a124119a <=( a124118a  and  a124115a );
 a124122a <=( A200  and  A199 );
 a124125a <=( (not A203)  and  A202 );
 a124126a <=( a124125a  and  a124122a );
 a124127a <=( a124126a  and  a124119a );
 a124130a <=( A266  and  A265 );
 a124133a <=( (not A269)  and  A268 );
 a124134a <=( a124133a  and  a124130a );
 a124137a <=( (not A299)  and  A298 );
 a124140a <=( A301  and  (not A300) );
 a124141a <=( a124140a  and  a124137a );
 a124142a <=( a124141a  and  a124134a );
 a124145a <=( A168  and  A169 );
 a124148a <=( A166  and  (not A167) );
 a124149a <=( a124148a  and  a124145a );
 a124152a <=( A200  and  A199 );
 a124155a <=( (not A203)  and  A202 );
 a124156a <=( a124155a  and  a124152a );
 a124157a <=( a124156a  and  a124149a );
 a124160a <=( A266  and  A265 );
 a124163a <=( (not A269)  and  A268 );
 a124164a <=( a124163a  and  a124160a );
 a124167a <=( (not A299)  and  A298 );
 a124170a <=( (not A302)  and  (not A300) );
 a124171a <=( a124170a  and  a124167a );
 a124172a <=( a124171a  and  a124164a );
 a124175a <=( A168  and  A169 );
 a124178a <=( A166  and  (not A167) );
 a124179a <=( a124178a  and  a124175a );
 a124182a <=( A200  and  A199 );
 a124185a <=( (not A203)  and  A202 );
 a124186a <=( a124185a  and  a124182a );
 a124187a <=( a124186a  and  a124179a );
 a124190a <=( A266  and  A265 );
 a124193a <=( (not A269)  and  A268 );
 a124194a <=( a124193a  and  a124190a );
 a124197a <=( A299  and  (not A298) );
 a124200a <=( A301  and  (not A300) );
 a124201a <=( a124200a  and  a124197a );
 a124202a <=( a124201a  and  a124194a );
 a124205a <=( A168  and  A169 );
 a124208a <=( A166  and  (not A167) );
 a124209a <=( a124208a  and  a124205a );
 a124212a <=( A200  and  A199 );
 a124215a <=( (not A203)  and  A202 );
 a124216a <=( a124215a  and  a124212a );
 a124217a <=( a124216a  and  a124209a );
 a124220a <=( A266  and  A265 );
 a124223a <=( (not A269)  and  A268 );
 a124224a <=( a124223a  and  a124220a );
 a124227a <=( A299  and  (not A298) );
 a124230a <=( (not A302)  and  (not A300) );
 a124231a <=( a124230a  and  a124227a );
 a124232a <=( a124231a  and  a124224a );
 a124235a <=( A168  and  A169 );
 a124238a <=( A166  and  (not A167) );
 a124239a <=( a124238a  and  a124235a );
 a124242a <=( A200  and  A199 );
 a124245a <=( (not A203)  and  A202 );
 a124246a <=( a124245a  and  a124242a );
 a124247a <=( a124246a  and  a124239a );
 a124250a <=( A266  and  (not A265) );
 a124253a <=( A269  and  (not A268) );
 a124254a <=( a124253a  and  a124250a );
 a124257a <=( A299  and  A298 );
 a124260a <=( (not A301)  and  (not A300) );
 a124261a <=( a124260a  and  a124257a );
 a124262a <=( a124261a  and  a124254a );
 a124265a <=( A168  and  A169 );
 a124268a <=( A166  and  (not A167) );
 a124269a <=( a124268a  and  a124265a );
 a124272a <=( A200  and  A199 );
 a124275a <=( (not A203)  and  A202 );
 a124276a <=( a124275a  and  a124272a );
 a124277a <=( a124276a  and  a124269a );
 a124280a <=( A266  and  (not A265) );
 a124283a <=( A269  and  (not A268) );
 a124284a <=( a124283a  and  a124280a );
 a124287a <=( A299  and  A298 );
 a124290a <=( A302  and  (not A300) );
 a124291a <=( a124290a  and  a124287a );
 a124292a <=( a124291a  and  a124284a );
 a124295a <=( A168  and  A169 );
 a124298a <=( A166  and  (not A167) );
 a124299a <=( a124298a  and  a124295a );
 a124302a <=( A200  and  A199 );
 a124305a <=( (not A203)  and  A202 );
 a124306a <=( a124305a  and  a124302a );
 a124307a <=( a124306a  and  a124299a );
 a124310a <=( A266  and  (not A265) );
 a124313a <=( A269  and  (not A268) );
 a124314a <=( a124313a  and  a124310a );
 a124317a <=( (not A299)  and  A298 );
 a124320a <=( A301  and  (not A300) );
 a124321a <=( a124320a  and  a124317a );
 a124322a <=( a124321a  and  a124314a );
 a124325a <=( A168  and  A169 );
 a124328a <=( A166  and  (not A167) );
 a124329a <=( a124328a  and  a124325a );
 a124332a <=( A200  and  A199 );
 a124335a <=( (not A203)  and  A202 );
 a124336a <=( a124335a  and  a124332a );
 a124337a <=( a124336a  and  a124329a );
 a124340a <=( A266  and  (not A265) );
 a124343a <=( A269  and  (not A268) );
 a124344a <=( a124343a  and  a124340a );
 a124347a <=( (not A299)  and  A298 );
 a124350a <=( (not A302)  and  (not A300) );
 a124351a <=( a124350a  and  a124347a );
 a124352a <=( a124351a  and  a124344a );
 a124355a <=( A168  and  A169 );
 a124358a <=( A166  and  (not A167) );
 a124359a <=( a124358a  and  a124355a );
 a124362a <=( A200  and  A199 );
 a124365a <=( (not A203)  and  A202 );
 a124366a <=( a124365a  and  a124362a );
 a124367a <=( a124366a  and  a124359a );
 a124370a <=( A266  and  (not A265) );
 a124373a <=( A269  and  (not A268) );
 a124374a <=( a124373a  and  a124370a );
 a124377a <=( A299  and  (not A298) );
 a124380a <=( A301  and  (not A300) );
 a124381a <=( a124380a  and  a124377a );
 a124382a <=( a124381a  and  a124374a );
 a124385a <=( A168  and  A169 );
 a124388a <=( A166  and  (not A167) );
 a124389a <=( a124388a  and  a124385a );
 a124392a <=( A200  and  A199 );
 a124395a <=( (not A203)  and  A202 );
 a124396a <=( a124395a  and  a124392a );
 a124397a <=( a124396a  and  a124389a );
 a124400a <=( A266  and  (not A265) );
 a124403a <=( A269  and  (not A268) );
 a124404a <=( a124403a  and  a124400a );
 a124407a <=( A299  and  (not A298) );
 a124410a <=( (not A302)  and  (not A300) );
 a124411a <=( a124410a  and  a124407a );
 a124412a <=( a124411a  and  a124404a );
 a124415a <=( A168  and  A169 );
 a124418a <=( A166  and  (not A167) );
 a124419a <=( a124418a  and  a124415a );
 a124422a <=( A200  and  A199 );
 a124425a <=( (not A203)  and  A202 );
 a124426a <=( a124425a  and  a124422a );
 a124427a <=( a124426a  and  a124419a );
 a124430a <=( (not A266)  and  A265 );
 a124433a <=( A269  and  (not A268) );
 a124434a <=( a124433a  and  a124430a );
 a124437a <=( A299  and  A298 );
 a124440a <=( (not A301)  and  (not A300) );
 a124441a <=( a124440a  and  a124437a );
 a124442a <=( a124441a  and  a124434a );
 a124445a <=( A168  and  A169 );
 a124448a <=( A166  and  (not A167) );
 a124449a <=( a124448a  and  a124445a );
 a124452a <=( A200  and  A199 );
 a124455a <=( (not A203)  and  A202 );
 a124456a <=( a124455a  and  a124452a );
 a124457a <=( a124456a  and  a124449a );
 a124460a <=( (not A266)  and  A265 );
 a124463a <=( A269  and  (not A268) );
 a124464a <=( a124463a  and  a124460a );
 a124467a <=( A299  and  A298 );
 a124470a <=( A302  and  (not A300) );
 a124471a <=( a124470a  and  a124467a );
 a124472a <=( a124471a  and  a124464a );
 a124475a <=( A168  and  A169 );
 a124478a <=( A166  and  (not A167) );
 a124479a <=( a124478a  and  a124475a );
 a124482a <=( A200  and  A199 );
 a124485a <=( (not A203)  and  A202 );
 a124486a <=( a124485a  and  a124482a );
 a124487a <=( a124486a  and  a124479a );
 a124490a <=( (not A266)  and  A265 );
 a124493a <=( A269  and  (not A268) );
 a124494a <=( a124493a  and  a124490a );
 a124497a <=( (not A299)  and  A298 );
 a124500a <=( A301  and  (not A300) );
 a124501a <=( a124500a  and  a124497a );
 a124502a <=( a124501a  and  a124494a );
 a124505a <=( A168  and  A169 );
 a124508a <=( A166  and  (not A167) );
 a124509a <=( a124508a  and  a124505a );
 a124512a <=( A200  and  A199 );
 a124515a <=( (not A203)  and  A202 );
 a124516a <=( a124515a  and  a124512a );
 a124517a <=( a124516a  and  a124509a );
 a124520a <=( (not A266)  and  A265 );
 a124523a <=( A269  and  (not A268) );
 a124524a <=( a124523a  and  a124520a );
 a124527a <=( (not A299)  and  A298 );
 a124530a <=( (not A302)  and  (not A300) );
 a124531a <=( a124530a  and  a124527a );
 a124532a <=( a124531a  and  a124524a );
 a124535a <=( A168  and  A169 );
 a124538a <=( A166  and  (not A167) );
 a124539a <=( a124538a  and  a124535a );
 a124542a <=( A200  and  A199 );
 a124545a <=( (not A203)  and  A202 );
 a124546a <=( a124545a  and  a124542a );
 a124547a <=( a124546a  and  a124539a );
 a124550a <=( (not A266)  and  A265 );
 a124553a <=( A269  and  (not A268) );
 a124554a <=( a124553a  and  a124550a );
 a124557a <=( A299  and  (not A298) );
 a124560a <=( A301  and  (not A300) );
 a124561a <=( a124560a  and  a124557a );
 a124562a <=( a124561a  and  a124554a );
 a124565a <=( A168  and  A169 );
 a124568a <=( A166  and  (not A167) );
 a124569a <=( a124568a  and  a124565a );
 a124572a <=( A200  and  A199 );
 a124575a <=( (not A203)  and  A202 );
 a124576a <=( a124575a  and  a124572a );
 a124577a <=( a124576a  and  a124569a );
 a124580a <=( (not A266)  and  A265 );
 a124583a <=( A269  and  (not A268) );
 a124584a <=( a124583a  and  a124580a );
 a124587a <=( A299  and  (not A298) );
 a124590a <=( (not A302)  and  (not A300) );
 a124591a <=( a124590a  and  a124587a );
 a124592a <=( a124591a  and  a124584a );
 a124595a <=( A168  and  A169 );
 a124598a <=( A166  and  (not A167) );
 a124599a <=( a124598a  and  a124595a );
 a124602a <=( A200  and  A199 );
 a124605a <=( (not A203)  and  A202 );
 a124606a <=( a124605a  and  a124602a );
 a124607a <=( a124606a  and  a124599a );
 a124610a <=( (not A266)  and  (not A265) );
 a124613a <=( (not A269)  and  A268 );
 a124614a <=( a124613a  and  a124610a );
 a124617a <=( A299  and  A298 );
 a124620a <=( (not A301)  and  (not A300) );
 a124621a <=( a124620a  and  a124617a );
 a124622a <=( a124621a  and  a124614a );
 a124625a <=( A168  and  A169 );
 a124628a <=( A166  and  (not A167) );
 a124629a <=( a124628a  and  a124625a );
 a124632a <=( A200  and  A199 );
 a124635a <=( (not A203)  and  A202 );
 a124636a <=( a124635a  and  a124632a );
 a124637a <=( a124636a  and  a124629a );
 a124640a <=( (not A266)  and  (not A265) );
 a124643a <=( (not A269)  and  A268 );
 a124644a <=( a124643a  and  a124640a );
 a124647a <=( A299  and  A298 );
 a124650a <=( A302  and  (not A300) );
 a124651a <=( a124650a  and  a124647a );
 a124652a <=( a124651a  and  a124644a );
 a124655a <=( A168  and  A169 );
 a124658a <=( A166  and  (not A167) );
 a124659a <=( a124658a  and  a124655a );
 a124662a <=( A200  and  A199 );
 a124665a <=( (not A203)  and  A202 );
 a124666a <=( a124665a  and  a124662a );
 a124667a <=( a124666a  and  a124659a );
 a124670a <=( (not A266)  and  (not A265) );
 a124673a <=( (not A269)  and  A268 );
 a124674a <=( a124673a  and  a124670a );
 a124677a <=( (not A299)  and  A298 );
 a124680a <=( A301  and  (not A300) );
 a124681a <=( a124680a  and  a124677a );
 a124682a <=( a124681a  and  a124674a );
 a124685a <=( A168  and  A169 );
 a124688a <=( A166  and  (not A167) );
 a124689a <=( a124688a  and  a124685a );
 a124692a <=( A200  and  A199 );
 a124695a <=( (not A203)  and  A202 );
 a124696a <=( a124695a  and  a124692a );
 a124697a <=( a124696a  and  a124689a );
 a124700a <=( (not A266)  and  (not A265) );
 a124703a <=( (not A269)  and  A268 );
 a124704a <=( a124703a  and  a124700a );
 a124707a <=( (not A299)  and  A298 );
 a124710a <=( (not A302)  and  (not A300) );
 a124711a <=( a124710a  and  a124707a );
 a124712a <=( a124711a  and  a124704a );
 a124715a <=( A168  and  A169 );
 a124718a <=( A166  and  (not A167) );
 a124719a <=( a124718a  and  a124715a );
 a124722a <=( A200  and  A199 );
 a124725a <=( (not A203)  and  A202 );
 a124726a <=( a124725a  and  a124722a );
 a124727a <=( a124726a  and  a124719a );
 a124730a <=( (not A266)  and  (not A265) );
 a124733a <=( (not A269)  and  A268 );
 a124734a <=( a124733a  and  a124730a );
 a124737a <=( A299  and  (not A298) );
 a124740a <=( A301  and  (not A300) );
 a124741a <=( a124740a  and  a124737a );
 a124742a <=( a124741a  and  a124734a );
 a124745a <=( A168  and  A169 );
 a124748a <=( A166  and  (not A167) );
 a124749a <=( a124748a  and  a124745a );
 a124752a <=( A200  and  A199 );
 a124755a <=( (not A203)  and  A202 );
 a124756a <=( a124755a  and  a124752a );
 a124757a <=( a124756a  and  a124749a );
 a124760a <=( (not A266)  and  (not A265) );
 a124763a <=( (not A269)  and  A268 );
 a124764a <=( a124763a  and  a124760a );
 a124767a <=( A299  and  (not A298) );
 a124770a <=( (not A302)  and  (not A300) );
 a124771a <=( a124770a  and  a124767a );
 a124772a <=( a124771a  and  a124764a );
 a124775a <=( A168  and  A169 );
 a124778a <=( A166  and  (not A167) );
 a124779a <=( a124778a  and  a124775a );
 a124782a <=( A200  and  A199 );
 a124785a <=( (not A202)  and  (not A201) );
 a124786a <=( a124785a  and  a124782a );
 a124787a <=( a124786a  and  a124779a );
 a124790a <=( A266  and  A265 );
 a124793a <=( (not A268)  and  (not A267) );
 a124794a <=( a124793a  and  a124790a );
 a124797a <=( A299  and  A298 );
 a124800a <=( (not A302)  and  A301 );
 a124801a <=( a124800a  and  a124797a );
 a124802a <=( a124801a  and  a124794a );
 a124805a <=( A168  and  A169 );
 a124808a <=( A166  and  (not A167) );
 a124809a <=( a124808a  and  a124805a );
 a124812a <=( A200  and  A199 );
 a124815a <=( (not A202)  and  (not A201) );
 a124816a <=( a124815a  and  a124812a );
 a124817a <=( a124816a  and  a124809a );
 a124820a <=( A266  and  A265 );
 a124823a <=( (not A268)  and  (not A267) );
 a124824a <=( a124823a  and  a124820a );
 a124827a <=( (not A299)  and  A298 );
 a124830a <=( A302  and  (not A301) );
 a124831a <=( a124830a  and  a124827a );
 a124832a <=( a124831a  and  a124824a );
 a124835a <=( A168  and  A169 );
 a124838a <=( A166  and  (not A167) );
 a124839a <=( a124838a  and  a124835a );
 a124842a <=( A200  and  A199 );
 a124845a <=( (not A202)  and  (not A201) );
 a124846a <=( a124845a  and  a124842a );
 a124847a <=( a124846a  and  a124839a );
 a124850a <=( A266  and  A265 );
 a124853a <=( (not A268)  and  (not A267) );
 a124854a <=( a124853a  and  a124850a );
 a124857a <=( A299  and  (not A298) );
 a124860a <=( A302  and  (not A301) );
 a124861a <=( a124860a  and  a124857a );
 a124862a <=( a124861a  and  a124854a );
 a124865a <=( A168  and  A169 );
 a124868a <=( A166  and  (not A167) );
 a124869a <=( a124868a  and  a124865a );
 a124872a <=( A200  and  A199 );
 a124875a <=( (not A202)  and  (not A201) );
 a124876a <=( a124875a  and  a124872a );
 a124877a <=( a124876a  and  a124869a );
 a124880a <=( A266  and  A265 );
 a124883a <=( (not A268)  and  (not A267) );
 a124884a <=( a124883a  and  a124880a );
 a124887a <=( (not A299)  and  (not A298) );
 a124890a <=( (not A302)  and  A301 );
 a124891a <=( a124890a  and  a124887a );
 a124892a <=( a124891a  and  a124884a );
 a124895a <=( A168  and  A169 );
 a124898a <=( A166  and  (not A167) );
 a124899a <=( a124898a  and  a124895a );
 a124902a <=( A200  and  A199 );
 a124905a <=( (not A202)  and  (not A201) );
 a124906a <=( a124905a  and  a124902a );
 a124907a <=( a124906a  and  a124899a );
 a124910a <=( A266  and  A265 );
 a124913a <=( A269  and  (not A267) );
 a124914a <=( a124913a  and  a124910a );
 a124917a <=( A299  and  A298 );
 a124920a <=( (not A302)  and  A301 );
 a124921a <=( a124920a  and  a124917a );
 a124922a <=( a124921a  and  a124914a );
 a124925a <=( A168  and  A169 );
 a124928a <=( A166  and  (not A167) );
 a124929a <=( a124928a  and  a124925a );
 a124932a <=( A200  and  A199 );
 a124935a <=( (not A202)  and  (not A201) );
 a124936a <=( a124935a  and  a124932a );
 a124937a <=( a124936a  and  a124929a );
 a124940a <=( A266  and  A265 );
 a124943a <=( A269  and  (not A267) );
 a124944a <=( a124943a  and  a124940a );
 a124947a <=( (not A299)  and  A298 );
 a124950a <=( A302  and  (not A301) );
 a124951a <=( a124950a  and  a124947a );
 a124952a <=( a124951a  and  a124944a );
 a124955a <=( A168  and  A169 );
 a124958a <=( A166  and  (not A167) );
 a124959a <=( a124958a  and  a124955a );
 a124962a <=( A200  and  A199 );
 a124965a <=( (not A202)  and  (not A201) );
 a124966a <=( a124965a  and  a124962a );
 a124967a <=( a124966a  and  a124959a );
 a124970a <=( A266  and  A265 );
 a124973a <=( A269  and  (not A267) );
 a124974a <=( a124973a  and  a124970a );
 a124977a <=( A299  and  (not A298) );
 a124980a <=( A302  and  (not A301) );
 a124981a <=( a124980a  and  a124977a );
 a124982a <=( a124981a  and  a124974a );
 a124985a <=( A168  and  A169 );
 a124988a <=( A166  and  (not A167) );
 a124989a <=( a124988a  and  a124985a );
 a124992a <=( A200  and  A199 );
 a124995a <=( (not A202)  and  (not A201) );
 a124996a <=( a124995a  and  a124992a );
 a124997a <=( a124996a  and  a124989a );
 a125000a <=( A266  and  A265 );
 a125003a <=( A269  and  (not A267) );
 a125004a <=( a125003a  and  a125000a );
 a125007a <=( (not A299)  and  (not A298) );
 a125010a <=( (not A302)  and  A301 );
 a125011a <=( a125010a  and  a125007a );
 a125012a <=( a125011a  and  a125004a );
 a125015a <=( A168  and  A169 );
 a125018a <=( A166  and  (not A167) );
 a125019a <=( a125018a  and  a125015a );
 a125022a <=( A200  and  A199 );
 a125025a <=( (not A202)  and  (not A201) );
 a125026a <=( a125025a  and  a125022a );
 a125027a <=( a125026a  and  a125019a );
 a125030a <=( A266  and  (not A265) );
 a125033a <=( A268  and  (not A267) );
 a125034a <=( a125033a  and  a125030a );
 a125037a <=( A299  and  A298 );
 a125040a <=( (not A302)  and  A301 );
 a125041a <=( a125040a  and  a125037a );
 a125042a <=( a125041a  and  a125034a );
 a125045a <=( A168  and  A169 );
 a125048a <=( A166  and  (not A167) );
 a125049a <=( a125048a  and  a125045a );
 a125052a <=( A200  and  A199 );
 a125055a <=( (not A202)  and  (not A201) );
 a125056a <=( a125055a  and  a125052a );
 a125057a <=( a125056a  and  a125049a );
 a125060a <=( A266  and  (not A265) );
 a125063a <=( A268  and  (not A267) );
 a125064a <=( a125063a  and  a125060a );
 a125067a <=( (not A299)  and  A298 );
 a125070a <=( A302  and  (not A301) );
 a125071a <=( a125070a  and  a125067a );
 a125072a <=( a125071a  and  a125064a );
 a125075a <=( A168  and  A169 );
 a125078a <=( A166  and  (not A167) );
 a125079a <=( a125078a  and  a125075a );
 a125082a <=( A200  and  A199 );
 a125085a <=( (not A202)  and  (not A201) );
 a125086a <=( a125085a  and  a125082a );
 a125087a <=( a125086a  and  a125079a );
 a125090a <=( A266  and  (not A265) );
 a125093a <=( A268  and  (not A267) );
 a125094a <=( a125093a  and  a125090a );
 a125097a <=( A299  and  (not A298) );
 a125100a <=( A302  and  (not A301) );
 a125101a <=( a125100a  and  a125097a );
 a125102a <=( a125101a  and  a125094a );
 a125105a <=( A168  and  A169 );
 a125108a <=( A166  and  (not A167) );
 a125109a <=( a125108a  and  a125105a );
 a125112a <=( A200  and  A199 );
 a125115a <=( (not A202)  and  (not A201) );
 a125116a <=( a125115a  and  a125112a );
 a125117a <=( a125116a  and  a125109a );
 a125120a <=( A266  and  (not A265) );
 a125123a <=( A268  and  (not A267) );
 a125124a <=( a125123a  and  a125120a );
 a125127a <=( (not A299)  and  (not A298) );
 a125130a <=( (not A302)  and  A301 );
 a125131a <=( a125130a  and  a125127a );
 a125132a <=( a125131a  and  a125124a );
 a125135a <=( A168  and  A169 );
 a125138a <=( A166  and  (not A167) );
 a125139a <=( a125138a  and  a125135a );
 a125142a <=( A200  and  A199 );
 a125145a <=( (not A202)  and  (not A201) );
 a125146a <=( a125145a  and  a125142a );
 a125147a <=( a125146a  and  a125139a );
 a125150a <=( A266  and  (not A265) );
 a125153a <=( (not A269)  and  (not A267) );
 a125154a <=( a125153a  and  a125150a );
 a125157a <=( A299  and  A298 );
 a125160a <=( (not A302)  and  A301 );
 a125161a <=( a125160a  and  a125157a );
 a125162a <=( a125161a  and  a125154a );
 a125165a <=( A168  and  A169 );
 a125168a <=( A166  and  (not A167) );
 a125169a <=( a125168a  and  a125165a );
 a125172a <=( A200  and  A199 );
 a125175a <=( (not A202)  and  (not A201) );
 a125176a <=( a125175a  and  a125172a );
 a125177a <=( a125176a  and  a125169a );
 a125180a <=( A266  and  (not A265) );
 a125183a <=( (not A269)  and  (not A267) );
 a125184a <=( a125183a  and  a125180a );
 a125187a <=( (not A299)  and  A298 );
 a125190a <=( A302  and  (not A301) );
 a125191a <=( a125190a  and  a125187a );
 a125192a <=( a125191a  and  a125184a );
 a125195a <=( A168  and  A169 );
 a125198a <=( A166  and  (not A167) );
 a125199a <=( a125198a  and  a125195a );
 a125202a <=( A200  and  A199 );
 a125205a <=( (not A202)  and  (not A201) );
 a125206a <=( a125205a  and  a125202a );
 a125207a <=( a125206a  and  a125199a );
 a125210a <=( A266  and  (not A265) );
 a125213a <=( (not A269)  and  (not A267) );
 a125214a <=( a125213a  and  a125210a );
 a125217a <=( A299  and  (not A298) );
 a125220a <=( A302  and  (not A301) );
 a125221a <=( a125220a  and  a125217a );
 a125222a <=( a125221a  and  a125214a );
 a125225a <=( A168  and  A169 );
 a125228a <=( A166  and  (not A167) );
 a125229a <=( a125228a  and  a125225a );
 a125232a <=( A200  and  A199 );
 a125235a <=( (not A202)  and  (not A201) );
 a125236a <=( a125235a  and  a125232a );
 a125237a <=( a125236a  and  a125229a );
 a125240a <=( A266  and  (not A265) );
 a125243a <=( (not A269)  and  (not A267) );
 a125244a <=( a125243a  and  a125240a );
 a125247a <=( (not A299)  and  (not A298) );
 a125250a <=( (not A302)  and  A301 );
 a125251a <=( a125250a  and  a125247a );
 a125252a <=( a125251a  and  a125244a );
 a125255a <=( A168  and  A169 );
 a125258a <=( A166  and  (not A167) );
 a125259a <=( a125258a  and  a125255a );
 a125262a <=( A200  and  A199 );
 a125265a <=( (not A202)  and  (not A201) );
 a125266a <=( a125265a  and  a125262a );
 a125267a <=( a125266a  and  a125259a );
 a125270a <=( (not A266)  and  A265 );
 a125273a <=( A268  and  (not A267) );
 a125274a <=( a125273a  and  a125270a );
 a125277a <=( A299  and  A298 );
 a125280a <=( (not A302)  and  A301 );
 a125281a <=( a125280a  and  a125277a );
 a125282a <=( a125281a  and  a125274a );
 a125285a <=( A168  and  A169 );
 a125288a <=( A166  and  (not A167) );
 a125289a <=( a125288a  and  a125285a );
 a125292a <=( A200  and  A199 );
 a125295a <=( (not A202)  and  (not A201) );
 a125296a <=( a125295a  and  a125292a );
 a125297a <=( a125296a  and  a125289a );
 a125300a <=( (not A266)  and  A265 );
 a125303a <=( A268  and  (not A267) );
 a125304a <=( a125303a  and  a125300a );
 a125307a <=( (not A299)  and  A298 );
 a125310a <=( A302  and  (not A301) );
 a125311a <=( a125310a  and  a125307a );
 a125312a <=( a125311a  and  a125304a );
 a125315a <=( A168  and  A169 );
 a125318a <=( A166  and  (not A167) );
 a125319a <=( a125318a  and  a125315a );
 a125322a <=( A200  and  A199 );
 a125325a <=( (not A202)  and  (not A201) );
 a125326a <=( a125325a  and  a125322a );
 a125327a <=( a125326a  and  a125319a );
 a125330a <=( (not A266)  and  A265 );
 a125333a <=( A268  and  (not A267) );
 a125334a <=( a125333a  and  a125330a );
 a125337a <=( A299  and  (not A298) );
 a125340a <=( A302  and  (not A301) );
 a125341a <=( a125340a  and  a125337a );
 a125342a <=( a125341a  and  a125334a );
 a125345a <=( A168  and  A169 );
 a125348a <=( A166  and  (not A167) );
 a125349a <=( a125348a  and  a125345a );
 a125352a <=( A200  and  A199 );
 a125355a <=( (not A202)  and  (not A201) );
 a125356a <=( a125355a  and  a125352a );
 a125357a <=( a125356a  and  a125349a );
 a125360a <=( (not A266)  and  A265 );
 a125363a <=( A268  and  (not A267) );
 a125364a <=( a125363a  and  a125360a );
 a125367a <=( (not A299)  and  (not A298) );
 a125370a <=( (not A302)  and  A301 );
 a125371a <=( a125370a  and  a125367a );
 a125372a <=( a125371a  and  a125364a );
 a125375a <=( A168  and  A169 );
 a125378a <=( A166  and  (not A167) );
 a125379a <=( a125378a  and  a125375a );
 a125382a <=( A200  and  A199 );
 a125385a <=( (not A202)  and  (not A201) );
 a125386a <=( a125385a  and  a125382a );
 a125387a <=( a125386a  and  a125379a );
 a125390a <=( (not A266)  and  A265 );
 a125393a <=( (not A269)  and  (not A267) );
 a125394a <=( a125393a  and  a125390a );
 a125397a <=( A299  and  A298 );
 a125400a <=( (not A302)  and  A301 );
 a125401a <=( a125400a  and  a125397a );
 a125402a <=( a125401a  and  a125394a );
 a125405a <=( A168  and  A169 );
 a125408a <=( A166  and  (not A167) );
 a125409a <=( a125408a  and  a125405a );
 a125412a <=( A200  and  A199 );
 a125415a <=( (not A202)  and  (not A201) );
 a125416a <=( a125415a  and  a125412a );
 a125417a <=( a125416a  and  a125409a );
 a125420a <=( (not A266)  and  A265 );
 a125423a <=( (not A269)  and  (not A267) );
 a125424a <=( a125423a  and  a125420a );
 a125427a <=( (not A299)  and  A298 );
 a125430a <=( A302  and  (not A301) );
 a125431a <=( a125430a  and  a125427a );
 a125432a <=( a125431a  and  a125424a );
 a125435a <=( A168  and  A169 );
 a125438a <=( A166  and  (not A167) );
 a125439a <=( a125438a  and  a125435a );
 a125442a <=( A200  and  A199 );
 a125445a <=( (not A202)  and  (not A201) );
 a125446a <=( a125445a  and  a125442a );
 a125447a <=( a125446a  and  a125439a );
 a125450a <=( (not A266)  and  A265 );
 a125453a <=( (not A269)  and  (not A267) );
 a125454a <=( a125453a  and  a125450a );
 a125457a <=( A299  and  (not A298) );
 a125460a <=( A302  and  (not A301) );
 a125461a <=( a125460a  and  a125457a );
 a125462a <=( a125461a  and  a125454a );
 a125465a <=( A168  and  A169 );
 a125468a <=( A166  and  (not A167) );
 a125469a <=( a125468a  and  a125465a );
 a125472a <=( A200  and  A199 );
 a125475a <=( (not A202)  and  (not A201) );
 a125476a <=( a125475a  and  a125472a );
 a125477a <=( a125476a  and  a125469a );
 a125480a <=( (not A266)  and  A265 );
 a125483a <=( (not A269)  and  (not A267) );
 a125484a <=( a125483a  and  a125480a );
 a125487a <=( (not A299)  and  (not A298) );
 a125490a <=( (not A302)  and  A301 );
 a125491a <=( a125490a  and  a125487a );
 a125492a <=( a125491a  and  a125484a );
 a125495a <=( A168  and  A169 );
 a125498a <=( A166  and  (not A167) );
 a125499a <=( a125498a  and  a125495a );
 a125502a <=( A200  and  A199 );
 a125505a <=( A203  and  (not A201) );
 a125506a <=( a125505a  and  a125502a );
 a125507a <=( a125506a  and  a125499a );
 a125510a <=( A266  and  A265 );
 a125513a <=( (not A268)  and  (not A267) );
 a125514a <=( a125513a  and  a125510a );
 a125517a <=( A299  and  A298 );
 a125520a <=( (not A302)  and  A301 );
 a125521a <=( a125520a  and  a125517a );
 a125522a <=( a125521a  and  a125514a );
 a125525a <=( A168  and  A169 );
 a125528a <=( A166  and  (not A167) );
 a125529a <=( a125528a  and  a125525a );
 a125532a <=( A200  and  A199 );
 a125535a <=( A203  and  (not A201) );
 a125536a <=( a125535a  and  a125532a );
 a125537a <=( a125536a  and  a125529a );
 a125540a <=( A266  and  A265 );
 a125543a <=( (not A268)  and  (not A267) );
 a125544a <=( a125543a  and  a125540a );
 a125547a <=( (not A299)  and  A298 );
 a125550a <=( A302  and  (not A301) );
 a125551a <=( a125550a  and  a125547a );
 a125552a <=( a125551a  and  a125544a );
 a125555a <=( A168  and  A169 );
 a125558a <=( A166  and  (not A167) );
 a125559a <=( a125558a  and  a125555a );
 a125562a <=( A200  and  A199 );
 a125565a <=( A203  and  (not A201) );
 a125566a <=( a125565a  and  a125562a );
 a125567a <=( a125566a  and  a125559a );
 a125570a <=( A266  and  A265 );
 a125573a <=( (not A268)  and  (not A267) );
 a125574a <=( a125573a  and  a125570a );
 a125577a <=( A299  and  (not A298) );
 a125580a <=( A302  and  (not A301) );
 a125581a <=( a125580a  and  a125577a );
 a125582a <=( a125581a  and  a125574a );
 a125585a <=( A168  and  A169 );
 a125588a <=( A166  and  (not A167) );
 a125589a <=( a125588a  and  a125585a );
 a125592a <=( A200  and  A199 );
 a125595a <=( A203  and  (not A201) );
 a125596a <=( a125595a  and  a125592a );
 a125597a <=( a125596a  and  a125589a );
 a125600a <=( A266  and  A265 );
 a125603a <=( (not A268)  and  (not A267) );
 a125604a <=( a125603a  and  a125600a );
 a125607a <=( (not A299)  and  (not A298) );
 a125610a <=( (not A302)  and  A301 );
 a125611a <=( a125610a  and  a125607a );
 a125612a <=( a125611a  and  a125604a );
 a125615a <=( A168  and  A169 );
 a125618a <=( A166  and  (not A167) );
 a125619a <=( a125618a  and  a125615a );
 a125622a <=( A200  and  A199 );
 a125625a <=( A203  and  (not A201) );
 a125626a <=( a125625a  and  a125622a );
 a125627a <=( a125626a  and  a125619a );
 a125630a <=( A266  and  A265 );
 a125633a <=( A269  and  (not A267) );
 a125634a <=( a125633a  and  a125630a );
 a125637a <=( A299  and  A298 );
 a125640a <=( (not A302)  and  A301 );
 a125641a <=( a125640a  and  a125637a );
 a125642a <=( a125641a  and  a125634a );
 a125645a <=( A168  and  A169 );
 a125648a <=( A166  and  (not A167) );
 a125649a <=( a125648a  and  a125645a );
 a125652a <=( A200  and  A199 );
 a125655a <=( A203  and  (not A201) );
 a125656a <=( a125655a  and  a125652a );
 a125657a <=( a125656a  and  a125649a );
 a125660a <=( A266  and  A265 );
 a125663a <=( A269  and  (not A267) );
 a125664a <=( a125663a  and  a125660a );
 a125667a <=( (not A299)  and  A298 );
 a125670a <=( A302  and  (not A301) );
 a125671a <=( a125670a  and  a125667a );
 a125672a <=( a125671a  and  a125664a );
 a125675a <=( A168  and  A169 );
 a125678a <=( A166  and  (not A167) );
 a125679a <=( a125678a  and  a125675a );
 a125682a <=( A200  and  A199 );
 a125685a <=( A203  and  (not A201) );
 a125686a <=( a125685a  and  a125682a );
 a125687a <=( a125686a  and  a125679a );
 a125690a <=( A266  and  A265 );
 a125693a <=( A269  and  (not A267) );
 a125694a <=( a125693a  and  a125690a );
 a125697a <=( A299  and  (not A298) );
 a125700a <=( A302  and  (not A301) );
 a125701a <=( a125700a  and  a125697a );
 a125702a <=( a125701a  and  a125694a );
 a125705a <=( A168  and  A169 );
 a125708a <=( A166  and  (not A167) );
 a125709a <=( a125708a  and  a125705a );
 a125712a <=( A200  and  A199 );
 a125715a <=( A203  and  (not A201) );
 a125716a <=( a125715a  and  a125712a );
 a125717a <=( a125716a  and  a125709a );
 a125720a <=( A266  and  A265 );
 a125723a <=( A269  and  (not A267) );
 a125724a <=( a125723a  and  a125720a );
 a125727a <=( (not A299)  and  (not A298) );
 a125730a <=( (not A302)  and  A301 );
 a125731a <=( a125730a  and  a125727a );
 a125732a <=( a125731a  and  a125724a );
 a125735a <=( A168  and  A169 );
 a125738a <=( A166  and  (not A167) );
 a125739a <=( a125738a  and  a125735a );
 a125742a <=( A200  and  A199 );
 a125745a <=( A203  and  (not A201) );
 a125746a <=( a125745a  and  a125742a );
 a125747a <=( a125746a  and  a125739a );
 a125750a <=( A266  and  (not A265) );
 a125753a <=( A268  and  (not A267) );
 a125754a <=( a125753a  and  a125750a );
 a125757a <=( A299  and  A298 );
 a125760a <=( (not A302)  and  A301 );
 a125761a <=( a125760a  and  a125757a );
 a125762a <=( a125761a  and  a125754a );
 a125765a <=( A168  and  A169 );
 a125768a <=( A166  and  (not A167) );
 a125769a <=( a125768a  and  a125765a );
 a125772a <=( A200  and  A199 );
 a125775a <=( A203  and  (not A201) );
 a125776a <=( a125775a  and  a125772a );
 a125777a <=( a125776a  and  a125769a );
 a125780a <=( A266  and  (not A265) );
 a125783a <=( A268  and  (not A267) );
 a125784a <=( a125783a  and  a125780a );
 a125787a <=( (not A299)  and  A298 );
 a125790a <=( A302  and  (not A301) );
 a125791a <=( a125790a  and  a125787a );
 a125792a <=( a125791a  and  a125784a );
 a125795a <=( A168  and  A169 );
 a125798a <=( A166  and  (not A167) );
 a125799a <=( a125798a  and  a125795a );
 a125802a <=( A200  and  A199 );
 a125805a <=( A203  and  (not A201) );
 a125806a <=( a125805a  and  a125802a );
 a125807a <=( a125806a  and  a125799a );
 a125810a <=( A266  and  (not A265) );
 a125813a <=( A268  and  (not A267) );
 a125814a <=( a125813a  and  a125810a );
 a125817a <=( A299  and  (not A298) );
 a125820a <=( A302  and  (not A301) );
 a125821a <=( a125820a  and  a125817a );
 a125822a <=( a125821a  and  a125814a );
 a125825a <=( A168  and  A169 );
 a125828a <=( A166  and  (not A167) );
 a125829a <=( a125828a  and  a125825a );
 a125832a <=( A200  and  A199 );
 a125835a <=( A203  and  (not A201) );
 a125836a <=( a125835a  and  a125832a );
 a125837a <=( a125836a  and  a125829a );
 a125840a <=( A266  and  (not A265) );
 a125843a <=( A268  and  (not A267) );
 a125844a <=( a125843a  and  a125840a );
 a125847a <=( (not A299)  and  (not A298) );
 a125850a <=( (not A302)  and  A301 );
 a125851a <=( a125850a  and  a125847a );
 a125852a <=( a125851a  and  a125844a );
 a125855a <=( A168  and  A169 );
 a125858a <=( A166  and  (not A167) );
 a125859a <=( a125858a  and  a125855a );
 a125862a <=( A200  and  A199 );
 a125865a <=( A203  and  (not A201) );
 a125866a <=( a125865a  and  a125862a );
 a125867a <=( a125866a  and  a125859a );
 a125870a <=( A266  and  (not A265) );
 a125873a <=( (not A269)  and  (not A267) );
 a125874a <=( a125873a  and  a125870a );
 a125877a <=( A299  and  A298 );
 a125880a <=( (not A302)  and  A301 );
 a125881a <=( a125880a  and  a125877a );
 a125882a <=( a125881a  and  a125874a );
 a125885a <=( A168  and  A169 );
 a125888a <=( A166  and  (not A167) );
 a125889a <=( a125888a  and  a125885a );
 a125892a <=( A200  and  A199 );
 a125895a <=( A203  and  (not A201) );
 a125896a <=( a125895a  and  a125892a );
 a125897a <=( a125896a  and  a125889a );
 a125900a <=( A266  and  (not A265) );
 a125903a <=( (not A269)  and  (not A267) );
 a125904a <=( a125903a  and  a125900a );
 a125907a <=( (not A299)  and  A298 );
 a125910a <=( A302  and  (not A301) );
 a125911a <=( a125910a  and  a125907a );
 a125912a <=( a125911a  and  a125904a );
 a125915a <=( A168  and  A169 );
 a125918a <=( A166  and  (not A167) );
 a125919a <=( a125918a  and  a125915a );
 a125922a <=( A200  and  A199 );
 a125925a <=( A203  and  (not A201) );
 a125926a <=( a125925a  and  a125922a );
 a125927a <=( a125926a  and  a125919a );
 a125930a <=( A266  and  (not A265) );
 a125933a <=( (not A269)  and  (not A267) );
 a125934a <=( a125933a  and  a125930a );
 a125937a <=( A299  and  (not A298) );
 a125940a <=( A302  and  (not A301) );
 a125941a <=( a125940a  and  a125937a );
 a125942a <=( a125941a  and  a125934a );
 a125945a <=( A168  and  A169 );
 a125948a <=( A166  and  (not A167) );
 a125949a <=( a125948a  and  a125945a );
 a125952a <=( A200  and  A199 );
 a125955a <=( A203  and  (not A201) );
 a125956a <=( a125955a  and  a125952a );
 a125957a <=( a125956a  and  a125949a );
 a125960a <=( A266  and  (not A265) );
 a125963a <=( (not A269)  and  (not A267) );
 a125964a <=( a125963a  and  a125960a );
 a125967a <=( (not A299)  and  (not A298) );
 a125970a <=( (not A302)  and  A301 );
 a125971a <=( a125970a  and  a125967a );
 a125972a <=( a125971a  and  a125964a );
 a125975a <=( A168  and  A169 );
 a125978a <=( A166  and  (not A167) );
 a125979a <=( a125978a  and  a125975a );
 a125982a <=( A200  and  A199 );
 a125985a <=( A203  and  (not A201) );
 a125986a <=( a125985a  and  a125982a );
 a125987a <=( a125986a  and  a125979a );
 a125990a <=( (not A266)  and  A265 );
 a125993a <=( A268  and  (not A267) );
 a125994a <=( a125993a  and  a125990a );
 a125997a <=( A299  and  A298 );
 a126000a <=( (not A302)  and  A301 );
 a126001a <=( a126000a  and  a125997a );
 a126002a <=( a126001a  and  a125994a );
 a126005a <=( A168  and  A169 );
 a126008a <=( A166  and  (not A167) );
 a126009a <=( a126008a  and  a126005a );
 a126012a <=( A200  and  A199 );
 a126015a <=( A203  and  (not A201) );
 a126016a <=( a126015a  and  a126012a );
 a126017a <=( a126016a  and  a126009a );
 a126020a <=( (not A266)  and  A265 );
 a126023a <=( A268  and  (not A267) );
 a126024a <=( a126023a  and  a126020a );
 a126027a <=( (not A299)  and  A298 );
 a126030a <=( A302  and  (not A301) );
 a126031a <=( a126030a  and  a126027a );
 a126032a <=( a126031a  and  a126024a );
 a126035a <=( A168  and  A169 );
 a126038a <=( A166  and  (not A167) );
 a126039a <=( a126038a  and  a126035a );
 a126042a <=( A200  and  A199 );
 a126045a <=( A203  and  (not A201) );
 a126046a <=( a126045a  and  a126042a );
 a126047a <=( a126046a  and  a126039a );
 a126050a <=( (not A266)  and  A265 );
 a126053a <=( A268  and  (not A267) );
 a126054a <=( a126053a  and  a126050a );
 a126057a <=( A299  and  (not A298) );
 a126060a <=( A302  and  (not A301) );
 a126061a <=( a126060a  and  a126057a );
 a126062a <=( a126061a  and  a126054a );
 a126065a <=( A168  and  A169 );
 a126068a <=( A166  and  (not A167) );
 a126069a <=( a126068a  and  a126065a );
 a126072a <=( A200  and  A199 );
 a126075a <=( A203  and  (not A201) );
 a126076a <=( a126075a  and  a126072a );
 a126077a <=( a126076a  and  a126069a );
 a126080a <=( (not A266)  and  A265 );
 a126083a <=( A268  and  (not A267) );
 a126084a <=( a126083a  and  a126080a );
 a126087a <=( (not A299)  and  (not A298) );
 a126090a <=( (not A302)  and  A301 );
 a126091a <=( a126090a  and  a126087a );
 a126092a <=( a126091a  and  a126084a );
 a126095a <=( A168  and  A169 );
 a126098a <=( A166  and  (not A167) );
 a126099a <=( a126098a  and  a126095a );
 a126102a <=( A200  and  A199 );
 a126105a <=( A203  and  (not A201) );
 a126106a <=( a126105a  and  a126102a );
 a126107a <=( a126106a  and  a126099a );
 a126110a <=( (not A266)  and  A265 );
 a126113a <=( (not A269)  and  (not A267) );
 a126114a <=( a126113a  and  a126110a );
 a126117a <=( A299  and  A298 );
 a126120a <=( (not A302)  and  A301 );
 a126121a <=( a126120a  and  a126117a );
 a126122a <=( a126121a  and  a126114a );
 a126125a <=( A168  and  A169 );
 a126128a <=( A166  and  (not A167) );
 a126129a <=( a126128a  and  a126125a );
 a126132a <=( A200  and  A199 );
 a126135a <=( A203  and  (not A201) );
 a126136a <=( a126135a  and  a126132a );
 a126137a <=( a126136a  and  a126129a );
 a126140a <=( (not A266)  and  A265 );
 a126143a <=( (not A269)  and  (not A267) );
 a126144a <=( a126143a  and  a126140a );
 a126147a <=( (not A299)  and  A298 );
 a126150a <=( A302  and  (not A301) );
 a126151a <=( a126150a  and  a126147a );
 a126152a <=( a126151a  and  a126144a );
 a126155a <=( A168  and  A169 );
 a126158a <=( A166  and  (not A167) );
 a126159a <=( a126158a  and  a126155a );
 a126162a <=( A200  and  A199 );
 a126165a <=( A203  and  (not A201) );
 a126166a <=( a126165a  and  a126162a );
 a126167a <=( a126166a  and  a126159a );
 a126170a <=( (not A266)  and  A265 );
 a126173a <=( (not A269)  and  (not A267) );
 a126174a <=( a126173a  and  a126170a );
 a126177a <=( A299  and  (not A298) );
 a126180a <=( A302  and  (not A301) );
 a126181a <=( a126180a  and  a126177a );
 a126182a <=( a126181a  and  a126174a );
 a126185a <=( A168  and  A169 );
 a126188a <=( A166  and  (not A167) );
 a126189a <=( a126188a  and  a126185a );
 a126192a <=( A200  and  A199 );
 a126195a <=( A203  and  (not A201) );
 a126196a <=( a126195a  and  a126192a );
 a126197a <=( a126196a  and  a126189a );
 a126200a <=( (not A266)  and  A265 );
 a126203a <=( (not A269)  and  (not A267) );
 a126204a <=( a126203a  and  a126200a );
 a126207a <=( (not A299)  and  (not A298) );
 a126210a <=( (not A302)  and  A301 );
 a126211a <=( a126210a  and  a126207a );
 a126212a <=( a126211a  and  a126204a );
 a126215a <=( A168  and  A169 );
 a126218a <=( A166  and  (not A167) );
 a126219a <=( a126218a  and  a126215a );
 a126222a <=( A200  and  (not A199) );
 a126225a <=( A203  and  (not A202) );
 a126226a <=( a126225a  and  a126222a );
 a126227a <=( a126226a  and  a126219a );
 a126230a <=( A266  and  A265 );
 a126233a <=( (not A269)  and  A268 );
 a126234a <=( a126233a  and  a126230a );
 a126237a <=( A299  and  A298 );
 a126240a <=( (not A301)  and  (not A300) );
 a126241a <=( a126240a  and  a126237a );
 a126242a <=( a126241a  and  a126234a );
 a126245a <=( A168  and  A169 );
 a126248a <=( A166  and  (not A167) );
 a126249a <=( a126248a  and  a126245a );
 a126252a <=( A200  and  (not A199) );
 a126255a <=( A203  and  (not A202) );
 a126256a <=( a126255a  and  a126252a );
 a126257a <=( a126256a  and  a126249a );
 a126260a <=( A266  and  A265 );
 a126263a <=( (not A269)  and  A268 );
 a126264a <=( a126263a  and  a126260a );
 a126267a <=( A299  and  A298 );
 a126270a <=( A302  and  (not A300) );
 a126271a <=( a126270a  and  a126267a );
 a126272a <=( a126271a  and  a126264a );
 a126275a <=( A168  and  A169 );
 a126278a <=( A166  and  (not A167) );
 a126279a <=( a126278a  and  a126275a );
 a126282a <=( A200  and  (not A199) );
 a126285a <=( A203  and  (not A202) );
 a126286a <=( a126285a  and  a126282a );
 a126287a <=( a126286a  and  a126279a );
 a126290a <=( A266  and  A265 );
 a126293a <=( (not A269)  and  A268 );
 a126294a <=( a126293a  and  a126290a );
 a126297a <=( (not A299)  and  A298 );
 a126300a <=( A301  and  (not A300) );
 a126301a <=( a126300a  and  a126297a );
 a126302a <=( a126301a  and  a126294a );
 a126305a <=( A168  and  A169 );
 a126308a <=( A166  and  (not A167) );
 a126309a <=( a126308a  and  a126305a );
 a126312a <=( A200  and  (not A199) );
 a126315a <=( A203  and  (not A202) );
 a126316a <=( a126315a  and  a126312a );
 a126317a <=( a126316a  and  a126309a );
 a126320a <=( A266  and  A265 );
 a126323a <=( (not A269)  and  A268 );
 a126324a <=( a126323a  and  a126320a );
 a126327a <=( (not A299)  and  A298 );
 a126330a <=( (not A302)  and  (not A300) );
 a126331a <=( a126330a  and  a126327a );
 a126332a <=( a126331a  and  a126324a );
 a126335a <=( A168  and  A169 );
 a126338a <=( A166  and  (not A167) );
 a126339a <=( a126338a  and  a126335a );
 a126342a <=( A200  and  (not A199) );
 a126345a <=( A203  and  (not A202) );
 a126346a <=( a126345a  and  a126342a );
 a126347a <=( a126346a  and  a126339a );
 a126350a <=( A266  and  A265 );
 a126353a <=( (not A269)  and  A268 );
 a126354a <=( a126353a  and  a126350a );
 a126357a <=( A299  and  (not A298) );
 a126360a <=( A301  and  (not A300) );
 a126361a <=( a126360a  and  a126357a );
 a126362a <=( a126361a  and  a126354a );
 a126365a <=( A168  and  A169 );
 a126368a <=( A166  and  (not A167) );
 a126369a <=( a126368a  and  a126365a );
 a126372a <=( A200  and  (not A199) );
 a126375a <=( A203  and  (not A202) );
 a126376a <=( a126375a  and  a126372a );
 a126377a <=( a126376a  and  a126369a );
 a126380a <=( A266  and  A265 );
 a126383a <=( (not A269)  and  A268 );
 a126384a <=( a126383a  and  a126380a );
 a126387a <=( A299  and  (not A298) );
 a126390a <=( (not A302)  and  (not A300) );
 a126391a <=( a126390a  and  a126387a );
 a126392a <=( a126391a  and  a126384a );
 a126395a <=( A168  and  A169 );
 a126398a <=( A166  and  (not A167) );
 a126399a <=( a126398a  and  a126395a );
 a126402a <=( A200  and  (not A199) );
 a126405a <=( A203  and  (not A202) );
 a126406a <=( a126405a  and  a126402a );
 a126407a <=( a126406a  and  a126399a );
 a126410a <=( A266  and  (not A265) );
 a126413a <=( A269  and  (not A268) );
 a126414a <=( a126413a  and  a126410a );
 a126417a <=( A299  and  A298 );
 a126420a <=( (not A301)  and  (not A300) );
 a126421a <=( a126420a  and  a126417a );
 a126422a <=( a126421a  and  a126414a );
 a126425a <=( A168  and  A169 );
 a126428a <=( A166  and  (not A167) );
 a126429a <=( a126428a  and  a126425a );
 a126432a <=( A200  and  (not A199) );
 a126435a <=( A203  and  (not A202) );
 a126436a <=( a126435a  and  a126432a );
 a126437a <=( a126436a  and  a126429a );
 a126440a <=( A266  and  (not A265) );
 a126443a <=( A269  and  (not A268) );
 a126444a <=( a126443a  and  a126440a );
 a126447a <=( A299  and  A298 );
 a126450a <=( A302  and  (not A300) );
 a126451a <=( a126450a  and  a126447a );
 a126452a <=( a126451a  and  a126444a );
 a126455a <=( A168  and  A169 );
 a126458a <=( A166  and  (not A167) );
 a126459a <=( a126458a  and  a126455a );
 a126462a <=( A200  and  (not A199) );
 a126465a <=( A203  and  (not A202) );
 a126466a <=( a126465a  and  a126462a );
 a126467a <=( a126466a  and  a126459a );
 a126470a <=( A266  and  (not A265) );
 a126473a <=( A269  and  (not A268) );
 a126474a <=( a126473a  and  a126470a );
 a126477a <=( (not A299)  and  A298 );
 a126480a <=( A301  and  (not A300) );
 a126481a <=( a126480a  and  a126477a );
 a126482a <=( a126481a  and  a126474a );
 a126485a <=( A168  and  A169 );
 a126488a <=( A166  and  (not A167) );
 a126489a <=( a126488a  and  a126485a );
 a126492a <=( A200  and  (not A199) );
 a126495a <=( A203  and  (not A202) );
 a126496a <=( a126495a  and  a126492a );
 a126497a <=( a126496a  and  a126489a );
 a126500a <=( A266  and  (not A265) );
 a126503a <=( A269  and  (not A268) );
 a126504a <=( a126503a  and  a126500a );
 a126507a <=( (not A299)  and  A298 );
 a126510a <=( (not A302)  and  (not A300) );
 a126511a <=( a126510a  and  a126507a );
 a126512a <=( a126511a  and  a126504a );
 a126515a <=( A168  and  A169 );
 a126518a <=( A166  and  (not A167) );
 a126519a <=( a126518a  and  a126515a );
 a126522a <=( A200  and  (not A199) );
 a126525a <=( A203  and  (not A202) );
 a126526a <=( a126525a  and  a126522a );
 a126527a <=( a126526a  and  a126519a );
 a126530a <=( A266  and  (not A265) );
 a126533a <=( A269  and  (not A268) );
 a126534a <=( a126533a  and  a126530a );
 a126537a <=( A299  and  (not A298) );
 a126540a <=( A301  and  (not A300) );
 a126541a <=( a126540a  and  a126537a );
 a126542a <=( a126541a  and  a126534a );
 a126545a <=( A168  and  A169 );
 a126548a <=( A166  and  (not A167) );
 a126549a <=( a126548a  and  a126545a );
 a126552a <=( A200  and  (not A199) );
 a126555a <=( A203  and  (not A202) );
 a126556a <=( a126555a  and  a126552a );
 a126557a <=( a126556a  and  a126549a );
 a126560a <=( A266  and  (not A265) );
 a126563a <=( A269  and  (not A268) );
 a126564a <=( a126563a  and  a126560a );
 a126567a <=( A299  and  (not A298) );
 a126570a <=( (not A302)  and  (not A300) );
 a126571a <=( a126570a  and  a126567a );
 a126572a <=( a126571a  and  a126564a );
 a126575a <=( A168  and  A169 );
 a126578a <=( A166  and  (not A167) );
 a126579a <=( a126578a  and  a126575a );
 a126582a <=( A200  and  (not A199) );
 a126585a <=( A203  and  (not A202) );
 a126586a <=( a126585a  and  a126582a );
 a126587a <=( a126586a  and  a126579a );
 a126590a <=( (not A266)  and  A265 );
 a126593a <=( A269  and  (not A268) );
 a126594a <=( a126593a  and  a126590a );
 a126597a <=( A299  and  A298 );
 a126600a <=( (not A301)  and  (not A300) );
 a126601a <=( a126600a  and  a126597a );
 a126602a <=( a126601a  and  a126594a );
 a126605a <=( A168  and  A169 );
 a126608a <=( A166  and  (not A167) );
 a126609a <=( a126608a  and  a126605a );
 a126612a <=( A200  and  (not A199) );
 a126615a <=( A203  and  (not A202) );
 a126616a <=( a126615a  and  a126612a );
 a126617a <=( a126616a  and  a126609a );
 a126620a <=( (not A266)  and  A265 );
 a126623a <=( A269  and  (not A268) );
 a126624a <=( a126623a  and  a126620a );
 a126627a <=( A299  and  A298 );
 a126630a <=( A302  and  (not A300) );
 a126631a <=( a126630a  and  a126627a );
 a126632a <=( a126631a  and  a126624a );
 a126635a <=( A168  and  A169 );
 a126638a <=( A166  and  (not A167) );
 a126639a <=( a126638a  and  a126635a );
 a126642a <=( A200  and  (not A199) );
 a126645a <=( A203  and  (not A202) );
 a126646a <=( a126645a  and  a126642a );
 a126647a <=( a126646a  and  a126639a );
 a126650a <=( (not A266)  and  A265 );
 a126653a <=( A269  and  (not A268) );
 a126654a <=( a126653a  and  a126650a );
 a126657a <=( (not A299)  and  A298 );
 a126660a <=( A301  and  (not A300) );
 a126661a <=( a126660a  and  a126657a );
 a126662a <=( a126661a  and  a126654a );
 a126665a <=( A168  and  A169 );
 a126668a <=( A166  and  (not A167) );
 a126669a <=( a126668a  and  a126665a );
 a126672a <=( A200  and  (not A199) );
 a126675a <=( A203  and  (not A202) );
 a126676a <=( a126675a  and  a126672a );
 a126677a <=( a126676a  and  a126669a );
 a126680a <=( (not A266)  and  A265 );
 a126683a <=( A269  and  (not A268) );
 a126684a <=( a126683a  and  a126680a );
 a126687a <=( (not A299)  and  A298 );
 a126690a <=( (not A302)  and  (not A300) );
 a126691a <=( a126690a  and  a126687a );
 a126692a <=( a126691a  and  a126684a );
 a126695a <=( A168  and  A169 );
 a126698a <=( A166  and  (not A167) );
 a126699a <=( a126698a  and  a126695a );
 a126702a <=( A200  and  (not A199) );
 a126705a <=( A203  and  (not A202) );
 a126706a <=( a126705a  and  a126702a );
 a126707a <=( a126706a  and  a126699a );
 a126710a <=( (not A266)  and  A265 );
 a126713a <=( A269  and  (not A268) );
 a126714a <=( a126713a  and  a126710a );
 a126717a <=( A299  and  (not A298) );
 a126720a <=( A301  and  (not A300) );
 a126721a <=( a126720a  and  a126717a );
 a126722a <=( a126721a  and  a126714a );
 a126725a <=( A168  and  A169 );
 a126728a <=( A166  and  (not A167) );
 a126729a <=( a126728a  and  a126725a );
 a126732a <=( A200  and  (not A199) );
 a126735a <=( A203  and  (not A202) );
 a126736a <=( a126735a  and  a126732a );
 a126737a <=( a126736a  and  a126729a );
 a126740a <=( (not A266)  and  A265 );
 a126743a <=( A269  and  (not A268) );
 a126744a <=( a126743a  and  a126740a );
 a126747a <=( A299  and  (not A298) );
 a126750a <=( (not A302)  and  (not A300) );
 a126751a <=( a126750a  and  a126747a );
 a126752a <=( a126751a  and  a126744a );
 a126755a <=( A168  and  A169 );
 a126758a <=( A166  and  (not A167) );
 a126759a <=( a126758a  and  a126755a );
 a126762a <=( A200  and  (not A199) );
 a126765a <=( A203  and  (not A202) );
 a126766a <=( a126765a  and  a126762a );
 a126767a <=( a126766a  and  a126759a );
 a126770a <=( (not A266)  and  (not A265) );
 a126773a <=( (not A269)  and  A268 );
 a126774a <=( a126773a  and  a126770a );
 a126777a <=( A299  and  A298 );
 a126780a <=( (not A301)  and  (not A300) );
 a126781a <=( a126780a  and  a126777a );
 a126782a <=( a126781a  and  a126774a );
 a126785a <=( A168  and  A169 );
 a126788a <=( A166  and  (not A167) );
 a126789a <=( a126788a  and  a126785a );
 a126792a <=( A200  and  (not A199) );
 a126795a <=( A203  and  (not A202) );
 a126796a <=( a126795a  and  a126792a );
 a126797a <=( a126796a  and  a126789a );
 a126800a <=( (not A266)  and  (not A265) );
 a126803a <=( (not A269)  and  A268 );
 a126804a <=( a126803a  and  a126800a );
 a126807a <=( A299  and  A298 );
 a126810a <=( A302  and  (not A300) );
 a126811a <=( a126810a  and  a126807a );
 a126812a <=( a126811a  and  a126804a );
 a126815a <=( A168  and  A169 );
 a126818a <=( A166  and  (not A167) );
 a126819a <=( a126818a  and  a126815a );
 a126822a <=( A200  and  (not A199) );
 a126825a <=( A203  and  (not A202) );
 a126826a <=( a126825a  and  a126822a );
 a126827a <=( a126826a  and  a126819a );
 a126830a <=( (not A266)  and  (not A265) );
 a126833a <=( (not A269)  and  A268 );
 a126834a <=( a126833a  and  a126830a );
 a126837a <=( (not A299)  and  A298 );
 a126840a <=( A301  and  (not A300) );
 a126841a <=( a126840a  and  a126837a );
 a126842a <=( a126841a  and  a126834a );
 a126845a <=( A168  and  A169 );
 a126848a <=( A166  and  (not A167) );
 a126849a <=( a126848a  and  a126845a );
 a126852a <=( A200  and  (not A199) );
 a126855a <=( A203  and  (not A202) );
 a126856a <=( a126855a  and  a126852a );
 a126857a <=( a126856a  and  a126849a );
 a126860a <=( (not A266)  and  (not A265) );
 a126863a <=( (not A269)  and  A268 );
 a126864a <=( a126863a  and  a126860a );
 a126867a <=( (not A299)  and  A298 );
 a126870a <=( (not A302)  and  (not A300) );
 a126871a <=( a126870a  and  a126867a );
 a126872a <=( a126871a  and  a126864a );
 a126875a <=( A168  and  A169 );
 a126878a <=( A166  and  (not A167) );
 a126879a <=( a126878a  and  a126875a );
 a126882a <=( A200  and  (not A199) );
 a126885a <=( A203  and  (not A202) );
 a126886a <=( a126885a  and  a126882a );
 a126887a <=( a126886a  and  a126879a );
 a126890a <=( (not A266)  and  (not A265) );
 a126893a <=( (not A269)  and  A268 );
 a126894a <=( a126893a  and  a126890a );
 a126897a <=( A299  and  (not A298) );
 a126900a <=( A301  and  (not A300) );
 a126901a <=( a126900a  and  a126897a );
 a126902a <=( a126901a  and  a126894a );
 a126905a <=( A168  and  A169 );
 a126908a <=( A166  and  (not A167) );
 a126909a <=( a126908a  and  a126905a );
 a126912a <=( A200  and  (not A199) );
 a126915a <=( A203  and  (not A202) );
 a126916a <=( a126915a  and  a126912a );
 a126917a <=( a126916a  and  a126909a );
 a126920a <=( (not A266)  and  (not A265) );
 a126923a <=( (not A269)  and  A268 );
 a126924a <=( a126923a  and  a126920a );
 a126927a <=( A299  and  (not A298) );
 a126930a <=( (not A302)  and  (not A300) );
 a126931a <=( a126930a  and  a126927a );
 a126932a <=( a126931a  and  a126924a );
 a126935a <=( A168  and  A169 );
 a126938a <=( A166  and  (not A167) );
 a126939a <=( a126938a  and  a126935a );
 a126942a <=( A200  and  (not A199) );
 a126945a <=( A202  and  (not A201) );
 a126946a <=( a126945a  and  a126942a );
 a126947a <=( a126946a  and  a126939a );
 a126950a <=( A266  and  A265 );
 a126953a <=( (not A268)  and  (not A267) );
 a126954a <=( a126953a  and  a126950a );
 a126957a <=( A299  and  A298 );
 a126960a <=( (not A302)  and  A301 );
 a126961a <=( a126960a  and  a126957a );
 a126962a <=( a126961a  and  a126954a );
 a126965a <=( A168  and  A169 );
 a126968a <=( A166  and  (not A167) );
 a126969a <=( a126968a  and  a126965a );
 a126972a <=( A200  and  (not A199) );
 a126975a <=( A202  and  (not A201) );
 a126976a <=( a126975a  and  a126972a );
 a126977a <=( a126976a  and  a126969a );
 a126980a <=( A266  and  A265 );
 a126983a <=( (not A268)  and  (not A267) );
 a126984a <=( a126983a  and  a126980a );
 a126987a <=( (not A299)  and  A298 );
 a126990a <=( A302  and  (not A301) );
 a126991a <=( a126990a  and  a126987a );
 a126992a <=( a126991a  and  a126984a );
 a126995a <=( A168  and  A169 );
 a126998a <=( A166  and  (not A167) );
 a126999a <=( a126998a  and  a126995a );
 a127002a <=( A200  and  (not A199) );
 a127005a <=( A202  and  (not A201) );
 a127006a <=( a127005a  and  a127002a );
 a127007a <=( a127006a  and  a126999a );
 a127010a <=( A266  and  A265 );
 a127013a <=( (not A268)  and  (not A267) );
 a127014a <=( a127013a  and  a127010a );
 a127017a <=( A299  and  (not A298) );
 a127020a <=( A302  and  (not A301) );
 a127021a <=( a127020a  and  a127017a );
 a127022a <=( a127021a  and  a127014a );
 a127025a <=( A168  and  A169 );
 a127028a <=( A166  and  (not A167) );
 a127029a <=( a127028a  and  a127025a );
 a127032a <=( A200  and  (not A199) );
 a127035a <=( A202  and  (not A201) );
 a127036a <=( a127035a  and  a127032a );
 a127037a <=( a127036a  and  a127029a );
 a127040a <=( A266  and  A265 );
 a127043a <=( (not A268)  and  (not A267) );
 a127044a <=( a127043a  and  a127040a );
 a127047a <=( (not A299)  and  (not A298) );
 a127050a <=( (not A302)  and  A301 );
 a127051a <=( a127050a  and  a127047a );
 a127052a <=( a127051a  and  a127044a );
 a127055a <=( A168  and  A169 );
 a127058a <=( A166  and  (not A167) );
 a127059a <=( a127058a  and  a127055a );
 a127062a <=( A200  and  (not A199) );
 a127065a <=( A202  and  (not A201) );
 a127066a <=( a127065a  and  a127062a );
 a127067a <=( a127066a  and  a127059a );
 a127070a <=( A266  and  A265 );
 a127073a <=( A269  and  (not A267) );
 a127074a <=( a127073a  and  a127070a );
 a127077a <=( A299  and  A298 );
 a127080a <=( (not A302)  and  A301 );
 a127081a <=( a127080a  and  a127077a );
 a127082a <=( a127081a  and  a127074a );
 a127085a <=( A168  and  A169 );
 a127088a <=( A166  and  (not A167) );
 a127089a <=( a127088a  and  a127085a );
 a127092a <=( A200  and  (not A199) );
 a127095a <=( A202  and  (not A201) );
 a127096a <=( a127095a  and  a127092a );
 a127097a <=( a127096a  and  a127089a );
 a127100a <=( A266  and  A265 );
 a127103a <=( A269  and  (not A267) );
 a127104a <=( a127103a  and  a127100a );
 a127107a <=( (not A299)  and  A298 );
 a127110a <=( A302  and  (not A301) );
 a127111a <=( a127110a  and  a127107a );
 a127112a <=( a127111a  and  a127104a );
 a127115a <=( A168  and  A169 );
 a127118a <=( A166  and  (not A167) );
 a127119a <=( a127118a  and  a127115a );
 a127122a <=( A200  and  (not A199) );
 a127125a <=( A202  and  (not A201) );
 a127126a <=( a127125a  and  a127122a );
 a127127a <=( a127126a  and  a127119a );
 a127130a <=( A266  and  A265 );
 a127133a <=( A269  and  (not A267) );
 a127134a <=( a127133a  and  a127130a );
 a127137a <=( A299  and  (not A298) );
 a127140a <=( A302  and  (not A301) );
 a127141a <=( a127140a  and  a127137a );
 a127142a <=( a127141a  and  a127134a );
 a127145a <=( A168  and  A169 );
 a127148a <=( A166  and  (not A167) );
 a127149a <=( a127148a  and  a127145a );
 a127152a <=( A200  and  (not A199) );
 a127155a <=( A202  and  (not A201) );
 a127156a <=( a127155a  and  a127152a );
 a127157a <=( a127156a  and  a127149a );
 a127160a <=( A266  and  A265 );
 a127163a <=( A269  and  (not A267) );
 a127164a <=( a127163a  and  a127160a );
 a127167a <=( (not A299)  and  (not A298) );
 a127170a <=( (not A302)  and  A301 );
 a127171a <=( a127170a  and  a127167a );
 a127172a <=( a127171a  and  a127164a );
 a127175a <=( A168  and  A169 );
 a127178a <=( A166  and  (not A167) );
 a127179a <=( a127178a  and  a127175a );
 a127182a <=( A200  and  (not A199) );
 a127185a <=( A202  and  (not A201) );
 a127186a <=( a127185a  and  a127182a );
 a127187a <=( a127186a  and  a127179a );
 a127190a <=( A266  and  (not A265) );
 a127193a <=( A268  and  (not A267) );
 a127194a <=( a127193a  and  a127190a );
 a127197a <=( A299  and  A298 );
 a127200a <=( (not A302)  and  A301 );
 a127201a <=( a127200a  and  a127197a );
 a127202a <=( a127201a  and  a127194a );
 a127205a <=( A168  and  A169 );
 a127208a <=( A166  and  (not A167) );
 a127209a <=( a127208a  and  a127205a );
 a127212a <=( A200  and  (not A199) );
 a127215a <=( A202  and  (not A201) );
 a127216a <=( a127215a  and  a127212a );
 a127217a <=( a127216a  and  a127209a );
 a127220a <=( A266  and  (not A265) );
 a127223a <=( A268  and  (not A267) );
 a127224a <=( a127223a  and  a127220a );
 a127227a <=( (not A299)  and  A298 );
 a127230a <=( A302  and  (not A301) );
 a127231a <=( a127230a  and  a127227a );
 a127232a <=( a127231a  and  a127224a );
 a127235a <=( A168  and  A169 );
 a127238a <=( A166  and  (not A167) );
 a127239a <=( a127238a  and  a127235a );
 a127242a <=( A200  and  (not A199) );
 a127245a <=( A202  and  (not A201) );
 a127246a <=( a127245a  and  a127242a );
 a127247a <=( a127246a  and  a127239a );
 a127250a <=( A266  and  (not A265) );
 a127253a <=( A268  and  (not A267) );
 a127254a <=( a127253a  and  a127250a );
 a127257a <=( A299  and  (not A298) );
 a127260a <=( A302  and  (not A301) );
 a127261a <=( a127260a  and  a127257a );
 a127262a <=( a127261a  and  a127254a );
 a127265a <=( A168  and  A169 );
 a127268a <=( A166  and  (not A167) );
 a127269a <=( a127268a  and  a127265a );
 a127272a <=( A200  and  (not A199) );
 a127275a <=( A202  and  (not A201) );
 a127276a <=( a127275a  and  a127272a );
 a127277a <=( a127276a  and  a127269a );
 a127280a <=( A266  and  (not A265) );
 a127283a <=( A268  and  (not A267) );
 a127284a <=( a127283a  and  a127280a );
 a127287a <=( (not A299)  and  (not A298) );
 a127290a <=( (not A302)  and  A301 );
 a127291a <=( a127290a  and  a127287a );
 a127292a <=( a127291a  and  a127284a );
 a127295a <=( A168  and  A169 );
 a127298a <=( A166  and  (not A167) );
 a127299a <=( a127298a  and  a127295a );
 a127302a <=( A200  and  (not A199) );
 a127305a <=( A202  and  (not A201) );
 a127306a <=( a127305a  and  a127302a );
 a127307a <=( a127306a  and  a127299a );
 a127310a <=( A266  and  (not A265) );
 a127313a <=( (not A269)  and  (not A267) );
 a127314a <=( a127313a  and  a127310a );
 a127317a <=( A299  and  A298 );
 a127320a <=( (not A302)  and  A301 );
 a127321a <=( a127320a  and  a127317a );
 a127322a <=( a127321a  and  a127314a );
 a127325a <=( A168  and  A169 );
 a127328a <=( A166  and  (not A167) );
 a127329a <=( a127328a  and  a127325a );
 a127332a <=( A200  and  (not A199) );
 a127335a <=( A202  and  (not A201) );
 a127336a <=( a127335a  and  a127332a );
 a127337a <=( a127336a  and  a127329a );
 a127340a <=( A266  and  (not A265) );
 a127343a <=( (not A269)  and  (not A267) );
 a127344a <=( a127343a  and  a127340a );
 a127347a <=( (not A299)  and  A298 );
 a127350a <=( A302  and  (not A301) );
 a127351a <=( a127350a  and  a127347a );
 a127352a <=( a127351a  and  a127344a );
 a127355a <=( A168  and  A169 );
 a127358a <=( A166  and  (not A167) );
 a127359a <=( a127358a  and  a127355a );
 a127362a <=( A200  and  (not A199) );
 a127365a <=( A202  and  (not A201) );
 a127366a <=( a127365a  and  a127362a );
 a127367a <=( a127366a  and  a127359a );
 a127370a <=( A266  and  (not A265) );
 a127373a <=( (not A269)  and  (not A267) );
 a127374a <=( a127373a  and  a127370a );
 a127377a <=( A299  and  (not A298) );
 a127380a <=( A302  and  (not A301) );
 a127381a <=( a127380a  and  a127377a );
 a127382a <=( a127381a  and  a127374a );
 a127385a <=( A168  and  A169 );
 a127388a <=( A166  and  (not A167) );
 a127389a <=( a127388a  and  a127385a );
 a127392a <=( A200  and  (not A199) );
 a127395a <=( A202  and  (not A201) );
 a127396a <=( a127395a  and  a127392a );
 a127397a <=( a127396a  and  a127389a );
 a127400a <=( A266  and  (not A265) );
 a127403a <=( (not A269)  and  (not A267) );
 a127404a <=( a127403a  and  a127400a );
 a127407a <=( (not A299)  and  (not A298) );
 a127410a <=( (not A302)  and  A301 );
 a127411a <=( a127410a  and  a127407a );
 a127412a <=( a127411a  and  a127404a );
 a127415a <=( A168  and  A169 );
 a127418a <=( A166  and  (not A167) );
 a127419a <=( a127418a  and  a127415a );
 a127422a <=( A200  and  (not A199) );
 a127425a <=( A202  and  (not A201) );
 a127426a <=( a127425a  and  a127422a );
 a127427a <=( a127426a  and  a127419a );
 a127430a <=( (not A266)  and  A265 );
 a127433a <=( A268  and  (not A267) );
 a127434a <=( a127433a  and  a127430a );
 a127437a <=( A299  and  A298 );
 a127440a <=( (not A302)  and  A301 );
 a127441a <=( a127440a  and  a127437a );
 a127442a <=( a127441a  and  a127434a );
 a127445a <=( A168  and  A169 );
 a127448a <=( A166  and  (not A167) );
 a127449a <=( a127448a  and  a127445a );
 a127452a <=( A200  and  (not A199) );
 a127455a <=( A202  and  (not A201) );
 a127456a <=( a127455a  and  a127452a );
 a127457a <=( a127456a  and  a127449a );
 a127460a <=( (not A266)  and  A265 );
 a127463a <=( A268  and  (not A267) );
 a127464a <=( a127463a  and  a127460a );
 a127467a <=( (not A299)  and  A298 );
 a127470a <=( A302  and  (not A301) );
 a127471a <=( a127470a  and  a127467a );
 a127472a <=( a127471a  and  a127464a );
 a127475a <=( A168  and  A169 );
 a127478a <=( A166  and  (not A167) );
 a127479a <=( a127478a  and  a127475a );
 a127482a <=( A200  and  (not A199) );
 a127485a <=( A202  and  (not A201) );
 a127486a <=( a127485a  and  a127482a );
 a127487a <=( a127486a  and  a127479a );
 a127490a <=( (not A266)  and  A265 );
 a127493a <=( A268  and  (not A267) );
 a127494a <=( a127493a  and  a127490a );
 a127497a <=( A299  and  (not A298) );
 a127500a <=( A302  and  (not A301) );
 a127501a <=( a127500a  and  a127497a );
 a127502a <=( a127501a  and  a127494a );
 a127505a <=( A168  and  A169 );
 a127508a <=( A166  and  (not A167) );
 a127509a <=( a127508a  and  a127505a );
 a127512a <=( A200  and  (not A199) );
 a127515a <=( A202  and  (not A201) );
 a127516a <=( a127515a  and  a127512a );
 a127517a <=( a127516a  and  a127509a );
 a127520a <=( (not A266)  and  A265 );
 a127523a <=( A268  and  (not A267) );
 a127524a <=( a127523a  and  a127520a );
 a127527a <=( (not A299)  and  (not A298) );
 a127530a <=( (not A302)  and  A301 );
 a127531a <=( a127530a  and  a127527a );
 a127532a <=( a127531a  and  a127524a );
 a127535a <=( A168  and  A169 );
 a127538a <=( A166  and  (not A167) );
 a127539a <=( a127538a  and  a127535a );
 a127542a <=( A200  and  (not A199) );
 a127545a <=( A202  and  (not A201) );
 a127546a <=( a127545a  and  a127542a );
 a127547a <=( a127546a  and  a127539a );
 a127550a <=( (not A266)  and  A265 );
 a127553a <=( (not A269)  and  (not A267) );
 a127554a <=( a127553a  and  a127550a );
 a127557a <=( A299  and  A298 );
 a127560a <=( (not A302)  and  A301 );
 a127561a <=( a127560a  and  a127557a );
 a127562a <=( a127561a  and  a127554a );
 a127565a <=( A168  and  A169 );
 a127568a <=( A166  and  (not A167) );
 a127569a <=( a127568a  and  a127565a );
 a127572a <=( A200  and  (not A199) );
 a127575a <=( A202  and  (not A201) );
 a127576a <=( a127575a  and  a127572a );
 a127577a <=( a127576a  and  a127569a );
 a127580a <=( (not A266)  and  A265 );
 a127583a <=( (not A269)  and  (not A267) );
 a127584a <=( a127583a  and  a127580a );
 a127587a <=( (not A299)  and  A298 );
 a127590a <=( A302  and  (not A301) );
 a127591a <=( a127590a  and  a127587a );
 a127592a <=( a127591a  and  a127584a );
 a127595a <=( A168  and  A169 );
 a127598a <=( A166  and  (not A167) );
 a127599a <=( a127598a  and  a127595a );
 a127602a <=( A200  and  (not A199) );
 a127605a <=( A202  and  (not A201) );
 a127606a <=( a127605a  and  a127602a );
 a127607a <=( a127606a  and  a127599a );
 a127610a <=( (not A266)  and  A265 );
 a127613a <=( (not A269)  and  (not A267) );
 a127614a <=( a127613a  and  a127610a );
 a127617a <=( A299  and  (not A298) );
 a127620a <=( A302  and  (not A301) );
 a127621a <=( a127620a  and  a127617a );
 a127622a <=( a127621a  and  a127614a );
 a127625a <=( A168  and  A169 );
 a127628a <=( A166  and  (not A167) );
 a127629a <=( a127628a  and  a127625a );
 a127632a <=( A200  and  (not A199) );
 a127635a <=( A202  and  (not A201) );
 a127636a <=( a127635a  and  a127632a );
 a127637a <=( a127636a  and  a127629a );
 a127640a <=( (not A266)  and  A265 );
 a127643a <=( (not A269)  and  (not A267) );
 a127644a <=( a127643a  and  a127640a );
 a127647a <=( (not A299)  and  (not A298) );
 a127650a <=( (not A302)  and  A301 );
 a127651a <=( a127650a  and  a127647a );
 a127652a <=( a127651a  and  a127644a );
 a127655a <=( A168  and  A169 );
 a127658a <=( A166  and  (not A167) );
 a127659a <=( a127658a  and  a127655a );
 a127662a <=( A200  and  (not A199) );
 a127665a <=( (not A203)  and  (not A201) );
 a127666a <=( a127665a  and  a127662a );
 a127667a <=( a127666a  and  a127659a );
 a127670a <=( A266  and  A265 );
 a127673a <=( (not A268)  and  (not A267) );
 a127674a <=( a127673a  and  a127670a );
 a127677a <=( A299  and  A298 );
 a127680a <=( (not A302)  and  A301 );
 a127681a <=( a127680a  and  a127677a );
 a127682a <=( a127681a  and  a127674a );
 a127685a <=( A168  and  A169 );
 a127688a <=( A166  and  (not A167) );
 a127689a <=( a127688a  and  a127685a );
 a127692a <=( A200  and  (not A199) );
 a127695a <=( (not A203)  and  (not A201) );
 a127696a <=( a127695a  and  a127692a );
 a127697a <=( a127696a  and  a127689a );
 a127700a <=( A266  and  A265 );
 a127703a <=( (not A268)  and  (not A267) );
 a127704a <=( a127703a  and  a127700a );
 a127707a <=( (not A299)  and  A298 );
 a127710a <=( A302  and  (not A301) );
 a127711a <=( a127710a  and  a127707a );
 a127712a <=( a127711a  and  a127704a );
 a127715a <=( A168  and  A169 );
 a127718a <=( A166  and  (not A167) );
 a127719a <=( a127718a  and  a127715a );
 a127722a <=( A200  and  (not A199) );
 a127725a <=( (not A203)  and  (not A201) );
 a127726a <=( a127725a  and  a127722a );
 a127727a <=( a127726a  and  a127719a );
 a127730a <=( A266  and  A265 );
 a127733a <=( (not A268)  and  (not A267) );
 a127734a <=( a127733a  and  a127730a );
 a127737a <=( A299  and  (not A298) );
 a127740a <=( A302  and  (not A301) );
 a127741a <=( a127740a  and  a127737a );
 a127742a <=( a127741a  and  a127734a );
 a127745a <=( A168  and  A169 );
 a127748a <=( A166  and  (not A167) );
 a127749a <=( a127748a  and  a127745a );
 a127752a <=( A200  and  (not A199) );
 a127755a <=( (not A203)  and  (not A201) );
 a127756a <=( a127755a  and  a127752a );
 a127757a <=( a127756a  and  a127749a );
 a127760a <=( A266  and  A265 );
 a127763a <=( (not A268)  and  (not A267) );
 a127764a <=( a127763a  and  a127760a );
 a127767a <=( (not A299)  and  (not A298) );
 a127770a <=( (not A302)  and  A301 );
 a127771a <=( a127770a  and  a127767a );
 a127772a <=( a127771a  and  a127764a );
 a127775a <=( A168  and  A169 );
 a127778a <=( A166  and  (not A167) );
 a127779a <=( a127778a  and  a127775a );
 a127782a <=( A200  and  (not A199) );
 a127785a <=( (not A203)  and  (not A201) );
 a127786a <=( a127785a  and  a127782a );
 a127787a <=( a127786a  and  a127779a );
 a127790a <=( A266  and  A265 );
 a127793a <=( A269  and  (not A267) );
 a127794a <=( a127793a  and  a127790a );
 a127797a <=( A299  and  A298 );
 a127800a <=( (not A302)  and  A301 );
 a127801a <=( a127800a  and  a127797a );
 a127802a <=( a127801a  and  a127794a );
 a127805a <=( A168  and  A169 );
 a127808a <=( A166  and  (not A167) );
 a127809a <=( a127808a  and  a127805a );
 a127812a <=( A200  and  (not A199) );
 a127815a <=( (not A203)  and  (not A201) );
 a127816a <=( a127815a  and  a127812a );
 a127817a <=( a127816a  and  a127809a );
 a127820a <=( A266  and  A265 );
 a127823a <=( A269  and  (not A267) );
 a127824a <=( a127823a  and  a127820a );
 a127827a <=( (not A299)  and  A298 );
 a127830a <=( A302  and  (not A301) );
 a127831a <=( a127830a  and  a127827a );
 a127832a <=( a127831a  and  a127824a );
 a127835a <=( A168  and  A169 );
 a127838a <=( A166  and  (not A167) );
 a127839a <=( a127838a  and  a127835a );
 a127842a <=( A200  and  (not A199) );
 a127845a <=( (not A203)  and  (not A201) );
 a127846a <=( a127845a  and  a127842a );
 a127847a <=( a127846a  and  a127839a );
 a127850a <=( A266  and  A265 );
 a127853a <=( A269  and  (not A267) );
 a127854a <=( a127853a  and  a127850a );
 a127857a <=( A299  and  (not A298) );
 a127860a <=( A302  and  (not A301) );
 a127861a <=( a127860a  and  a127857a );
 a127862a <=( a127861a  and  a127854a );
 a127865a <=( A168  and  A169 );
 a127868a <=( A166  and  (not A167) );
 a127869a <=( a127868a  and  a127865a );
 a127872a <=( A200  and  (not A199) );
 a127875a <=( (not A203)  and  (not A201) );
 a127876a <=( a127875a  and  a127872a );
 a127877a <=( a127876a  and  a127869a );
 a127880a <=( A266  and  A265 );
 a127883a <=( A269  and  (not A267) );
 a127884a <=( a127883a  and  a127880a );
 a127887a <=( (not A299)  and  (not A298) );
 a127890a <=( (not A302)  and  A301 );
 a127891a <=( a127890a  and  a127887a );
 a127892a <=( a127891a  and  a127884a );
 a127895a <=( A168  and  A169 );
 a127898a <=( A166  and  (not A167) );
 a127899a <=( a127898a  and  a127895a );
 a127902a <=( A200  and  (not A199) );
 a127905a <=( (not A203)  and  (not A201) );
 a127906a <=( a127905a  and  a127902a );
 a127907a <=( a127906a  and  a127899a );
 a127910a <=( A266  and  (not A265) );
 a127913a <=( A268  and  (not A267) );
 a127914a <=( a127913a  and  a127910a );
 a127917a <=( A299  and  A298 );
 a127920a <=( (not A302)  and  A301 );
 a127921a <=( a127920a  and  a127917a );
 a127922a <=( a127921a  and  a127914a );
 a127925a <=( A168  and  A169 );
 a127928a <=( A166  and  (not A167) );
 a127929a <=( a127928a  and  a127925a );
 a127932a <=( A200  and  (not A199) );
 a127935a <=( (not A203)  and  (not A201) );
 a127936a <=( a127935a  and  a127932a );
 a127937a <=( a127936a  and  a127929a );
 a127940a <=( A266  and  (not A265) );
 a127943a <=( A268  and  (not A267) );
 a127944a <=( a127943a  and  a127940a );
 a127947a <=( (not A299)  and  A298 );
 a127950a <=( A302  and  (not A301) );
 a127951a <=( a127950a  and  a127947a );
 a127952a <=( a127951a  and  a127944a );
 a127955a <=( A168  and  A169 );
 a127958a <=( A166  and  (not A167) );
 a127959a <=( a127958a  and  a127955a );
 a127962a <=( A200  and  (not A199) );
 a127965a <=( (not A203)  and  (not A201) );
 a127966a <=( a127965a  and  a127962a );
 a127967a <=( a127966a  and  a127959a );
 a127970a <=( A266  and  (not A265) );
 a127973a <=( A268  and  (not A267) );
 a127974a <=( a127973a  and  a127970a );
 a127977a <=( A299  and  (not A298) );
 a127980a <=( A302  and  (not A301) );
 a127981a <=( a127980a  and  a127977a );
 a127982a <=( a127981a  and  a127974a );
 a127985a <=( A168  and  A169 );
 a127988a <=( A166  and  (not A167) );
 a127989a <=( a127988a  and  a127985a );
 a127992a <=( A200  and  (not A199) );
 a127995a <=( (not A203)  and  (not A201) );
 a127996a <=( a127995a  and  a127992a );
 a127997a <=( a127996a  and  a127989a );
 a128000a <=( A266  and  (not A265) );
 a128003a <=( A268  and  (not A267) );
 a128004a <=( a128003a  and  a128000a );
 a128007a <=( (not A299)  and  (not A298) );
 a128010a <=( (not A302)  and  A301 );
 a128011a <=( a128010a  and  a128007a );
 a128012a <=( a128011a  and  a128004a );
 a128015a <=( A168  and  A169 );
 a128018a <=( A166  and  (not A167) );
 a128019a <=( a128018a  and  a128015a );
 a128022a <=( A200  and  (not A199) );
 a128025a <=( (not A203)  and  (not A201) );
 a128026a <=( a128025a  and  a128022a );
 a128027a <=( a128026a  and  a128019a );
 a128030a <=( A266  and  (not A265) );
 a128033a <=( (not A269)  and  (not A267) );
 a128034a <=( a128033a  and  a128030a );
 a128037a <=( A299  and  A298 );
 a128040a <=( (not A302)  and  A301 );
 a128041a <=( a128040a  and  a128037a );
 a128042a <=( a128041a  and  a128034a );
 a128045a <=( A168  and  A169 );
 a128048a <=( A166  and  (not A167) );
 a128049a <=( a128048a  and  a128045a );
 a128052a <=( A200  and  (not A199) );
 a128055a <=( (not A203)  and  (not A201) );
 a128056a <=( a128055a  and  a128052a );
 a128057a <=( a128056a  and  a128049a );
 a128060a <=( A266  and  (not A265) );
 a128063a <=( (not A269)  and  (not A267) );
 a128064a <=( a128063a  and  a128060a );
 a128067a <=( (not A299)  and  A298 );
 a128070a <=( A302  and  (not A301) );
 a128071a <=( a128070a  and  a128067a );
 a128072a <=( a128071a  and  a128064a );
 a128075a <=( A168  and  A169 );
 a128078a <=( A166  and  (not A167) );
 a128079a <=( a128078a  and  a128075a );
 a128082a <=( A200  and  (not A199) );
 a128085a <=( (not A203)  and  (not A201) );
 a128086a <=( a128085a  and  a128082a );
 a128087a <=( a128086a  and  a128079a );
 a128090a <=( A266  and  (not A265) );
 a128093a <=( (not A269)  and  (not A267) );
 a128094a <=( a128093a  and  a128090a );
 a128097a <=( A299  and  (not A298) );
 a128100a <=( A302  and  (not A301) );
 a128101a <=( a128100a  and  a128097a );
 a128102a <=( a128101a  and  a128094a );
 a128105a <=( A168  and  A169 );
 a128108a <=( A166  and  (not A167) );
 a128109a <=( a128108a  and  a128105a );
 a128112a <=( A200  and  (not A199) );
 a128115a <=( (not A203)  and  (not A201) );
 a128116a <=( a128115a  and  a128112a );
 a128117a <=( a128116a  and  a128109a );
 a128120a <=( A266  and  (not A265) );
 a128123a <=( (not A269)  and  (not A267) );
 a128124a <=( a128123a  and  a128120a );
 a128127a <=( (not A299)  and  (not A298) );
 a128130a <=( (not A302)  and  A301 );
 a128131a <=( a128130a  and  a128127a );
 a128132a <=( a128131a  and  a128124a );
 a128135a <=( A168  and  A169 );
 a128138a <=( A166  and  (not A167) );
 a128139a <=( a128138a  and  a128135a );
 a128142a <=( A200  and  (not A199) );
 a128145a <=( (not A203)  and  (not A201) );
 a128146a <=( a128145a  and  a128142a );
 a128147a <=( a128146a  and  a128139a );
 a128150a <=( (not A266)  and  A265 );
 a128153a <=( A268  and  (not A267) );
 a128154a <=( a128153a  and  a128150a );
 a128157a <=( A299  and  A298 );
 a128160a <=( (not A302)  and  A301 );
 a128161a <=( a128160a  and  a128157a );
 a128162a <=( a128161a  and  a128154a );
 a128165a <=( A168  and  A169 );
 a128168a <=( A166  and  (not A167) );
 a128169a <=( a128168a  and  a128165a );
 a128172a <=( A200  and  (not A199) );
 a128175a <=( (not A203)  and  (not A201) );
 a128176a <=( a128175a  and  a128172a );
 a128177a <=( a128176a  and  a128169a );
 a128180a <=( (not A266)  and  A265 );
 a128183a <=( A268  and  (not A267) );
 a128184a <=( a128183a  and  a128180a );
 a128187a <=( (not A299)  and  A298 );
 a128190a <=( A302  and  (not A301) );
 a128191a <=( a128190a  and  a128187a );
 a128192a <=( a128191a  and  a128184a );
 a128195a <=( A168  and  A169 );
 a128198a <=( A166  and  (not A167) );
 a128199a <=( a128198a  and  a128195a );
 a128202a <=( A200  and  (not A199) );
 a128205a <=( (not A203)  and  (not A201) );
 a128206a <=( a128205a  and  a128202a );
 a128207a <=( a128206a  and  a128199a );
 a128210a <=( (not A266)  and  A265 );
 a128213a <=( A268  and  (not A267) );
 a128214a <=( a128213a  and  a128210a );
 a128217a <=( A299  and  (not A298) );
 a128220a <=( A302  and  (not A301) );
 a128221a <=( a128220a  and  a128217a );
 a128222a <=( a128221a  and  a128214a );
 a128225a <=( A168  and  A169 );
 a128228a <=( A166  and  (not A167) );
 a128229a <=( a128228a  and  a128225a );
 a128232a <=( A200  and  (not A199) );
 a128235a <=( (not A203)  and  (not A201) );
 a128236a <=( a128235a  and  a128232a );
 a128237a <=( a128236a  and  a128229a );
 a128240a <=( (not A266)  and  A265 );
 a128243a <=( A268  and  (not A267) );
 a128244a <=( a128243a  and  a128240a );
 a128247a <=( (not A299)  and  (not A298) );
 a128250a <=( (not A302)  and  A301 );
 a128251a <=( a128250a  and  a128247a );
 a128252a <=( a128251a  and  a128244a );
 a128255a <=( A168  and  A169 );
 a128258a <=( A166  and  (not A167) );
 a128259a <=( a128258a  and  a128255a );
 a128262a <=( A200  and  (not A199) );
 a128265a <=( (not A203)  and  (not A201) );
 a128266a <=( a128265a  and  a128262a );
 a128267a <=( a128266a  and  a128259a );
 a128270a <=( (not A266)  and  A265 );
 a128273a <=( (not A269)  and  (not A267) );
 a128274a <=( a128273a  and  a128270a );
 a128277a <=( A299  and  A298 );
 a128280a <=( (not A302)  and  A301 );
 a128281a <=( a128280a  and  a128277a );
 a128282a <=( a128281a  and  a128274a );
 a128285a <=( A168  and  A169 );
 a128288a <=( A166  and  (not A167) );
 a128289a <=( a128288a  and  a128285a );
 a128292a <=( A200  and  (not A199) );
 a128295a <=( (not A203)  and  (not A201) );
 a128296a <=( a128295a  and  a128292a );
 a128297a <=( a128296a  and  a128289a );
 a128300a <=( (not A266)  and  A265 );
 a128303a <=( (not A269)  and  (not A267) );
 a128304a <=( a128303a  and  a128300a );
 a128307a <=( (not A299)  and  A298 );
 a128310a <=( A302  and  (not A301) );
 a128311a <=( a128310a  and  a128307a );
 a128312a <=( a128311a  and  a128304a );
 a128315a <=( A168  and  A169 );
 a128318a <=( A166  and  (not A167) );
 a128319a <=( a128318a  and  a128315a );
 a128322a <=( A200  and  (not A199) );
 a128325a <=( (not A203)  and  (not A201) );
 a128326a <=( a128325a  and  a128322a );
 a128327a <=( a128326a  and  a128319a );
 a128330a <=( (not A266)  and  A265 );
 a128333a <=( (not A269)  and  (not A267) );
 a128334a <=( a128333a  and  a128330a );
 a128337a <=( A299  and  (not A298) );
 a128340a <=( A302  and  (not A301) );
 a128341a <=( a128340a  and  a128337a );
 a128342a <=( a128341a  and  a128334a );
 a128345a <=( A168  and  A169 );
 a128348a <=( A166  and  (not A167) );
 a128349a <=( a128348a  and  a128345a );
 a128352a <=( A200  and  (not A199) );
 a128355a <=( (not A203)  and  (not A201) );
 a128356a <=( a128355a  and  a128352a );
 a128357a <=( a128356a  and  a128349a );
 a128360a <=( (not A266)  and  A265 );
 a128363a <=( (not A269)  and  (not A267) );
 a128364a <=( a128363a  and  a128360a );
 a128367a <=( (not A299)  and  (not A298) );
 a128370a <=( (not A302)  and  A301 );
 a128371a <=( a128370a  and  a128367a );
 a128372a <=( a128371a  and  a128364a );
 a128375a <=( A168  and  A169 );
 a128378a <=( A166  and  (not A167) );
 a128379a <=( a128378a  and  a128375a );
 a128382a <=( (not A200)  and  A199 );
 a128385a <=( A203  and  (not A202) );
 a128386a <=( a128385a  and  a128382a );
 a128387a <=( a128386a  and  a128379a );
 a128390a <=( A266  and  A265 );
 a128393a <=( (not A269)  and  A268 );
 a128394a <=( a128393a  and  a128390a );
 a128397a <=( A299  and  A298 );
 a128400a <=( (not A301)  and  (not A300) );
 a128401a <=( a128400a  and  a128397a );
 a128402a <=( a128401a  and  a128394a );
 a128405a <=( A168  and  A169 );
 a128408a <=( A166  and  (not A167) );
 a128409a <=( a128408a  and  a128405a );
 a128412a <=( (not A200)  and  A199 );
 a128415a <=( A203  and  (not A202) );
 a128416a <=( a128415a  and  a128412a );
 a128417a <=( a128416a  and  a128409a );
 a128420a <=( A266  and  A265 );
 a128423a <=( (not A269)  and  A268 );
 a128424a <=( a128423a  and  a128420a );
 a128427a <=( A299  and  A298 );
 a128430a <=( A302  and  (not A300) );
 a128431a <=( a128430a  and  a128427a );
 a128432a <=( a128431a  and  a128424a );
 a128435a <=( A168  and  A169 );
 a128438a <=( A166  and  (not A167) );
 a128439a <=( a128438a  and  a128435a );
 a128442a <=( (not A200)  and  A199 );
 a128445a <=( A203  and  (not A202) );
 a128446a <=( a128445a  and  a128442a );
 a128447a <=( a128446a  and  a128439a );
 a128450a <=( A266  and  A265 );
 a128453a <=( (not A269)  and  A268 );
 a128454a <=( a128453a  and  a128450a );
 a128457a <=( (not A299)  and  A298 );
 a128460a <=( A301  and  (not A300) );
 a128461a <=( a128460a  and  a128457a );
 a128462a <=( a128461a  and  a128454a );
 a128465a <=( A168  and  A169 );
 a128468a <=( A166  and  (not A167) );
 a128469a <=( a128468a  and  a128465a );
 a128472a <=( (not A200)  and  A199 );
 a128475a <=( A203  and  (not A202) );
 a128476a <=( a128475a  and  a128472a );
 a128477a <=( a128476a  and  a128469a );
 a128480a <=( A266  and  A265 );
 a128483a <=( (not A269)  and  A268 );
 a128484a <=( a128483a  and  a128480a );
 a128487a <=( (not A299)  and  A298 );
 a128490a <=( (not A302)  and  (not A300) );
 a128491a <=( a128490a  and  a128487a );
 a128492a <=( a128491a  and  a128484a );
 a128495a <=( A168  and  A169 );
 a128498a <=( A166  and  (not A167) );
 a128499a <=( a128498a  and  a128495a );
 a128502a <=( (not A200)  and  A199 );
 a128505a <=( A203  and  (not A202) );
 a128506a <=( a128505a  and  a128502a );
 a128507a <=( a128506a  and  a128499a );
 a128510a <=( A266  and  A265 );
 a128513a <=( (not A269)  and  A268 );
 a128514a <=( a128513a  and  a128510a );
 a128517a <=( A299  and  (not A298) );
 a128520a <=( A301  and  (not A300) );
 a128521a <=( a128520a  and  a128517a );
 a128522a <=( a128521a  and  a128514a );
 a128525a <=( A168  and  A169 );
 a128528a <=( A166  and  (not A167) );
 a128529a <=( a128528a  and  a128525a );
 a128532a <=( (not A200)  and  A199 );
 a128535a <=( A203  and  (not A202) );
 a128536a <=( a128535a  and  a128532a );
 a128537a <=( a128536a  and  a128529a );
 a128540a <=( A266  and  A265 );
 a128543a <=( (not A269)  and  A268 );
 a128544a <=( a128543a  and  a128540a );
 a128547a <=( A299  and  (not A298) );
 a128550a <=( (not A302)  and  (not A300) );
 a128551a <=( a128550a  and  a128547a );
 a128552a <=( a128551a  and  a128544a );
 a128555a <=( A168  and  A169 );
 a128558a <=( A166  and  (not A167) );
 a128559a <=( a128558a  and  a128555a );
 a128562a <=( (not A200)  and  A199 );
 a128565a <=( A203  and  (not A202) );
 a128566a <=( a128565a  and  a128562a );
 a128567a <=( a128566a  and  a128559a );
 a128570a <=( A266  and  (not A265) );
 a128573a <=( A269  and  (not A268) );
 a128574a <=( a128573a  and  a128570a );
 a128577a <=( A299  and  A298 );
 a128580a <=( (not A301)  and  (not A300) );
 a128581a <=( a128580a  and  a128577a );
 a128582a <=( a128581a  and  a128574a );
 a128585a <=( A168  and  A169 );
 a128588a <=( A166  and  (not A167) );
 a128589a <=( a128588a  and  a128585a );
 a128592a <=( (not A200)  and  A199 );
 a128595a <=( A203  and  (not A202) );
 a128596a <=( a128595a  and  a128592a );
 a128597a <=( a128596a  and  a128589a );
 a128600a <=( A266  and  (not A265) );
 a128603a <=( A269  and  (not A268) );
 a128604a <=( a128603a  and  a128600a );
 a128607a <=( A299  and  A298 );
 a128610a <=( A302  and  (not A300) );
 a128611a <=( a128610a  and  a128607a );
 a128612a <=( a128611a  and  a128604a );
 a128615a <=( A168  and  A169 );
 a128618a <=( A166  and  (not A167) );
 a128619a <=( a128618a  and  a128615a );
 a128622a <=( (not A200)  and  A199 );
 a128625a <=( A203  and  (not A202) );
 a128626a <=( a128625a  and  a128622a );
 a128627a <=( a128626a  and  a128619a );
 a128630a <=( A266  and  (not A265) );
 a128633a <=( A269  and  (not A268) );
 a128634a <=( a128633a  and  a128630a );
 a128637a <=( (not A299)  and  A298 );
 a128640a <=( A301  and  (not A300) );
 a128641a <=( a128640a  and  a128637a );
 a128642a <=( a128641a  and  a128634a );
 a128645a <=( A168  and  A169 );
 a128648a <=( A166  and  (not A167) );
 a128649a <=( a128648a  and  a128645a );
 a128652a <=( (not A200)  and  A199 );
 a128655a <=( A203  and  (not A202) );
 a128656a <=( a128655a  and  a128652a );
 a128657a <=( a128656a  and  a128649a );
 a128660a <=( A266  and  (not A265) );
 a128663a <=( A269  and  (not A268) );
 a128664a <=( a128663a  and  a128660a );
 a128667a <=( (not A299)  and  A298 );
 a128670a <=( (not A302)  and  (not A300) );
 a128671a <=( a128670a  and  a128667a );
 a128672a <=( a128671a  and  a128664a );
 a128675a <=( A168  and  A169 );
 a128678a <=( A166  and  (not A167) );
 a128679a <=( a128678a  and  a128675a );
 a128682a <=( (not A200)  and  A199 );
 a128685a <=( A203  and  (not A202) );
 a128686a <=( a128685a  and  a128682a );
 a128687a <=( a128686a  and  a128679a );
 a128690a <=( A266  and  (not A265) );
 a128693a <=( A269  and  (not A268) );
 a128694a <=( a128693a  and  a128690a );
 a128697a <=( A299  and  (not A298) );
 a128700a <=( A301  and  (not A300) );
 a128701a <=( a128700a  and  a128697a );
 a128702a <=( a128701a  and  a128694a );
 a128705a <=( A168  and  A169 );
 a128708a <=( A166  and  (not A167) );
 a128709a <=( a128708a  and  a128705a );
 a128712a <=( (not A200)  and  A199 );
 a128715a <=( A203  and  (not A202) );
 a128716a <=( a128715a  and  a128712a );
 a128717a <=( a128716a  and  a128709a );
 a128720a <=( A266  and  (not A265) );
 a128723a <=( A269  and  (not A268) );
 a128724a <=( a128723a  and  a128720a );
 a128727a <=( A299  and  (not A298) );
 a128730a <=( (not A302)  and  (not A300) );
 a128731a <=( a128730a  and  a128727a );
 a128732a <=( a128731a  and  a128724a );
 a128735a <=( A168  and  A169 );
 a128738a <=( A166  and  (not A167) );
 a128739a <=( a128738a  and  a128735a );
 a128742a <=( (not A200)  and  A199 );
 a128745a <=( A203  and  (not A202) );
 a128746a <=( a128745a  and  a128742a );
 a128747a <=( a128746a  and  a128739a );
 a128750a <=( (not A266)  and  A265 );
 a128753a <=( A269  and  (not A268) );
 a128754a <=( a128753a  and  a128750a );
 a128757a <=( A299  and  A298 );
 a128760a <=( (not A301)  and  (not A300) );
 a128761a <=( a128760a  and  a128757a );
 a128762a <=( a128761a  and  a128754a );
 a128765a <=( A168  and  A169 );
 a128768a <=( A166  and  (not A167) );
 a128769a <=( a128768a  and  a128765a );
 a128772a <=( (not A200)  and  A199 );
 a128775a <=( A203  and  (not A202) );
 a128776a <=( a128775a  and  a128772a );
 a128777a <=( a128776a  and  a128769a );
 a128780a <=( (not A266)  and  A265 );
 a128783a <=( A269  and  (not A268) );
 a128784a <=( a128783a  and  a128780a );
 a128787a <=( A299  and  A298 );
 a128790a <=( A302  and  (not A300) );
 a128791a <=( a128790a  and  a128787a );
 a128792a <=( a128791a  and  a128784a );
 a128795a <=( A168  and  A169 );
 a128798a <=( A166  and  (not A167) );
 a128799a <=( a128798a  and  a128795a );
 a128802a <=( (not A200)  and  A199 );
 a128805a <=( A203  and  (not A202) );
 a128806a <=( a128805a  and  a128802a );
 a128807a <=( a128806a  and  a128799a );
 a128810a <=( (not A266)  and  A265 );
 a128813a <=( A269  and  (not A268) );
 a128814a <=( a128813a  and  a128810a );
 a128817a <=( (not A299)  and  A298 );
 a128820a <=( A301  and  (not A300) );
 a128821a <=( a128820a  and  a128817a );
 a128822a <=( a128821a  and  a128814a );
 a128825a <=( A168  and  A169 );
 a128828a <=( A166  and  (not A167) );
 a128829a <=( a128828a  and  a128825a );
 a128832a <=( (not A200)  and  A199 );
 a128835a <=( A203  and  (not A202) );
 a128836a <=( a128835a  and  a128832a );
 a128837a <=( a128836a  and  a128829a );
 a128840a <=( (not A266)  and  A265 );
 a128843a <=( A269  and  (not A268) );
 a128844a <=( a128843a  and  a128840a );
 a128847a <=( (not A299)  and  A298 );
 a128850a <=( (not A302)  and  (not A300) );
 a128851a <=( a128850a  and  a128847a );
 a128852a <=( a128851a  and  a128844a );
 a128855a <=( A168  and  A169 );
 a128858a <=( A166  and  (not A167) );
 a128859a <=( a128858a  and  a128855a );
 a128862a <=( (not A200)  and  A199 );
 a128865a <=( A203  and  (not A202) );
 a128866a <=( a128865a  and  a128862a );
 a128867a <=( a128866a  and  a128859a );
 a128870a <=( (not A266)  and  A265 );
 a128873a <=( A269  and  (not A268) );
 a128874a <=( a128873a  and  a128870a );
 a128877a <=( A299  and  (not A298) );
 a128880a <=( A301  and  (not A300) );
 a128881a <=( a128880a  and  a128877a );
 a128882a <=( a128881a  and  a128874a );
 a128885a <=( A168  and  A169 );
 a128888a <=( A166  and  (not A167) );
 a128889a <=( a128888a  and  a128885a );
 a128892a <=( (not A200)  and  A199 );
 a128895a <=( A203  and  (not A202) );
 a128896a <=( a128895a  and  a128892a );
 a128897a <=( a128896a  and  a128889a );
 a128900a <=( (not A266)  and  A265 );
 a128903a <=( A269  and  (not A268) );
 a128904a <=( a128903a  and  a128900a );
 a128907a <=( A299  and  (not A298) );
 a128910a <=( (not A302)  and  (not A300) );
 a128911a <=( a128910a  and  a128907a );
 a128912a <=( a128911a  and  a128904a );
 a128915a <=( A168  and  A169 );
 a128918a <=( A166  and  (not A167) );
 a128919a <=( a128918a  and  a128915a );
 a128922a <=( (not A200)  and  A199 );
 a128925a <=( A203  and  (not A202) );
 a128926a <=( a128925a  and  a128922a );
 a128927a <=( a128926a  and  a128919a );
 a128930a <=( (not A266)  and  (not A265) );
 a128933a <=( (not A269)  and  A268 );
 a128934a <=( a128933a  and  a128930a );
 a128937a <=( A299  and  A298 );
 a128940a <=( (not A301)  and  (not A300) );
 a128941a <=( a128940a  and  a128937a );
 a128942a <=( a128941a  and  a128934a );
 a128945a <=( A168  and  A169 );
 a128948a <=( A166  and  (not A167) );
 a128949a <=( a128948a  and  a128945a );
 a128952a <=( (not A200)  and  A199 );
 a128955a <=( A203  and  (not A202) );
 a128956a <=( a128955a  and  a128952a );
 a128957a <=( a128956a  and  a128949a );
 a128960a <=( (not A266)  and  (not A265) );
 a128963a <=( (not A269)  and  A268 );
 a128964a <=( a128963a  and  a128960a );
 a128967a <=( A299  and  A298 );
 a128970a <=( A302  and  (not A300) );
 a128971a <=( a128970a  and  a128967a );
 a128972a <=( a128971a  and  a128964a );
 a128975a <=( A168  and  A169 );
 a128978a <=( A166  and  (not A167) );
 a128979a <=( a128978a  and  a128975a );
 a128982a <=( (not A200)  and  A199 );
 a128985a <=( A203  and  (not A202) );
 a128986a <=( a128985a  and  a128982a );
 a128987a <=( a128986a  and  a128979a );
 a128990a <=( (not A266)  and  (not A265) );
 a128993a <=( (not A269)  and  A268 );
 a128994a <=( a128993a  and  a128990a );
 a128997a <=( (not A299)  and  A298 );
 a129000a <=( A301  and  (not A300) );
 a129001a <=( a129000a  and  a128997a );
 a129002a <=( a129001a  and  a128994a );
 a129005a <=( A168  and  A169 );
 a129008a <=( A166  and  (not A167) );
 a129009a <=( a129008a  and  a129005a );
 a129012a <=( (not A200)  and  A199 );
 a129015a <=( A203  and  (not A202) );
 a129016a <=( a129015a  and  a129012a );
 a129017a <=( a129016a  and  a129009a );
 a129020a <=( (not A266)  and  (not A265) );
 a129023a <=( (not A269)  and  A268 );
 a129024a <=( a129023a  and  a129020a );
 a129027a <=( (not A299)  and  A298 );
 a129030a <=( (not A302)  and  (not A300) );
 a129031a <=( a129030a  and  a129027a );
 a129032a <=( a129031a  and  a129024a );
 a129035a <=( A168  and  A169 );
 a129038a <=( A166  and  (not A167) );
 a129039a <=( a129038a  and  a129035a );
 a129042a <=( (not A200)  and  A199 );
 a129045a <=( A203  and  (not A202) );
 a129046a <=( a129045a  and  a129042a );
 a129047a <=( a129046a  and  a129039a );
 a129050a <=( (not A266)  and  (not A265) );
 a129053a <=( (not A269)  and  A268 );
 a129054a <=( a129053a  and  a129050a );
 a129057a <=( A299  and  (not A298) );
 a129060a <=( A301  and  (not A300) );
 a129061a <=( a129060a  and  a129057a );
 a129062a <=( a129061a  and  a129054a );
 a129065a <=( A168  and  A169 );
 a129068a <=( A166  and  (not A167) );
 a129069a <=( a129068a  and  a129065a );
 a129072a <=( (not A200)  and  A199 );
 a129075a <=( A203  and  (not A202) );
 a129076a <=( a129075a  and  a129072a );
 a129077a <=( a129076a  and  a129069a );
 a129080a <=( (not A266)  and  (not A265) );
 a129083a <=( (not A269)  and  A268 );
 a129084a <=( a129083a  and  a129080a );
 a129087a <=( A299  and  (not A298) );
 a129090a <=( (not A302)  and  (not A300) );
 a129091a <=( a129090a  and  a129087a );
 a129092a <=( a129091a  and  a129084a );
 a129095a <=( A168  and  A169 );
 a129098a <=( A166  and  (not A167) );
 a129099a <=( a129098a  and  a129095a );
 a129102a <=( (not A200)  and  A199 );
 a129105a <=( A202  and  (not A201) );
 a129106a <=( a129105a  and  a129102a );
 a129107a <=( a129106a  and  a129099a );
 a129110a <=( A266  and  A265 );
 a129113a <=( (not A268)  and  (not A267) );
 a129114a <=( a129113a  and  a129110a );
 a129117a <=( A299  and  A298 );
 a129120a <=( (not A302)  and  A301 );
 a129121a <=( a129120a  and  a129117a );
 a129122a <=( a129121a  and  a129114a );
 a129125a <=( A168  and  A169 );
 a129128a <=( A166  and  (not A167) );
 a129129a <=( a129128a  and  a129125a );
 a129132a <=( (not A200)  and  A199 );
 a129135a <=( A202  and  (not A201) );
 a129136a <=( a129135a  and  a129132a );
 a129137a <=( a129136a  and  a129129a );
 a129140a <=( A266  and  A265 );
 a129143a <=( (not A268)  and  (not A267) );
 a129144a <=( a129143a  and  a129140a );
 a129147a <=( (not A299)  and  A298 );
 a129150a <=( A302  and  (not A301) );
 a129151a <=( a129150a  and  a129147a );
 a129152a <=( a129151a  and  a129144a );
 a129155a <=( A168  and  A169 );
 a129158a <=( A166  and  (not A167) );
 a129159a <=( a129158a  and  a129155a );
 a129162a <=( (not A200)  and  A199 );
 a129165a <=( A202  and  (not A201) );
 a129166a <=( a129165a  and  a129162a );
 a129167a <=( a129166a  and  a129159a );
 a129170a <=( A266  and  A265 );
 a129173a <=( (not A268)  and  (not A267) );
 a129174a <=( a129173a  and  a129170a );
 a129177a <=( A299  and  (not A298) );
 a129180a <=( A302  and  (not A301) );
 a129181a <=( a129180a  and  a129177a );
 a129182a <=( a129181a  and  a129174a );
 a129185a <=( A168  and  A169 );
 a129188a <=( A166  and  (not A167) );
 a129189a <=( a129188a  and  a129185a );
 a129192a <=( (not A200)  and  A199 );
 a129195a <=( A202  and  (not A201) );
 a129196a <=( a129195a  and  a129192a );
 a129197a <=( a129196a  and  a129189a );
 a129200a <=( A266  and  A265 );
 a129203a <=( (not A268)  and  (not A267) );
 a129204a <=( a129203a  and  a129200a );
 a129207a <=( (not A299)  and  (not A298) );
 a129210a <=( (not A302)  and  A301 );
 a129211a <=( a129210a  and  a129207a );
 a129212a <=( a129211a  and  a129204a );
 a129215a <=( A168  and  A169 );
 a129218a <=( A166  and  (not A167) );
 a129219a <=( a129218a  and  a129215a );
 a129222a <=( (not A200)  and  A199 );
 a129225a <=( A202  and  (not A201) );
 a129226a <=( a129225a  and  a129222a );
 a129227a <=( a129226a  and  a129219a );
 a129230a <=( A266  and  A265 );
 a129233a <=( A269  and  (not A267) );
 a129234a <=( a129233a  and  a129230a );
 a129237a <=( A299  and  A298 );
 a129240a <=( (not A302)  and  A301 );
 a129241a <=( a129240a  and  a129237a );
 a129242a <=( a129241a  and  a129234a );
 a129245a <=( A168  and  A169 );
 a129248a <=( A166  and  (not A167) );
 a129249a <=( a129248a  and  a129245a );
 a129252a <=( (not A200)  and  A199 );
 a129255a <=( A202  and  (not A201) );
 a129256a <=( a129255a  and  a129252a );
 a129257a <=( a129256a  and  a129249a );
 a129260a <=( A266  and  A265 );
 a129263a <=( A269  and  (not A267) );
 a129264a <=( a129263a  and  a129260a );
 a129267a <=( (not A299)  and  A298 );
 a129270a <=( A302  and  (not A301) );
 a129271a <=( a129270a  and  a129267a );
 a129272a <=( a129271a  and  a129264a );
 a129275a <=( A168  and  A169 );
 a129278a <=( A166  and  (not A167) );
 a129279a <=( a129278a  and  a129275a );
 a129282a <=( (not A200)  and  A199 );
 a129285a <=( A202  and  (not A201) );
 a129286a <=( a129285a  and  a129282a );
 a129287a <=( a129286a  and  a129279a );
 a129290a <=( A266  and  A265 );
 a129293a <=( A269  and  (not A267) );
 a129294a <=( a129293a  and  a129290a );
 a129297a <=( A299  and  (not A298) );
 a129300a <=( A302  and  (not A301) );
 a129301a <=( a129300a  and  a129297a );
 a129302a <=( a129301a  and  a129294a );
 a129305a <=( A168  and  A169 );
 a129308a <=( A166  and  (not A167) );
 a129309a <=( a129308a  and  a129305a );
 a129312a <=( (not A200)  and  A199 );
 a129315a <=( A202  and  (not A201) );
 a129316a <=( a129315a  and  a129312a );
 a129317a <=( a129316a  and  a129309a );
 a129320a <=( A266  and  A265 );
 a129323a <=( A269  and  (not A267) );
 a129324a <=( a129323a  and  a129320a );
 a129327a <=( (not A299)  and  (not A298) );
 a129330a <=( (not A302)  and  A301 );
 a129331a <=( a129330a  and  a129327a );
 a129332a <=( a129331a  and  a129324a );
 a129335a <=( A168  and  A169 );
 a129338a <=( A166  and  (not A167) );
 a129339a <=( a129338a  and  a129335a );
 a129342a <=( (not A200)  and  A199 );
 a129345a <=( A202  and  (not A201) );
 a129346a <=( a129345a  and  a129342a );
 a129347a <=( a129346a  and  a129339a );
 a129350a <=( A266  and  (not A265) );
 a129353a <=( A268  and  (not A267) );
 a129354a <=( a129353a  and  a129350a );
 a129357a <=( A299  and  A298 );
 a129360a <=( (not A302)  and  A301 );
 a129361a <=( a129360a  and  a129357a );
 a129362a <=( a129361a  and  a129354a );
 a129365a <=( A168  and  A169 );
 a129368a <=( A166  and  (not A167) );
 a129369a <=( a129368a  and  a129365a );
 a129372a <=( (not A200)  and  A199 );
 a129375a <=( A202  and  (not A201) );
 a129376a <=( a129375a  and  a129372a );
 a129377a <=( a129376a  and  a129369a );
 a129380a <=( A266  and  (not A265) );
 a129383a <=( A268  and  (not A267) );
 a129384a <=( a129383a  and  a129380a );
 a129387a <=( (not A299)  and  A298 );
 a129390a <=( A302  and  (not A301) );
 a129391a <=( a129390a  and  a129387a );
 a129392a <=( a129391a  and  a129384a );
 a129395a <=( A168  and  A169 );
 a129398a <=( A166  and  (not A167) );
 a129399a <=( a129398a  and  a129395a );
 a129402a <=( (not A200)  and  A199 );
 a129405a <=( A202  and  (not A201) );
 a129406a <=( a129405a  and  a129402a );
 a129407a <=( a129406a  and  a129399a );
 a129410a <=( A266  and  (not A265) );
 a129413a <=( A268  and  (not A267) );
 a129414a <=( a129413a  and  a129410a );
 a129417a <=( A299  and  (not A298) );
 a129420a <=( A302  and  (not A301) );
 a129421a <=( a129420a  and  a129417a );
 a129422a <=( a129421a  and  a129414a );
 a129425a <=( A168  and  A169 );
 a129428a <=( A166  and  (not A167) );
 a129429a <=( a129428a  and  a129425a );
 a129432a <=( (not A200)  and  A199 );
 a129435a <=( A202  and  (not A201) );
 a129436a <=( a129435a  and  a129432a );
 a129437a <=( a129436a  and  a129429a );
 a129440a <=( A266  and  (not A265) );
 a129443a <=( A268  and  (not A267) );
 a129444a <=( a129443a  and  a129440a );
 a129447a <=( (not A299)  and  (not A298) );
 a129450a <=( (not A302)  and  A301 );
 a129451a <=( a129450a  and  a129447a );
 a129452a <=( a129451a  and  a129444a );
 a129455a <=( A168  and  A169 );
 a129458a <=( A166  and  (not A167) );
 a129459a <=( a129458a  and  a129455a );
 a129462a <=( (not A200)  and  A199 );
 a129465a <=( A202  and  (not A201) );
 a129466a <=( a129465a  and  a129462a );
 a129467a <=( a129466a  and  a129459a );
 a129470a <=( A266  and  (not A265) );
 a129473a <=( (not A269)  and  (not A267) );
 a129474a <=( a129473a  and  a129470a );
 a129477a <=( A299  and  A298 );
 a129480a <=( (not A302)  and  A301 );
 a129481a <=( a129480a  and  a129477a );
 a129482a <=( a129481a  and  a129474a );
 a129485a <=( A168  and  A169 );
 a129488a <=( A166  and  (not A167) );
 a129489a <=( a129488a  and  a129485a );
 a129492a <=( (not A200)  and  A199 );
 a129495a <=( A202  and  (not A201) );
 a129496a <=( a129495a  and  a129492a );
 a129497a <=( a129496a  and  a129489a );
 a129500a <=( A266  and  (not A265) );
 a129503a <=( (not A269)  and  (not A267) );
 a129504a <=( a129503a  and  a129500a );
 a129507a <=( (not A299)  and  A298 );
 a129510a <=( A302  and  (not A301) );
 a129511a <=( a129510a  and  a129507a );
 a129512a <=( a129511a  and  a129504a );
 a129515a <=( A168  and  A169 );
 a129518a <=( A166  and  (not A167) );
 a129519a <=( a129518a  and  a129515a );
 a129522a <=( (not A200)  and  A199 );
 a129525a <=( A202  and  (not A201) );
 a129526a <=( a129525a  and  a129522a );
 a129527a <=( a129526a  and  a129519a );
 a129530a <=( A266  and  (not A265) );
 a129533a <=( (not A269)  and  (not A267) );
 a129534a <=( a129533a  and  a129530a );
 a129537a <=( A299  and  (not A298) );
 a129540a <=( A302  and  (not A301) );
 a129541a <=( a129540a  and  a129537a );
 a129542a <=( a129541a  and  a129534a );
 a129545a <=( A168  and  A169 );
 a129548a <=( A166  and  (not A167) );
 a129549a <=( a129548a  and  a129545a );
 a129552a <=( (not A200)  and  A199 );
 a129555a <=( A202  and  (not A201) );
 a129556a <=( a129555a  and  a129552a );
 a129557a <=( a129556a  and  a129549a );
 a129560a <=( A266  and  (not A265) );
 a129563a <=( (not A269)  and  (not A267) );
 a129564a <=( a129563a  and  a129560a );
 a129567a <=( (not A299)  and  (not A298) );
 a129570a <=( (not A302)  and  A301 );
 a129571a <=( a129570a  and  a129567a );
 a129572a <=( a129571a  and  a129564a );
 a129575a <=( A168  and  A169 );
 a129578a <=( A166  and  (not A167) );
 a129579a <=( a129578a  and  a129575a );
 a129582a <=( (not A200)  and  A199 );
 a129585a <=( A202  and  (not A201) );
 a129586a <=( a129585a  and  a129582a );
 a129587a <=( a129586a  and  a129579a );
 a129590a <=( (not A266)  and  A265 );
 a129593a <=( A268  and  (not A267) );
 a129594a <=( a129593a  and  a129590a );
 a129597a <=( A299  and  A298 );
 a129600a <=( (not A302)  and  A301 );
 a129601a <=( a129600a  and  a129597a );
 a129602a <=( a129601a  and  a129594a );
 a129605a <=( A168  and  A169 );
 a129608a <=( A166  and  (not A167) );
 a129609a <=( a129608a  and  a129605a );
 a129612a <=( (not A200)  and  A199 );
 a129615a <=( A202  and  (not A201) );
 a129616a <=( a129615a  and  a129612a );
 a129617a <=( a129616a  and  a129609a );
 a129620a <=( (not A266)  and  A265 );
 a129623a <=( A268  and  (not A267) );
 a129624a <=( a129623a  and  a129620a );
 a129627a <=( (not A299)  and  A298 );
 a129630a <=( A302  and  (not A301) );
 a129631a <=( a129630a  and  a129627a );
 a129632a <=( a129631a  and  a129624a );
 a129635a <=( A168  and  A169 );
 a129638a <=( A166  and  (not A167) );
 a129639a <=( a129638a  and  a129635a );
 a129642a <=( (not A200)  and  A199 );
 a129645a <=( A202  and  (not A201) );
 a129646a <=( a129645a  and  a129642a );
 a129647a <=( a129646a  and  a129639a );
 a129650a <=( (not A266)  and  A265 );
 a129653a <=( A268  and  (not A267) );
 a129654a <=( a129653a  and  a129650a );
 a129657a <=( A299  and  (not A298) );
 a129660a <=( A302  and  (not A301) );
 a129661a <=( a129660a  and  a129657a );
 a129662a <=( a129661a  and  a129654a );
 a129665a <=( A168  and  A169 );
 a129668a <=( A166  and  (not A167) );
 a129669a <=( a129668a  and  a129665a );
 a129672a <=( (not A200)  and  A199 );
 a129675a <=( A202  and  (not A201) );
 a129676a <=( a129675a  and  a129672a );
 a129677a <=( a129676a  and  a129669a );
 a129680a <=( (not A266)  and  A265 );
 a129683a <=( A268  and  (not A267) );
 a129684a <=( a129683a  and  a129680a );
 a129687a <=( (not A299)  and  (not A298) );
 a129690a <=( (not A302)  and  A301 );
 a129691a <=( a129690a  and  a129687a );
 a129692a <=( a129691a  and  a129684a );
 a129695a <=( A168  and  A169 );
 a129698a <=( A166  and  (not A167) );
 a129699a <=( a129698a  and  a129695a );
 a129702a <=( (not A200)  and  A199 );
 a129705a <=( A202  and  (not A201) );
 a129706a <=( a129705a  and  a129702a );
 a129707a <=( a129706a  and  a129699a );
 a129710a <=( (not A266)  and  A265 );
 a129713a <=( (not A269)  and  (not A267) );
 a129714a <=( a129713a  and  a129710a );
 a129717a <=( A299  and  A298 );
 a129720a <=( (not A302)  and  A301 );
 a129721a <=( a129720a  and  a129717a );
 a129722a <=( a129721a  and  a129714a );
 a129725a <=( A168  and  A169 );
 a129728a <=( A166  and  (not A167) );
 a129729a <=( a129728a  and  a129725a );
 a129732a <=( (not A200)  and  A199 );
 a129735a <=( A202  and  (not A201) );
 a129736a <=( a129735a  and  a129732a );
 a129737a <=( a129736a  and  a129729a );
 a129740a <=( (not A266)  and  A265 );
 a129743a <=( (not A269)  and  (not A267) );
 a129744a <=( a129743a  and  a129740a );
 a129747a <=( (not A299)  and  A298 );
 a129750a <=( A302  and  (not A301) );
 a129751a <=( a129750a  and  a129747a );
 a129752a <=( a129751a  and  a129744a );
 a129755a <=( A168  and  A169 );
 a129758a <=( A166  and  (not A167) );
 a129759a <=( a129758a  and  a129755a );
 a129762a <=( (not A200)  and  A199 );
 a129765a <=( A202  and  (not A201) );
 a129766a <=( a129765a  and  a129762a );
 a129767a <=( a129766a  and  a129759a );
 a129770a <=( (not A266)  and  A265 );
 a129773a <=( (not A269)  and  (not A267) );
 a129774a <=( a129773a  and  a129770a );
 a129777a <=( A299  and  (not A298) );
 a129780a <=( A302  and  (not A301) );
 a129781a <=( a129780a  and  a129777a );
 a129782a <=( a129781a  and  a129774a );
 a129785a <=( A168  and  A169 );
 a129788a <=( A166  and  (not A167) );
 a129789a <=( a129788a  and  a129785a );
 a129792a <=( (not A200)  and  A199 );
 a129795a <=( A202  and  (not A201) );
 a129796a <=( a129795a  and  a129792a );
 a129797a <=( a129796a  and  a129789a );
 a129800a <=( (not A266)  and  A265 );
 a129803a <=( (not A269)  and  (not A267) );
 a129804a <=( a129803a  and  a129800a );
 a129807a <=( (not A299)  and  (not A298) );
 a129810a <=( (not A302)  and  A301 );
 a129811a <=( a129810a  and  a129807a );
 a129812a <=( a129811a  and  a129804a );
 a129815a <=( A168  and  A169 );
 a129818a <=( A166  and  (not A167) );
 a129819a <=( a129818a  and  a129815a );
 a129822a <=( (not A200)  and  A199 );
 a129825a <=( (not A203)  and  (not A201) );
 a129826a <=( a129825a  and  a129822a );
 a129827a <=( a129826a  and  a129819a );
 a129830a <=( A266  and  A265 );
 a129833a <=( (not A268)  and  (not A267) );
 a129834a <=( a129833a  and  a129830a );
 a129837a <=( A299  and  A298 );
 a129840a <=( (not A302)  and  A301 );
 a129841a <=( a129840a  and  a129837a );
 a129842a <=( a129841a  and  a129834a );
 a129845a <=( A168  and  A169 );
 a129848a <=( A166  and  (not A167) );
 a129849a <=( a129848a  and  a129845a );
 a129852a <=( (not A200)  and  A199 );
 a129855a <=( (not A203)  and  (not A201) );
 a129856a <=( a129855a  and  a129852a );
 a129857a <=( a129856a  and  a129849a );
 a129860a <=( A266  and  A265 );
 a129863a <=( (not A268)  and  (not A267) );
 a129864a <=( a129863a  and  a129860a );
 a129867a <=( (not A299)  and  A298 );
 a129870a <=( A302  and  (not A301) );
 a129871a <=( a129870a  and  a129867a );
 a129872a <=( a129871a  and  a129864a );
 a129875a <=( A168  and  A169 );
 a129878a <=( A166  and  (not A167) );
 a129879a <=( a129878a  and  a129875a );
 a129882a <=( (not A200)  and  A199 );
 a129885a <=( (not A203)  and  (not A201) );
 a129886a <=( a129885a  and  a129882a );
 a129887a <=( a129886a  and  a129879a );
 a129890a <=( A266  and  A265 );
 a129893a <=( (not A268)  and  (not A267) );
 a129894a <=( a129893a  and  a129890a );
 a129897a <=( A299  and  (not A298) );
 a129900a <=( A302  and  (not A301) );
 a129901a <=( a129900a  and  a129897a );
 a129902a <=( a129901a  and  a129894a );
 a129905a <=( A168  and  A169 );
 a129908a <=( A166  and  (not A167) );
 a129909a <=( a129908a  and  a129905a );
 a129912a <=( (not A200)  and  A199 );
 a129915a <=( (not A203)  and  (not A201) );
 a129916a <=( a129915a  and  a129912a );
 a129917a <=( a129916a  and  a129909a );
 a129920a <=( A266  and  A265 );
 a129923a <=( (not A268)  and  (not A267) );
 a129924a <=( a129923a  and  a129920a );
 a129927a <=( (not A299)  and  (not A298) );
 a129930a <=( (not A302)  and  A301 );
 a129931a <=( a129930a  and  a129927a );
 a129932a <=( a129931a  and  a129924a );
 a129935a <=( A168  and  A169 );
 a129938a <=( A166  and  (not A167) );
 a129939a <=( a129938a  and  a129935a );
 a129942a <=( (not A200)  and  A199 );
 a129945a <=( (not A203)  and  (not A201) );
 a129946a <=( a129945a  and  a129942a );
 a129947a <=( a129946a  and  a129939a );
 a129950a <=( A266  and  A265 );
 a129953a <=( A269  and  (not A267) );
 a129954a <=( a129953a  and  a129950a );
 a129957a <=( A299  and  A298 );
 a129960a <=( (not A302)  and  A301 );
 a129961a <=( a129960a  and  a129957a );
 a129962a <=( a129961a  and  a129954a );
 a129965a <=( A168  and  A169 );
 a129968a <=( A166  and  (not A167) );
 a129969a <=( a129968a  and  a129965a );
 a129972a <=( (not A200)  and  A199 );
 a129975a <=( (not A203)  and  (not A201) );
 a129976a <=( a129975a  and  a129972a );
 a129977a <=( a129976a  and  a129969a );
 a129980a <=( A266  and  A265 );
 a129983a <=( A269  and  (not A267) );
 a129984a <=( a129983a  and  a129980a );
 a129987a <=( (not A299)  and  A298 );
 a129990a <=( A302  and  (not A301) );
 a129991a <=( a129990a  and  a129987a );
 a129992a <=( a129991a  and  a129984a );
 a129995a <=( A168  and  A169 );
 a129998a <=( A166  and  (not A167) );
 a129999a <=( a129998a  and  a129995a );
 a130002a <=( (not A200)  and  A199 );
 a130005a <=( (not A203)  and  (not A201) );
 a130006a <=( a130005a  and  a130002a );
 a130007a <=( a130006a  and  a129999a );
 a130010a <=( A266  and  A265 );
 a130013a <=( A269  and  (not A267) );
 a130014a <=( a130013a  and  a130010a );
 a130017a <=( A299  and  (not A298) );
 a130020a <=( A302  and  (not A301) );
 a130021a <=( a130020a  and  a130017a );
 a130022a <=( a130021a  and  a130014a );
 a130025a <=( A168  and  A169 );
 a130028a <=( A166  and  (not A167) );
 a130029a <=( a130028a  and  a130025a );
 a130032a <=( (not A200)  and  A199 );
 a130035a <=( (not A203)  and  (not A201) );
 a130036a <=( a130035a  and  a130032a );
 a130037a <=( a130036a  and  a130029a );
 a130040a <=( A266  and  A265 );
 a130043a <=( A269  and  (not A267) );
 a130044a <=( a130043a  and  a130040a );
 a130047a <=( (not A299)  and  (not A298) );
 a130050a <=( (not A302)  and  A301 );
 a130051a <=( a130050a  and  a130047a );
 a130052a <=( a130051a  and  a130044a );
 a130055a <=( A168  and  A169 );
 a130058a <=( A166  and  (not A167) );
 a130059a <=( a130058a  and  a130055a );
 a130062a <=( (not A200)  and  A199 );
 a130065a <=( (not A203)  and  (not A201) );
 a130066a <=( a130065a  and  a130062a );
 a130067a <=( a130066a  and  a130059a );
 a130070a <=( A266  and  (not A265) );
 a130073a <=( A268  and  (not A267) );
 a130074a <=( a130073a  and  a130070a );
 a130077a <=( A299  and  A298 );
 a130080a <=( (not A302)  and  A301 );
 a130081a <=( a130080a  and  a130077a );
 a130082a <=( a130081a  and  a130074a );
 a130085a <=( A168  and  A169 );
 a130088a <=( A166  and  (not A167) );
 a130089a <=( a130088a  and  a130085a );
 a130092a <=( (not A200)  and  A199 );
 a130095a <=( (not A203)  and  (not A201) );
 a130096a <=( a130095a  and  a130092a );
 a130097a <=( a130096a  and  a130089a );
 a130100a <=( A266  and  (not A265) );
 a130103a <=( A268  and  (not A267) );
 a130104a <=( a130103a  and  a130100a );
 a130107a <=( (not A299)  and  A298 );
 a130110a <=( A302  and  (not A301) );
 a130111a <=( a130110a  and  a130107a );
 a130112a <=( a130111a  and  a130104a );
 a130115a <=( A168  and  A169 );
 a130118a <=( A166  and  (not A167) );
 a130119a <=( a130118a  and  a130115a );
 a130122a <=( (not A200)  and  A199 );
 a130125a <=( (not A203)  and  (not A201) );
 a130126a <=( a130125a  and  a130122a );
 a130127a <=( a130126a  and  a130119a );
 a130130a <=( A266  and  (not A265) );
 a130133a <=( A268  and  (not A267) );
 a130134a <=( a130133a  and  a130130a );
 a130137a <=( A299  and  (not A298) );
 a130140a <=( A302  and  (not A301) );
 a130141a <=( a130140a  and  a130137a );
 a130142a <=( a130141a  and  a130134a );
 a130145a <=( A168  and  A169 );
 a130148a <=( A166  and  (not A167) );
 a130149a <=( a130148a  and  a130145a );
 a130152a <=( (not A200)  and  A199 );
 a130155a <=( (not A203)  and  (not A201) );
 a130156a <=( a130155a  and  a130152a );
 a130157a <=( a130156a  and  a130149a );
 a130160a <=( A266  and  (not A265) );
 a130163a <=( A268  and  (not A267) );
 a130164a <=( a130163a  and  a130160a );
 a130167a <=( (not A299)  and  (not A298) );
 a130170a <=( (not A302)  and  A301 );
 a130171a <=( a130170a  and  a130167a );
 a130172a <=( a130171a  and  a130164a );
 a130175a <=( A168  and  A169 );
 a130178a <=( A166  and  (not A167) );
 a130179a <=( a130178a  and  a130175a );
 a130182a <=( (not A200)  and  A199 );
 a130185a <=( (not A203)  and  (not A201) );
 a130186a <=( a130185a  and  a130182a );
 a130187a <=( a130186a  and  a130179a );
 a130190a <=( A266  and  (not A265) );
 a130193a <=( (not A269)  and  (not A267) );
 a130194a <=( a130193a  and  a130190a );
 a130197a <=( A299  and  A298 );
 a130200a <=( (not A302)  and  A301 );
 a130201a <=( a130200a  and  a130197a );
 a130202a <=( a130201a  and  a130194a );
 a130205a <=( A168  and  A169 );
 a130208a <=( A166  and  (not A167) );
 a130209a <=( a130208a  and  a130205a );
 a130212a <=( (not A200)  and  A199 );
 a130215a <=( (not A203)  and  (not A201) );
 a130216a <=( a130215a  and  a130212a );
 a130217a <=( a130216a  and  a130209a );
 a130220a <=( A266  and  (not A265) );
 a130223a <=( (not A269)  and  (not A267) );
 a130224a <=( a130223a  and  a130220a );
 a130227a <=( (not A299)  and  A298 );
 a130230a <=( A302  and  (not A301) );
 a130231a <=( a130230a  and  a130227a );
 a130232a <=( a130231a  and  a130224a );
 a130235a <=( A168  and  A169 );
 a130238a <=( A166  and  (not A167) );
 a130239a <=( a130238a  and  a130235a );
 a130242a <=( (not A200)  and  A199 );
 a130245a <=( (not A203)  and  (not A201) );
 a130246a <=( a130245a  and  a130242a );
 a130247a <=( a130246a  and  a130239a );
 a130250a <=( A266  and  (not A265) );
 a130253a <=( (not A269)  and  (not A267) );
 a130254a <=( a130253a  and  a130250a );
 a130257a <=( A299  and  (not A298) );
 a130260a <=( A302  and  (not A301) );
 a130261a <=( a130260a  and  a130257a );
 a130262a <=( a130261a  and  a130254a );
 a130265a <=( A168  and  A169 );
 a130268a <=( A166  and  (not A167) );
 a130269a <=( a130268a  and  a130265a );
 a130272a <=( (not A200)  and  A199 );
 a130275a <=( (not A203)  and  (not A201) );
 a130276a <=( a130275a  and  a130272a );
 a130277a <=( a130276a  and  a130269a );
 a130280a <=( A266  and  (not A265) );
 a130283a <=( (not A269)  and  (not A267) );
 a130284a <=( a130283a  and  a130280a );
 a130287a <=( (not A299)  and  (not A298) );
 a130290a <=( (not A302)  and  A301 );
 a130291a <=( a130290a  and  a130287a );
 a130292a <=( a130291a  and  a130284a );
 a130295a <=( A168  and  A169 );
 a130298a <=( A166  and  (not A167) );
 a130299a <=( a130298a  and  a130295a );
 a130302a <=( (not A200)  and  A199 );
 a130305a <=( (not A203)  and  (not A201) );
 a130306a <=( a130305a  and  a130302a );
 a130307a <=( a130306a  and  a130299a );
 a130310a <=( (not A266)  and  A265 );
 a130313a <=( A268  and  (not A267) );
 a130314a <=( a130313a  and  a130310a );
 a130317a <=( A299  and  A298 );
 a130320a <=( (not A302)  and  A301 );
 a130321a <=( a130320a  and  a130317a );
 a130322a <=( a130321a  and  a130314a );
 a130325a <=( A168  and  A169 );
 a130328a <=( A166  and  (not A167) );
 a130329a <=( a130328a  and  a130325a );
 a130332a <=( (not A200)  and  A199 );
 a130335a <=( (not A203)  and  (not A201) );
 a130336a <=( a130335a  and  a130332a );
 a130337a <=( a130336a  and  a130329a );
 a130340a <=( (not A266)  and  A265 );
 a130343a <=( A268  and  (not A267) );
 a130344a <=( a130343a  and  a130340a );
 a130347a <=( (not A299)  and  A298 );
 a130350a <=( A302  and  (not A301) );
 a130351a <=( a130350a  and  a130347a );
 a130352a <=( a130351a  and  a130344a );
 a130355a <=( A168  and  A169 );
 a130358a <=( A166  and  (not A167) );
 a130359a <=( a130358a  and  a130355a );
 a130362a <=( (not A200)  and  A199 );
 a130365a <=( (not A203)  and  (not A201) );
 a130366a <=( a130365a  and  a130362a );
 a130367a <=( a130366a  and  a130359a );
 a130370a <=( (not A266)  and  A265 );
 a130373a <=( A268  and  (not A267) );
 a130374a <=( a130373a  and  a130370a );
 a130377a <=( A299  and  (not A298) );
 a130380a <=( A302  and  (not A301) );
 a130381a <=( a130380a  and  a130377a );
 a130382a <=( a130381a  and  a130374a );
 a130385a <=( A168  and  A169 );
 a130388a <=( A166  and  (not A167) );
 a130389a <=( a130388a  and  a130385a );
 a130392a <=( (not A200)  and  A199 );
 a130395a <=( (not A203)  and  (not A201) );
 a130396a <=( a130395a  and  a130392a );
 a130397a <=( a130396a  and  a130389a );
 a130400a <=( (not A266)  and  A265 );
 a130403a <=( A268  and  (not A267) );
 a130404a <=( a130403a  and  a130400a );
 a130407a <=( (not A299)  and  (not A298) );
 a130410a <=( (not A302)  and  A301 );
 a130411a <=( a130410a  and  a130407a );
 a130412a <=( a130411a  and  a130404a );
 a130415a <=( A168  and  A169 );
 a130418a <=( A166  and  (not A167) );
 a130419a <=( a130418a  and  a130415a );
 a130422a <=( (not A200)  and  A199 );
 a130425a <=( (not A203)  and  (not A201) );
 a130426a <=( a130425a  and  a130422a );
 a130427a <=( a130426a  and  a130419a );
 a130430a <=( (not A266)  and  A265 );
 a130433a <=( (not A269)  and  (not A267) );
 a130434a <=( a130433a  and  a130430a );
 a130437a <=( A299  and  A298 );
 a130440a <=( (not A302)  and  A301 );
 a130441a <=( a130440a  and  a130437a );
 a130442a <=( a130441a  and  a130434a );
 a130445a <=( A168  and  A169 );
 a130448a <=( A166  and  (not A167) );
 a130449a <=( a130448a  and  a130445a );
 a130452a <=( (not A200)  and  A199 );
 a130455a <=( (not A203)  and  (not A201) );
 a130456a <=( a130455a  and  a130452a );
 a130457a <=( a130456a  and  a130449a );
 a130460a <=( (not A266)  and  A265 );
 a130463a <=( (not A269)  and  (not A267) );
 a130464a <=( a130463a  and  a130460a );
 a130467a <=( (not A299)  and  A298 );
 a130470a <=( A302  and  (not A301) );
 a130471a <=( a130470a  and  a130467a );
 a130472a <=( a130471a  and  a130464a );
 a130475a <=( A168  and  A169 );
 a130478a <=( A166  and  (not A167) );
 a130479a <=( a130478a  and  a130475a );
 a130482a <=( (not A200)  and  A199 );
 a130485a <=( (not A203)  and  (not A201) );
 a130486a <=( a130485a  and  a130482a );
 a130487a <=( a130486a  and  a130479a );
 a130490a <=( (not A266)  and  A265 );
 a130493a <=( (not A269)  and  (not A267) );
 a130494a <=( a130493a  and  a130490a );
 a130497a <=( A299  and  (not A298) );
 a130500a <=( A302  and  (not A301) );
 a130501a <=( a130500a  and  a130497a );
 a130502a <=( a130501a  and  a130494a );
 a130505a <=( A168  and  A169 );
 a130508a <=( A166  and  (not A167) );
 a130509a <=( a130508a  and  a130505a );
 a130512a <=( (not A200)  and  A199 );
 a130515a <=( (not A203)  and  (not A201) );
 a130516a <=( a130515a  and  a130512a );
 a130517a <=( a130516a  and  a130509a );
 a130520a <=( (not A266)  and  A265 );
 a130523a <=( (not A269)  and  (not A267) );
 a130524a <=( a130523a  and  a130520a );
 a130527a <=( (not A299)  and  (not A298) );
 a130530a <=( (not A302)  and  A301 );
 a130531a <=( a130530a  and  a130527a );
 a130532a <=( a130531a  and  a130524a );
 a130535a <=( A168  and  A169 );
 a130538a <=( A166  and  (not A167) );
 a130539a <=( a130538a  and  a130535a );
 a130542a <=( (not A200)  and  (not A199) );
 a130545a <=( (not A203)  and  A202 );
 a130546a <=( a130545a  and  a130542a );
 a130547a <=( a130546a  and  a130539a );
 a130550a <=( A266  and  A265 );
 a130553a <=( (not A269)  and  A268 );
 a130554a <=( a130553a  and  a130550a );
 a130557a <=( A299  and  A298 );
 a130560a <=( (not A301)  and  (not A300) );
 a130561a <=( a130560a  and  a130557a );
 a130562a <=( a130561a  and  a130554a );
 a130565a <=( A168  and  A169 );
 a130568a <=( A166  and  (not A167) );
 a130569a <=( a130568a  and  a130565a );
 a130572a <=( (not A200)  and  (not A199) );
 a130575a <=( (not A203)  and  A202 );
 a130576a <=( a130575a  and  a130572a );
 a130577a <=( a130576a  and  a130569a );
 a130580a <=( A266  and  A265 );
 a130583a <=( (not A269)  and  A268 );
 a130584a <=( a130583a  and  a130580a );
 a130587a <=( A299  and  A298 );
 a130590a <=( A302  and  (not A300) );
 a130591a <=( a130590a  and  a130587a );
 a130592a <=( a130591a  and  a130584a );
 a130595a <=( A168  and  A169 );
 a130598a <=( A166  and  (not A167) );
 a130599a <=( a130598a  and  a130595a );
 a130602a <=( (not A200)  and  (not A199) );
 a130605a <=( (not A203)  and  A202 );
 a130606a <=( a130605a  and  a130602a );
 a130607a <=( a130606a  and  a130599a );
 a130610a <=( A266  and  A265 );
 a130613a <=( (not A269)  and  A268 );
 a130614a <=( a130613a  and  a130610a );
 a130617a <=( (not A299)  and  A298 );
 a130620a <=( A301  and  (not A300) );
 a130621a <=( a130620a  and  a130617a );
 a130622a <=( a130621a  and  a130614a );
 a130625a <=( A168  and  A169 );
 a130628a <=( A166  and  (not A167) );
 a130629a <=( a130628a  and  a130625a );
 a130632a <=( (not A200)  and  (not A199) );
 a130635a <=( (not A203)  and  A202 );
 a130636a <=( a130635a  and  a130632a );
 a130637a <=( a130636a  and  a130629a );
 a130640a <=( A266  and  A265 );
 a130643a <=( (not A269)  and  A268 );
 a130644a <=( a130643a  and  a130640a );
 a130647a <=( (not A299)  and  A298 );
 a130650a <=( (not A302)  and  (not A300) );
 a130651a <=( a130650a  and  a130647a );
 a130652a <=( a130651a  and  a130644a );
 a130655a <=( A168  and  A169 );
 a130658a <=( A166  and  (not A167) );
 a130659a <=( a130658a  and  a130655a );
 a130662a <=( (not A200)  and  (not A199) );
 a130665a <=( (not A203)  and  A202 );
 a130666a <=( a130665a  and  a130662a );
 a130667a <=( a130666a  and  a130659a );
 a130670a <=( A266  and  A265 );
 a130673a <=( (not A269)  and  A268 );
 a130674a <=( a130673a  and  a130670a );
 a130677a <=( A299  and  (not A298) );
 a130680a <=( A301  and  (not A300) );
 a130681a <=( a130680a  and  a130677a );
 a130682a <=( a130681a  and  a130674a );
 a130685a <=( A168  and  A169 );
 a130688a <=( A166  and  (not A167) );
 a130689a <=( a130688a  and  a130685a );
 a130692a <=( (not A200)  and  (not A199) );
 a130695a <=( (not A203)  and  A202 );
 a130696a <=( a130695a  and  a130692a );
 a130697a <=( a130696a  and  a130689a );
 a130700a <=( A266  and  A265 );
 a130703a <=( (not A269)  and  A268 );
 a130704a <=( a130703a  and  a130700a );
 a130707a <=( A299  and  (not A298) );
 a130710a <=( (not A302)  and  (not A300) );
 a130711a <=( a130710a  and  a130707a );
 a130712a <=( a130711a  and  a130704a );
 a130715a <=( A168  and  A169 );
 a130718a <=( A166  and  (not A167) );
 a130719a <=( a130718a  and  a130715a );
 a130722a <=( (not A200)  and  (not A199) );
 a130725a <=( (not A203)  and  A202 );
 a130726a <=( a130725a  and  a130722a );
 a130727a <=( a130726a  and  a130719a );
 a130730a <=( A266  and  (not A265) );
 a130733a <=( A269  and  (not A268) );
 a130734a <=( a130733a  and  a130730a );
 a130737a <=( A299  and  A298 );
 a130740a <=( (not A301)  and  (not A300) );
 a130741a <=( a130740a  and  a130737a );
 a130742a <=( a130741a  and  a130734a );
 a130745a <=( A168  and  A169 );
 a130748a <=( A166  and  (not A167) );
 a130749a <=( a130748a  and  a130745a );
 a130752a <=( (not A200)  and  (not A199) );
 a130755a <=( (not A203)  and  A202 );
 a130756a <=( a130755a  and  a130752a );
 a130757a <=( a130756a  and  a130749a );
 a130760a <=( A266  and  (not A265) );
 a130763a <=( A269  and  (not A268) );
 a130764a <=( a130763a  and  a130760a );
 a130767a <=( A299  and  A298 );
 a130770a <=( A302  and  (not A300) );
 a130771a <=( a130770a  and  a130767a );
 a130772a <=( a130771a  and  a130764a );
 a130775a <=( A168  and  A169 );
 a130778a <=( A166  and  (not A167) );
 a130779a <=( a130778a  and  a130775a );
 a130782a <=( (not A200)  and  (not A199) );
 a130785a <=( (not A203)  and  A202 );
 a130786a <=( a130785a  and  a130782a );
 a130787a <=( a130786a  and  a130779a );
 a130790a <=( A266  and  (not A265) );
 a130793a <=( A269  and  (not A268) );
 a130794a <=( a130793a  and  a130790a );
 a130797a <=( (not A299)  and  A298 );
 a130800a <=( A301  and  (not A300) );
 a130801a <=( a130800a  and  a130797a );
 a130802a <=( a130801a  and  a130794a );
 a130805a <=( A168  and  A169 );
 a130808a <=( A166  and  (not A167) );
 a130809a <=( a130808a  and  a130805a );
 a130812a <=( (not A200)  and  (not A199) );
 a130815a <=( (not A203)  and  A202 );
 a130816a <=( a130815a  and  a130812a );
 a130817a <=( a130816a  and  a130809a );
 a130820a <=( A266  and  (not A265) );
 a130823a <=( A269  and  (not A268) );
 a130824a <=( a130823a  and  a130820a );
 a130827a <=( (not A299)  and  A298 );
 a130830a <=( (not A302)  and  (not A300) );
 a130831a <=( a130830a  and  a130827a );
 a130832a <=( a130831a  and  a130824a );
 a130835a <=( A168  and  A169 );
 a130838a <=( A166  and  (not A167) );
 a130839a <=( a130838a  and  a130835a );
 a130842a <=( (not A200)  and  (not A199) );
 a130845a <=( (not A203)  and  A202 );
 a130846a <=( a130845a  and  a130842a );
 a130847a <=( a130846a  and  a130839a );
 a130850a <=( A266  and  (not A265) );
 a130853a <=( A269  and  (not A268) );
 a130854a <=( a130853a  and  a130850a );
 a130857a <=( A299  and  (not A298) );
 a130860a <=( A301  and  (not A300) );
 a130861a <=( a130860a  and  a130857a );
 a130862a <=( a130861a  and  a130854a );
 a130865a <=( A168  and  A169 );
 a130868a <=( A166  and  (not A167) );
 a130869a <=( a130868a  and  a130865a );
 a130872a <=( (not A200)  and  (not A199) );
 a130875a <=( (not A203)  and  A202 );
 a130876a <=( a130875a  and  a130872a );
 a130877a <=( a130876a  and  a130869a );
 a130880a <=( A266  and  (not A265) );
 a130883a <=( A269  and  (not A268) );
 a130884a <=( a130883a  and  a130880a );
 a130887a <=( A299  and  (not A298) );
 a130890a <=( (not A302)  and  (not A300) );
 a130891a <=( a130890a  and  a130887a );
 a130892a <=( a130891a  and  a130884a );
 a130895a <=( A168  and  A169 );
 a130898a <=( A166  and  (not A167) );
 a130899a <=( a130898a  and  a130895a );
 a130902a <=( (not A200)  and  (not A199) );
 a130905a <=( (not A203)  and  A202 );
 a130906a <=( a130905a  and  a130902a );
 a130907a <=( a130906a  and  a130899a );
 a130910a <=( (not A266)  and  A265 );
 a130913a <=( A269  and  (not A268) );
 a130914a <=( a130913a  and  a130910a );
 a130917a <=( A299  and  A298 );
 a130920a <=( (not A301)  and  (not A300) );
 a130921a <=( a130920a  and  a130917a );
 a130922a <=( a130921a  and  a130914a );
 a130925a <=( A168  and  A169 );
 a130928a <=( A166  and  (not A167) );
 a130929a <=( a130928a  and  a130925a );
 a130932a <=( (not A200)  and  (not A199) );
 a130935a <=( (not A203)  and  A202 );
 a130936a <=( a130935a  and  a130932a );
 a130937a <=( a130936a  and  a130929a );
 a130940a <=( (not A266)  and  A265 );
 a130943a <=( A269  and  (not A268) );
 a130944a <=( a130943a  and  a130940a );
 a130947a <=( A299  and  A298 );
 a130950a <=( A302  and  (not A300) );
 a130951a <=( a130950a  and  a130947a );
 a130952a <=( a130951a  and  a130944a );
 a130955a <=( A168  and  A169 );
 a130958a <=( A166  and  (not A167) );
 a130959a <=( a130958a  and  a130955a );
 a130962a <=( (not A200)  and  (not A199) );
 a130965a <=( (not A203)  and  A202 );
 a130966a <=( a130965a  and  a130962a );
 a130967a <=( a130966a  and  a130959a );
 a130970a <=( (not A266)  and  A265 );
 a130973a <=( A269  and  (not A268) );
 a130974a <=( a130973a  and  a130970a );
 a130977a <=( (not A299)  and  A298 );
 a130980a <=( A301  and  (not A300) );
 a130981a <=( a130980a  and  a130977a );
 a130982a <=( a130981a  and  a130974a );
 a130985a <=( A168  and  A169 );
 a130988a <=( A166  and  (not A167) );
 a130989a <=( a130988a  and  a130985a );
 a130992a <=( (not A200)  and  (not A199) );
 a130995a <=( (not A203)  and  A202 );
 a130996a <=( a130995a  and  a130992a );
 a130997a <=( a130996a  and  a130989a );
 a131000a <=( (not A266)  and  A265 );
 a131003a <=( A269  and  (not A268) );
 a131004a <=( a131003a  and  a131000a );
 a131007a <=( (not A299)  and  A298 );
 a131010a <=( (not A302)  and  (not A300) );
 a131011a <=( a131010a  and  a131007a );
 a131012a <=( a131011a  and  a131004a );
 a131015a <=( A168  and  A169 );
 a131018a <=( A166  and  (not A167) );
 a131019a <=( a131018a  and  a131015a );
 a131022a <=( (not A200)  and  (not A199) );
 a131025a <=( (not A203)  and  A202 );
 a131026a <=( a131025a  and  a131022a );
 a131027a <=( a131026a  and  a131019a );
 a131030a <=( (not A266)  and  A265 );
 a131033a <=( A269  and  (not A268) );
 a131034a <=( a131033a  and  a131030a );
 a131037a <=( A299  and  (not A298) );
 a131040a <=( A301  and  (not A300) );
 a131041a <=( a131040a  and  a131037a );
 a131042a <=( a131041a  and  a131034a );
 a131045a <=( A168  and  A169 );
 a131048a <=( A166  and  (not A167) );
 a131049a <=( a131048a  and  a131045a );
 a131052a <=( (not A200)  and  (not A199) );
 a131055a <=( (not A203)  and  A202 );
 a131056a <=( a131055a  and  a131052a );
 a131057a <=( a131056a  and  a131049a );
 a131060a <=( (not A266)  and  A265 );
 a131063a <=( A269  and  (not A268) );
 a131064a <=( a131063a  and  a131060a );
 a131067a <=( A299  and  (not A298) );
 a131070a <=( (not A302)  and  (not A300) );
 a131071a <=( a131070a  and  a131067a );
 a131072a <=( a131071a  and  a131064a );
 a131075a <=( A168  and  A169 );
 a131078a <=( A166  and  (not A167) );
 a131079a <=( a131078a  and  a131075a );
 a131082a <=( (not A200)  and  (not A199) );
 a131085a <=( (not A203)  and  A202 );
 a131086a <=( a131085a  and  a131082a );
 a131087a <=( a131086a  and  a131079a );
 a131090a <=( (not A266)  and  (not A265) );
 a131093a <=( (not A269)  and  A268 );
 a131094a <=( a131093a  and  a131090a );
 a131097a <=( A299  and  A298 );
 a131100a <=( (not A301)  and  (not A300) );
 a131101a <=( a131100a  and  a131097a );
 a131102a <=( a131101a  and  a131094a );
 a131105a <=( A168  and  A169 );
 a131108a <=( A166  and  (not A167) );
 a131109a <=( a131108a  and  a131105a );
 a131112a <=( (not A200)  and  (not A199) );
 a131115a <=( (not A203)  and  A202 );
 a131116a <=( a131115a  and  a131112a );
 a131117a <=( a131116a  and  a131109a );
 a131120a <=( (not A266)  and  (not A265) );
 a131123a <=( (not A269)  and  A268 );
 a131124a <=( a131123a  and  a131120a );
 a131127a <=( A299  and  A298 );
 a131130a <=( A302  and  (not A300) );
 a131131a <=( a131130a  and  a131127a );
 a131132a <=( a131131a  and  a131124a );
 a131135a <=( A168  and  A169 );
 a131138a <=( A166  and  (not A167) );
 a131139a <=( a131138a  and  a131135a );
 a131142a <=( (not A200)  and  (not A199) );
 a131145a <=( (not A203)  and  A202 );
 a131146a <=( a131145a  and  a131142a );
 a131147a <=( a131146a  and  a131139a );
 a131150a <=( (not A266)  and  (not A265) );
 a131153a <=( (not A269)  and  A268 );
 a131154a <=( a131153a  and  a131150a );
 a131157a <=( (not A299)  and  A298 );
 a131160a <=( A301  and  (not A300) );
 a131161a <=( a131160a  and  a131157a );
 a131162a <=( a131161a  and  a131154a );
 a131165a <=( A168  and  A169 );
 a131168a <=( A166  and  (not A167) );
 a131169a <=( a131168a  and  a131165a );
 a131172a <=( (not A200)  and  (not A199) );
 a131175a <=( (not A203)  and  A202 );
 a131176a <=( a131175a  and  a131172a );
 a131177a <=( a131176a  and  a131169a );
 a131180a <=( (not A266)  and  (not A265) );
 a131183a <=( (not A269)  and  A268 );
 a131184a <=( a131183a  and  a131180a );
 a131187a <=( (not A299)  and  A298 );
 a131190a <=( (not A302)  and  (not A300) );
 a131191a <=( a131190a  and  a131187a );
 a131192a <=( a131191a  and  a131184a );
 a131195a <=( A168  and  A169 );
 a131198a <=( A166  and  (not A167) );
 a131199a <=( a131198a  and  a131195a );
 a131202a <=( (not A200)  and  (not A199) );
 a131205a <=( (not A203)  and  A202 );
 a131206a <=( a131205a  and  a131202a );
 a131207a <=( a131206a  and  a131199a );
 a131210a <=( (not A266)  and  (not A265) );
 a131213a <=( (not A269)  and  A268 );
 a131214a <=( a131213a  and  a131210a );
 a131217a <=( A299  and  (not A298) );
 a131220a <=( A301  and  (not A300) );
 a131221a <=( a131220a  and  a131217a );
 a131222a <=( a131221a  and  a131214a );
 a131225a <=( A168  and  A169 );
 a131228a <=( A166  and  (not A167) );
 a131229a <=( a131228a  and  a131225a );
 a131232a <=( (not A200)  and  (not A199) );
 a131235a <=( (not A203)  and  A202 );
 a131236a <=( a131235a  and  a131232a );
 a131237a <=( a131236a  and  a131229a );
 a131240a <=( (not A266)  and  (not A265) );
 a131243a <=( (not A269)  and  A268 );
 a131244a <=( a131243a  and  a131240a );
 a131247a <=( A299  and  (not A298) );
 a131250a <=( (not A302)  and  (not A300) );
 a131251a <=( a131250a  and  a131247a );
 a131252a <=( a131251a  and  a131244a );


end x25_19x_behav;
