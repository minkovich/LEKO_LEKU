Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_14x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A73: buffer std_logic
);
end x25_14x;

architecture x25_14x_behav of x25_14x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1014a,a1015a,a1018a,a1021a,a1022a,a1023a,a1026a,a1029a,a1030a,a1033a,a1036a,a1037a,a1038a,a1039a,a1042a,a1045a,a1046a,a1049a,a1052a,a1053a,a1054a,a1057a,a1060a,a1061a,a1064a,a1067a,a1068a,a1069a,a1070a,a1071a,a1074a,a1077a,a1078a,a1081a,a1084a,a1085a,a1086a,a1089a,a1092a,a1093a,a1096a,a1099a,a1100a,a1101a,a1102a,a1105a,a1108a,a1109a,a1112a,a1115a,a1116a,a1117a,a1120a,a1123a,a1124a,a1127a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1139a,a1140a,a1143a,a1146a,a1147a,a1148a,a1151a,a1154a,a1155a,a1158a,a1161a,a1162a,a1163a,a1164a,a1167a,a1170a,a1171a,a1174a,a1177a,a1178a,a1179a,a1182a,a1185a,a1186a,a1189a,a1192a,a1193a,a1194a,a1195a,a1196a,a1199a,a1202a,a1203a,a1206a,a1209a,a1210a,a1211a,a1214a,a1217a,a1218a,a1221a,a1224a,a1225a,a1226a,a1227a,a1230a,a1233a,a1234a,a1237a,a1240a,a1241a,a1242a,a1245a,a1248a,a1249a,a1252a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1265a,a1266a,a1269a,a1272a,a1273a,a1274a,a1277a,a1280a,a1281a,a1284a,a1287a,a1288a,a1289a,a1290a,a1293a,a1296a,a1297a,a1300a,a1303a,a1304a,a1305a,a1308a,a1311a,a1312a,a1315a,a1318a,a1319a,a1320a,a1321a,a1322a,a1325a,a1328a,a1329a,a1332a,a1335a,a1336a,a1337a,a1340a,a1343a,a1344a,a1347a,a1350a,a1351a,a1352a,a1353a,a1356a,a1359a,a1360a,a1363a,a1366a,a1367a,a1368a,a1371a,a1374a,a1375a,a1378a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1390a,a1391a,a1394a,a1397a,a1398a,a1399a,a1402a,a1405a,a1406a,a1409a,a1412a,a1413a,a1414a,a1415a,a1418a,a1421a,a1422a,a1425a,a1428a,a1429a,a1430a,a1433a,a1436a,a1437a,a1440a,a1443a,a1444a,a1445a,a1446a,a1447a,a1450a,a1453a,a1454a,a1457a,a1460a,a1461a,a1462a,a1465a,a1468a,a1469a,a1472a,a1475a,a1476a,a1477a,a1478a,a1481a,a1484a,a1485a,a1488a,a1491a,a1492a,a1493a,a1496a,a1499a,a1500a,a1503a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1517a,a1518a,a1521a,a1524a,a1525a,a1526a,a1529a,a1532a,a1533a,a1536a,a1539a,a1540a,a1541a,a1542a,a1545a,a1548a,a1549a,a1552a,a1555a,a1556a,a1557a,a1560a,a1563a,a1564a,a1567a,a1570a,a1571a,a1572a,a1573a,a1574a,a1577a,a1580a,a1581a,a1584a,a1587a,a1588a,a1589a,a1592a,a1595a,a1596a,a1599a,a1602a,a1603a,a1604a,a1605a,a1608a,a1611a,a1612a,a1615a,a1618a,a1619a,a1620a,a1623a,a1626a,a1627a,a1630a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1642a,a1643a,a1646a,a1649a,a1650a,a1651a,a1654a,a1657a,a1658a,a1661a,a1664a,a1665a,a1666a,a1667a,a1670a,a1673a,a1674a,a1677a,a1680a,a1681a,a1682a,a1685a,a1688a,a1689a,a1692a,a1695a,a1696a,a1697a,a1698a,a1699a,a1702a,a1705a,a1706a,a1709a,a1712a,a1713a,a1714a,a1717a,a1720a,a1721a,a1724a,a1727a,a1728a,a1729a,a1730a,a1733a,a1736a,a1737a,a1740a,a1743a,a1744a,a1745a,a1748a,a1751a,a1752a,a1755a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1768a,a1769a,a1772a,a1775a,a1776a,a1777a,a1780a,a1783a,a1784a,a1787a,a1790a,a1791a,a1792a,a1793a,a1796a,a1799a,a1800a,a1803a,a1806a,a1807a,a1808a,a1811a,a1814a,a1815a,a1818a,a1821a,a1822a,a1823a,a1824a,a1825a,a1828a,a1831a,a1832a,a1835a,a1838a,a1839a,a1840a,a1843a,a1846a,a1847a,a1850a,a1853a,a1854a,a1855a,a1856a,a1859a,a1862a,a1863a,a1866a,a1869a,a1870a,a1871a,a1874a,a1877a,a1878a,a1881a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1892a,a1895a,a1896a,a1899a,a1902a,a1903a,a1904a,a1907a,a1910a,a1911a,a1914a,a1917a,a1918a,a1919a,a1920a,a1923a,a1926a,a1927a,a1930a,a1933a,a1934a,a1935a,a1938a,a1941a,a1942a,a1945a,a1948a,a1949a,a1950a,a1951a,a1952a,a1955a,a1958a,a1959a,a1962a,a1965a,a1966a,a1967a,a1970a,a1973a,a1974a,a1977a,a1980a,a1981a,a1982a,a1983a,a1986a,a1989a,a1990a,a1993a,a1996a,a1997a,a1998a,a2001a,a2004a,a2005a,a2008a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2023a,a2024a,a2027a,a2030a,a2031a,a2032a,a2035a,a2038a,a2039a,a2042a,a2045a,a2046a,a2047a,a2048a,a2051a,a2054a,a2055a,a2058a,a2061a,a2062a,a2063a,a2066a,a2069a,a2070a,a2073a,a2076a,a2077a,a2078a,a2079a,a2080a,a2083a,a2086a,a2087a,a2090a,a2093a,a2094a,a2095a,a2098a,a2101a,a2102a,a2105a,a2108a,a2109a,a2110a,a2111a,a2114a,a2117a,a2118a,a2121a,a2124a,a2125a,a2126a,a2129a,a2132a,a2133a,a2136a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2148a,a2149a,a2152a,a2155a,a2156a,a2157a,a2160a,a2163a,a2164a,a2167a,a2170a,a2171a,a2172a,a2173a,a2176a,a2179a,a2180a,a2183a,a2186a,a2187a,a2188a,a2191a,a2194a,a2195a,a2198a,a2201a,a2202a,a2203a,a2204a,a2205a,a2208a,a2211a,a2212a,a2215a,a2218a,a2219a,a2220a,a2223a,a2226a,a2227a,a2230a,a2233a,a2234a,a2235a,a2236a,a2239a,a2242a,a2243a,a2246a,a2249a,a2250a,a2251a,a2254a,a2257a,a2258a,a2261a,a2264a,a2265a,a2266a,a2267a,a2268a,a2269a,a2270a,a2274a,a2275a,a2278a,a2281a,a2282a,a2283a,a2286a,a2289a,a2290a,a2293a,a2296a,a2297a,a2298a,a2299a,a2302a,a2305a,a2306a,a2309a,a2312a,a2313a,a2314a,a2317a,a2320a,a2321a,a2324a,a2327a,a2328a,a2329a,a2330a,a2331a,a2334a,a2337a,a2338a,a2341a,a2344a,a2345a,a2346a,a2349a,a2352a,a2353a,a2356a,a2359a,a2360a,a2361a,a2362a,a2365a,a2368a,a2369a,a2372a,a2375a,a2376a,a2377a,a2380a,a2383a,a2384a,a2387a,a2390a,a2391a,a2392a,a2393a,a2394a,a2395a,a2399a,a2400a,a2403a,a2406a,a2407a,a2408a,a2411a,a2414a,a2415a,a2418a,a2421a,a2422a,a2423a,a2424a,a2427a,a2430a,a2431a,a2434a,a2437a,a2438a,a2439a,a2442a,a2445a,a2446a,a2449a,a2452a,a2453a,a2454a,a2455a,a2456a,a2459a,a2462a,a2463a,a2466a,a2469a,a2470a,a2471a,a2474a,a2477a,a2478a,a2481a,a2484a,a2485a,a2486a,a2487a,a2490a,a2493a,a2494a,a2497a,a2500a,a2501a,a2502a,a2505a,a2508a,a2509a,a2512a,a2515a,a2516a,a2517a,a2518a,a2519a,a2520a,a2521a,a2522a,a2526a,a2527a,a2530a,a2533a,a2534a,a2535a,a2538a,a2541a,a2542a,a2545a,a2548a,a2549a,a2550a,a2551a,a2554a,a2557a,a2558a,a2561a,a2564a,a2565a,a2566a,a2569a,a2572a,a2573a,a2576a,a2579a,a2580a,a2581a,a2582a,a2583a,a2586a,a2589a,a2590a,a2593a,a2596a,a2597a,a2598a,a2601a,a2604a,a2605a,a2608a,a2611a,a2612a,a2613a,a2614a,a2617a,a2620a,a2621a,a2624a,a2627a,a2628a,a2629a,a2632a,a2635a,a2636a,a2639a,a2642a,a2643a,a2644a,a2645a,a2646a,a2647a,a2651a,a2652a,a2655a,a2658a,a2659a,a2660a,a2663a,a2666a,a2667a,a2670a,a2673a,a2674a,a2675a,a2676a,a2679a,a2682a,a2683a,a2686a,a2689a,a2690a,a2691a,a2694a,a2697a,a2698a,a2701a,a2704a,a2705a,a2706a,a2707a,a2708a,a2711a,a2714a,a2715a,a2718a,a2721a,a2722a,a2723a,a2726a,a2729a,a2730a,a2733a,a2736a,a2737a,a2738a,a2739a,a2742a,a2745a,a2746a,a2749a,a2752a,a2753a,a2754a,a2757a,a2760a,a2761a,a2764a,a2767a,a2768a,a2769a,a2770a,a2771a,a2772a,a2773a,a2777a,a2778a,a2781a,a2784a,a2785a,a2786a,a2789a,a2792a,a2793a,a2796a,a2799a,a2800a,a2801a,a2802a,a2805a,a2808a,a2809a,a2812a,a2815a,a2816a,a2817a,a2820a,a2823a,a2824a,a2827a,a2830a,a2831a,a2832a,a2833a,a2834a,a2837a,a2840a,a2841a,a2844a,a2847a,a2848a,a2849a,a2852a,a2855a,a2856a,a2859a,a2862a,a2863a,a2864a,a2865a,a2868a,a2871a,a2872a,a2875a,a2878a,a2879a,a2880a,a2883a,a2886a,a2887a,a2890a,a2893a,a2894a,a2895a,a2896a,a2897a,a2898a,a2901a,a2904a,a2905a,a2908a,a2911a,a2912a,a2913a,a2916a,a2919a,a2920a,a2923a,a2926a,a2927a,a2928a,a2929a,a2932a,a2935a,a2936a,a2939a,a2942a,a2943a,a2944a,a2947a,a2950a,a2951a,a2954a,a2957a,a2958a,a2959a,a2960a,a2961a,a2964a,a2967a,a2968a,a2971a,a2974a,a2975a,a2976a,a2979a,a2982a,a2983a,a2986a,a2989a,a2990a,a2991a,a2992a,a2995a,a2998a,a2999a,a3002a,a3005a,a3006a,a3007a,a3010a,a3013a,a3014a,a3017a,a3020a,a3021a,a3022a,a3023a,a3024a,a3025a,a3026a,a3027a,a3028a,a3036a,a3040a,a3044a,a3048a,a3052a,a3056a,a3060a,a3064a,a3067a,a3070a,a3073a,a3076a,a3079a,a3082a,a3085a,a3088a,a3091a,a3094a,a3097a,a3100a,a3103a,a3106a,a3109a,a3112a,a3115a,a3118a,a3121a,a3124a,a3127a,a3130a,a3133a,a3136a,a3139a,a3142a,a3145a,a3148a,a3151a,a3154a,a3157a,a3160a,a3163a,a3167a,a3168a,a3171a,a3175a,a3176a,a3179a,a3183a,a3184a,a3187a,a3191a,a3192a,a3195a,a3199a,a3200a,a3203a,a3207a,a3208a,a3211a,a3215a,a3216a,a3219a,a3223a,a3224a,a3227a,a3231a,a3232a,a3235a,a3239a,a3240a,a3243a,a3247a,a3248a,a3251a,a3255a,a3256a,a3259a,a3263a,a3264a,a3267a,a3271a,a3272a,a3275a,a3279a,a3280a,a3283a,a3287a,a3288a,a3292a,a3293a,a3297a,a3298a,a3302a,a3303a,a3307a,a3308a,a3312a,a3313a,a3317a,a3318a,a3322a,a3323a,a3327a,a3328a,a3332a,a3333a,a3337a,a3338a,a3342a,a3343a,a3347a,a3348a,a3352a,a3353a,a3357a,a3358a,a3362a,a3363a,a3367a,a3368a,a3372a,a3373a,a3377a,a3378a,a3382a,a3383a,a3387a,a3388a,a3392a,a3393a,a3396a,a3399a,a3400a,a3404a,a3405a,a3408a,a3411a,a3412a,a3416a,a3417a,a3420a,a3423a,a3424a,a3428a,a3429a,a3432a,a3435a,a3436a,a3440a,a3441a,a3444a,a3447a,a3448a,a3452a,a3453a,a3456a,a3459a,a3460a,a3464a,a3465a,a3468a,a3471a,a3472a,a3476a,a3477a,a3480a,a3483a,a3484a,a3488a,a3489a,a3492a,a3495a,a3496a,a3500a,a3501a,a3504a,a3507a,a3508a,a3512a,a3513a,a3516a,a3519a,a3520a,a3524a,a3525a,a3528a,a3531a,a3532a,a3536a,a3537a,a3540a,a3543a,a3544a,a3547a,a3550a,a3551a,a3554a,a3557a,a3558a,a3561a,a3564a,a3565a,a3568a,a3571a,a3572a,a3575a,a3578a,a3579a,a3582a,a3585a,a3586a,a3589a,a3592a,a3593a,a3596a,a3599a,a3600a,a3603a,a3606a,a3607a,a3610a,a3613a,a3614a,a3617a,a3620a,a3621a,a3624a,a3627a,a3628a,a3631a,a3634a,a3635a,a3638a,a3641a,a3642a,a3645a,a3648a,a3649a,a3652a,a3655a,a3656a,a3659a,a3662a,a3663a,a3666a,a3669a,a3670a,a3673a,a3676a,a3677a,a3680a,a3683a,a3684a,a3687a,a3690a,a3691a,a3694a,a3697a,a3698a,a3701a,a3704a,a3705a,a3708a,a3711a,a3712a,a3715a,a3718a,a3719a,a3722a,a3725a,a3726a,a3729a,a3732a,a3733a,a3736a,a3739a,a3740a,a3743a,a3746a,a3747a,a3750a,a3753a,a3754a,a3757a,a3760a,a3761a,a3764a,a3767a,a3768a,a3771a,a3774a,a3775a,a3778a,a3781a,a3782a,a3785a,a3788a,a3789a,a3792a,a3795a,a3796a,a3799a,a3802a,a3803a,a3806a,a3809a,a3810a,a3813a,a3816a,a3817a,a3820a,a3823a,a3824a,a3827a,a3830a,a3831a,a3834a,a3837a,a3838a,a3841a,a3844a,a3845a,a3848a,a3851a,a3852a,a3855a,a3858a,a3859a,a3862a,a3865a,a3866a,a3869a,a3872a,a3873a,a3876a,a3879a,a3880a,a3883a,a3886a,a3887a,a3890a,a3893a,a3894a,a3897a,a3900a,a3901a,a3904a,a3907a,a3908a,a3911a,a3914a,a3915a,a3918a,a3921a,a3922a,a3925a,a3928a,a3929a,a3932a,a3935a,a3936a,a3939a,a3942a,a3943a,a3946a,a3949a,a3950a,a3953a,a3956a,a3957a,a3960a,a3963a,a3964a,a3967a,a3970a,a3971a,a3974a,a3977a,a3978a,a3981a,a3984a,a3985a,a3988a,a3991a,a3992a,a3995a,a3998a,a3999a,a4002a,a4005a,a4006a,a4009a,a4012a,a4013a,a4016a,a4019a,a4020a,a4023a,a4026a,a4027a,a4030a,a4033a,a4034a,a4037a,a4040a,a4041a,a4044a,a4047a,a4048a,a4051a,a4054a,a4055a,a4058a,a4061a,a4062a,a4065a,a4068a,a4069a,a4072a,a4075a,a4076a,a4079a,a4082a,a4083a,a4086a,a4089a,a4090a,a4093a,a4096a,a4097a,a4100a,a4103a,a4104a,a4107a,a4110a,a4111a,a4114a,a4117a,a4118a,a4121a,a4124a,a4125a,a4128a,a4131a,a4132a,a4135a,a4138a,a4139a,a4142a,a4145a,a4146a,a4149a,a4152a,a4153a,a4156a,a4159a,a4160a,a4163a,a4166a,a4167a,a4170a,a4173a,a4174a,a4177a,a4180a,a4181a,a4184a,a4187a,a4188a,a4191a,a4194a,a4195a,a4198a,a4201a,a4202a,a4205a,a4208a,a4209a,a4212a,a4215a,a4216a,a4219a,a4222a,a4223a,a4226a,a4229a,a4230a,a4233a,a4236a,a4237a,a4240a,a4243a,a4244a,a4247a,a4250a,a4251a,a4254a,a4258a,a4259a,a4260a,a4263a,a4266a,a4267a,a4270a,a4274a,a4275a,a4276a,a4279a,a4282a,a4283a,a4286a,a4290a,a4291a,a4292a,a4295a,a4298a,a4299a,a4302a,a4306a,a4307a,a4308a,a4311a,a4314a,a4315a,a4318a,a4322a,a4323a,a4324a,a4327a,a4330a,a4331a,a4334a,a4338a,a4339a,a4340a,a4343a,a4346a,a4347a,a4350a,a4354a,a4355a,a4356a,a4359a,a4362a,a4363a,a4366a,a4370a,a4371a,a4372a,a4375a,a4378a,a4379a,a4382a,a4386a,a4387a,a4388a,a4391a,a4394a,a4395a,a4398a,a4402a,a4403a,a4404a,a4407a,a4410a,a4411a,a4414a,a4418a,a4419a,a4420a,a4423a,a4426a,a4427a,a4430a,a4434a,a4435a,a4436a,a4439a,a4442a,a4443a,a4446a,a4450a,a4451a,a4452a,a4455a,a4458a,a4459a,a4462a,a4466a,a4467a,a4468a,a4471a,a4474a,a4475a,a4478a,a4482a,a4483a,a4484a,a4487a,a4490a,a4491a,a4494a,a4498a,a4499a,a4500a,a4503a,a4506a,a4507a,a4510a,a4514a,a4515a,a4516a,a4519a,a4522a,a4523a,a4526a,a4530a,a4531a,a4532a,a4535a,a4538a,a4539a,a4542a,a4546a,a4547a,a4548a,a4551a,a4554a,a4555a,a4558a,a4562a,a4563a,a4564a,a4567a,a4570a,a4571a,a4574a,a4578a,a4579a,a4580a,a4583a,a4586a,a4587a,a4590a,a4594a,a4595a,a4596a,a4599a,a4602a,a4603a,a4606a,a4610a,a4611a,a4612a,a4615a,a4618a,a4619a,a4622a,a4626a,a4627a,a4628a,a4631a,a4634a,a4635a,a4638a,a4642a,a4643a,a4644a,a4647a,a4650a,a4651a,a4654a,a4658a,a4659a,a4660a,a4663a,a4666a,a4667a,a4670a,a4674a,a4675a,a4676a,a4679a,a4682a,a4683a,a4686a,a4690a,a4691a,a4692a,a4695a,a4698a,a4699a,a4702a,a4706a,a4707a,a4708a,a4711a,a4714a,a4715a,a4718a,a4722a,a4723a,a4724a,a4727a,a4730a,a4731a,a4734a,a4738a,a4739a,a4740a,a4743a,a4746a,a4747a,a4750a,a4754a,a4755a,a4756a,a4759a,a4762a,a4763a,a4766a,a4770a,a4771a,a4772a,a4775a,a4778a,a4779a,a4782a,a4786a,a4787a,a4788a,a4791a,a4794a,a4795a,a4798a,a4802a,a4803a,a4804a,a4807a,a4810a,a4811a,a4814a,a4818a,a4819a,a4820a,a4823a,a4826a,a4827a,a4830a,a4834a,a4835a,a4836a,a4839a,a4842a,a4843a,a4846a,a4850a,a4851a,a4852a,a4855a,a4858a,a4859a,a4862a,a4866a,a4867a,a4868a,a4871a,a4874a,a4875a,a4878a,a4882a,a4883a,a4884a,a4887a,a4890a,a4891a,a4894a,a4898a,a4899a,a4900a,a4903a,a4906a,a4907a,a4910a,a4914a,a4915a,a4916a,a4919a,a4922a,a4923a,a4926a,a4930a,a4931a,a4932a,a4935a,a4938a,a4939a,a4942a,a4946a,a4947a,a4948a,a4951a,a4954a,a4955a,a4958a,a4962a,a4963a,a4964a,a4967a,a4970a,a4971a,a4974a,a4978a,a4979a,a4980a,a4983a,a4986a,a4987a,a4990a,a4994a,a4995a,a4996a,a4999a,a5002a,a5003a,a5006a,a5010a,a5011a,a5012a,a5015a,a5018a,a5019a,a5022a,a5026a,a5027a,a5028a,a5031a,a5034a,a5035a,a5038a,a5042a,a5043a,a5044a,a5047a,a5050a,a5051a,a5054a,a5058a,a5059a,a5060a,a5063a,a5066a,a5067a,a5070a,a5074a,a5075a,a5076a,a5079a,a5082a,a5083a,a5086a,a5090a,a5091a,a5092a,a5095a,a5098a,a5099a,a5102a,a5106a,a5107a,a5108a,a5111a,a5114a,a5115a,a5118a,a5122a,a5123a,a5124a,a5127a,a5130a,a5131a,a5134a,a5138a,a5139a,a5140a,a5143a,a5146a,a5147a,a5150a,a5154a,a5155a,a5156a,a5159a,a5162a,a5163a,a5166a,a5170a,a5171a,a5172a,a5175a,a5178a,a5179a,a5182a,a5186a,a5187a,a5188a,a5191a,a5194a,a5195a,a5198a,a5202a,a5203a,a5204a,a5207a,a5210a,a5211a,a5214a,a5218a,a5219a,a5220a,a5223a,a5226a,a5227a,a5230a,a5234a,a5235a,a5236a,a5239a,a5242a,a5243a,a5246a,a5250a,a5251a,a5252a,a5255a,a5258a,a5259a,a5262a,a5266a,a5267a,a5268a,a5271a,a5274a,a5275a,a5278a,a5282a,a5283a,a5284a,a5287a,a5290a,a5291a,a5294a,a5298a,a5299a,a5300a,a5303a,a5306a,a5307a,a5310a,a5314a,a5315a,a5316a,a5319a,a5322a,a5323a,a5326a,a5330a,a5331a,a5332a,a5335a,a5338a,a5339a,a5342a,a5346a,a5347a,a5348a,a5351a,a5354a,a5355a,a5358a,a5362a,a5363a,a5364a,a5367a,a5370a,a5371a,a5374a,a5378a,a5379a,a5380a,a5383a,a5386a,a5387a,a5390a,a5394a,a5395a,a5396a,a5399a,a5402a,a5403a,a5406a,a5410a,a5411a,a5412a,a5415a,a5418a,a5419a,a5422a,a5426a,a5427a,a5428a,a5431a,a5434a,a5435a,a5438a,a5442a,a5443a,a5444a,a5447a,a5450a,a5451a,a5454a,a5458a,a5459a,a5460a,a5463a,a5466a,a5467a,a5470a,a5474a,a5475a,a5476a,a5479a,a5482a,a5483a,a5486a,a5490a,a5491a,a5492a,a5495a,a5498a,a5499a,a5502a,a5506a,a5507a,a5508a,a5511a,a5514a,a5515a,a5518a,a5522a,a5523a,a5524a,a5527a,a5530a,a5531a,a5534a,a5538a,a5539a,a5540a,a5543a,a5546a,a5547a,a5550a,a5554a,a5555a,a5556a,a5559a,a5562a,a5563a,a5566a,a5570a,a5571a,a5572a,a5575a,a5578a,a5579a,a5582a,a5586a,a5587a,a5588a,a5591a,a5594a,a5595a,a5598a,a5602a,a5603a,a5604a,a5607a,a5610a,a5611a,a5614a,a5618a,a5619a,a5620a,a5623a,a5626a,a5627a,a5630a,a5634a,a5635a,a5636a,a5639a,a5642a,a5643a,a5646a,a5650a,a5651a,a5652a,a5655a,a5658a,a5659a,a5662a,a5666a,a5667a,a5668a,a5671a,a5674a,a5675a,a5678a,a5682a,a5683a,a5684a,a5687a,a5690a,a5691a,a5694a,a5698a,a5699a,a5700a,a5703a,a5706a,a5707a,a5710a,a5714a,a5715a,a5716a,a5719a,a5722a,a5723a,a5726a,a5730a,a5731a,a5732a,a5735a,a5738a,a5739a,a5742a,a5746a,a5747a,a5748a,a5751a,a5754a,a5755a,a5758a,a5762a,a5763a,a5764a,a5767a,a5770a,a5771a,a5774a,a5778a,a5779a,a5780a,a5783a,a5786a,a5787a,a5790a,a5794a,a5795a,a5796a,a5799a,a5802a,a5803a,a5806a,a5810a,a5811a,a5812a,a5815a,a5818a,a5819a,a5822a,a5826a,a5827a,a5828a,a5831a,a5834a,a5835a,a5838a,a5842a,a5843a,a5844a,a5847a,a5850a,a5851a,a5854a,a5858a,a5859a,a5860a,a5863a,a5866a,a5867a,a5870a,a5874a,a5875a,a5876a,a5879a,a5882a,a5883a,a5886a,a5890a,a5891a,a5892a,a5895a,a5898a,a5899a,a5902a,a5906a,a5907a,a5908a,a5911a,a5914a,a5915a,a5918a,a5922a,a5923a,a5924a,a5927a,a5930a,a5931a,a5934a,a5938a,a5939a,a5940a,a5943a,a5946a,a5947a,a5950a,a5954a,a5955a,a5956a,a5959a,a5962a,a5963a,a5966a,a5970a,a5971a,a5972a,a5975a,a5978a,a5979a,a5982a,a5986a,a5987a,a5988a,a5991a,a5994a,a5995a,a5998a,a6002a,a6003a,a6004a,a6007a,a6010a,a6011a,a6014a,a6018a,a6019a,a6020a,a6023a,a6026a,a6027a,a6030a,a6034a,a6035a,a6036a,a6039a,a6042a,a6043a,a6046a,a6050a,a6051a,a6052a,a6055a,a6058a,a6059a,a6062a,a6066a,a6067a,a6068a,a6071a,a6074a,a6075a,a6078a,a6082a,a6083a,a6084a,a6087a,a6090a,a6091a,a6094a,a6098a,a6099a,a6100a,a6103a,a6106a,a6107a,a6110a,a6114a,a6115a,a6116a,a6119a,a6122a,a6123a,a6126a,a6130a,a6131a,a6132a,a6135a,a6138a,a6139a,a6142a,a6146a,a6147a,a6148a,a6151a,a6154a,a6155a,a6158a,a6162a,a6163a,a6164a,a6167a,a6170a,a6171a,a6174a,a6178a,a6179a,a6180a,a6183a,a6186a,a6187a,a6190a,a6194a,a6195a,a6196a,a6199a,a6203a,a6204a,a6205a,a6208a,a6212a,a6213a,a6214a,a6217a,a6221a,a6222a,a6223a,a6226a,a6230a,a6231a,a6232a,a6235a,a6239a,a6240a,a6241a,a6244a,a6248a,a6249a,a6250a,a6253a,a6257a,a6258a,a6259a,a6262a,a6266a,a6267a,a6268a,a6271a,a6275a,a6276a,a6277a,a6280a,a6284a,a6285a,a6286a,a6289a,a6293a,a6294a,a6295a,a6298a,a6302a,a6303a,a6304a,a6307a,a6311a,a6312a,a6313a,a6316a,a6320a,a6321a,a6322a,a6325a,a6329a,a6330a,a6331a,a6334a,a6338a,a6339a,a6340a,a6343a,a6347a,a6348a,a6349a,a6352a,a6356a,a6357a,a6358a,a6361a,a6365a,a6366a,a6367a,a6370a,a6374a,a6375a,a6376a,a6379a,a6383a,a6384a,a6385a,a6388a,a6392a,a6393a,a6394a,a6397a,a6401a,a6402a,a6403a,a6406a,a6410a,a6411a,a6412a,a6415a,a6419a,a6420a,a6421a,a6424a,a6428a,a6429a,a6430a,a6433a,a6437a,a6438a,a6439a,a6442a,a6446a,a6447a,a6448a,a6451a,a6455a,a6456a,a6457a,a6460a,a6464a,a6465a,a6466a,a6469a,a6473a,a6474a,a6475a,a6478a,a6482a,a6483a,a6484a,a6487a,a6491a,a6492a,a6493a,a6496a,a6500a,a6501a,a6502a,a6505a,a6509a,a6510a,a6511a,a6514a,a6518a,a6519a,a6520a,a6523a,a6527a,a6528a,a6529a,a6532a,a6536a,a6537a,a6538a,a6541a,a6545a,a6546a,a6547a,a6550a,a6554a,a6555a,a6556a,a6559a,a6563a,a6564a,a6565a,a6568a,a6572a,a6573a,a6574a,a6577a,a6581a,a6582a,a6583a,a6586a,a6590a,a6591a,a6592a,a6595a,a6599a,a6600a,a6601a,a6604a,a6608a,a6609a,a6610a,a6613a,a6617a,a6618a,a6619a,a6622a,a6626a,a6627a,a6628a,a6631a,a6635a,a6636a,a6637a,a6640a,a6644a,a6645a,a6646a,a6649a,a6653a,a6654a,a6655a,a6658a,a6662a,a6663a,a6664a,a6667a,a6671a,a6672a,a6673a,a6676a,a6680a,a6681a,a6682a,a6685a,a6689a,a6690a,a6691a,a6694a,a6698a,a6699a,a6700a,a6703a,a6707a,a6708a,a6709a,a6712a,a6716a,a6717a,a6718a,a6721a,a6725a,a6726a,a6727a,a6730a,a6734a,a6735a,a6736a,a6739a,a6743a,a6744a,a6745a,a6748a,a6752a,a6753a,a6754a,a6757a,a6761a,a6762a,a6763a,a6766a,a6770a,a6771a,a6772a,a6775a,a6779a,a6780a,a6781a,a6784a,a6788a,a6789a,a6790a,a6793a,a6797a,a6798a,a6799a,a6802a,a6806a,a6807a,a6808a,a6811a,a6815a,a6816a,a6817a,a6820a,a6824a,a6825a,a6826a,a6829a,a6833a,a6834a,a6835a,a6838a,a6842a,a6843a,a6844a,a6847a,a6851a,a6852a,a6853a,a6856a,a6860a,a6861a,a6862a,a6865a,a6869a,a6870a,a6871a,a6874a,a6878a,a6879a,a6880a,a6883a,a6887a,a6888a,a6889a,a6892a,a6896a,a6897a,a6898a,a6901a,a6905a,a6906a,a6907a,a6910a,a6914a,a6915a,a6916a,a6919a,a6923a,a6924a,a6925a,a6928a,a6932a,a6933a,a6934a,a6937a,a6941a,a6942a,a6943a,a6946a,a6950a,a6951a,a6952a,a6955a,a6959a,a6960a,a6961a,a6964a,a6968a,a6969a,a6970a,a6973a,a6977a,a6978a,a6979a,a6982a,a6986a,a6987a,a6988a,a6991a,a6995a,a6996a,a6997a,a7000a,a7004a,a7005a,a7006a,a7009a,a7013a,a7014a,a7015a,a7018a,a7022a,a7023a,a7024a,a7027a,a7031a,a7032a,a7033a,a7036a,a7040a,a7041a,a7042a,a7045a,a7049a,a7050a,a7051a,a7054a,a7058a,a7059a,a7060a,a7063a,a7067a,a7068a,a7069a,a7072a,a7076a,a7077a,a7078a,a7081a,a7085a,a7086a,a7087a,a7090a,a7094a,a7095a,a7096a,a7099a,a7103a,a7104a,a7105a,a7108a,a7112a,a7113a,a7114a,a7117a,a7121a,a7122a,a7123a,a7126a,a7130a,a7131a,a7132a,a7135a,a7139a,a7140a,a7141a,a7144a,a7148a,a7149a,a7150a,a7153a,a7157a,a7158a,a7159a,a7162a,a7166a,a7167a,a7168a,a7171a,a7175a,a7176a,a7177a,a7180a,a7184a,a7185a,a7186a,a7189a,a7193a,a7194a,a7195a,a7198a,a7202a,a7203a,a7204a,a7207a,a7211a,a7212a,a7213a,a7216a,a7220a,a7221a,a7222a,a7225a,a7229a,a7230a,a7231a,a7234a,a7238a,a7239a,a7240a,a7243a,a7247a,a7248a,a7249a,a7252a,a7256a,a7257a,a7258a,a7261a,a7265a,a7266a,a7267a,a7270a,a7274a,a7275a,a7276a,a7279a,a7283a,a7284a,a7285a,a7288a,a7292a,a7293a,a7294a,a7297a,a7301a,a7302a,a7303a,a7306a,a7310a,a7311a,a7312a,a7315a,a7319a,a7320a,a7321a,a7324a,a7328a,a7329a,a7330a,a7333a,a7337a,a7338a,a7339a,a7342a,a7346a,a7347a,a7348a,a7351a,a7355a,a7356a,a7357a,a7360a,a7364a,a7365a,a7366a,a7369a,a7373a,a7374a,a7375a,a7378a,a7382a,a7383a,a7384a,a7387a,a7391a,a7392a,a7393a,a7396a,a7400a,a7401a,a7402a,a7405a,a7409a,a7410a,a7411a,a7414a,a7418a,a7419a,a7420a,a7423a,a7427a,a7428a,a7429a,a7432a,a7436a,a7437a,a7438a,a7441a,a7445a,a7446a,a7447a,a7450a,a7454a,a7455a,a7456a,a7459a,a7463a,a7464a,a7465a,a7468a,a7472a,a7473a,a7474a,a7477a,a7481a,a7482a,a7483a,a7486a,a7490a,a7491a,a7492a,a7495a,a7499a,a7500a,a7501a,a7504a,a7508a,a7509a,a7510a,a7513a,a7517a,a7518a,a7519a,a7522a,a7526a,a7527a,a7528a,a7531a,a7535a,a7536a,a7537a,a7540a,a7544a,a7545a,a7546a,a7549a,a7553a,a7554a,a7555a,a7558a,a7562a,a7563a,a7564a,a7567a,a7571a,a7572a,a7573a,a7576a,a7580a,a7581a,a7582a,a7585a,a7589a,a7590a,a7591a,a7594a,a7598a,a7599a,a7600a,a7603a,a7607a,a7608a,a7609a,a7612a,a7616a,a7617a,a7618a,a7621a,a7625a,a7626a,a7627a,a7630a,a7634a,a7635a,a7636a,a7639a,a7643a,a7644a,a7645a,a7648a,a7652a,a7653a,a7654a,a7657a,a7661a,a7662a,a7663a,a7666a,a7670a,a7671a,a7672a,a7675a,a7679a,a7680a,a7681a,a7684a,a7688a,a7689a,a7690a,a7693a,a7697a,a7698a,a7699a,a7702a,a7706a,a7707a,a7708a,a7711a,a7715a,a7716a,a7717a,a7720a,a7724a,a7725a,a7726a,a7729a,a7733a,a7734a,a7735a,a7738a,a7742a,a7743a,a7744a,a7747a,a7751a,a7752a,a7753a,a7756a,a7760a,a7761a,a7762a,a7765a,a7769a,a7770a,a7771a,a7774a,a7778a,a7779a,a7780a,a7783a,a7787a,a7788a,a7789a,a7792a,a7796a,a7797a,a7798a,a7801a,a7805a,a7806a,a7807a,a7810a,a7814a,a7815a,a7816a,a7819a,a7823a,a7824a,a7825a,a7828a,a7832a,a7833a,a7834a,a7837a,a7841a,a7842a,a7843a,a7846a,a7850a,a7851a,a7852a,a7855a,a7859a,a7860a,a7861a,a7864a,a7868a,a7869a,a7870a,a7873a,a7877a,a7878a,a7879a,a7882a,a7886a,a7887a,a7888a,a7891a,a7895a,a7896a,a7897a,a7900a,a7904a,a7905a,a7906a,a7909a,a7913a,a7914a,a7915a,a7918a,a7922a,a7923a,a7924a,a7927a,a7931a,a7932a,a7933a,a7936a,a7940a,a7941a,a7942a,a7945a,a7949a,a7950a,a7951a,a7954a,a7958a,a7959a,a7960a,a7963a,a7967a,a7968a,a7969a,a7972a,a7976a,a7977a,a7978a,a7981a,a7985a,a7986a,a7987a,a7990a,a7994a,a7995a,a7996a,a7999a,a8003a,a8004a,a8005a,a8008a,a8012a,a8013a,a8014a,a8017a,a8021a,a8022a,a8023a,a8026a,a8030a,a8031a,a8032a,a8035a,a8039a,a8040a,a8041a,a8044a,a8048a,a8049a,a8050a,a8053a,a8057a,a8058a,a8059a,a8062a,a8066a,a8067a,a8068a,a8071a,a8075a,a8076a,a8077a,a8080a,a8084a,a8085a,a8086a,a8089a,a8093a,a8094a,a8095a,a8098a,a8102a,a8103a,a8104a,a8107a,a8111a,a8112a,a8113a,a8116a,a8120a,a8121a,a8122a,a8125a,a8129a,a8130a,a8131a,a8134a,a8138a,a8139a,a8140a,a8143a,a8147a,a8148a,a8149a,a8152a,a8156a,a8157a,a8158a,a8161a,a8165a,a8166a,a8167a,a8170a,a8174a,a8175a,a8176a,a8179a,a8183a,a8184a,a8185a,a8188a,a8192a,a8193a,a8194a,a8197a,a8201a,a8202a,a8203a,a8206a,a8210a,a8211a,a8212a,a8215a,a8219a,a8220a,a8221a,a8224a,a8228a,a8229a,a8230a,a8233a,a8237a,a8238a,a8239a,a8242a,a8246a,a8247a,a8248a,a8251a,a8255a,a8256a,a8257a,a8260a,a8264a,a8265a,a8266a,a8269a,a8273a,a8274a,a8275a,a8278a,a8282a,a8283a,a8284a,a8287a,a8291a,a8292a,a8293a,a8296a,a8300a,a8301a,a8302a,a8305a,a8309a,a8310a,a8311a,a8314a,a8318a,a8319a,a8320a,a8323a,a8327a,a8328a,a8329a,a8332a,a8336a,a8337a,a8338a,a8341a,a8345a,a8346a,a8347a,a8350a,a8354a,a8355a,a8356a,a8359a,a8363a,a8364a,a8365a,a8368a,a8372a,a8373a,a8374a,a8377a,a8381a,a8382a,a8383a,a8386a,a8390a,a8391a,a8392a,a8395a,a8399a,a8400a,a8401a,a8404a,a8408a,a8409a,a8410a,a8413a,a8417a,a8418a,a8419a,a8422a,a8426a,a8427a,a8428a,a8431a,a8435a,a8436a,a8437a,a8440a,a8444a,a8445a,a8446a,a8449a,a8453a,a8454a,a8455a,a8458a,a8462a,a8463a,a8464a,a8467a,a8471a,a8472a,a8473a,a8476a,a8480a,a8481a,a8482a,a8485a,a8489a,a8490a,a8491a,a8494a,a8498a,a8499a,a8500a,a8503a,a8507a,a8508a,a8509a,a8512a,a8516a,a8517a,a8518a,a8521a,a8525a,a8526a,a8527a,a8530a,a8534a,a8535a,a8536a,a8539a,a8543a,a8544a,a8545a,a8548a,a8552a,a8553a,a8554a,a8557a,a8561a,a8562a,a8563a,a8566a,a8570a,a8571a,a8572a,a8575a,a8579a,a8580a,a8581a,a8584a,a8588a,a8589a,a8590a,a8593a,a8597a,a8598a,a8599a,a8602a,a8606a,a8607a,a8608a,a8611a,a8615a,a8616a,a8617a,a8620a,a8624a,a8625a,a8626a,a8629a,a8633a,a8634a,a8635a,a8638a,a8642a,a8643a,a8644a,a8647a,a8651a,a8652a,a8653a,a8656a,a8660a,a8661a,a8662a,a8665a,a8669a,a8670a,a8671a,a8674a,a8678a,a8679a,a8680a,a8683a,a8687a,a8688a,a8689a,a8692a,a8696a,a8697a,a8698a,a8701a,a8705a,a8706a,a8707a,a8710a,a8714a,a8715a,a8716a,a8719a,a8723a,a8724a,a8725a,a8728a,a8732a,a8733a,a8734a,a8737a,a8741a,a8742a,a8743a,a8746a,a8750a,a8751a,a8752a,a8755a,a8759a,a8760a,a8761a,a8764a,a8768a,a8769a,a8770a,a8773a,a8777a,a8778a,a8779a,a8782a,a8786a,a8787a,a8788a,a8791a,a8795a,a8796a,a8797a,a8800a,a8804a,a8805a,a8806a,a8809a,a8813a,a8814a,a8815a,a8818a,a8822a,a8823a,a8824a,a8827a,a8831a,a8832a,a8833a,a8836a,a8840a,a8841a,a8842a,a8845a,a8849a,a8850a,a8851a,a8854a,a8858a,a8859a,a8860a,a8863a,a8867a,a8868a,a8869a,a8872a,a8876a,a8877a,a8878a,a8881a,a8885a,a8886a,a8887a,a8890a,a8894a,a8895a,a8896a,a8899a,a8903a,a8904a,a8905a,a8908a,a8912a,a8913a,a8914a,a8917a,a8921a,a8922a,a8923a,a8926a,a8930a,a8931a,a8932a,a8935a,a8939a,a8940a,a8941a,a8944a,a8948a,a8949a,a8950a,a8953a,a8957a,a8958a,a8959a,a8962a,a8966a,a8967a,a8968a,a8971a,a8975a,a8976a,a8977a,a8980a,a8984a,a8985a,a8986a,a8989a,a8993a,a8994a,a8995a,a8998a,a9002a,a9003a,a9004a,a9007a,a9011a,a9012a,a9013a,a9016a,a9020a,a9021a,a9022a,a9025a,a9029a,a9030a,a9031a,a9034a,a9038a,a9039a,a9040a,a9043a,a9047a,a9048a,a9049a,a9052a,a9056a,a9057a,a9058a,a9061a,a9065a,a9066a,a9067a,a9070a,a9074a,a9075a,a9076a,a9079a,a9083a,a9084a,a9085a,a9088a,a9092a,a9093a,a9094a,a9097a,a9101a,a9102a,a9103a,a9106a,a9110a,a9111a,a9112a,a9115a,a9119a,a9120a,a9121a,a9124a,a9128a,a9129a,a9130a,a9133a,a9137a,a9138a,a9139a,a9142a,a9146a,a9147a,a9148a,a9151a,a9155a,a9156a,a9157a,a9160a,a9164a,a9165a,a9166a,a9169a,a9173a,a9174a,a9175a,a9178a,a9182a,a9183a,a9184a,a9187a,a9191a,a9192a,a9193a,a9196a,a9200a,a9201a,a9202a,a9205a,a9209a,a9210a,a9211a,a9214a,a9218a,a9219a,a9220a,a9223a,a9227a,a9228a,a9229a,a9232a,a9236a,a9237a,a9238a,a9241a,a9245a,a9246a,a9247a,a9250a,a9254a,a9255a,a9256a,a9259a,a9263a,a9264a,a9265a,a9268a,a9272a,a9273a,a9274a,a9277a,a9281a,a9282a,a9283a,a9286a,a9290a,a9291a,a9292a,a9295a,a9299a,a9300a,a9301a,a9304a,a9308a,a9309a,a9310a,a9313a,a9317a,a9318a,a9319a,a9322a,a9326a,a9327a,a9328a,a9331a,a9335a,a9336a,a9337a,a9340a,a9344a,a9345a,a9346a,a9349a,a9353a,a9354a,a9355a,a9358a,a9362a,a9363a,a9364a,a9367a,a9371a,a9372a,a9373a,a9376a,a9380a,a9381a,a9382a,a9385a,a9389a,a9390a,a9391a,a9394a,a9398a,a9399a,a9400a,a9403a,a9407a,a9408a,a9409a,a9412a,a9416a,a9417a,a9418a,a9421a,a9425a,a9426a,a9427a,a9430a,a9434a,a9435a,a9436a,a9439a,a9443a,a9444a,a9445a,a9448a,a9452a,a9453a,a9454a,a9457a,a9461a,a9462a,a9463a,a9466a,a9470a,a9471a,a9472a,a9475a,a9479a,a9480a,a9481a,a9484a,a9488a,a9489a,a9490a,a9493a,a9497a,a9498a,a9499a,a9502a,a9506a,a9507a,a9508a,a9511a,a9515a,a9516a,a9517a,a9520a,a9524a,a9525a,a9526a,a9529a,a9533a,a9534a,a9535a,a9538a,a9542a,a9543a,a9544a,a9547a,a9551a,a9552a,a9553a,a9556a,a9560a,a9561a,a9562a,a9565a,a9569a,a9570a,a9571a,a9574a,a9578a,a9579a,a9580a,a9583a,a9587a,a9588a,a9589a,a9592a,a9596a,a9597a,a9598a,a9601a,a9605a,a9606a,a9607a,a9610a,a9614a,a9615a,a9616a,a9619a,a9623a,a9624a,a9625a,a9628a,a9632a,a9633a,a9634a,a9637a,a9641a,a9642a,a9643a,a9646a,a9650a,a9651a,a9652a,a9655a,a9659a,a9660a,a9661a,a9664a,a9668a,a9669a,a9670a,a9673a,a9677a,a9678a,a9679a,a9682a,a9686a,a9687a,a9688a,a9691a,a9695a,a9696a,a9697a,a9700a,a9704a,a9705a,a9706a,a9709a,a9713a,a9714a,a9715a,a9718a,a9722a,a9723a,a9724a,a9727a,a9731a,a9732a,a9733a,a9736a,a9740a,a9741a,a9742a,a9745a,a9749a,a9750a,a9751a,a9754a,a9758a,a9759a,a9760a,a9763a,a9767a,a9768a,a9769a,a9772a,a9776a,a9777a,a9778a,a9781a,a9785a,a9786a,a9787a,a9790a,a9794a,a9795a,a9796a,a9799a,a9803a,a9804a,a9805a,a9808a,a9812a,a9813a,a9814a,a9817a,a9821a,a9822a,a9823a,a9826a,a9830a,a9831a,a9832a,a9835a,a9839a,a9840a,a9841a,a9844a,a9848a,a9849a,a9850a,a9853a,a9857a,a9858a,a9859a,a9862a,a9866a,a9867a,a9868a,a9871a,a9875a,a9876a,a9877a,a9880a,a9884a,a9885a,a9886a,a9889a,a9893a,a9894a,a9895a,a9898a,a9902a,a9903a,a9904a,a9907a,a9911a,a9912a,a9913a,a9916a,a9920a,a9921a,a9922a,a9925a,a9929a,a9930a,a9931a,a9934a,a9938a,a9939a,a9940a,a9943a,a9947a,a9948a,a9949a,a9952a,a9956a,a9957a,a9958a,a9961a,a9965a,a9966a,a9967a,a9970a,a9974a,a9975a,a9976a,a9979a,a9983a,a9984a,a9985a,a9989a,a9990a,a9994a,a9995a,a9996a,a9999a,a10003a,a10004a,a10005a,a10009a,a10010a,a10014a,a10015a,a10016a,a10019a,a10023a,a10024a,a10025a,a10029a,a10030a,a10034a,a10035a,a10036a,a10039a,a10043a,a10044a,a10045a,a10049a,a10050a,a10054a,a10055a,a10056a,a10059a,a10063a,a10064a,a10065a,a10069a,a10070a,a10074a,a10075a,a10076a,a10079a,a10083a,a10084a,a10085a,a10089a,a10090a,a10094a,a10095a,a10096a,a10099a,a10103a,a10104a,a10105a,a10109a,a10110a,a10114a,a10115a,a10116a,a10119a,a10123a,a10124a,a10125a,a10129a,a10130a,a10134a,a10135a,a10136a,a10139a,a10143a,a10144a,a10145a,a10149a,a10150a,a10154a,a10155a,a10156a,a10159a,a10163a,a10164a,a10165a,a10169a,a10170a,a10174a,a10175a,a10176a,a10179a,a10183a,a10184a,a10185a,a10189a,a10190a,a10194a,a10195a,a10196a,a10199a,a10203a,a10204a,a10205a,a10209a,a10210a,a10214a,a10215a,a10216a,a10219a,a10223a,a10224a,a10225a,a10229a,a10230a,a10234a,a10235a,a10236a,a10239a,a10243a,a10244a,a10245a,a10249a,a10250a,a10254a,a10255a,a10256a,a10259a,a10263a,a10264a,a10265a,a10269a,a10270a,a10274a,a10275a,a10276a,a10279a,a10283a,a10284a,a10285a,a10289a,a10290a,a10294a,a10295a,a10296a,a10299a,a10303a,a10304a,a10305a,a10309a,a10310a,a10314a,a10315a,a10316a,a10319a,a10323a,a10324a,a10325a,a10329a,a10330a,a10334a,a10335a,a10336a,a10339a,a10343a,a10344a,a10345a,a10349a,a10350a,a10354a,a10355a,a10356a,a10359a,a10363a,a10364a,a10365a,a10369a,a10370a,a10374a,a10375a,a10376a,a10379a,a10383a,a10384a,a10385a,a10389a,a10390a,a10394a,a10395a,a10396a,a10399a,a10403a,a10404a,a10405a,a10409a,a10410a,a10414a,a10415a,a10416a,a10419a,a10423a,a10424a,a10425a,a10429a,a10430a,a10434a,a10435a,a10436a,a10439a,a10443a,a10444a,a10445a,a10449a,a10450a,a10454a,a10455a,a10456a,a10459a,a10463a,a10464a,a10465a,a10469a,a10470a,a10474a,a10475a,a10476a,a10479a,a10483a,a10484a,a10485a,a10489a,a10490a,a10494a,a10495a,a10496a,a10499a,a10503a,a10504a,a10505a,a10509a,a10510a,a10514a,a10515a,a10516a,a10519a,a10523a,a10524a,a10525a,a10529a,a10530a,a10534a,a10535a,a10536a,a10539a,a10543a,a10544a,a10545a,a10549a,a10550a,a10554a,a10555a,a10556a,a10559a,a10563a,a10564a,a10565a,a10569a,a10570a,a10574a,a10575a,a10576a,a10579a,a10583a,a10584a,a10585a,a10589a,a10590a,a10594a,a10595a,a10596a,a10599a,a10603a,a10604a,a10605a,a10609a,a10610a,a10614a,a10615a,a10616a,a10619a,a10623a,a10624a,a10625a,a10629a,a10630a,a10634a,a10635a,a10636a,a10639a,a10643a,a10644a,a10645a,a10649a,a10650a,a10654a,a10655a,a10656a,a10659a,a10663a,a10664a,a10665a,a10669a,a10670a,a10674a,a10675a,a10676a,a10679a,a10683a,a10684a,a10685a,a10689a,a10690a,a10694a,a10695a,a10696a,a10699a,a10703a,a10704a,a10705a,a10709a,a10710a,a10714a,a10715a,a10716a,a10719a,a10723a,a10724a,a10725a,a10729a,a10730a,a10734a,a10735a,a10736a,a10739a,a10743a,a10744a,a10745a,a10749a,a10750a,a10754a,a10755a,a10756a,a10759a,a10763a,a10764a,a10765a,a10769a,a10770a,a10774a,a10775a,a10776a,a10779a,a10783a,a10784a,a10785a,a10789a,a10790a,a10794a,a10795a,a10796a,a10799a,a10803a,a10804a,a10805a,a10809a,a10810a,a10814a,a10815a,a10816a,a10819a,a10823a,a10824a,a10825a,a10829a,a10830a,a10834a,a10835a,a10836a,a10839a,a10843a,a10844a,a10845a,a10849a,a10850a,a10854a,a10855a,a10856a,a10859a,a10863a,a10864a,a10865a,a10869a,a10870a,a10874a,a10875a,a10876a,a10879a,a10883a,a10884a,a10885a,a10889a,a10890a,a10894a,a10895a,a10896a,a10899a,a10903a,a10904a,a10905a,a10909a,a10910a,a10914a,a10915a,a10916a,a10919a,a10923a,a10924a,a10925a,a10929a,a10930a,a10934a,a10935a,a10936a,a10939a,a10943a,a10944a,a10945a,a10949a,a10950a,a10954a,a10955a,a10956a,a10959a,a10963a,a10964a,a10965a,a10969a,a10970a,a10974a,a10975a,a10976a,a10979a,a10983a,a10984a,a10985a,a10989a,a10990a,a10994a,a10995a,a10996a,a10999a,a11003a,a11004a,a11005a,a11009a,a11010a,a11014a,a11015a,a11016a,a11019a,a11023a,a11024a,a11025a,a11029a,a11030a,a11034a,a11035a,a11036a,a11039a,a11043a,a11044a,a11045a,a11049a,a11050a,a11054a,a11055a,a11056a,a11059a,a11063a,a11064a,a11065a,a11069a,a11070a,a11074a,a11075a,a11076a,a11079a,a11083a,a11084a,a11085a,a11089a,a11090a,a11094a,a11095a,a11096a,a11099a,a11103a,a11104a,a11105a,a11109a,a11110a,a11114a,a11115a,a11116a,a11119a,a11123a,a11124a,a11125a,a11129a,a11130a,a11134a,a11135a,a11136a,a11139a,a11143a,a11144a,a11145a,a11149a,a11150a,a11154a,a11155a,a11156a,a11159a,a11163a,a11164a,a11165a,a11169a,a11170a,a11174a,a11175a,a11176a,a11179a,a11183a,a11184a,a11185a,a11189a,a11190a,a11194a,a11195a,a11196a,a11199a,a11203a,a11204a,a11205a,a11209a,a11210a,a11214a,a11215a,a11216a,a11219a,a11223a,a11224a,a11225a,a11229a,a11230a,a11234a,a11235a,a11236a,a11239a,a11243a,a11244a,a11245a,a11249a,a11250a,a11254a,a11255a,a11256a,a11259a,a11263a,a11264a,a11265a,a11269a,a11270a,a11274a,a11275a,a11276a,a11279a,a11283a,a11284a,a11285a,a11289a,a11290a,a11294a,a11295a,a11296a,a11299a,a11303a,a11304a,a11305a,a11309a,a11310a,a11314a,a11315a,a11316a,a11319a,a11323a,a11324a,a11325a,a11329a,a11330a,a11334a,a11335a,a11336a,a11339a,a11343a,a11344a,a11345a,a11349a,a11350a,a11354a,a11355a,a11356a,a11359a,a11363a,a11364a,a11365a,a11369a,a11370a,a11374a,a11375a,a11376a,a11379a,a11383a,a11384a,a11385a,a11389a,a11390a,a11394a,a11395a,a11396a,a11399a,a11403a,a11404a,a11405a,a11409a,a11410a,a11414a,a11415a,a11416a,a11419a,a11423a,a11424a,a11425a,a11429a,a11430a,a11434a,a11435a,a11436a,a11439a,a11443a,a11444a,a11445a,a11449a,a11450a,a11454a,a11455a,a11456a,a11459a,a11463a,a11464a,a11465a,a11469a,a11470a,a11474a,a11475a,a11476a,a11479a,a11483a,a11484a,a11485a,a11489a,a11490a,a11494a,a11495a,a11496a,a11499a,a11503a,a11504a,a11505a,a11509a,a11510a,a11514a,a11515a,a11516a,a11519a,a11523a,a11524a,a11525a,a11529a,a11530a,a11534a,a11535a,a11536a,a11539a,a11543a,a11544a,a11545a,a11549a,a11550a,a11554a,a11555a,a11556a,a11559a,a11563a,a11564a,a11565a,a11569a,a11570a,a11574a,a11575a,a11576a,a11579a,a11583a,a11584a,a11585a,a11589a,a11590a,a11594a,a11595a,a11596a,a11599a,a11603a,a11604a,a11605a,a11609a,a11610a,a11614a,a11615a,a11616a,a11619a,a11623a,a11624a,a11625a,a11629a,a11630a,a11634a,a11635a,a11636a,a11639a,a11643a,a11644a,a11645a,a11649a,a11650a,a11654a,a11655a,a11656a,a11659a,a11663a,a11664a,a11665a,a11669a,a11670a,a11674a,a11675a,a11676a,a11679a,a11683a,a11684a,a11685a,a11689a,a11690a,a11694a,a11695a,a11696a,a11699a,a11703a,a11704a,a11705a,a11709a,a11710a,a11714a,a11715a,a11716a,a11719a,a11723a,a11724a,a11725a,a11729a,a11730a,a11734a,a11735a,a11736a,a11739a,a11743a,a11744a,a11745a,a11749a,a11750a,a11754a,a11755a,a11756a,a11759a,a11763a,a11764a,a11765a,a11769a,a11770a,a11774a,a11775a,a11776a,a11779a,a11783a,a11784a,a11785a,a11789a,a11790a,a11794a,a11795a,a11796a,a11799a,a11803a,a11804a,a11805a,a11809a,a11810a,a11814a,a11815a,a11816a,a11819a,a11823a,a11824a,a11825a,a11829a,a11830a,a11834a,a11835a,a11836a,a11839a,a11843a,a11844a,a11845a,a11849a,a11850a,a11854a,a11855a,a11856a,a11859a,a11863a,a11864a,a11865a,a11869a,a11870a,a11874a,a11875a,a11876a,a11879a,a11883a,a11884a,a11885a,a11889a,a11890a,a11894a,a11895a,a11896a,a11899a,a11903a,a11904a,a11905a,a11909a,a11910a,a11914a,a11915a,a11916a,a11919a,a11923a,a11924a,a11925a,a11929a,a11930a,a11934a,a11935a,a11936a,a11939a,a11943a,a11944a,a11945a,a11949a,a11950a,a11954a,a11955a,a11956a,a11959a,a11963a,a11964a,a11965a,a11969a,a11970a,a11974a,a11975a,a11976a,a11979a,a11983a,a11984a,a11985a,a11989a,a11990a,a11994a,a11995a,a11996a,a11999a,a12003a,a12004a,a12005a,a12009a,a12010a,a12014a,a12015a,a12016a,a12019a,a12023a,a12024a,a12025a,a12029a,a12030a,a12034a,a12035a,a12036a,a12039a,a12043a,a12044a,a12045a,a12049a,a12050a,a12054a,a12055a,a12056a,a12059a,a12063a,a12064a,a12065a,a12069a,a12070a,a12074a,a12075a,a12076a,a12079a,a12083a,a12084a,a12085a,a12089a,a12090a,a12094a,a12095a,a12096a,a12099a,a12103a,a12104a,a12105a,a12109a,a12110a,a12114a,a12115a,a12116a,a12119a,a12123a,a12124a,a12125a,a12129a,a12130a,a12134a,a12135a,a12136a,a12139a,a12143a,a12144a,a12145a,a12149a,a12150a,a12154a,a12155a,a12156a,a12159a,a12163a,a12164a,a12165a,a12169a,a12170a,a12174a,a12175a,a12176a,a12179a,a12183a,a12184a,a12185a,a12189a,a12190a,a12194a,a12195a,a12196a,a12199a,a12203a,a12204a,a12205a,a12209a,a12210a,a12214a,a12215a,a12216a,a12219a,a12223a,a12224a,a12225a,a12229a,a12230a,a12234a,a12235a,a12236a,a12239a,a12243a,a12244a,a12245a,a12249a,a12250a,a12254a,a12255a,a12256a,a12259a,a12263a,a12264a,a12265a,a12269a,a12270a,a12274a,a12275a,a12276a,a12279a,a12283a,a12284a,a12285a,a12289a,a12290a,a12294a,a12295a,a12296a,a12299a,a12303a,a12304a,a12305a,a12309a,a12310a,a12314a,a12315a,a12316a,a12319a,a12323a,a12324a,a12325a,a12329a,a12330a,a12334a,a12335a,a12336a,a12339a,a12343a,a12344a,a12345a,a12349a,a12350a,a12354a,a12355a,a12356a,a12359a,a12363a,a12364a,a12365a,a12369a,a12370a,a12374a,a12375a,a12376a,a12379a,a12383a,a12384a,a12385a,a12389a,a12390a,a12394a,a12395a,a12396a,a12399a,a12403a,a12404a,a12405a,a12409a,a12410a,a12414a,a12415a,a12416a,a12419a,a12423a,a12424a,a12425a,a12429a,a12430a,a12434a,a12435a,a12436a,a12439a,a12443a,a12444a,a12445a,a12449a,a12450a,a12454a,a12455a,a12456a,a12459a,a12463a,a12464a,a12465a,a12469a,a12470a,a12474a,a12475a,a12476a,a12479a,a12483a,a12484a,a12485a,a12489a,a12490a,a12494a,a12495a,a12496a,a12499a,a12503a,a12504a,a12505a,a12509a,a12510a,a12514a,a12515a,a12516a,a12519a,a12523a,a12524a,a12525a,a12529a,a12530a,a12534a,a12535a,a12536a,a12539a,a12543a,a12544a,a12545a,a12549a,a12550a,a12554a,a12555a,a12556a,a12559a,a12563a,a12564a,a12565a,a12569a,a12570a,a12574a,a12575a,a12576a,a12579a,a12583a,a12584a,a12585a,a12589a,a12590a,a12594a,a12595a,a12596a,a12599a,a12603a,a12604a,a12605a,a12609a,a12610a,a12614a,a12615a,a12616a,a12619a,a12623a,a12624a,a12625a,a12629a,a12630a,a12634a,a12635a,a12636a,a12639a,a12643a,a12644a,a12645a,a12649a,a12650a,a12654a,a12655a,a12656a,a12659a,a12663a,a12664a,a12665a,a12669a,a12670a,a12674a,a12675a,a12676a,a12679a,a12683a,a12684a,a12685a,a12689a,a12690a,a12694a,a12695a,a12696a,a12699a,a12703a,a12704a,a12705a,a12709a,a12710a,a12714a,a12715a,a12716a,a12719a,a12723a,a12724a,a12725a,a12729a,a12730a,a12734a,a12735a,a12736a,a12739a,a12743a,a12744a,a12745a,a12749a,a12750a,a12754a,a12755a,a12756a,a12759a,a12763a,a12764a,a12765a,a12769a,a12770a,a12774a,a12775a,a12776a,a12779a,a12783a,a12784a,a12785a,a12789a,a12790a,a12794a,a12795a,a12796a,a12799a,a12803a,a12804a,a12805a,a12809a,a12810a,a12814a,a12815a,a12816a,a12819a,a12823a,a12824a,a12825a,a12829a,a12830a,a12834a,a12835a,a12836a,a12839a,a12843a,a12844a,a12845a,a12849a,a12850a,a12854a,a12855a,a12856a,a12859a,a12863a,a12864a,a12865a,a12869a,a12870a,a12874a,a12875a,a12876a,a12879a,a12883a,a12884a,a12885a,a12889a,a12890a,a12894a,a12895a,a12896a,a12899a,a12903a,a12904a,a12905a,a12909a,a12910a,a12914a,a12915a,a12916a,a12919a,a12923a,a12924a,a12925a,a12929a,a12930a,a12934a,a12935a,a12936a,a12939a,a12943a,a12944a,a12945a,a12949a,a12950a,a12954a,a12955a,a12956a,a12959a,a12963a,a12964a,a12965a,a12969a,a12970a,a12974a,a12975a,a12976a,a12979a,a12983a,a12984a,a12985a,a12989a,a12990a,a12994a,a12995a,a12996a,a12999a,a13003a,a13004a,a13005a,a13009a,a13010a,a13014a,a13015a,a13016a,a13019a,a13023a,a13024a,a13025a,a13029a,a13030a,a13034a,a13035a,a13036a,a13039a,a13043a,a13044a,a13045a,a13049a,a13050a,a13054a,a13055a,a13056a,a13059a,a13063a,a13064a,a13065a,a13069a,a13070a,a13074a,a13075a,a13076a,a13079a,a13083a,a13084a,a13085a,a13089a,a13090a,a13094a,a13095a,a13096a,a13099a,a13103a,a13104a,a13105a,a13109a,a13110a,a13114a,a13115a,a13116a,a13119a,a13123a,a13124a,a13125a,a13129a,a13130a,a13134a,a13135a,a13136a,a13139a,a13143a,a13144a,a13145a,a13149a,a13150a,a13154a,a13155a,a13156a,a13159a,a13163a,a13164a,a13165a,a13169a,a13170a,a13174a,a13175a,a13176a,a13179a,a13183a,a13184a,a13185a,a13189a,a13190a,a13194a,a13195a,a13196a,a13199a,a13203a,a13204a,a13205a,a13209a,a13210a,a13214a,a13215a,a13216a,a13219a,a13223a,a13224a,a13225a,a13229a,a13230a,a13234a,a13235a,a13236a,a13239a,a13243a,a13244a,a13245a,a13249a,a13250a,a13254a,a13255a,a13256a,a13259a,a13263a,a13264a,a13265a,a13269a,a13270a,a13274a,a13275a,a13276a,a13279a,a13283a,a13284a,a13285a,a13289a,a13290a,a13294a,a13295a,a13296a,a13299a,a13303a,a13304a,a13305a,a13309a,a13310a,a13314a,a13315a,a13316a,a13319a,a13323a,a13324a,a13325a,a13329a,a13330a,a13334a,a13335a,a13336a,a13339a,a13343a,a13344a,a13345a,a13349a,a13350a,a13354a,a13355a,a13356a,a13359a,a13363a,a13364a,a13365a,a13369a,a13370a,a13374a,a13375a,a13376a,a13379a,a13383a,a13384a,a13385a,a13389a,a13390a,a13394a,a13395a,a13396a,a13399a,a13403a,a13404a,a13405a,a13409a,a13410a,a13414a,a13415a,a13416a,a13419a,a13423a,a13424a,a13425a,a13429a,a13430a,a13434a,a13435a,a13436a,a13439a,a13443a,a13444a,a13445a,a13449a,a13450a,a13454a,a13455a,a13456a,a13459a,a13463a,a13464a,a13465a,a13469a,a13470a,a13474a,a13475a,a13476a,a13479a,a13483a,a13484a,a13485a,a13489a,a13490a,a13494a,a13495a,a13496a,a13499a,a13503a,a13504a,a13505a,a13509a,a13510a,a13514a,a13515a,a13516a,a13519a,a13523a,a13524a,a13525a,a13529a,a13530a,a13534a,a13535a,a13536a,a13539a,a13543a,a13544a,a13545a,a13549a,a13550a,a13554a,a13555a,a13556a,a13559a,a13563a,a13564a,a13565a,a13569a,a13570a,a13574a,a13575a,a13576a,a13579a,a13583a,a13584a,a13585a,a13589a,a13590a,a13594a,a13595a,a13596a,a13599a,a13603a,a13604a,a13605a,a13609a,a13610a,a13614a,a13615a,a13616a,a13619a,a13623a,a13624a,a13625a,a13629a,a13630a,a13634a,a13635a,a13636a,a13639a,a13643a,a13644a,a13645a,a13649a,a13650a,a13654a,a13655a,a13656a,a13659a,a13663a,a13664a,a13665a,a13669a,a13670a,a13674a,a13675a,a13676a,a13679a,a13683a,a13684a,a13685a,a13689a,a13690a,a13694a,a13695a,a13696a,a13699a,a13703a,a13704a,a13705a,a13709a,a13710a,a13714a,a13715a,a13716a,a13719a,a13723a,a13724a,a13725a,a13729a,a13730a,a13734a,a13735a,a13736a,a13739a,a13743a,a13744a,a13745a,a13749a,a13750a,a13754a,a13755a,a13756a,a13759a,a13763a,a13764a,a13765a,a13769a,a13770a,a13774a,a13775a,a13776a,a13779a,a13783a,a13784a,a13785a,a13789a,a13790a,a13794a,a13795a,a13796a,a13799a,a13803a,a13804a,a13805a,a13809a,a13810a,a13814a,a13815a,a13816a,a13819a,a13823a,a13824a,a13825a,a13829a,a13830a,a13834a,a13835a,a13836a,a13839a,a13843a,a13844a,a13845a,a13849a,a13850a,a13854a,a13855a,a13856a,a13859a,a13863a,a13864a,a13865a,a13869a,a13870a,a13874a,a13875a,a13876a,a13879a,a13883a,a13884a,a13885a,a13889a,a13890a,a13894a,a13895a,a13896a,a13899a,a13903a,a13904a,a13905a,a13909a,a13910a,a13914a,a13915a,a13916a,a13919a,a13923a,a13924a,a13925a,a13929a,a13930a,a13934a,a13935a,a13936a,a13939a,a13943a,a13944a,a13945a,a13949a,a13950a,a13954a,a13955a,a13956a,a13959a,a13963a,a13964a,a13965a,a13969a,a13970a,a13974a,a13975a,a13976a,a13979a,a13983a,a13984a,a13985a,a13989a,a13990a,a13994a,a13995a,a13996a,a13999a,a14003a,a14004a,a14005a,a14009a,a14010a,a14014a,a14015a,a14016a,a14019a,a14023a,a14024a,a14025a,a14029a,a14030a,a14034a,a14035a,a14036a,a14039a,a14043a,a14044a,a14045a,a14049a,a14050a,a14054a,a14055a,a14056a,a14059a,a14063a,a14064a,a14065a,a14069a,a14070a,a14074a,a14075a,a14076a,a14079a,a14083a,a14084a,a14085a,a14089a,a14090a,a14094a,a14095a,a14096a,a14099a,a14103a,a14104a,a14105a,a14109a,a14110a,a14114a,a14115a,a14116a,a14119a,a14123a,a14124a,a14125a,a14129a,a14130a,a14134a,a14135a,a14136a,a14139a,a14143a,a14144a,a14145a,a14149a,a14150a,a14154a,a14155a,a14156a,a14159a,a14163a,a14164a,a14165a,a14169a,a14170a,a14174a,a14175a,a14176a,a14179a,a14183a,a14184a,a14185a,a14189a,a14190a,a14194a,a14195a,a14196a,a14199a,a14203a,a14204a,a14205a,a14209a,a14210a,a14214a,a14215a,a14216a,a14219a,a14223a,a14224a,a14225a,a14229a,a14230a,a14234a,a14235a,a14236a,a14239a,a14243a,a14244a,a14245a,a14249a,a14250a,a14254a,a14255a,a14256a,a14259a,a14263a,a14264a,a14265a,a14269a,a14270a,a14274a,a14275a,a14276a,a14279a,a14283a,a14284a,a14285a,a14289a,a14290a,a14294a,a14295a,a14296a,a14299a,a14303a,a14304a,a14305a,a14309a,a14310a,a14314a,a14315a,a14316a,a14319a,a14323a,a14324a,a14325a,a14329a,a14330a,a14334a,a14335a,a14336a,a14339a,a14343a,a14344a,a14345a,a14349a,a14350a,a14354a,a14355a,a14356a,a14359a,a14363a,a14364a,a14365a,a14369a,a14370a,a14374a,a14375a,a14376a,a14379a,a14383a,a14384a,a14385a,a14389a,a14390a,a14394a,a14395a,a14396a,a14399a,a14403a,a14404a,a14405a,a14409a,a14410a,a14414a,a14415a,a14416a,a14419a,a14423a,a14424a,a14425a,a14429a,a14430a,a14434a,a14435a,a14436a,a14439a,a14443a,a14444a,a14445a,a14449a,a14450a,a14454a,a14455a,a14456a,a14459a,a14463a,a14464a,a14465a,a14469a,a14470a,a14474a,a14475a,a14476a,a14479a,a14483a,a14484a,a14485a,a14489a,a14490a,a14494a,a14495a,a14496a,a14499a,a14503a,a14504a,a14505a,a14509a,a14510a,a14514a,a14515a,a14516a,a14519a,a14523a,a14524a,a14525a,a14529a,a14530a,a14534a,a14535a,a14536a,a14539a,a14543a,a14544a,a14545a,a14549a,a14550a,a14554a,a14555a,a14556a,a14559a,a14563a,a14564a,a14565a,a14569a,a14570a,a14574a,a14575a,a14576a,a14579a,a14583a,a14584a,a14585a,a14589a,a14590a,a14594a,a14595a,a14596a,a14599a,a14603a,a14604a,a14605a,a14609a,a14610a,a14614a,a14615a,a14616a,a14619a,a14623a,a14624a,a14625a,a14629a,a14630a,a14634a,a14635a,a14636a,a14639a,a14643a,a14644a,a14645a,a14649a,a14650a,a14654a,a14655a,a14656a,a14659a,a14663a,a14664a,a14665a,a14669a,a14670a,a14674a,a14675a,a14676a,a14679a,a14683a,a14684a,a14685a,a14689a,a14690a,a14694a,a14695a,a14696a,a14699a,a14703a,a14704a,a14705a,a14709a,a14710a,a14714a,a14715a,a14716a,a14719a,a14723a,a14724a,a14725a,a14729a,a14730a,a14734a,a14735a,a14736a,a14739a,a14743a,a14744a,a14745a,a14749a,a14750a,a14754a,a14755a,a14756a,a14759a,a14763a,a14764a,a14765a,a14769a,a14770a,a14774a,a14775a,a14776a,a14779a,a14783a,a14784a,a14785a,a14789a,a14790a,a14794a,a14795a,a14796a,a14799a,a14803a,a14804a,a14805a,a14809a,a14810a,a14814a,a14815a,a14816a,a14819a,a14823a,a14824a,a14825a,a14829a,a14830a,a14834a,a14835a,a14836a,a14839a,a14843a,a14844a,a14845a,a14849a,a14850a,a14854a,a14855a,a14856a,a14859a,a14863a,a14864a,a14865a,a14869a,a14870a,a14874a,a14875a,a14876a,a14879a,a14883a,a14884a,a14885a,a14889a,a14890a,a14894a,a14895a,a14896a,a14899a,a14903a,a14904a,a14905a,a14909a,a14910a,a14914a,a14915a,a14916a,a14919a,a14923a,a14924a,a14925a,a14929a,a14930a,a14934a,a14935a,a14936a,a14940a,a14941a,a14945a,a14946a,a14947a,a14951a,a14952a,a14956a,a14957a,a14958a,a14962a,a14963a,a14967a,a14968a,a14969a,a14973a,a14974a,a14978a,a14979a,a14980a,a14984a,a14985a,a14989a,a14990a,a14991a,a14995a,a14996a,a15000a,a15001a,a15002a,a15006a,a15007a,a15011a,a15012a,a15013a,a15017a,a15018a,a15022a,a15023a,a15024a,a15028a,a15029a,a15033a,a15034a,a15035a,a15039a,a15040a,a15044a,a15045a,a15046a,a15050a,a15051a,a15055a,a15056a,a15057a,a15061a,a15062a,a15066a,a15067a,a15068a,a15072a,a15073a,a15077a,a15078a,a15079a,a15083a,a15084a,a15088a,a15089a,a15090a,a15094a,a15095a,a15099a,a15100a,a15101a,a15105a,a15106a,a15110a,a15111a,a15112a,a15116a,a15117a,a15121a,a15122a,a15123a,a15127a,a15128a,a15132a,a15133a,a15134a,a15138a,a15139a,a15143a,a15144a,a15145a,a15149a,a15150a,a15154a,a15155a,a15156a,a15160a,a15161a,a15165a,a15166a,a15167a,a15171a,a15172a,a15176a,a15177a,a15178a,a15182a,a15183a,a15187a,a15188a,a15189a,a15193a,a15194a,a15198a,a15199a,a15200a,a15204a,a15205a,a15209a,a15210a,a15211a,a15215a,a15216a,a15220a,a15221a,a15222a,a15226a,a15227a,a15231a,a15232a,a15233a,a15237a,a15238a,a15242a,a15243a,a15244a,a15248a,a15249a,a15253a,a15254a,a15255a,a15259a,a15260a,a15264a,a15265a,a15266a,a15270a,a15271a,a15275a,a15276a,a15277a,a15281a,a15282a,a15286a,a15287a,a15288a,a15292a,a15293a,a15297a,a15298a,a15299a,a15303a,a15304a,a15308a,a15309a,a15310a,a15314a,a15315a,a15319a,a15320a,a15321a,a15325a,a15326a,a15330a,a15331a,a15332a,a15336a,a15337a,a15341a,a15342a,a15343a,a15347a,a15348a,a15352a,a15353a,a15354a,a15358a,a15359a,a15363a,a15364a,a15365a,a15369a,a15370a,a15374a,a15375a,a15376a,a15380a,a15381a,a15385a,a15386a,a15387a,a15391a,a15392a,a15396a,a15397a,a15398a,a15402a,a15403a,a15407a,a15408a,a15409a,a15413a,a15414a,a15418a,a15419a,a15420a,a15424a,a15425a,a15429a,a15430a,a15431a,a15435a,a15436a,a15440a,a15441a,a15442a,a15446a,a15447a,a15451a,a15452a,a15453a,a15457a,a15458a,a15462a,a15463a,a15464a,a15468a,a15469a,a15473a,a15474a,a15475a,a15479a,a15480a,a15484a,a15485a,a15486a,a15490a,a15491a,a15495a,a15496a,a15497a,a15501a,a15502a,a15506a,a15507a,a15508a,a15512a,a15513a,a15517a,a15518a,a15519a,a15523a,a15524a,a15528a,a15529a,a15530a,a15534a,a15535a,a15539a,a15540a,a15541a,a15545a,a15546a,a15550a,a15551a,a15552a,a15556a,a15557a,a15561a,a15562a,a15563a,a15567a,a15568a,a15572a,a15573a,a15574a,a15578a,a15579a,a15583a,a15584a,a15585a,a15589a,a15590a,a15594a,a15595a,a15596a,a15600a,a15601a,a15605a,a15606a,a15607a,a15611a,a15612a,a15616a,a15617a,a15618a,a15622a,a15623a,a15627a,a15628a,a15629a,a15633a,a15634a,a15638a,a15639a,a15640a,a15644a,a15645a,a15649a,a15650a,a15651a,a15655a,a15656a,a15660a,a15661a,a15662a,a15666a,a15667a,a15671a,a15672a,a15673a,a15677a,a15678a,a15682a,a15683a,a15684a,a15688a,a15689a,a15693a,a15694a,a15695a,a15699a,a15700a,a15704a,a15705a,a15706a,a15710a,a15711a,a15715a,a15716a,a15717a,a15721a,a15722a,a15726a,a15727a,a15728a,a15732a,a15733a,a15737a,a15738a,a15739a,a15743a,a15744a,a15748a,a15749a,a15750a,a15754a,a15755a,a15759a,a15760a,a15761a,a15765a,a15766a,a15770a,a15771a,a15772a,a15776a,a15777a,a15781a,a15782a,a15783a,a15787a,a15788a,a15792a,a15793a,a15794a,a15798a,a15799a,a15803a,a15804a,a15805a,a15809a,a15810a,a15814a,a15815a,a15816a,a15820a,a15821a,a15825a,a15826a,a15827a,a15831a,a15832a,a15836a,a15837a,a15838a,a15842a,a15843a,a15847a,a15848a,a15849a,a15853a,a15854a,a15858a,a15859a,a15860a,a15864a,a15865a,a15869a,a15870a,a15871a,a15875a,a15876a,a15880a,a15881a,a15882a,a15886a,a15887a,a15891a,a15892a,a15893a,a15897a,a15898a,a15902a,a15903a,a15904a,a15908a,a15909a,a15913a,a15914a,a15915a,a15919a,a15920a,a15924a,a15925a,a15926a,a15930a,a15931a,a15935a,a15936a,a15937a,a15941a,a15942a,a15946a,a15947a,a15948a,a15952a,a15953a,a15957a,a15958a,a15959a,a15963a,a15964a,a15968a,a15969a,a15970a,a15974a,a15975a,a15979a,a15980a,a15981a,a15985a,a15986a,a15990a,a15991a,a15992a,a15996a,a15997a,a16001a,a16002a,a16003a,a16007a,a16008a,a16012a,a16013a,a16014a,a16018a,a16019a,a16023a,a16024a,a16025a,a16029a,a16030a,a16034a,a16035a,a16036a,a16040a,a16041a,a16045a,a16046a,a16047a,a16051a,a16052a,a16056a,a16057a,a16058a,a16062a,a16063a,a16067a,a16068a,a16069a,a16073a,a16074a,a16078a,a16079a,a16080a,a16084a,a16085a,a16089a,a16090a,a16091a,a16095a,a16096a,a16100a,a16101a,a16102a,a16106a,a16107a,a16111a,a16112a,a16113a,a16117a,a16118a,a16122a,a16123a,a16124a,a16128a,a16129a,a16133a,a16134a,a16135a,a16139a,a16140a,a16144a,a16145a,a16146a,a16150a,a16151a,a16155a,a16156a,a16157a,a16161a,a16162a,a16166a,a16167a,a16168a,a16172a,a16173a,a16177a,a16178a,a16179a,a16183a,a16184a,a16188a,a16189a,a16190a,a16194a,a16195a,a16199a,a16200a,a16201a,a16205a,a16206a,a16210a,a16211a,a16212a,a16216a,a16217a,a16221a,a16222a,a16223a,a16227a,a16228a,a16232a,a16233a,a16234a,a16238a,a16239a,a16243a,a16244a,a16245a,a16249a,a16250a,a16254a,a16255a,a16256a,a16260a,a16261a,a16265a,a16266a,a16267a,a16271a,a16272a,a16276a,a16277a,a16278a,a16282a,a16283a,a16287a,a16288a,a16289a,a16293a,a16294a,a16298a,a16299a,a16300a,a16304a,a16305a,a16309a,a16310a,a16311a,a16315a,a16316a,a16320a,a16321a,a16322a,a16326a,a16327a,a16331a,a16332a,a16333a,a16337a,a16338a,a16342a,a16343a,a16344a,a16348a,a16349a,a16353a,a16354a,a16355a,a16359a,a16360a,a16364a,a16365a,a16366a,a16370a,a16371a,a16375a,a16376a,a16377a,a16381a,a16382a,a16386a,a16387a,a16388a,a16392a,a16393a,a16397a,a16398a,a16399a,a16403a,a16404a,a16408a,a16409a,a16410a,a16414a,a16415a,a16419a,a16420a,a16421a,a16425a,a16426a,a16430a,a16431a,a16432a,a16436a,a16437a,a16441a,a16442a,a16443a,a16447a,a16448a,a16452a,a16453a,a16454a,a16458a,a16459a,a16463a,a16464a,a16465a,a16469a,a16470a,a16474a,a16475a,a16476a,a16480a,a16481a,a16485a,a16486a,a16487a,a16491a,a16492a,a16496a,a16497a,a16498a,a16502a,a16503a,a16507a,a16508a,a16509a,a16513a,a16514a,a16518a,a16519a,a16520a,a16524a,a16525a,a16529a,a16530a,a16531a,a16535a,a16536a,a16540a,a16541a,a16542a,a16546a,a16547a,a16551a,a16552a,a16553a,a16557a,a16558a,a16562a,a16563a,a16564a,a16568a,a16569a,a16573a,a16574a,a16575a,a16579a,a16580a,a16584a,a16585a,a16586a,a16590a,a16591a,a16595a,a16596a,a16597a,a16601a,a16602a,a16606a,a16607a,a16608a,a16612a,a16613a,a16617a,a16618a,a16619a,a16623a,a16624a,a16628a,a16629a,a16630a,a16634a,a16635a,a16639a,a16640a,a16641a,a16645a,a16646a,a16650a,a16651a,a16652a,a16656a,a16657a,a16661a,a16662a,a16663a,a16667a,a16668a,a16672a,a16673a,a16674a,a16678a,a16679a,a16683a,a16684a,a16685a,a16689a,a16690a,a16694a,a16695a,a16696a,a16700a,a16701a,a16705a,a16706a,a16707a,a16711a,a16712a,a16716a,a16717a,a16718a,a16722a,a16723a,a16727a,a16728a,a16729a,a16733a,a16734a,a16738a,a16739a,a16740a,a16744a,a16745a,a16749a,a16750a,a16751a,a16755a,a16756a,a16760a,a16761a,a16762a,a16766a,a16767a,a16771a,a16772a,a16773a,a16777a,a16778a,a16782a,a16783a,a16784a,a16788a,a16789a,a16793a,a16794a,a16795a,a16799a,a16800a,a16804a,a16805a,a16806a,a16810a,a16811a,a16815a,a16816a,a16817a,a16821a,a16822a,a16826a,a16827a,a16828a,a16832a,a16833a,a16837a,a16838a,a16839a,a16843a,a16844a,a16848a,a16849a,a16850a,a16854a,a16855a,a16859a,a16860a,a16861a,a16865a,a16866a,a16870a,a16871a,a16872a,a16876a,a16877a,a16881a,a16882a,a16883a,a16887a,a16888a,a16892a,a16893a,a16894a,a16898a,a16899a,a16903a,a16904a,a16905a,a16909a,a16910a,a16914a,a16915a,a16916a,a16920a,a16921a,a16925a,a16926a,a16927a,a16931a,a16932a,a16936a,a16937a,a16938a,a16942a,a16943a,a16947a,a16948a,a16949a,a16953a,a16954a,a16958a,a16959a,a16960a,a16964a,a16965a,a16969a,a16970a,a16971a,a16975a,a16976a,a16980a,a16981a,a16982a,a16986a,a16987a,a16991a,a16992a,a16993a,a16997a,a16998a,a17002a,a17003a,a17004a,a17008a,a17009a,a17013a,a17014a,a17015a,a17019a,a17020a,a17024a,a17025a,a17026a,a17030a,a17031a,a17035a,a17036a,a17037a,a17041a,a17042a,a17046a,a17047a,a17048a,a17052a,a17053a,a17057a,a17058a,a17059a,a17063a,a17064a,a17068a,a17069a,a17070a,a17074a,a17075a,a17079a,a17080a,a17081a,a17085a,a17086a,a17090a,a17091a,a17092a,a17096a,a17097a,a17101a,a17102a,a17103a,a17107a,a17108a,a17112a,a17113a,a17114a,a17118a,a17119a,a17123a,a17124a,a17125a,a17129a,a17130a,a17134a,a17135a,a17136a,a17140a,a17141a,a17145a,a17146a,a17147a,a17151a,a17152a,a17156a,a17157a,a17158a,a17162a,a17163a,a17167a,a17168a,a17169a,a17173a,a17174a,a17178a,a17179a,a17180a,a17184a,a17185a,a17189a,a17190a,a17191a,a17195a,a17196a,a17200a,a17201a,a17202a,a17206a,a17207a,a17211a,a17212a,a17213a,a17217a,a17218a,a17222a,a17223a,a17224a,a17228a,a17229a,a17233a,a17234a,a17235a,a17239a,a17240a,a17244a,a17245a,a17246a,a17250a,a17251a,a17255a,a17256a,a17257a,a17261a,a17262a,a17266a,a17267a,a17268a,a17272a,a17273a,a17277a,a17278a,a17279a,a17283a,a17284a,a17288a,a17289a,a17290a,a17294a,a17295a,a17299a,a17300a,a17301a,a17305a,a17306a,a17310a,a17311a,a17312a,a17316a,a17317a,a17321a,a17322a,a17323a,a17327a,a17328a,a17332a,a17333a,a17334a,a17338a,a17339a,a17343a,a17344a,a17345a,a17349a,a17350a,a17354a,a17355a,a17356a,a17360a,a17361a,a17365a,a17366a,a17367a,a17371a,a17372a,a17376a,a17377a,a17378a,a17382a,a17383a,a17387a,a17388a,a17389a,a17393a,a17394a,a17398a,a17399a,a17400a,a17404a,a17405a,a17409a,a17410a,a17411a,a17415a,a17416a,a17420a,a17421a,a17422a,a17426a,a17427a,a17431a,a17432a,a17433a,a17437a,a17438a,a17442a,a17443a,a17444a,a17448a,a17449a,a17453a,a17454a,a17455a,a17459a,a17460a,a17464a,a17465a,a17466a,a17470a,a17471a,a17475a,a17476a,a17477a,a17481a,a17482a,a17486a,a17487a,a17488a,a17492a,a17493a,a17497a,a17498a,a17499a,a17503a,a17504a,a17508a,a17509a,a17510a,a17514a,a17515a,a17519a,a17520a,a17521a,a17525a,a17526a,a17530a,a17531a,a17532a,a17536a,a17537a,a17541a,a17542a,a17543a,a17547a,a17548a,a17552a,a17553a,a17554a,a17558a,a17559a,a17563a,a17564a,a17565a,a17569a,a17570a,a17574a,a17575a,a17576a,a17580a,a17581a,a17585a,a17586a,a17587a,a17591a,a17592a,a17596a,a17597a,a17598a,a17602a,a17603a,a17607a,a17608a,a17609a,a17613a,a17614a,a17618a,a17619a,a17620a,a17624a,a17625a,a17629a,a17630a,a17631a,a17635a,a17636a,a17640a,a17641a,a17642a,a17646a,a17647a,a17651a,a17652a,a17653a,a17657a,a17658a,a17662a,a17663a,a17664a,a17668a,a17669a,a17673a,a17674a,a17675a,a17679a,a17680a,a17684a,a17685a,a17686a,a17690a,a17691a,a17695a,a17696a,a17697a,a17701a,a17702a,a17706a,a17707a,a17708a,a17712a,a17713a,a17717a,a17718a,a17719a,a17723a,a17724a,a17728a,a17729a,a17730a,a17734a,a17735a,a17739a,a17740a,a17741a,a17745a,a17746a,a17750a,a17751a,a17752a,a17756a,a17757a,a17761a,a17762a,a17763a,a17767a,a17768a,a17772a,a17773a,a17774a,a17778a,a17779a,a17783a,a17784a,a17785a,a17789a,a17790a,a17794a,a17795a,a17796a,a17800a,a17801a,a17805a,a17806a,a17807a,a17811a,a17812a,a17816a,a17817a,a17818a,a17822a,a17823a,a17827a,a17828a,a17829a,a17833a,a17834a,a17838a,a17839a,a17840a,a17844a,a17845a,a17849a,a17850a,a17851a,a17855a,a17856a,a17860a,a17861a,a17862a,a17866a,a17867a,a17871a,a17872a,a17873a,a17877a,a17878a,a17882a,a17883a,a17884a,a17888a,a17889a,a17893a,a17894a,a17895a,a17899a,a17900a,a17904a,a17905a,a17906a,a17910a,a17911a,a17915a,a17916a,a17917a,a17921a,a17922a,a17926a,a17927a,a17928a,a17932a,a17933a,a17937a,a17938a,a17939a,a17943a,a17944a,a17948a,a17949a,a17950a,a17954a,a17955a,a17959a,a17960a,a17961a,a17965a,a17966a,a17970a,a17971a,a17972a,a17976a,a17977a,a17981a,a17982a,a17983a,a17987a,a17988a,a17992a,a17993a,a17994a,a17998a,a17999a,a18003a,a18004a,a18005a,a18009a,a18010a,a18014a,a18015a,a18016a,a18020a,a18021a,a18025a,a18026a,a18027a,a18031a,a18032a,a18036a,a18037a,a18038a,a18042a,a18043a,a18047a,a18048a,a18049a,a18053a,a18054a,a18058a,a18059a,a18060a,a18064a,a18065a,a18069a,a18070a,a18071a,a18075a,a18076a,a18080a,a18081a,a18082a,a18086a,a18087a,a18091a,a18092a,a18093a,a18097a,a18098a,a18102a,a18103a,a18104a,a18108a,a18109a,a18113a,a18114a,a18115a,a18119a,a18120a,a18124a,a18125a,a18126a,a18130a,a18131a,a18135a,a18136a,a18137a,a18141a,a18142a,a18146a,a18147a,a18148a,a18152a,a18153a,a18157a,a18158a,a18159a,a18163a,a18164a,a18168a,a18169a,a18170a,a18174a,a18175a,a18179a,a18180a,a18181a,a18185a,a18186a,a18190a,a18191a,a18192a,a18196a,a18197a,a18201a,a18202a,a18203a,a18207a,a18208a,a18212a,a18213a,a18214a,a18218a,a18219a,a18223a,a18224a,a18225a,a18229a,a18230a,a18234a,a18235a,a18236a,a18240a,a18241a,a18245a,a18246a,a18247a,a18251a,a18252a,a18256a,a18257a,a18258a,a18262a,a18263a,a18267a,a18268a,a18269a,a18273a,a18274a,a18278a,a18279a,a18280a,a18284a,a18285a,a18289a,a18290a,a18291a,a18295a,a18296a,a18300a,a18301a,a18302a,a18306a,a18307a,a18311a,a18312a,a18313a,a18317a,a18318a,a18322a,a18323a,a18324a,a18328a,a18329a,a18333a,a18334a,a18335a,a18339a,a18340a,a18344a,a18345a,a18346a,a18350a,a18351a,a18355a,a18356a,a18357a,a18361a,a18362a,a18366a,a18367a,a18368a,a18372a,a18373a,a18377a,a18378a,a18379a,a18383a,a18384a,a18388a,a18389a,a18390a,a18394a,a18395a,a18399a,a18400a,a18401a,a18405a,a18406a,a18410a,a18411a,a18412a,a18416a,a18417a,a18421a,a18422a,a18423a,a18427a,a18428a,a18432a,a18433a,a18434a,a18438a,a18439a,a18443a,a18444a,a18445a,a18449a,a18450a,a18454a,a18455a,a18456a,a18460a,a18461a,a18465a,a18466a,a18467a,a18471a,a18472a,a18476a,a18477a,a18478a,a18482a,a18483a,a18487a,a18488a,a18489a,a18493a,a18494a,a18498a,a18499a,a18500a,a18504a,a18505a,a18509a,a18510a,a18511a,a18515a,a18516a,a18520a,a18521a,a18522a,a18526a,a18527a,a18531a,a18532a,a18533a,a18537a,a18538a,a18542a,a18543a,a18544a,a18548a,a18549a,a18553a,a18554a,a18555a,a18559a,a18560a,a18564a,a18565a,a18566a,a18570a,a18571a,a18575a,a18576a,a18577a,a18581a,a18582a,a18586a,a18587a,a18588a,a18592a,a18593a,a18597a,a18598a,a18599a,a18603a,a18604a,a18608a,a18609a,a18610a,a18614a,a18615a,a18619a,a18620a,a18621a,a18625a,a18626a,a18630a,a18631a,a18632a,a18636a,a18637a,a18641a,a18642a,a18643a,a18647a,a18648a,a18652a,a18653a,a18654a,a18658a,a18659a,a18663a,a18664a,a18665a,a18669a,a18670a,a18674a,a18675a,a18676a,a18680a,a18681a,a18685a,a18686a,a18687a,a18691a,a18692a,a18696a,a18697a,a18698a,a18702a,a18703a,a18707a,a18708a,a18709a,a18713a,a18714a,a18718a,a18719a,a18720a,a18724a,a18725a,a18729a,a18730a,a18731a,a18735a,a18736a,a18740a,a18741a,a18742a,a18746a,a18747a,a18751a,a18752a,a18753a,a18757a,a18758a,a18762a,a18763a,a18764a,a18768a,a18769a,a18773a,a18774a,a18775a,a18779a,a18780a,a18784a,a18785a,a18786a,a18790a,a18791a,a18795a,a18796a,a18797a,a18801a,a18802a,a18806a,a18807a,a18808a,a18812a,a18813a,a18817a,a18818a,a18819a,a18823a,a18824a,a18828a,a18829a,a18830a,a18834a,a18835a,a18839a,a18840a,a18841a,a18845a,a18846a,a18850a,a18851a,a18852a,a18856a,a18857a,a18861a,a18862a,a18863a,a18867a,a18868a,a18872a,a18873a,a18874a,a18878a,a18879a,a18883a,a18884a,a18885a,a18889a,a18890a,a18894a,a18895a,a18896a,a18900a,a18901a,a18905a,a18906a,a18907a,a18911a,a18912a,a18916a,a18917a,a18918a,a18922a,a18923a,a18927a,a18928a,a18929a,a18933a,a18934a,a18938a,a18939a,a18940a,a18944a,a18945a,a18949a,a18950a,a18951a,a18955a,a18956a,a18960a,a18961a,a18962a,a18966a,a18967a,a18971a,a18972a,a18973a,a18977a,a18978a,a18982a,a18983a,a18984a,a18988a,a18989a,a18993a,a18994a,a18995a,a18999a,a19000a,a19004a,a19005a,a19006a,a19010a,a19011a,a19015a,a19016a,a19017a,a19021a,a19022a,a19026a,a19027a,a19028a,a19032a,a19033a,a19037a,a19038a,a19039a,a19043a,a19044a,a19048a,a19049a,a19050a,a19054a,a19055a,a19059a,a19060a,a19061a,a19065a,a19066a,a19070a,a19071a,a19072a,a19076a,a19077a,a19081a,a19082a,a19083a,a19087a,a19088a,a19092a,a19093a,a19094a,a19098a,a19099a,a19103a,a19104a,a19105a,a19109a,a19110a,a19114a,a19115a,a19116a,a19120a,a19121a,a19125a,a19126a,a19127a,a19131a,a19132a,a19136a,a19137a,a19138a,a19142a,a19143a,a19147a,a19148a,a19149a,a19153a,a19154a,a19158a,a19159a,a19160a,a19164a,a19165a,a19169a,a19170a,a19171a,a19175a,a19176a,a19180a,a19181a,a19182a,a19186a,a19187a,a19191a,a19192a,a19193a,a19197a,a19198a,a19202a,a19203a,a19204a,a19208a,a19209a,a19213a,a19214a,a19215a,a19219a,a19220a,a19224a,a19225a,a19226a,a19230a,a19231a,a19235a,a19236a,a19237a,a19241a,a19242a,a19246a,a19247a,a19248a,a19252a,a19253a,a19257a,a19258a,a19259a,a19263a,a19264a,a19268a,a19269a,a19270a,a19274a,a19275a,a19279a,a19280a,a19281a,a19285a,a19286a,a19290a,a19291a,a19292a,a19296a,a19297a,a19301a,a19302a,a19303a,a19307a,a19308a,a19311a,a19314a,a19315a,a19316a,a19320a,a19321a,a19325a,a19326a,a19327a,a19331a,a19332a,a19335a,a19338a,a19339a,a19340a,a19344a,a19345a,a19349a,a19350a,a19351a,a19355a,a19356a,a19359a,a19362a,a19363a,a19364a,a19368a,a19369a,a19373a,a19374a,a19375a,a19379a,a19380a,a19383a,a19386a,a19387a,a19388a,a19392a,a19393a,a19397a,a19398a,a19399a,a19403a,a19404a,a19407a,a19410a,a19411a,a19412a,a19416a,a19417a,a19421a,a19422a,a19423a,a19427a,a19428a,a19431a,a19434a,a19435a,a19436a,a19440a,a19441a,a19445a,a19446a,a19447a,a19451a,a19452a,a19455a,a19458a,a19459a,a19460a,a19464a,a19465a,a19469a,a19470a,a19471a,a19475a,a19476a,a19479a,a19482a,a19483a,a19484a,a19488a,a19489a,a19493a,a19494a,a19495a,a19499a,a19500a,a19503a,a19506a,a19507a,a19508a,a19512a,a19513a,a19517a,a19518a,a19519a,a19523a,a19524a,a19527a,a19530a,a19531a,a19532a,a19536a,a19537a,a19541a,a19542a,a19543a,a19547a,a19548a,a19551a,a19554a,a19555a,a19556a,a19560a,a19561a,a19565a,a19566a,a19567a,a19571a,a19572a,a19575a,a19578a,a19579a,a19580a,a19584a,a19585a,a19589a,a19590a,a19591a,a19595a,a19596a,a19599a,a19602a,a19603a,a19604a,a19608a,a19609a,a19613a,a19614a,a19615a,a19619a,a19620a,a19623a,a19626a,a19627a,a19628a,a19632a,a19633a,a19637a,a19638a,a19639a,a19643a,a19644a,a19647a,a19650a,a19651a,a19652a,a19656a,a19657a,a19661a,a19662a,a19663a,a19667a,a19668a,a19671a,a19674a,a19675a,a19676a,a19680a,a19681a,a19685a,a19686a,a19687a,a19691a,a19692a,a19695a,a19698a,a19699a,a19700a,a19704a,a19705a,a19709a,a19710a,a19711a,a19715a,a19716a,a19719a,a19722a,a19723a,a19724a,a19728a,a19729a,a19733a,a19734a,a19735a,a19739a,a19740a,a19743a,a19746a,a19747a,a19748a,a19752a,a19753a,a19757a,a19758a,a19759a,a19763a,a19764a,a19767a,a19770a,a19771a,a19772a,a19776a,a19777a,a19781a,a19782a,a19783a,a19787a,a19788a,a19791a,a19794a,a19795a,a19796a,a19800a,a19801a,a19805a,a19806a,a19807a,a19811a,a19812a,a19815a,a19818a,a19819a,a19820a,a19824a,a19825a,a19829a,a19830a,a19831a,a19835a,a19836a,a19839a,a19842a,a19843a,a19844a,a19848a,a19849a,a19853a,a19854a,a19855a,a19859a,a19860a,a19863a,a19866a,a19867a,a19868a,a19872a,a19873a,a19877a,a19878a,a19879a,a19883a,a19884a,a19887a,a19890a,a19891a,a19892a,a19896a,a19897a,a19901a,a19902a,a19903a,a19907a,a19908a,a19911a,a19914a,a19915a,a19916a,a19920a,a19921a,a19925a,a19926a,a19927a,a19931a,a19932a,a19935a,a19938a,a19939a,a19940a,a19944a,a19945a,a19949a,a19950a,a19951a,a19955a,a19956a,a19959a,a19962a,a19963a,a19964a,a19968a,a19969a,a19973a,a19974a,a19975a,a19979a,a19980a,a19983a,a19986a,a19987a,a19988a,a19992a,a19993a,a19997a,a19998a,a19999a,a20003a,a20004a,a20007a,a20010a,a20011a,a20012a,a20016a,a20017a,a20021a,a20022a,a20023a,a20027a,a20028a,a20031a,a20034a,a20035a,a20036a,a20040a,a20041a,a20045a,a20046a,a20047a,a20051a,a20052a,a20055a,a20058a,a20059a,a20060a,a20064a,a20065a,a20069a,a20070a,a20071a,a20075a,a20076a,a20079a,a20082a,a20083a,a20084a,a20088a,a20089a,a20093a,a20094a,a20095a,a20099a,a20100a,a20103a,a20106a,a20107a,a20108a,a20112a,a20113a,a20117a,a20118a,a20119a,a20123a,a20124a,a20127a,a20130a,a20131a,a20132a,a20136a,a20137a,a20141a,a20142a,a20143a,a20147a,a20148a,a20151a,a20154a,a20155a,a20156a,a20160a,a20161a,a20165a,a20166a,a20167a,a20171a,a20172a,a20175a,a20178a,a20179a,a20180a,a20184a,a20185a,a20189a,a20190a,a20191a,a20195a,a20196a,a20199a,a20202a,a20203a,a20204a,a20208a,a20209a,a20213a,a20214a,a20215a,a20219a,a20220a,a20223a,a20226a,a20227a,a20228a,a20232a,a20233a,a20237a,a20238a,a20239a,a20243a,a20244a,a20247a,a20250a,a20251a,a20252a,a20256a,a20257a,a20261a,a20262a,a20263a,a20267a,a20268a,a20271a,a20274a,a20275a,a20276a,a20280a,a20281a,a20285a,a20286a,a20287a,a20291a,a20292a,a20295a,a20298a,a20299a,a20300a,a20304a,a20305a,a20309a,a20310a,a20311a,a20315a,a20316a,a20319a,a20322a,a20323a,a20324a,a20328a,a20329a,a20333a,a20334a,a20335a,a20339a,a20340a,a20343a,a20346a,a20347a,a20348a,a20352a,a20353a,a20357a,a20358a,a20359a,a20363a,a20364a,a20367a,a20370a,a20371a,a20372a,a20376a,a20377a,a20381a,a20382a,a20383a,a20387a,a20388a,a20391a,a20394a,a20395a,a20396a,a20400a,a20401a,a20405a,a20406a,a20407a,a20411a,a20412a,a20415a,a20418a,a20419a,a20420a,a20424a,a20425a,a20429a,a20430a,a20431a,a20435a,a20436a,a20439a,a20442a,a20443a,a20444a,a20448a,a20449a,a20453a,a20454a,a20455a,a20459a,a20460a,a20463a,a20466a,a20467a,a20468a,a20472a,a20473a,a20477a,a20478a,a20479a,a20483a,a20484a,a20487a,a20490a,a20491a,a20492a,a20496a,a20497a,a20501a,a20502a,a20503a,a20507a,a20508a,a20511a,a20514a,a20515a,a20516a,a20520a,a20521a,a20525a,a20526a,a20527a,a20531a,a20532a,a20535a,a20538a,a20539a,a20540a,a20544a,a20545a,a20549a,a20550a,a20551a,a20555a,a20556a,a20559a,a20562a,a20563a,a20564a,a20568a,a20569a,a20573a,a20574a,a20575a,a20579a,a20580a,a20583a,a20586a,a20587a,a20588a,a20592a,a20593a,a20597a,a20598a,a20599a,a20603a,a20604a,a20607a,a20610a,a20611a,a20612a,a20616a,a20617a,a20621a,a20622a,a20623a,a20627a,a20628a,a20631a,a20634a,a20635a,a20636a,a20640a,a20641a,a20645a,a20646a,a20647a,a20651a,a20652a,a20655a,a20658a,a20659a,a20660a,a20664a,a20665a,a20669a,a20670a,a20671a,a20675a,a20676a,a20679a,a20682a,a20683a,a20684a,a20688a,a20689a,a20693a,a20694a,a20695a,a20699a,a20700a,a20703a,a20706a,a20707a,a20708a,a20712a,a20713a,a20717a,a20718a,a20719a,a20723a,a20724a,a20727a,a20730a,a20731a,a20732a,a20736a,a20737a,a20741a,a20742a,a20743a,a20747a,a20748a,a20751a,a20754a,a20755a,a20756a,a20760a,a20761a,a20765a,a20766a,a20767a,a20771a,a20772a,a20775a,a20778a,a20779a,a20780a,a20784a,a20785a,a20789a,a20790a,a20791a,a20795a,a20796a,a20799a,a20802a,a20803a,a20804a,a20808a,a20809a,a20813a,a20814a,a20815a,a20819a,a20820a,a20823a,a20826a,a20827a,a20828a,a20832a,a20833a,a20837a,a20838a,a20839a,a20843a,a20844a,a20847a,a20850a,a20851a,a20852a,a20856a,a20857a,a20861a,a20862a,a20863a,a20867a,a20868a,a20871a,a20874a,a20875a,a20876a,a20880a,a20881a,a20885a,a20886a,a20887a,a20891a,a20892a,a20895a,a20898a,a20899a,a20900a,a20904a,a20905a,a20909a,a20910a,a20911a,a20915a,a20916a,a20919a,a20922a,a20923a,a20924a,a20928a,a20929a,a20933a,a20934a,a20935a,a20939a,a20940a,a20943a,a20946a,a20947a,a20948a,a20952a,a20953a,a20957a,a20958a,a20959a,a20963a,a20964a,a20967a,a20970a,a20971a,a20972a,a20976a,a20977a,a20981a,a20982a,a20983a,a20987a,a20988a,a20991a,a20994a,a20995a,a20996a,a21000a,a21001a,a21005a,a21006a,a21007a,a21011a,a21012a,a21015a,a21018a,a21019a,a21020a,a21024a,a21025a,a21029a,a21030a,a21031a,a21035a,a21036a,a21039a,a21042a,a21043a,a21044a,a21048a,a21049a,a21053a,a21054a,a21055a,a21059a,a21060a,a21063a,a21066a,a21067a,a21068a,a21072a,a21073a,a21077a,a21078a,a21079a,a21083a,a21084a,a21087a,a21090a,a21091a,a21092a,a21096a,a21097a,a21101a,a21102a,a21103a,a21107a,a21108a,a21111a,a21114a,a21115a,a21116a,a21120a,a21121a,a21125a,a21126a,a21127a,a21131a,a21132a,a21135a,a21138a,a21139a,a21140a,a21144a,a21145a,a21149a,a21150a,a21151a,a21155a,a21156a,a21159a,a21162a,a21163a,a21164a,a21168a,a21169a,a21173a,a21174a,a21175a,a21179a,a21180a,a21183a,a21186a,a21187a,a21188a,a21192a,a21193a,a21197a,a21198a,a21199a,a21203a,a21204a,a21207a,a21210a,a21211a,a21212a,a21216a,a21217a,a21221a,a21222a,a21223a,a21227a,a21228a,a21231a,a21234a,a21235a,a21236a,a21240a,a21241a,a21245a,a21246a,a21247a,a21251a,a21252a,a21255a,a21258a,a21259a,a21260a,a21264a,a21265a,a21269a,a21270a,a21271a,a21275a,a21276a,a21279a,a21282a,a21283a,a21284a,a21288a,a21289a,a21293a,a21294a,a21295a,a21299a,a21300a,a21303a,a21306a,a21307a,a21308a,a21312a,a21313a,a21317a,a21318a,a21319a,a21323a,a21324a,a21327a,a21330a,a21331a,a21332a,a21336a,a21337a,a21341a,a21342a,a21343a,a21347a,a21348a,a21351a,a21354a,a21355a,a21356a,a21360a,a21361a,a21365a,a21366a,a21367a,a21371a,a21372a,a21375a,a21378a,a21379a,a21380a,a21384a,a21385a,a21389a,a21390a,a21391a,a21395a,a21396a,a21399a,a21402a,a21403a,a21404a,a21408a,a21409a,a21413a,a21414a,a21415a,a21419a,a21420a,a21423a,a21426a,a21427a,a21428a,a21432a,a21433a,a21437a,a21438a,a21439a,a21443a,a21444a,a21447a,a21450a,a21451a,a21452a,a21456a,a21457a,a21461a,a21462a,a21463a,a21467a,a21468a,a21471a,a21474a,a21475a,a21476a,a21480a,a21481a,a21485a,a21486a,a21487a,a21491a,a21492a,a21495a,a21498a,a21499a,a21500a,a21504a,a21505a,a21509a,a21510a,a21511a,a21515a,a21516a,a21519a,a21522a,a21523a,a21524a,a21528a,a21529a,a21532a,a21535a,a21536a,a21537a,a21541a,a21542a,a21545a,a21548a,a21549a,a21550a,a21554a,a21555a,a21558a,a21561a,a21562a,a21563a,a21567a,a21568a,a21571a,a21574a,a21575a,a21576a,a21580a,a21581a,a21584a,a21587a,a21588a,a21589a,a21593a,a21594a,a21597a,a21600a,a21601a,a21602a,a21606a,a21607a,a21610a,a21613a,a21614a,a21615a,a21619a,a21620a,a21623a,a21626a,a21627a,a21628a,a21632a,a21633a,a21636a,a21639a,a21640a,a21641a,a21645a,a21646a,a21649a,a21652a,a21653a,a21654a,a21658a,a21659a,a21662a,a21665a,a21666a,a21667a,a21671a,a21672a,a21675a,a21678a,a21679a,a21680a,a21684a,a21685a,a21688a,a21691a,a21692a,a21693a,a21697a,a21698a,a21701a,a21704a,a21705a,a21706a,a21710a,a21711a,a21714a,a21717a,a21718a,a21719a,a21723a,a21724a,a21727a,a21730a,a21731a,a21732a,a21736a,a21737a,a21740a,a21743a,a21744a,a21745a,a21749a,a21750a,a21753a,a21756a,a21757a,a21758a,a21762a,a21763a,a21766a,a21769a,a21770a,a21771a,a21775a,a21776a,a21779a,a21782a,a21783a,a21784a,a21788a,a21789a,a21792a,a21795a,a21796a,a21797a,a21801a,a21802a,a21805a,a21808a,a21809a,a21810a,a21814a,a21815a,a21818a,a21821a,a21822a,a21823a,a21827a,a21828a,a21831a,a21834a,a21835a,a21836a,a21840a,a21841a,a21844a,a21847a,a21848a,a21849a,a21853a,a21854a,a21857a,a21860a,a21861a,a21862a,a21866a,a21867a,a21870a,a21873a,a21874a,a21875a,a21879a,a21880a,a21883a,a21886a,a21887a,a21888a,a21892a,a21893a,a21896a,a21899a,a21900a,a21901a,a21905a,a21906a,a21909a,a21912a,a21913a,a21914a,a21918a,a21919a,a21922a,a21925a,a21926a,a21927a,a21931a,a21932a,a21935a,a21938a,a21939a,a21940a,a21944a,a21945a,a21948a,a21951a,a21952a,a21953a,a21957a,a21958a,a21961a,a21964a,a21965a,a21966a,a21970a,a21971a,a21974a,a21977a,a21978a,a21979a,a21983a,a21984a,a21987a,a21990a,a21991a,a21992a,a21996a,a21997a,a22000a,a22003a,a22004a,a22005a,a22009a,a22010a,a22013a,a22016a,a22017a,a22018a,a22022a,a22023a,a22026a,a22029a,a22030a,a22031a,a22035a,a22036a,a22039a,a22042a,a22043a,a22044a,a22048a,a22049a,a22052a,a22055a,a22056a,a22057a,a22061a,a22062a,a22065a,a22068a,a22069a,a22070a,a22074a,a22075a,a22078a,a22081a,a22082a,a22083a,a22087a,a22088a,a22091a,a22094a,a22095a,a22096a,a22100a,a22101a,a22104a,a22107a,a22108a,a22109a,a22112a,a22115a,a22116a,a22119a,a22122a,a22123a,a22124a,a22128a,a22129a,a22132a,a22135a,a22136a,a22137a,a22140a,a22143a,a22144a,a22147a,a22150a,a22151a,a22152a: std_logic;
begin

A73 <=( a3028a ) or ( a2019a );
 a1a <=( a22152a  and  a22137a );
 a2a <=( a22124a  and  a22109a );
 a3a <=( a22096a  and  a22083a );
 a4a <=( a22070a  and  a22057a );
 a5a <=( a22044a  and  a22031a );
 a6a <=( a22018a  and  a22005a );
 a7a <=( a21992a  and  a21979a );
 a8a <=( a21966a  and  a21953a );
 a9a <=( a21940a  and  a21927a );
 a10a <=( a21914a  and  a21901a );
 a11a <=( a21888a  and  a21875a );
 a12a <=( a21862a  and  a21849a );
 a13a <=( a21836a  and  a21823a );
 a14a <=( a21810a  and  a21797a );
 a15a <=( a21784a  and  a21771a );
 a16a <=( a21758a  and  a21745a );
 a17a <=( a21732a  and  a21719a );
 a18a <=( a21706a  and  a21693a );
 a19a <=( a21680a  and  a21667a );
 a20a <=( a21654a  and  a21641a );
 a21a <=( a21628a  and  a21615a );
 a22a <=( a21602a  and  a21589a );
 a23a <=( a21576a  and  a21563a );
 a24a <=( a21550a  and  a21537a );
 a25a <=( a21524a  and  a21511a );
 a26a <=( a21500a  and  a21487a );
 a27a <=( a21476a  and  a21463a );
 a28a <=( a21452a  and  a21439a );
 a29a <=( a21428a  and  a21415a );
 a30a <=( a21404a  and  a21391a );
 a31a <=( a21380a  and  a21367a );
 a32a <=( a21356a  and  a21343a );
 a33a <=( a21332a  and  a21319a );
 a34a <=( a21308a  and  a21295a );
 a35a <=( a21284a  and  a21271a );
 a36a <=( a21260a  and  a21247a );
 a37a <=( a21236a  and  a21223a );
 a38a <=( a21212a  and  a21199a );
 a39a <=( a21188a  and  a21175a );
 a40a <=( a21164a  and  a21151a );
 a41a <=( a21140a  and  a21127a );
 a42a <=( a21116a  and  a21103a );
 a43a <=( a21092a  and  a21079a );
 a44a <=( a21068a  and  a21055a );
 a45a <=( a21044a  and  a21031a );
 a46a <=( a21020a  and  a21007a );
 a47a <=( a20996a  and  a20983a );
 a48a <=( a20972a  and  a20959a );
 a49a <=( a20948a  and  a20935a );
 a50a <=( a20924a  and  a20911a );
 a51a <=( a20900a  and  a20887a );
 a52a <=( a20876a  and  a20863a );
 a53a <=( a20852a  and  a20839a );
 a54a <=( a20828a  and  a20815a );
 a55a <=( a20804a  and  a20791a );
 a56a <=( a20780a  and  a20767a );
 a57a <=( a20756a  and  a20743a );
 a58a <=( a20732a  and  a20719a );
 a59a <=( a20708a  and  a20695a );
 a60a <=( a20684a  and  a20671a );
 a61a <=( a20660a  and  a20647a );
 a62a <=( a20636a  and  a20623a );
 a63a <=( a20612a  and  a20599a );
 a64a <=( a20588a  and  a20575a );
 a65a <=( a20564a  and  a20551a );
 a66a <=( a20540a  and  a20527a );
 a67a <=( a20516a  and  a20503a );
 a68a <=( a20492a  and  a20479a );
 a69a <=( a20468a  and  a20455a );
 a70a <=( a20444a  and  a20431a );
 a71a <=( a20420a  and  a20407a );
 a72a <=( a20396a  and  a20383a );
 a73a <=( a20372a  and  a20359a );
 a74a <=( a20348a  and  a20335a );
 a75a <=( a20324a  and  a20311a );
 a76a <=( a20300a  and  a20287a );
 a77a <=( a20276a  and  a20263a );
 a78a <=( a20252a  and  a20239a );
 a79a <=( a20228a  and  a20215a );
 a80a <=( a20204a  and  a20191a );
 a81a <=( a20180a  and  a20167a );
 a82a <=( a20156a  and  a20143a );
 a83a <=( a20132a  and  a20119a );
 a84a <=( a20108a  and  a20095a );
 a85a <=( a20084a  and  a20071a );
 a86a <=( a20060a  and  a20047a );
 a87a <=( a20036a  and  a20023a );
 a88a <=( a20012a  and  a19999a );
 a89a <=( a19988a  and  a19975a );
 a90a <=( a19964a  and  a19951a );
 a91a <=( a19940a  and  a19927a );
 a92a <=( a19916a  and  a19903a );
 a93a <=( a19892a  and  a19879a );
 a94a <=( a19868a  and  a19855a );
 a95a <=( a19844a  and  a19831a );
 a96a <=( a19820a  and  a19807a );
 a97a <=( a19796a  and  a19783a );
 a98a <=( a19772a  and  a19759a );
 a99a <=( a19748a  and  a19735a );
 a100a <=( a19724a  and  a19711a );
 a101a <=( a19700a  and  a19687a );
 a102a <=( a19676a  and  a19663a );
 a103a <=( a19652a  and  a19639a );
 a104a <=( a19628a  and  a19615a );
 a105a <=( a19604a  and  a19591a );
 a106a <=( a19580a  and  a19567a );
 a107a <=( a19556a  and  a19543a );
 a108a <=( a19532a  and  a19519a );
 a109a <=( a19508a  and  a19495a );
 a110a <=( a19484a  and  a19471a );
 a111a <=( a19460a  and  a19447a );
 a112a <=( a19436a  and  a19423a );
 a113a <=( a19412a  and  a19399a );
 a114a <=( a19388a  and  a19375a );
 a115a <=( a19364a  and  a19351a );
 a116a <=( a19340a  and  a19327a );
 a117a <=( a19316a  and  a19303a );
 a118a <=( a19292a  and  a19281a );
 a119a <=( a19270a  and  a19259a );
 a120a <=( a19248a  and  a19237a );
 a121a <=( a19226a  and  a19215a );
 a122a <=( a19204a  and  a19193a );
 a123a <=( a19182a  and  a19171a );
 a124a <=( a19160a  and  a19149a );
 a125a <=( a19138a  and  a19127a );
 a126a <=( a19116a  and  a19105a );
 a127a <=( a19094a  and  a19083a );
 a128a <=( a19072a  and  a19061a );
 a129a <=( a19050a  and  a19039a );
 a130a <=( a19028a  and  a19017a );
 a131a <=( a19006a  and  a18995a );
 a132a <=( a18984a  and  a18973a );
 a133a <=( a18962a  and  a18951a );
 a134a <=( a18940a  and  a18929a );
 a135a <=( a18918a  and  a18907a );
 a136a <=( a18896a  and  a18885a );
 a137a <=( a18874a  and  a18863a );
 a138a <=( a18852a  and  a18841a );
 a139a <=( a18830a  and  a18819a );
 a140a <=( a18808a  and  a18797a );
 a141a <=( a18786a  and  a18775a );
 a142a <=( a18764a  and  a18753a );
 a143a <=( a18742a  and  a18731a );
 a144a <=( a18720a  and  a18709a );
 a145a <=( a18698a  and  a18687a );
 a146a <=( a18676a  and  a18665a );
 a147a <=( a18654a  and  a18643a );
 a148a <=( a18632a  and  a18621a );
 a149a <=( a18610a  and  a18599a );
 a150a <=( a18588a  and  a18577a );
 a151a <=( a18566a  and  a18555a );
 a152a <=( a18544a  and  a18533a );
 a153a <=( a18522a  and  a18511a );
 a154a <=( a18500a  and  a18489a );
 a155a <=( a18478a  and  a18467a );
 a156a <=( a18456a  and  a18445a );
 a157a <=( a18434a  and  a18423a );
 a158a <=( a18412a  and  a18401a );
 a159a <=( a18390a  and  a18379a );
 a160a <=( a18368a  and  a18357a );
 a161a <=( a18346a  and  a18335a );
 a162a <=( a18324a  and  a18313a );
 a163a <=( a18302a  and  a18291a );
 a164a <=( a18280a  and  a18269a );
 a165a <=( a18258a  and  a18247a );
 a166a <=( a18236a  and  a18225a );
 a167a <=( a18214a  and  a18203a );
 a168a <=( a18192a  and  a18181a );
 a169a <=( a18170a  and  a18159a );
 a170a <=( a18148a  and  a18137a );
 a171a <=( a18126a  and  a18115a );
 a172a <=( a18104a  and  a18093a );
 a173a <=( a18082a  and  a18071a );
 a174a <=( a18060a  and  a18049a );
 a175a <=( a18038a  and  a18027a );
 a176a <=( a18016a  and  a18005a );
 a177a <=( a17994a  and  a17983a );
 a178a <=( a17972a  and  a17961a );
 a179a <=( a17950a  and  a17939a );
 a180a <=( a17928a  and  a17917a );
 a181a <=( a17906a  and  a17895a );
 a182a <=( a17884a  and  a17873a );
 a183a <=( a17862a  and  a17851a );
 a184a <=( a17840a  and  a17829a );
 a185a <=( a17818a  and  a17807a );
 a186a <=( a17796a  and  a17785a );
 a187a <=( a17774a  and  a17763a );
 a188a <=( a17752a  and  a17741a );
 a189a <=( a17730a  and  a17719a );
 a190a <=( a17708a  and  a17697a );
 a191a <=( a17686a  and  a17675a );
 a192a <=( a17664a  and  a17653a );
 a193a <=( a17642a  and  a17631a );
 a194a <=( a17620a  and  a17609a );
 a195a <=( a17598a  and  a17587a );
 a196a <=( a17576a  and  a17565a );
 a197a <=( a17554a  and  a17543a );
 a198a <=( a17532a  and  a17521a );
 a199a <=( a17510a  and  a17499a );
 a200a <=( a17488a  and  a17477a );
 a201a <=( a17466a  and  a17455a );
 a202a <=( a17444a  and  a17433a );
 a203a <=( a17422a  and  a17411a );
 a204a <=( a17400a  and  a17389a );
 a205a <=( a17378a  and  a17367a );
 a206a <=( a17356a  and  a17345a );
 a207a <=( a17334a  and  a17323a );
 a208a <=( a17312a  and  a17301a );
 a209a <=( a17290a  and  a17279a );
 a210a <=( a17268a  and  a17257a );
 a211a <=( a17246a  and  a17235a );
 a212a <=( a17224a  and  a17213a );
 a213a <=( a17202a  and  a17191a );
 a214a <=( a17180a  and  a17169a );
 a215a <=( a17158a  and  a17147a );
 a216a <=( a17136a  and  a17125a );
 a217a <=( a17114a  and  a17103a );
 a218a <=( a17092a  and  a17081a );
 a219a <=( a17070a  and  a17059a );
 a220a <=( a17048a  and  a17037a );
 a221a <=( a17026a  and  a17015a );
 a222a <=( a17004a  and  a16993a );
 a223a <=( a16982a  and  a16971a );
 a224a <=( a16960a  and  a16949a );
 a225a <=( a16938a  and  a16927a );
 a226a <=( a16916a  and  a16905a );
 a227a <=( a16894a  and  a16883a );
 a228a <=( a16872a  and  a16861a );
 a229a <=( a16850a  and  a16839a );
 a230a <=( a16828a  and  a16817a );
 a231a <=( a16806a  and  a16795a );
 a232a <=( a16784a  and  a16773a );
 a233a <=( a16762a  and  a16751a );
 a234a <=( a16740a  and  a16729a );
 a235a <=( a16718a  and  a16707a );
 a236a <=( a16696a  and  a16685a );
 a237a <=( a16674a  and  a16663a );
 a238a <=( a16652a  and  a16641a );
 a239a <=( a16630a  and  a16619a );
 a240a <=( a16608a  and  a16597a );
 a241a <=( a16586a  and  a16575a );
 a242a <=( a16564a  and  a16553a );
 a243a <=( a16542a  and  a16531a );
 a244a <=( a16520a  and  a16509a );
 a245a <=( a16498a  and  a16487a );
 a246a <=( a16476a  and  a16465a );
 a247a <=( a16454a  and  a16443a );
 a248a <=( a16432a  and  a16421a );
 a249a <=( a16410a  and  a16399a );
 a250a <=( a16388a  and  a16377a );
 a251a <=( a16366a  and  a16355a );
 a252a <=( a16344a  and  a16333a );
 a253a <=( a16322a  and  a16311a );
 a254a <=( a16300a  and  a16289a );
 a255a <=( a16278a  and  a16267a );
 a256a <=( a16256a  and  a16245a );
 a257a <=( a16234a  and  a16223a );
 a258a <=( a16212a  and  a16201a );
 a259a <=( a16190a  and  a16179a );
 a260a <=( a16168a  and  a16157a );
 a261a <=( a16146a  and  a16135a );
 a262a <=( a16124a  and  a16113a );
 a263a <=( a16102a  and  a16091a );
 a264a <=( a16080a  and  a16069a );
 a265a <=( a16058a  and  a16047a );
 a266a <=( a16036a  and  a16025a );
 a267a <=( a16014a  and  a16003a );
 a268a <=( a15992a  and  a15981a );
 a269a <=( a15970a  and  a15959a );
 a270a <=( a15948a  and  a15937a );
 a271a <=( a15926a  and  a15915a );
 a272a <=( a15904a  and  a15893a );
 a273a <=( a15882a  and  a15871a );
 a274a <=( a15860a  and  a15849a );
 a275a <=( a15838a  and  a15827a );
 a276a <=( a15816a  and  a15805a );
 a277a <=( a15794a  and  a15783a );
 a278a <=( a15772a  and  a15761a );
 a279a <=( a15750a  and  a15739a );
 a280a <=( a15728a  and  a15717a );
 a281a <=( a15706a  and  a15695a );
 a282a <=( a15684a  and  a15673a );
 a283a <=( a15662a  and  a15651a );
 a284a <=( a15640a  and  a15629a );
 a285a <=( a15618a  and  a15607a );
 a286a <=( a15596a  and  a15585a );
 a287a <=( a15574a  and  a15563a );
 a288a <=( a15552a  and  a15541a );
 a289a <=( a15530a  and  a15519a );
 a290a <=( a15508a  and  a15497a );
 a291a <=( a15486a  and  a15475a );
 a292a <=( a15464a  and  a15453a );
 a293a <=( a15442a  and  a15431a );
 a294a <=( a15420a  and  a15409a );
 a295a <=( a15398a  and  a15387a );
 a296a <=( a15376a  and  a15365a );
 a297a <=( a15354a  and  a15343a );
 a298a <=( a15332a  and  a15321a );
 a299a <=( a15310a  and  a15299a );
 a300a <=( a15288a  and  a15277a );
 a301a <=( a15266a  and  a15255a );
 a302a <=( a15244a  and  a15233a );
 a303a <=( a15222a  and  a15211a );
 a304a <=( a15200a  and  a15189a );
 a305a <=( a15178a  and  a15167a );
 a306a <=( a15156a  and  a15145a );
 a307a <=( a15134a  and  a15123a );
 a308a <=( a15112a  and  a15101a );
 a309a <=( a15090a  and  a15079a );
 a310a <=( a15068a  and  a15057a );
 a311a <=( a15046a  and  a15035a );
 a312a <=( a15024a  and  a15013a );
 a313a <=( a15002a  and  a14991a );
 a314a <=( a14980a  and  a14969a );
 a315a <=( a14958a  and  a14947a );
 a316a <=( a14936a  and  a14925a );
 a317a <=( a14916a  and  a14905a );
 a318a <=( a14896a  and  a14885a );
 a319a <=( a14876a  and  a14865a );
 a320a <=( a14856a  and  a14845a );
 a321a <=( a14836a  and  a14825a );
 a322a <=( a14816a  and  a14805a );
 a323a <=( a14796a  and  a14785a );
 a324a <=( a14776a  and  a14765a );
 a325a <=( a14756a  and  a14745a );
 a326a <=( a14736a  and  a14725a );
 a327a <=( a14716a  and  a14705a );
 a328a <=( a14696a  and  a14685a );
 a329a <=( a14676a  and  a14665a );
 a330a <=( a14656a  and  a14645a );
 a331a <=( a14636a  and  a14625a );
 a332a <=( a14616a  and  a14605a );
 a333a <=( a14596a  and  a14585a );
 a334a <=( a14576a  and  a14565a );
 a335a <=( a14556a  and  a14545a );
 a336a <=( a14536a  and  a14525a );
 a337a <=( a14516a  and  a14505a );
 a338a <=( a14496a  and  a14485a );
 a339a <=( a14476a  and  a14465a );
 a340a <=( a14456a  and  a14445a );
 a341a <=( a14436a  and  a14425a );
 a342a <=( a14416a  and  a14405a );
 a343a <=( a14396a  and  a14385a );
 a344a <=( a14376a  and  a14365a );
 a345a <=( a14356a  and  a14345a );
 a346a <=( a14336a  and  a14325a );
 a347a <=( a14316a  and  a14305a );
 a348a <=( a14296a  and  a14285a );
 a349a <=( a14276a  and  a14265a );
 a350a <=( a14256a  and  a14245a );
 a351a <=( a14236a  and  a14225a );
 a352a <=( a14216a  and  a14205a );
 a353a <=( a14196a  and  a14185a );
 a354a <=( a14176a  and  a14165a );
 a355a <=( a14156a  and  a14145a );
 a356a <=( a14136a  and  a14125a );
 a357a <=( a14116a  and  a14105a );
 a358a <=( a14096a  and  a14085a );
 a359a <=( a14076a  and  a14065a );
 a360a <=( a14056a  and  a14045a );
 a361a <=( a14036a  and  a14025a );
 a362a <=( a14016a  and  a14005a );
 a363a <=( a13996a  and  a13985a );
 a364a <=( a13976a  and  a13965a );
 a365a <=( a13956a  and  a13945a );
 a366a <=( a13936a  and  a13925a );
 a367a <=( a13916a  and  a13905a );
 a368a <=( a13896a  and  a13885a );
 a369a <=( a13876a  and  a13865a );
 a370a <=( a13856a  and  a13845a );
 a371a <=( a13836a  and  a13825a );
 a372a <=( a13816a  and  a13805a );
 a373a <=( a13796a  and  a13785a );
 a374a <=( a13776a  and  a13765a );
 a375a <=( a13756a  and  a13745a );
 a376a <=( a13736a  and  a13725a );
 a377a <=( a13716a  and  a13705a );
 a378a <=( a13696a  and  a13685a );
 a379a <=( a13676a  and  a13665a );
 a380a <=( a13656a  and  a13645a );
 a381a <=( a13636a  and  a13625a );
 a382a <=( a13616a  and  a13605a );
 a383a <=( a13596a  and  a13585a );
 a384a <=( a13576a  and  a13565a );
 a385a <=( a13556a  and  a13545a );
 a386a <=( a13536a  and  a13525a );
 a387a <=( a13516a  and  a13505a );
 a388a <=( a13496a  and  a13485a );
 a389a <=( a13476a  and  a13465a );
 a390a <=( a13456a  and  a13445a );
 a391a <=( a13436a  and  a13425a );
 a392a <=( a13416a  and  a13405a );
 a393a <=( a13396a  and  a13385a );
 a394a <=( a13376a  and  a13365a );
 a395a <=( a13356a  and  a13345a );
 a396a <=( a13336a  and  a13325a );
 a397a <=( a13316a  and  a13305a );
 a398a <=( a13296a  and  a13285a );
 a399a <=( a13276a  and  a13265a );
 a400a <=( a13256a  and  a13245a );
 a401a <=( a13236a  and  a13225a );
 a402a <=( a13216a  and  a13205a );
 a403a <=( a13196a  and  a13185a );
 a404a <=( a13176a  and  a13165a );
 a405a <=( a13156a  and  a13145a );
 a406a <=( a13136a  and  a13125a );
 a407a <=( a13116a  and  a13105a );
 a408a <=( a13096a  and  a13085a );
 a409a <=( a13076a  and  a13065a );
 a410a <=( a13056a  and  a13045a );
 a411a <=( a13036a  and  a13025a );
 a412a <=( a13016a  and  a13005a );
 a413a <=( a12996a  and  a12985a );
 a414a <=( a12976a  and  a12965a );
 a415a <=( a12956a  and  a12945a );
 a416a <=( a12936a  and  a12925a );
 a417a <=( a12916a  and  a12905a );
 a418a <=( a12896a  and  a12885a );
 a419a <=( a12876a  and  a12865a );
 a420a <=( a12856a  and  a12845a );
 a421a <=( a12836a  and  a12825a );
 a422a <=( a12816a  and  a12805a );
 a423a <=( a12796a  and  a12785a );
 a424a <=( a12776a  and  a12765a );
 a425a <=( a12756a  and  a12745a );
 a426a <=( a12736a  and  a12725a );
 a427a <=( a12716a  and  a12705a );
 a428a <=( a12696a  and  a12685a );
 a429a <=( a12676a  and  a12665a );
 a430a <=( a12656a  and  a12645a );
 a431a <=( a12636a  and  a12625a );
 a432a <=( a12616a  and  a12605a );
 a433a <=( a12596a  and  a12585a );
 a434a <=( a12576a  and  a12565a );
 a435a <=( a12556a  and  a12545a );
 a436a <=( a12536a  and  a12525a );
 a437a <=( a12516a  and  a12505a );
 a438a <=( a12496a  and  a12485a );
 a439a <=( a12476a  and  a12465a );
 a440a <=( a12456a  and  a12445a );
 a441a <=( a12436a  and  a12425a );
 a442a <=( a12416a  and  a12405a );
 a443a <=( a12396a  and  a12385a );
 a444a <=( a12376a  and  a12365a );
 a445a <=( a12356a  and  a12345a );
 a446a <=( a12336a  and  a12325a );
 a447a <=( a12316a  and  a12305a );
 a448a <=( a12296a  and  a12285a );
 a449a <=( a12276a  and  a12265a );
 a450a <=( a12256a  and  a12245a );
 a451a <=( a12236a  and  a12225a );
 a452a <=( a12216a  and  a12205a );
 a453a <=( a12196a  and  a12185a );
 a454a <=( a12176a  and  a12165a );
 a455a <=( a12156a  and  a12145a );
 a456a <=( a12136a  and  a12125a );
 a457a <=( a12116a  and  a12105a );
 a458a <=( a12096a  and  a12085a );
 a459a <=( a12076a  and  a12065a );
 a460a <=( a12056a  and  a12045a );
 a461a <=( a12036a  and  a12025a );
 a462a <=( a12016a  and  a12005a );
 a463a <=( a11996a  and  a11985a );
 a464a <=( a11976a  and  a11965a );
 a465a <=( a11956a  and  a11945a );
 a466a <=( a11936a  and  a11925a );
 a467a <=( a11916a  and  a11905a );
 a468a <=( a11896a  and  a11885a );
 a469a <=( a11876a  and  a11865a );
 a470a <=( a11856a  and  a11845a );
 a471a <=( a11836a  and  a11825a );
 a472a <=( a11816a  and  a11805a );
 a473a <=( a11796a  and  a11785a );
 a474a <=( a11776a  and  a11765a );
 a475a <=( a11756a  and  a11745a );
 a476a <=( a11736a  and  a11725a );
 a477a <=( a11716a  and  a11705a );
 a478a <=( a11696a  and  a11685a );
 a479a <=( a11676a  and  a11665a );
 a480a <=( a11656a  and  a11645a );
 a481a <=( a11636a  and  a11625a );
 a482a <=( a11616a  and  a11605a );
 a483a <=( a11596a  and  a11585a );
 a484a <=( a11576a  and  a11565a );
 a485a <=( a11556a  and  a11545a );
 a486a <=( a11536a  and  a11525a );
 a487a <=( a11516a  and  a11505a );
 a488a <=( a11496a  and  a11485a );
 a489a <=( a11476a  and  a11465a );
 a490a <=( a11456a  and  a11445a );
 a491a <=( a11436a  and  a11425a );
 a492a <=( a11416a  and  a11405a );
 a493a <=( a11396a  and  a11385a );
 a494a <=( a11376a  and  a11365a );
 a495a <=( a11356a  and  a11345a );
 a496a <=( a11336a  and  a11325a );
 a497a <=( a11316a  and  a11305a );
 a498a <=( a11296a  and  a11285a );
 a499a <=( a11276a  and  a11265a );
 a500a <=( a11256a  and  a11245a );
 a501a <=( a11236a  and  a11225a );
 a502a <=( a11216a  and  a11205a );
 a503a <=( a11196a  and  a11185a );
 a504a <=( a11176a  and  a11165a );
 a505a <=( a11156a  and  a11145a );
 a506a <=( a11136a  and  a11125a );
 a507a <=( a11116a  and  a11105a );
 a508a <=( a11096a  and  a11085a );
 a509a <=( a11076a  and  a11065a );
 a510a <=( a11056a  and  a11045a );
 a511a <=( a11036a  and  a11025a );
 a512a <=( a11016a  and  a11005a );
 a513a <=( a10996a  and  a10985a );
 a514a <=( a10976a  and  a10965a );
 a515a <=( a10956a  and  a10945a );
 a516a <=( a10936a  and  a10925a );
 a517a <=( a10916a  and  a10905a );
 a518a <=( a10896a  and  a10885a );
 a519a <=( a10876a  and  a10865a );
 a520a <=( a10856a  and  a10845a );
 a521a <=( a10836a  and  a10825a );
 a522a <=( a10816a  and  a10805a );
 a523a <=( a10796a  and  a10785a );
 a524a <=( a10776a  and  a10765a );
 a525a <=( a10756a  and  a10745a );
 a526a <=( a10736a  and  a10725a );
 a527a <=( a10716a  and  a10705a );
 a528a <=( a10696a  and  a10685a );
 a529a <=( a10676a  and  a10665a );
 a530a <=( a10656a  and  a10645a );
 a531a <=( a10636a  and  a10625a );
 a532a <=( a10616a  and  a10605a );
 a533a <=( a10596a  and  a10585a );
 a534a <=( a10576a  and  a10565a );
 a535a <=( a10556a  and  a10545a );
 a536a <=( a10536a  and  a10525a );
 a537a <=( a10516a  and  a10505a );
 a538a <=( a10496a  and  a10485a );
 a539a <=( a10476a  and  a10465a );
 a540a <=( a10456a  and  a10445a );
 a541a <=( a10436a  and  a10425a );
 a542a <=( a10416a  and  a10405a );
 a543a <=( a10396a  and  a10385a );
 a544a <=( a10376a  and  a10365a );
 a545a <=( a10356a  and  a10345a );
 a546a <=( a10336a  and  a10325a );
 a547a <=( a10316a  and  a10305a );
 a548a <=( a10296a  and  a10285a );
 a549a <=( a10276a  and  a10265a );
 a550a <=( a10256a  and  a10245a );
 a551a <=( a10236a  and  a10225a );
 a552a <=( a10216a  and  a10205a );
 a553a <=( a10196a  and  a10185a );
 a554a <=( a10176a  and  a10165a );
 a555a <=( a10156a  and  a10145a );
 a556a <=( a10136a  and  a10125a );
 a557a <=( a10116a  and  a10105a );
 a558a <=( a10096a  and  a10085a );
 a559a <=( a10076a  and  a10065a );
 a560a <=( a10056a  and  a10045a );
 a561a <=( a10036a  and  a10025a );
 a562a <=( a10016a  and  a10005a );
 a563a <=( a9996a  and  a9985a );
 a564a <=( a9976a  and  a9967a );
 a565a <=( a9958a  and  a9949a );
 a566a <=( a9940a  and  a9931a );
 a567a <=( a9922a  and  a9913a );
 a568a <=( a9904a  and  a9895a );
 a569a <=( a9886a  and  a9877a );
 a570a <=( a9868a  and  a9859a );
 a571a <=( a9850a  and  a9841a );
 a572a <=( a9832a  and  a9823a );
 a573a <=( a9814a  and  a9805a );
 a574a <=( a9796a  and  a9787a );
 a575a <=( a9778a  and  a9769a );
 a576a <=( a9760a  and  a9751a );
 a577a <=( a9742a  and  a9733a );
 a578a <=( a9724a  and  a9715a );
 a579a <=( a9706a  and  a9697a );
 a580a <=( a9688a  and  a9679a );
 a581a <=( a9670a  and  a9661a );
 a582a <=( a9652a  and  a9643a );
 a583a <=( a9634a  and  a9625a );
 a584a <=( a9616a  and  a9607a );
 a585a <=( a9598a  and  a9589a );
 a586a <=( a9580a  and  a9571a );
 a587a <=( a9562a  and  a9553a );
 a588a <=( a9544a  and  a9535a );
 a589a <=( a9526a  and  a9517a );
 a590a <=( a9508a  and  a9499a );
 a591a <=( a9490a  and  a9481a );
 a592a <=( a9472a  and  a9463a );
 a593a <=( a9454a  and  a9445a );
 a594a <=( a9436a  and  a9427a );
 a595a <=( a9418a  and  a9409a );
 a596a <=( a9400a  and  a9391a );
 a597a <=( a9382a  and  a9373a );
 a598a <=( a9364a  and  a9355a );
 a599a <=( a9346a  and  a9337a );
 a600a <=( a9328a  and  a9319a );
 a601a <=( a9310a  and  a9301a );
 a602a <=( a9292a  and  a9283a );
 a603a <=( a9274a  and  a9265a );
 a604a <=( a9256a  and  a9247a );
 a605a <=( a9238a  and  a9229a );
 a606a <=( a9220a  and  a9211a );
 a607a <=( a9202a  and  a9193a );
 a608a <=( a9184a  and  a9175a );
 a609a <=( a9166a  and  a9157a );
 a610a <=( a9148a  and  a9139a );
 a611a <=( a9130a  and  a9121a );
 a612a <=( a9112a  and  a9103a );
 a613a <=( a9094a  and  a9085a );
 a614a <=( a9076a  and  a9067a );
 a615a <=( a9058a  and  a9049a );
 a616a <=( a9040a  and  a9031a );
 a617a <=( a9022a  and  a9013a );
 a618a <=( a9004a  and  a8995a );
 a619a <=( a8986a  and  a8977a );
 a620a <=( a8968a  and  a8959a );
 a621a <=( a8950a  and  a8941a );
 a622a <=( a8932a  and  a8923a );
 a623a <=( a8914a  and  a8905a );
 a624a <=( a8896a  and  a8887a );
 a625a <=( a8878a  and  a8869a );
 a626a <=( a8860a  and  a8851a );
 a627a <=( a8842a  and  a8833a );
 a628a <=( a8824a  and  a8815a );
 a629a <=( a8806a  and  a8797a );
 a630a <=( a8788a  and  a8779a );
 a631a <=( a8770a  and  a8761a );
 a632a <=( a8752a  and  a8743a );
 a633a <=( a8734a  and  a8725a );
 a634a <=( a8716a  and  a8707a );
 a635a <=( a8698a  and  a8689a );
 a636a <=( a8680a  and  a8671a );
 a637a <=( a8662a  and  a8653a );
 a638a <=( a8644a  and  a8635a );
 a639a <=( a8626a  and  a8617a );
 a640a <=( a8608a  and  a8599a );
 a641a <=( a8590a  and  a8581a );
 a642a <=( a8572a  and  a8563a );
 a643a <=( a8554a  and  a8545a );
 a644a <=( a8536a  and  a8527a );
 a645a <=( a8518a  and  a8509a );
 a646a <=( a8500a  and  a8491a );
 a647a <=( a8482a  and  a8473a );
 a648a <=( a8464a  and  a8455a );
 a649a <=( a8446a  and  a8437a );
 a650a <=( a8428a  and  a8419a );
 a651a <=( a8410a  and  a8401a );
 a652a <=( a8392a  and  a8383a );
 a653a <=( a8374a  and  a8365a );
 a654a <=( a8356a  and  a8347a );
 a655a <=( a8338a  and  a8329a );
 a656a <=( a8320a  and  a8311a );
 a657a <=( a8302a  and  a8293a );
 a658a <=( a8284a  and  a8275a );
 a659a <=( a8266a  and  a8257a );
 a660a <=( a8248a  and  a8239a );
 a661a <=( a8230a  and  a8221a );
 a662a <=( a8212a  and  a8203a );
 a663a <=( a8194a  and  a8185a );
 a664a <=( a8176a  and  a8167a );
 a665a <=( a8158a  and  a8149a );
 a666a <=( a8140a  and  a8131a );
 a667a <=( a8122a  and  a8113a );
 a668a <=( a8104a  and  a8095a );
 a669a <=( a8086a  and  a8077a );
 a670a <=( a8068a  and  a8059a );
 a671a <=( a8050a  and  a8041a );
 a672a <=( a8032a  and  a8023a );
 a673a <=( a8014a  and  a8005a );
 a674a <=( a7996a  and  a7987a );
 a675a <=( a7978a  and  a7969a );
 a676a <=( a7960a  and  a7951a );
 a677a <=( a7942a  and  a7933a );
 a678a <=( a7924a  and  a7915a );
 a679a <=( a7906a  and  a7897a );
 a680a <=( a7888a  and  a7879a );
 a681a <=( a7870a  and  a7861a );
 a682a <=( a7852a  and  a7843a );
 a683a <=( a7834a  and  a7825a );
 a684a <=( a7816a  and  a7807a );
 a685a <=( a7798a  and  a7789a );
 a686a <=( a7780a  and  a7771a );
 a687a <=( a7762a  and  a7753a );
 a688a <=( a7744a  and  a7735a );
 a689a <=( a7726a  and  a7717a );
 a690a <=( a7708a  and  a7699a );
 a691a <=( a7690a  and  a7681a );
 a692a <=( a7672a  and  a7663a );
 a693a <=( a7654a  and  a7645a );
 a694a <=( a7636a  and  a7627a );
 a695a <=( a7618a  and  a7609a );
 a696a <=( a7600a  and  a7591a );
 a697a <=( a7582a  and  a7573a );
 a698a <=( a7564a  and  a7555a );
 a699a <=( a7546a  and  a7537a );
 a700a <=( a7528a  and  a7519a );
 a701a <=( a7510a  and  a7501a );
 a702a <=( a7492a  and  a7483a );
 a703a <=( a7474a  and  a7465a );
 a704a <=( a7456a  and  a7447a );
 a705a <=( a7438a  and  a7429a );
 a706a <=( a7420a  and  a7411a );
 a707a <=( a7402a  and  a7393a );
 a708a <=( a7384a  and  a7375a );
 a709a <=( a7366a  and  a7357a );
 a710a <=( a7348a  and  a7339a );
 a711a <=( a7330a  and  a7321a );
 a712a <=( a7312a  and  a7303a );
 a713a <=( a7294a  and  a7285a );
 a714a <=( a7276a  and  a7267a );
 a715a <=( a7258a  and  a7249a );
 a716a <=( a7240a  and  a7231a );
 a717a <=( a7222a  and  a7213a );
 a718a <=( a7204a  and  a7195a );
 a719a <=( a7186a  and  a7177a );
 a720a <=( a7168a  and  a7159a );
 a721a <=( a7150a  and  a7141a );
 a722a <=( a7132a  and  a7123a );
 a723a <=( a7114a  and  a7105a );
 a724a <=( a7096a  and  a7087a );
 a725a <=( a7078a  and  a7069a );
 a726a <=( a7060a  and  a7051a );
 a727a <=( a7042a  and  a7033a );
 a728a <=( a7024a  and  a7015a );
 a729a <=( a7006a  and  a6997a );
 a730a <=( a6988a  and  a6979a );
 a731a <=( a6970a  and  a6961a );
 a732a <=( a6952a  and  a6943a );
 a733a <=( a6934a  and  a6925a );
 a734a <=( a6916a  and  a6907a );
 a735a <=( a6898a  and  a6889a );
 a736a <=( a6880a  and  a6871a );
 a737a <=( a6862a  and  a6853a );
 a738a <=( a6844a  and  a6835a );
 a739a <=( a6826a  and  a6817a );
 a740a <=( a6808a  and  a6799a );
 a741a <=( a6790a  and  a6781a );
 a742a <=( a6772a  and  a6763a );
 a743a <=( a6754a  and  a6745a );
 a744a <=( a6736a  and  a6727a );
 a745a <=( a6718a  and  a6709a );
 a746a <=( a6700a  and  a6691a );
 a747a <=( a6682a  and  a6673a );
 a748a <=( a6664a  and  a6655a );
 a749a <=( a6646a  and  a6637a );
 a750a <=( a6628a  and  a6619a );
 a751a <=( a6610a  and  a6601a );
 a752a <=( a6592a  and  a6583a );
 a753a <=( a6574a  and  a6565a );
 a754a <=( a6556a  and  a6547a );
 a755a <=( a6538a  and  a6529a );
 a756a <=( a6520a  and  a6511a );
 a757a <=( a6502a  and  a6493a );
 a758a <=( a6484a  and  a6475a );
 a759a <=( a6466a  and  a6457a );
 a760a <=( a6448a  and  a6439a );
 a761a <=( a6430a  and  a6421a );
 a762a <=( a6412a  and  a6403a );
 a763a <=( a6394a  and  a6385a );
 a764a <=( a6376a  and  a6367a );
 a765a <=( a6358a  and  a6349a );
 a766a <=( a6340a  and  a6331a );
 a767a <=( a6322a  and  a6313a );
 a768a <=( a6304a  and  a6295a );
 a769a <=( a6286a  and  a6277a );
 a770a <=( a6268a  and  a6259a );
 a771a <=( a6250a  and  a6241a );
 a772a <=( a6232a  and  a6223a );
 a773a <=( a6214a  and  a6205a );
 a774a <=( a6196a  and  a6187a );
 a775a <=( a6180a  and  a6171a );
 a776a <=( a6164a  and  a6155a );
 a777a <=( a6148a  and  a6139a );
 a778a <=( a6132a  and  a6123a );
 a779a <=( a6116a  and  a6107a );
 a780a <=( a6100a  and  a6091a );
 a781a <=( a6084a  and  a6075a );
 a782a <=( a6068a  and  a6059a );
 a783a <=( a6052a  and  a6043a );
 a784a <=( a6036a  and  a6027a );
 a785a <=( a6020a  and  a6011a );
 a786a <=( a6004a  and  a5995a );
 a787a <=( a5988a  and  a5979a );
 a788a <=( a5972a  and  a5963a );
 a789a <=( a5956a  and  a5947a );
 a790a <=( a5940a  and  a5931a );
 a791a <=( a5924a  and  a5915a );
 a792a <=( a5908a  and  a5899a );
 a793a <=( a5892a  and  a5883a );
 a794a <=( a5876a  and  a5867a );
 a795a <=( a5860a  and  a5851a );
 a796a <=( a5844a  and  a5835a );
 a797a <=( a5828a  and  a5819a );
 a798a <=( a5812a  and  a5803a );
 a799a <=( a5796a  and  a5787a );
 a800a <=( a5780a  and  a5771a );
 a801a <=( a5764a  and  a5755a );
 a802a <=( a5748a  and  a5739a );
 a803a <=( a5732a  and  a5723a );
 a804a <=( a5716a  and  a5707a );
 a805a <=( a5700a  and  a5691a );
 a806a <=( a5684a  and  a5675a );
 a807a <=( a5668a  and  a5659a );
 a808a <=( a5652a  and  a5643a );
 a809a <=( a5636a  and  a5627a );
 a810a <=( a5620a  and  a5611a );
 a811a <=( a5604a  and  a5595a );
 a812a <=( a5588a  and  a5579a );
 a813a <=( a5572a  and  a5563a );
 a814a <=( a5556a  and  a5547a );
 a815a <=( a5540a  and  a5531a );
 a816a <=( a5524a  and  a5515a );
 a817a <=( a5508a  and  a5499a );
 a818a <=( a5492a  and  a5483a );
 a819a <=( a5476a  and  a5467a );
 a820a <=( a5460a  and  a5451a );
 a821a <=( a5444a  and  a5435a );
 a822a <=( a5428a  and  a5419a );
 a823a <=( a5412a  and  a5403a );
 a824a <=( a5396a  and  a5387a );
 a825a <=( a5380a  and  a5371a );
 a826a <=( a5364a  and  a5355a );
 a827a <=( a5348a  and  a5339a );
 a828a <=( a5332a  and  a5323a );
 a829a <=( a5316a  and  a5307a );
 a830a <=( a5300a  and  a5291a );
 a831a <=( a5284a  and  a5275a );
 a832a <=( a5268a  and  a5259a );
 a833a <=( a5252a  and  a5243a );
 a834a <=( a5236a  and  a5227a );
 a835a <=( a5220a  and  a5211a );
 a836a <=( a5204a  and  a5195a );
 a837a <=( a5188a  and  a5179a );
 a838a <=( a5172a  and  a5163a );
 a839a <=( a5156a  and  a5147a );
 a840a <=( a5140a  and  a5131a );
 a841a <=( a5124a  and  a5115a );
 a842a <=( a5108a  and  a5099a );
 a843a <=( a5092a  and  a5083a );
 a844a <=( a5076a  and  a5067a );
 a845a <=( a5060a  and  a5051a );
 a846a <=( a5044a  and  a5035a );
 a847a <=( a5028a  and  a5019a );
 a848a <=( a5012a  and  a5003a );
 a849a <=( a4996a  and  a4987a );
 a850a <=( a4980a  and  a4971a );
 a851a <=( a4964a  and  a4955a );
 a852a <=( a4948a  and  a4939a );
 a853a <=( a4932a  and  a4923a );
 a854a <=( a4916a  and  a4907a );
 a855a <=( a4900a  and  a4891a );
 a856a <=( a4884a  and  a4875a );
 a857a <=( a4868a  and  a4859a );
 a858a <=( a4852a  and  a4843a );
 a859a <=( a4836a  and  a4827a );
 a860a <=( a4820a  and  a4811a );
 a861a <=( a4804a  and  a4795a );
 a862a <=( a4788a  and  a4779a );
 a863a <=( a4772a  and  a4763a );
 a864a <=( a4756a  and  a4747a );
 a865a <=( a4740a  and  a4731a );
 a866a <=( a4724a  and  a4715a );
 a867a <=( a4708a  and  a4699a );
 a868a <=( a4692a  and  a4683a );
 a869a <=( a4676a  and  a4667a );
 a870a <=( a4660a  and  a4651a );
 a871a <=( a4644a  and  a4635a );
 a872a <=( a4628a  and  a4619a );
 a873a <=( a4612a  and  a4603a );
 a874a <=( a4596a  and  a4587a );
 a875a <=( a4580a  and  a4571a );
 a876a <=( a4564a  and  a4555a );
 a877a <=( a4548a  and  a4539a );
 a878a <=( a4532a  and  a4523a );
 a879a <=( a4516a  and  a4507a );
 a880a <=( a4500a  and  a4491a );
 a881a <=( a4484a  and  a4475a );
 a882a <=( a4468a  and  a4459a );
 a883a <=( a4452a  and  a4443a );
 a884a <=( a4436a  and  a4427a );
 a885a <=( a4420a  and  a4411a );
 a886a <=( a4404a  and  a4395a );
 a887a <=( a4388a  and  a4379a );
 a888a <=( a4372a  and  a4363a );
 a889a <=( a4356a  and  a4347a );
 a890a <=( a4340a  and  a4331a );
 a891a <=( a4324a  and  a4315a );
 a892a <=( a4308a  and  a4299a );
 a893a <=( a4292a  and  a4283a );
 a894a <=( a4276a  and  a4267a );
 a895a <=( a4260a  and  a4251a );
 a896a <=( a4244a  and  a4237a );
 a897a <=( a4230a  and  a4223a );
 a898a <=( a4216a  and  a4209a );
 a899a <=( a4202a  and  a4195a );
 a900a <=( a4188a  and  a4181a );
 a901a <=( a4174a  and  a4167a );
 a902a <=( a4160a  and  a4153a );
 a903a <=( a4146a  and  a4139a );
 a904a <=( a4132a  and  a4125a );
 a905a <=( a4118a  and  a4111a );
 a906a <=( a4104a  and  a4097a );
 a907a <=( a4090a  and  a4083a );
 a908a <=( a4076a  and  a4069a );
 a909a <=( a4062a  and  a4055a );
 a910a <=( a4048a  and  a4041a );
 a911a <=( a4034a  and  a4027a );
 a912a <=( a4020a  and  a4013a );
 a913a <=( a4006a  and  a3999a );
 a914a <=( a3992a  and  a3985a );
 a915a <=( a3978a  and  a3971a );
 a916a <=( a3964a  and  a3957a );
 a917a <=( a3950a  and  a3943a );
 a918a <=( a3936a  and  a3929a );
 a919a <=( a3922a  and  a3915a );
 a920a <=( a3908a  and  a3901a );
 a921a <=( a3894a  and  a3887a );
 a922a <=( a3880a  and  a3873a );
 a923a <=( a3866a  and  a3859a );
 a924a <=( a3852a  and  a3845a );
 a925a <=( a3838a  and  a3831a );
 a926a <=( a3824a  and  a3817a );
 a927a <=( a3810a  and  a3803a );
 a928a <=( a3796a  and  a3789a );
 a929a <=( a3782a  and  a3775a );
 a930a <=( a3768a  and  a3761a );
 a931a <=( a3754a  and  a3747a );
 a932a <=( a3740a  and  a3733a );
 a933a <=( a3726a  and  a3719a );
 a934a <=( a3712a  and  a3705a );
 a935a <=( a3698a  and  a3691a );
 a936a <=( a3684a  and  a3677a );
 a937a <=( a3670a  and  a3663a );
 a938a <=( a3656a  and  a3649a );
 a939a <=( a3642a  and  a3635a );
 a940a <=( a3628a  and  a3621a );
 a941a <=( a3614a  and  a3607a );
 a942a <=( a3600a  and  a3593a );
 a943a <=( a3586a  and  a3579a );
 a944a <=( a3572a  and  a3565a );
 a945a <=( a3558a  and  a3551a );
 a946a <=( a3544a  and  a3537a );
 a947a <=( a3532a  and  a3525a );
 a948a <=( a3520a  and  a3513a );
 a949a <=( a3508a  and  a3501a );
 a950a <=( a3496a  and  a3489a );
 a951a <=( a3484a  and  a3477a );
 a952a <=( a3472a  and  a3465a );
 a953a <=( a3460a  and  a3453a );
 a954a <=( a3448a  and  a3441a );
 a955a <=( a3436a  and  a3429a );
 a956a <=( a3424a  and  a3417a );
 a957a <=( a3412a  and  a3405a );
 a958a <=( a3400a  and  a3393a );
 a959a <=( a3388a  and  a3383a );
 a960a <=( a3378a  and  a3373a );
 a961a <=( a3368a  and  a3363a );
 a962a <=( a3358a  and  a3353a );
 a963a <=( a3348a  and  a3343a );
 a964a <=( a3338a  and  a3333a );
 a965a <=( a3328a  and  a3323a );
 a966a <=( a3318a  and  a3313a );
 a967a <=( a3308a  and  a3303a );
 a968a <=( a3298a  and  a3293a );
 a969a <=( a3288a  and  a3283a );
 a970a <=( a3280a  and  a3275a );
 a971a <=( a3272a  and  a3267a );
 a972a <=( a3264a  and  a3259a );
 a973a <=( a3256a  and  a3251a );
 a974a <=( a3248a  and  a3243a );
 a975a <=( a3240a  and  a3235a );
 a976a <=( a3232a  and  a3227a );
 a977a <=( a3224a  and  a3219a );
 a978a <=( a3216a  and  a3211a );
 a979a <=( a3208a  and  a3203a );
 a980a <=( a3200a  and  a3195a );
 a981a <=( a3192a  and  a3187a );
 a982a <=( a3184a  and  a3179a );
 a983a <=( a3176a  and  a3171a );
 a984a <=( a3168a  and  a3163a );
 a985a <=( a3160a  and  a3157a );
 a986a <=( a3154a  and  a3151a );
 a987a <=( a3148a  and  a3145a );
 a988a <=( a3142a  and  a3139a );
 a989a <=( a3136a  and  a3133a );
 a990a <=( a3130a  and  a3127a );
 a991a <=( a3124a  and  a3121a );
 a992a <=( a3118a  and  a3115a );
 a993a <=( a3112a  and  a3109a );
 a994a <=( a3106a  and  a3103a );
 a995a <=( a3100a  and  a3097a );
 a996a <=( a3094a  and  a3091a );
 a997a <=( a3088a  and  a3085a );
 a998a <=( a3082a  and  a3079a );
 a999a <=( a3076a  and  a3073a );
 a1000a <=( a3070a  and  a3067a );
 a1001a <=( A169  and  a3064a );
 a1002a <=( A169  and  a3060a );
 a1003a <=( A168  and  a3056a );
 a1004a <=( A168  and  a3052a );
 a1005a <=( A200  and  a3048a );
 a1006a <=( A199  and  a3044a );
 a1007a <=( A202  and  a3040a );
 a1008a <=( A202  and  a3036a );
 a1009a <=( A235  and  A169 );
 a1010a <=( A235  and  A202 );
 a1014a <=( a1008a ) or ( a1009a );
 a1015a <=( a1010a ) or ( a1014a );
 a1018a <=( a1006a ) or ( a1007a );
 a1021a <=( a1004a ) or ( a1005a );
 a1022a <=( a1021a ) or ( a1018a );
 a1023a <=( a1022a ) or ( a1015a );
 a1026a <=( a1002a ) or ( a1003a );
 a1029a <=( a1000a ) or ( a1001a );
 a1030a <=( a1029a ) or ( a1026a );
 a1033a <=( a998a ) or ( a999a );
 a1036a <=( a996a ) or ( a997a );
 a1037a <=( a1036a ) or ( a1033a );
 a1038a <=( a1037a ) or ( a1030a );
 a1039a <=( a1038a ) or ( a1023a );
 a1042a <=( a994a ) or ( a995a );
 a1045a <=( a992a ) or ( a993a );
 a1046a <=( a1045a ) or ( a1042a );
 a1049a <=( a990a ) or ( a991a );
 a1052a <=( a988a ) or ( a989a );
 a1053a <=( a1052a ) or ( a1049a );
 a1054a <=( a1053a ) or ( a1046a );
 a1057a <=( a986a ) or ( a987a );
 a1060a <=( a984a ) or ( a985a );
 a1061a <=( a1060a ) or ( a1057a );
 a1064a <=( a982a ) or ( a983a );
 a1067a <=( a980a ) or ( a981a );
 a1068a <=( a1067a ) or ( a1064a );
 a1069a <=( a1068a ) or ( a1061a );
 a1070a <=( a1069a ) or ( a1054a );
 a1071a <=( a1070a ) or ( a1039a );
 a1074a <=( a978a ) or ( a979a );
 a1077a <=( a976a ) or ( a977a );
 a1078a <=( a1077a ) or ( a1074a );
 a1081a <=( a974a ) or ( a975a );
 a1084a <=( a972a ) or ( a973a );
 a1085a <=( a1084a ) or ( a1081a );
 a1086a <=( a1085a ) or ( a1078a );
 a1089a <=( a970a ) or ( a971a );
 a1092a <=( a968a ) or ( a969a );
 a1093a <=( a1092a ) or ( a1089a );
 a1096a <=( a966a ) or ( a967a );
 a1099a <=( a964a ) or ( a965a );
 a1100a <=( a1099a ) or ( a1096a );
 a1101a <=( a1100a ) or ( a1093a );
 a1102a <=( a1101a ) or ( a1086a );
 a1105a <=( a962a ) or ( a963a );
 a1108a <=( a960a ) or ( a961a );
 a1109a <=( a1108a ) or ( a1105a );
 a1112a <=( a958a ) or ( a959a );
 a1115a <=( a956a ) or ( a957a );
 a1116a <=( a1115a ) or ( a1112a );
 a1117a <=( a1116a ) or ( a1109a );
 a1120a <=( a954a ) or ( a955a );
 a1123a <=( a952a ) or ( a953a );
 a1124a <=( a1123a ) or ( a1120a );
 a1127a <=( a950a ) or ( a951a );
 a1130a <=( a948a ) or ( a949a );
 a1131a <=( a1130a ) or ( a1127a );
 a1132a <=( a1131a ) or ( a1124a );
 a1133a <=( a1132a ) or ( a1117a );
 a1134a <=( a1133a ) or ( a1102a );
 a1135a <=( a1134a ) or ( a1071a );
 a1139a <=( a945a ) or ( a946a );
 a1140a <=( a947a ) or ( a1139a );
 a1143a <=( a943a ) or ( a944a );
 a1146a <=( a941a ) or ( a942a );
 a1147a <=( a1146a ) or ( a1143a );
 a1148a <=( a1147a ) or ( a1140a );
 a1151a <=( a939a ) or ( a940a );
 a1154a <=( a937a ) or ( a938a );
 a1155a <=( a1154a ) or ( a1151a );
 a1158a <=( a935a ) or ( a936a );
 a1161a <=( a933a ) or ( a934a );
 a1162a <=( a1161a ) or ( a1158a );
 a1163a <=( a1162a ) or ( a1155a );
 a1164a <=( a1163a ) or ( a1148a );
 a1167a <=( a931a ) or ( a932a );
 a1170a <=( a929a ) or ( a930a );
 a1171a <=( a1170a ) or ( a1167a );
 a1174a <=( a927a ) or ( a928a );
 a1177a <=( a925a ) or ( a926a );
 a1178a <=( a1177a ) or ( a1174a );
 a1179a <=( a1178a ) or ( a1171a );
 a1182a <=( a923a ) or ( a924a );
 a1185a <=( a921a ) or ( a922a );
 a1186a <=( a1185a ) or ( a1182a );
 a1189a <=( a919a ) or ( a920a );
 a1192a <=( a917a ) or ( a918a );
 a1193a <=( a1192a ) or ( a1189a );
 a1194a <=( a1193a ) or ( a1186a );
 a1195a <=( a1194a ) or ( a1179a );
 a1196a <=( a1195a ) or ( a1164a );
 a1199a <=( a915a ) or ( a916a );
 a1202a <=( a913a ) or ( a914a );
 a1203a <=( a1202a ) or ( a1199a );
 a1206a <=( a911a ) or ( a912a );
 a1209a <=( a909a ) or ( a910a );
 a1210a <=( a1209a ) or ( a1206a );
 a1211a <=( a1210a ) or ( a1203a );
 a1214a <=( a907a ) or ( a908a );
 a1217a <=( a905a ) or ( a906a );
 a1218a <=( a1217a ) or ( a1214a );
 a1221a <=( a903a ) or ( a904a );
 a1224a <=( a901a ) or ( a902a );
 a1225a <=( a1224a ) or ( a1221a );
 a1226a <=( a1225a ) or ( a1218a );
 a1227a <=( a1226a ) or ( a1211a );
 a1230a <=( a899a ) or ( a900a );
 a1233a <=( a897a ) or ( a898a );
 a1234a <=( a1233a ) or ( a1230a );
 a1237a <=( a895a ) or ( a896a );
 a1240a <=( a893a ) or ( a894a );
 a1241a <=( a1240a ) or ( a1237a );
 a1242a <=( a1241a ) or ( a1234a );
 a1245a <=( a891a ) or ( a892a );
 a1248a <=( a889a ) or ( a890a );
 a1249a <=( a1248a ) or ( a1245a );
 a1252a <=( a887a ) or ( a888a );
 a1255a <=( a885a ) or ( a886a );
 a1256a <=( a1255a ) or ( a1252a );
 a1257a <=( a1256a ) or ( a1249a );
 a1258a <=( a1257a ) or ( a1242a );
 a1259a <=( a1258a ) or ( a1227a );
 a1260a <=( a1259a ) or ( a1196a );
 a1261a <=( a1260a ) or ( a1135a );
 a1265a <=( a882a ) or ( a883a );
 a1266a <=( a884a ) or ( a1265a );
 a1269a <=( a880a ) or ( a881a );
 a1272a <=( a878a ) or ( a879a );
 a1273a <=( a1272a ) or ( a1269a );
 a1274a <=( a1273a ) or ( a1266a );
 a1277a <=( a876a ) or ( a877a );
 a1280a <=( a874a ) or ( a875a );
 a1281a <=( a1280a ) or ( a1277a );
 a1284a <=( a872a ) or ( a873a );
 a1287a <=( a870a ) or ( a871a );
 a1288a <=( a1287a ) or ( a1284a );
 a1289a <=( a1288a ) or ( a1281a );
 a1290a <=( a1289a ) or ( a1274a );
 a1293a <=( a868a ) or ( a869a );
 a1296a <=( a866a ) or ( a867a );
 a1297a <=( a1296a ) or ( a1293a );
 a1300a <=( a864a ) or ( a865a );
 a1303a <=( a862a ) or ( a863a );
 a1304a <=( a1303a ) or ( a1300a );
 a1305a <=( a1304a ) or ( a1297a );
 a1308a <=( a860a ) or ( a861a );
 a1311a <=( a858a ) or ( a859a );
 a1312a <=( a1311a ) or ( a1308a );
 a1315a <=( a856a ) or ( a857a );
 a1318a <=( a854a ) or ( a855a );
 a1319a <=( a1318a ) or ( a1315a );
 a1320a <=( a1319a ) or ( a1312a );
 a1321a <=( a1320a ) or ( a1305a );
 a1322a <=( a1321a ) or ( a1290a );
 a1325a <=( a852a ) or ( a853a );
 a1328a <=( a850a ) or ( a851a );
 a1329a <=( a1328a ) or ( a1325a );
 a1332a <=( a848a ) or ( a849a );
 a1335a <=( a846a ) or ( a847a );
 a1336a <=( a1335a ) or ( a1332a );
 a1337a <=( a1336a ) or ( a1329a );
 a1340a <=( a844a ) or ( a845a );
 a1343a <=( a842a ) or ( a843a );
 a1344a <=( a1343a ) or ( a1340a );
 a1347a <=( a840a ) or ( a841a );
 a1350a <=( a838a ) or ( a839a );
 a1351a <=( a1350a ) or ( a1347a );
 a1352a <=( a1351a ) or ( a1344a );
 a1353a <=( a1352a ) or ( a1337a );
 a1356a <=( a836a ) or ( a837a );
 a1359a <=( a834a ) or ( a835a );
 a1360a <=( a1359a ) or ( a1356a );
 a1363a <=( a832a ) or ( a833a );
 a1366a <=( a830a ) or ( a831a );
 a1367a <=( a1366a ) or ( a1363a );
 a1368a <=( a1367a ) or ( a1360a );
 a1371a <=( a828a ) or ( a829a );
 a1374a <=( a826a ) or ( a827a );
 a1375a <=( a1374a ) or ( a1371a );
 a1378a <=( a824a ) or ( a825a );
 a1381a <=( a822a ) or ( a823a );
 a1382a <=( a1381a ) or ( a1378a );
 a1383a <=( a1382a ) or ( a1375a );
 a1384a <=( a1383a ) or ( a1368a );
 a1385a <=( a1384a ) or ( a1353a );
 a1386a <=( a1385a ) or ( a1322a );
 a1390a <=( a819a ) or ( a820a );
 a1391a <=( a821a ) or ( a1390a );
 a1394a <=( a817a ) or ( a818a );
 a1397a <=( a815a ) or ( a816a );
 a1398a <=( a1397a ) or ( a1394a );
 a1399a <=( a1398a ) or ( a1391a );
 a1402a <=( a813a ) or ( a814a );
 a1405a <=( a811a ) or ( a812a );
 a1406a <=( a1405a ) or ( a1402a );
 a1409a <=( a809a ) or ( a810a );
 a1412a <=( a807a ) or ( a808a );
 a1413a <=( a1412a ) or ( a1409a );
 a1414a <=( a1413a ) or ( a1406a );
 a1415a <=( a1414a ) or ( a1399a );
 a1418a <=( a805a ) or ( a806a );
 a1421a <=( a803a ) or ( a804a );
 a1422a <=( a1421a ) or ( a1418a );
 a1425a <=( a801a ) or ( a802a );
 a1428a <=( a799a ) or ( a800a );
 a1429a <=( a1428a ) or ( a1425a );
 a1430a <=( a1429a ) or ( a1422a );
 a1433a <=( a797a ) or ( a798a );
 a1436a <=( a795a ) or ( a796a );
 a1437a <=( a1436a ) or ( a1433a );
 a1440a <=( a793a ) or ( a794a );
 a1443a <=( a791a ) or ( a792a );
 a1444a <=( a1443a ) or ( a1440a );
 a1445a <=( a1444a ) or ( a1437a );
 a1446a <=( a1445a ) or ( a1430a );
 a1447a <=( a1446a ) or ( a1415a );
 a1450a <=( a789a ) or ( a790a );
 a1453a <=( a787a ) or ( a788a );
 a1454a <=( a1453a ) or ( a1450a );
 a1457a <=( a785a ) or ( a786a );
 a1460a <=( a783a ) or ( a784a );
 a1461a <=( a1460a ) or ( a1457a );
 a1462a <=( a1461a ) or ( a1454a );
 a1465a <=( a781a ) or ( a782a );
 a1468a <=( a779a ) or ( a780a );
 a1469a <=( a1468a ) or ( a1465a );
 a1472a <=( a777a ) or ( a778a );
 a1475a <=( a775a ) or ( a776a );
 a1476a <=( a1475a ) or ( a1472a );
 a1477a <=( a1476a ) or ( a1469a );
 a1478a <=( a1477a ) or ( a1462a );
 a1481a <=( a773a ) or ( a774a );
 a1484a <=( a771a ) or ( a772a );
 a1485a <=( a1484a ) or ( a1481a );
 a1488a <=( a769a ) or ( a770a );
 a1491a <=( a767a ) or ( a768a );
 a1492a <=( a1491a ) or ( a1488a );
 a1493a <=( a1492a ) or ( a1485a );
 a1496a <=( a765a ) or ( a766a );
 a1499a <=( a763a ) or ( a764a );
 a1500a <=( a1499a ) or ( a1496a );
 a1503a <=( a761a ) or ( a762a );
 a1506a <=( a759a ) or ( a760a );
 a1507a <=( a1506a ) or ( a1503a );
 a1508a <=( a1507a ) or ( a1500a );
 a1509a <=( a1508a ) or ( a1493a );
 a1510a <=( a1509a ) or ( a1478a );
 a1511a <=( a1510a ) or ( a1447a );
 a1512a <=( a1511a ) or ( a1386a );
 a1513a <=( a1512a ) or ( a1261a );
 a1517a <=( a756a ) or ( a757a );
 a1518a <=( a758a ) or ( a1517a );
 a1521a <=( a754a ) or ( a755a );
 a1524a <=( a752a ) or ( a753a );
 a1525a <=( a1524a ) or ( a1521a );
 a1526a <=( a1525a ) or ( a1518a );
 a1529a <=( a750a ) or ( a751a );
 a1532a <=( a748a ) or ( a749a );
 a1533a <=( a1532a ) or ( a1529a );
 a1536a <=( a746a ) or ( a747a );
 a1539a <=( a744a ) or ( a745a );
 a1540a <=( a1539a ) or ( a1536a );
 a1541a <=( a1540a ) or ( a1533a );
 a1542a <=( a1541a ) or ( a1526a );
 a1545a <=( a742a ) or ( a743a );
 a1548a <=( a740a ) or ( a741a );
 a1549a <=( a1548a ) or ( a1545a );
 a1552a <=( a738a ) or ( a739a );
 a1555a <=( a736a ) or ( a737a );
 a1556a <=( a1555a ) or ( a1552a );
 a1557a <=( a1556a ) or ( a1549a );
 a1560a <=( a734a ) or ( a735a );
 a1563a <=( a732a ) or ( a733a );
 a1564a <=( a1563a ) or ( a1560a );
 a1567a <=( a730a ) or ( a731a );
 a1570a <=( a728a ) or ( a729a );
 a1571a <=( a1570a ) or ( a1567a );
 a1572a <=( a1571a ) or ( a1564a );
 a1573a <=( a1572a ) or ( a1557a );
 a1574a <=( a1573a ) or ( a1542a );
 a1577a <=( a726a ) or ( a727a );
 a1580a <=( a724a ) or ( a725a );
 a1581a <=( a1580a ) or ( a1577a );
 a1584a <=( a722a ) or ( a723a );
 a1587a <=( a720a ) or ( a721a );
 a1588a <=( a1587a ) or ( a1584a );
 a1589a <=( a1588a ) or ( a1581a );
 a1592a <=( a718a ) or ( a719a );
 a1595a <=( a716a ) or ( a717a );
 a1596a <=( a1595a ) or ( a1592a );
 a1599a <=( a714a ) or ( a715a );
 a1602a <=( a712a ) or ( a713a );
 a1603a <=( a1602a ) or ( a1599a );
 a1604a <=( a1603a ) or ( a1596a );
 a1605a <=( a1604a ) or ( a1589a );
 a1608a <=( a710a ) or ( a711a );
 a1611a <=( a708a ) or ( a709a );
 a1612a <=( a1611a ) or ( a1608a );
 a1615a <=( a706a ) or ( a707a );
 a1618a <=( a704a ) or ( a705a );
 a1619a <=( a1618a ) or ( a1615a );
 a1620a <=( a1619a ) or ( a1612a );
 a1623a <=( a702a ) or ( a703a );
 a1626a <=( a700a ) or ( a701a );
 a1627a <=( a1626a ) or ( a1623a );
 a1630a <=( a698a ) or ( a699a );
 a1633a <=( a696a ) or ( a697a );
 a1634a <=( a1633a ) or ( a1630a );
 a1635a <=( a1634a ) or ( a1627a );
 a1636a <=( a1635a ) or ( a1620a );
 a1637a <=( a1636a ) or ( a1605a );
 a1638a <=( a1637a ) or ( a1574a );
 a1642a <=( a693a ) or ( a694a );
 a1643a <=( a695a ) or ( a1642a );
 a1646a <=( a691a ) or ( a692a );
 a1649a <=( a689a ) or ( a690a );
 a1650a <=( a1649a ) or ( a1646a );
 a1651a <=( a1650a ) or ( a1643a );
 a1654a <=( a687a ) or ( a688a );
 a1657a <=( a685a ) or ( a686a );
 a1658a <=( a1657a ) or ( a1654a );
 a1661a <=( a683a ) or ( a684a );
 a1664a <=( a681a ) or ( a682a );
 a1665a <=( a1664a ) or ( a1661a );
 a1666a <=( a1665a ) or ( a1658a );
 a1667a <=( a1666a ) or ( a1651a );
 a1670a <=( a679a ) or ( a680a );
 a1673a <=( a677a ) or ( a678a );
 a1674a <=( a1673a ) or ( a1670a );
 a1677a <=( a675a ) or ( a676a );
 a1680a <=( a673a ) or ( a674a );
 a1681a <=( a1680a ) or ( a1677a );
 a1682a <=( a1681a ) or ( a1674a );
 a1685a <=( a671a ) or ( a672a );
 a1688a <=( a669a ) or ( a670a );
 a1689a <=( a1688a ) or ( a1685a );
 a1692a <=( a667a ) or ( a668a );
 a1695a <=( a665a ) or ( a666a );
 a1696a <=( a1695a ) or ( a1692a );
 a1697a <=( a1696a ) or ( a1689a );
 a1698a <=( a1697a ) or ( a1682a );
 a1699a <=( a1698a ) or ( a1667a );
 a1702a <=( a663a ) or ( a664a );
 a1705a <=( a661a ) or ( a662a );
 a1706a <=( a1705a ) or ( a1702a );
 a1709a <=( a659a ) or ( a660a );
 a1712a <=( a657a ) or ( a658a );
 a1713a <=( a1712a ) or ( a1709a );
 a1714a <=( a1713a ) or ( a1706a );
 a1717a <=( a655a ) or ( a656a );
 a1720a <=( a653a ) or ( a654a );
 a1721a <=( a1720a ) or ( a1717a );
 a1724a <=( a651a ) or ( a652a );
 a1727a <=( a649a ) or ( a650a );
 a1728a <=( a1727a ) or ( a1724a );
 a1729a <=( a1728a ) or ( a1721a );
 a1730a <=( a1729a ) or ( a1714a );
 a1733a <=( a647a ) or ( a648a );
 a1736a <=( a645a ) or ( a646a );
 a1737a <=( a1736a ) or ( a1733a );
 a1740a <=( a643a ) or ( a644a );
 a1743a <=( a641a ) or ( a642a );
 a1744a <=( a1743a ) or ( a1740a );
 a1745a <=( a1744a ) or ( a1737a );
 a1748a <=( a639a ) or ( a640a );
 a1751a <=( a637a ) or ( a638a );
 a1752a <=( a1751a ) or ( a1748a );
 a1755a <=( a635a ) or ( a636a );
 a1758a <=( a633a ) or ( a634a );
 a1759a <=( a1758a ) or ( a1755a );
 a1760a <=( a1759a ) or ( a1752a );
 a1761a <=( a1760a ) or ( a1745a );
 a1762a <=( a1761a ) or ( a1730a );
 a1763a <=( a1762a ) or ( a1699a );
 a1764a <=( a1763a ) or ( a1638a );
 a1768a <=( a630a ) or ( a631a );
 a1769a <=( a632a ) or ( a1768a );
 a1772a <=( a628a ) or ( a629a );
 a1775a <=( a626a ) or ( a627a );
 a1776a <=( a1775a ) or ( a1772a );
 a1777a <=( a1776a ) or ( a1769a );
 a1780a <=( a624a ) or ( a625a );
 a1783a <=( a622a ) or ( a623a );
 a1784a <=( a1783a ) or ( a1780a );
 a1787a <=( a620a ) or ( a621a );
 a1790a <=( a618a ) or ( a619a );
 a1791a <=( a1790a ) or ( a1787a );
 a1792a <=( a1791a ) or ( a1784a );
 a1793a <=( a1792a ) or ( a1777a );
 a1796a <=( a616a ) or ( a617a );
 a1799a <=( a614a ) or ( a615a );
 a1800a <=( a1799a ) or ( a1796a );
 a1803a <=( a612a ) or ( a613a );
 a1806a <=( a610a ) or ( a611a );
 a1807a <=( a1806a ) or ( a1803a );
 a1808a <=( a1807a ) or ( a1800a );
 a1811a <=( a608a ) or ( a609a );
 a1814a <=( a606a ) or ( a607a );
 a1815a <=( a1814a ) or ( a1811a );
 a1818a <=( a604a ) or ( a605a );
 a1821a <=( a602a ) or ( a603a );
 a1822a <=( a1821a ) or ( a1818a );
 a1823a <=( a1822a ) or ( a1815a );
 a1824a <=( a1823a ) or ( a1808a );
 a1825a <=( a1824a ) or ( a1793a );
 a1828a <=( a600a ) or ( a601a );
 a1831a <=( a598a ) or ( a599a );
 a1832a <=( a1831a ) or ( a1828a );
 a1835a <=( a596a ) or ( a597a );
 a1838a <=( a594a ) or ( a595a );
 a1839a <=( a1838a ) or ( a1835a );
 a1840a <=( a1839a ) or ( a1832a );
 a1843a <=( a592a ) or ( a593a );
 a1846a <=( a590a ) or ( a591a );
 a1847a <=( a1846a ) or ( a1843a );
 a1850a <=( a588a ) or ( a589a );
 a1853a <=( a586a ) or ( a587a );
 a1854a <=( a1853a ) or ( a1850a );
 a1855a <=( a1854a ) or ( a1847a );
 a1856a <=( a1855a ) or ( a1840a );
 a1859a <=( a584a ) or ( a585a );
 a1862a <=( a582a ) or ( a583a );
 a1863a <=( a1862a ) or ( a1859a );
 a1866a <=( a580a ) or ( a581a );
 a1869a <=( a578a ) or ( a579a );
 a1870a <=( a1869a ) or ( a1866a );
 a1871a <=( a1870a ) or ( a1863a );
 a1874a <=( a576a ) or ( a577a );
 a1877a <=( a574a ) or ( a575a );
 a1878a <=( a1877a ) or ( a1874a );
 a1881a <=( a572a ) or ( a573a );
 a1884a <=( a570a ) or ( a571a );
 a1885a <=( a1884a ) or ( a1881a );
 a1886a <=( a1885a ) or ( a1878a );
 a1887a <=( a1886a ) or ( a1871a );
 a1888a <=( a1887a ) or ( a1856a );
 a1889a <=( a1888a ) or ( a1825a );
 a1892a <=( a568a ) or ( a569a );
 a1895a <=( a566a ) or ( a567a );
 a1896a <=( a1895a ) or ( a1892a );
 a1899a <=( a564a ) or ( a565a );
 a1902a <=( a562a ) or ( a563a );
 a1903a <=( a1902a ) or ( a1899a );
 a1904a <=( a1903a ) or ( a1896a );
 a1907a <=( a560a ) or ( a561a );
 a1910a <=( a558a ) or ( a559a );
 a1911a <=( a1910a ) or ( a1907a );
 a1914a <=( a556a ) or ( a557a );
 a1917a <=( a554a ) or ( a555a );
 a1918a <=( a1917a ) or ( a1914a );
 a1919a <=( a1918a ) or ( a1911a );
 a1920a <=( a1919a ) or ( a1904a );
 a1923a <=( a552a ) or ( a553a );
 a1926a <=( a550a ) or ( a551a );
 a1927a <=( a1926a ) or ( a1923a );
 a1930a <=( a548a ) or ( a549a );
 a1933a <=( a546a ) or ( a547a );
 a1934a <=( a1933a ) or ( a1930a );
 a1935a <=( a1934a ) or ( a1927a );
 a1938a <=( a544a ) or ( a545a );
 a1941a <=( a542a ) or ( a543a );
 a1942a <=( a1941a ) or ( a1938a );
 a1945a <=( a540a ) or ( a541a );
 a1948a <=( a538a ) or ( a539a );
 a1949a <=( a1948a ) or ( a1945a );
 a1950a <=( a1949a ) or ( a1942a );
 a1951a <=( a1950a ) or ( a1935a );
 a1952a <=( a1951a ) or ( a1920a );
 a1955a <=( a536a ) or ( a537a );
 a1958a <=( a534a ) or ( a535a );
 a1959a <=( a1958a ) or ( a1955a );
 a1962a <=( a532a ) or ( a533a );
 a1965a <=( a530a ) or ( a531a );
 a1966a <=( a1965a ) or ( a1962a );
 a1967a <=( a1966a ) or ( a1959a );
 a1970a <=( a528a ) or ( a529a );
 a1973a <=( a526a ) or ( a527a );
 a1974a <=( a1973a ) or ( a1970a );
 a1977a <=( a524a ) or ( a525a );
 a1980a <=( a522a ) or ( a523a );
 a1981a <=( a1980a ) or ( a1977a );
 a1982a <=( a1981a ) or ( a1974a );
 a1983a <=( a1982a ) or ( a1967a );
 a1986a <=( a520a ) or ( a521a );
 a1989a <=( a518a ) or ( a519a );
 a1990a <=( a1989a ) or ( a1986a );
 a1993a <=( a516a ) or ( a517a );
 a1996a <=( a514a ) or ( a515a );
 a1997a <=( a1996a ) or ( a1993a );
 a1998a <=( a1997a ) or ( a1990a );
 a2001a <=( a512a ) or ( a513a );
 a2004a <=( a510a ) or ( a511a );
 a2005a <=( a2004a ) or ( a2001a );
 a2008a <=( a508a ) or ( a509a );
 a2011a <=( a506a ) or ( a507a );
 a2012a <=( a2011a ) or ( a2008a );
 a2013a <=( a2012a ) or ( a2005a );
 a2014a <=( a2013a ) or ( a1998a );
 a2015a <=( a2014a ) or ( a1983a );
 a2016a <=( a2015a ) or ( a1952a );
 a2017a <=( a2016a ) or ( a1889a );
 a2018a <=( a2017a ) or ( a1764a );
 a2019a <=( a2018a ) or ( a1513a );
 a2023a <=( a503a ) or ( a504a );
 a2024a <=( a505a ) or ( a2023a );
 a2027a <=( a501a ) or ( a502a );
 a2030a <=( a499a ) or ( a500a );
 a2031a <=( a2030a ) or ( a2027a );
 a2032a <=( a2031a ) or ( a2024a );
 a2035a <=( a497a ) or ( a498a );
 a2038a <=( a495a ) or ( a496a );
 a2039a <=( a2038a ) or ( a2035a );
 a2042a <=( a493a ) or ( a494a );
 a2045a <=( a491a ) or ( a492a );
 a2046a <=( a2045a ) or ( a2042a );
 a2047a <=( a2046a ) or ( a2039a );
 a2048a <=( a2047a ) or ( a2032a );
 a2051a <=( a489a ) or ( a490a );
 a2054a <=( a487a ) or ( a488a );
 a2055a <=( a2054a ) or ( a2051a );
 a2058a <=( a485a ) or ( a486a );
 a2061a <=( a483a ) or ( a484a );
 a2062a <=( a2061a ) or ( a2058a );
 a2063a <=( a2062a ) or ( a2055a );
 a2066a <=( a481a ) or ( a482a );
 a2069a <=( a479a ) or ( a480a );
 a2070a <=( a2069a ) or ( a2066a );
 a2073a <=( a477a ) or ( a478a );
 a2076a <=( a475a ) or ( a476a );
 a2077a <=( a2076a ) or ( a2073a );
 a2078a <=( a2077a ) or ( a2070a );
 a2079a <=( a2078a ) or ( a2063a );
 a2080a <=( a2079a ) or ( a2048a );
 a2083a <=( a473a ) or ( a474a );
 a2086a <=( a471a ) or ( a472a );
 a2087a <=( a2086a ) or ( a2083a );
 a2090a <=( a469a ) or ( a470a );
 a2093a <=( a467a ) or ( a468a );
 a2094a <=( a2093a ) or ( a2090a );
 a2095a <=( a2094a ) or ( a2087a );
 a2098a <=( a465a ) or ( a466a );
 a2101a <=( a463a ) or ( a464a );
 a2102a <=( a2101a ) or ( a2098a );
 a2105a <=( a461a ) or ( a462a );
 a2108a <=( a459a ) or ( a460a );
 a2109a <=( a2108a ) or ( a2105a );
 a2110a <=( a2109a ) or ( a2102a );
 a2111a <=( a2110a ) or ( a2095a );
 a2114a <=( a457a ) or ( a458a );
 a2117a <=( a455a ) or ( a456a );
 a2118a <=( a2117a ) or ( a2114a );
 a2121a <=( a453a ) or ( a454a );
 a2124a <=( a451a ) or ( a452a );
 a2125a <=( a2124a ) or ( a2121a );
 a2126a <=( a2125a ) or ( a2118a );
 a2129a <=( a449a ) or ( a450a );
 a2132a <=( a447a ) or ( a448a );
 a2133a <=( a2132a ) or ( a2129a );
 a2136a <=( a445a ) or ( a446a );
 a2139a <=( a443a ) or ( a444a );
 a2140a <=( a2139a ) or ( a2136a );
 a2141a <=( a2140a ) or ( a2133a );
 a2142a <=( a2141a ) or ( a2126a );
 a2143a <=( a2142a ) or ( a2111a );
 a2144a <=( a2143a ) or ( a2080a );
 a2148a <=( a440a ) or ( a441a );
 a2149a <=( a442a ) or ( a2148a );
 a2152a <=( a438a ) or ( a439a );
 a2155a <=( a436a ) or ( a437a );
 a2156a <=( a2155a ) or ( a2152a );
 a2157a <=( a2156a ) or ( a2149a );
 a2160a <=( a434a ) or ( a435a );
 a2163a <=( a432a ) or ( a433a );
 a2164a <=( a2163a ) or ( a2160a );
 a2167a <=( a430a ) or ( a431a );
 a2170a <=( a428a ) or ( a429a );
 a2171a <=( a2170a ) or ( a2167a );
 a2172a <=( a2171a ) or ( a2164a );
 a2173a <=( a2172a ) or ( a2157a );
 a2176a <=( a426a ) or ( a427a );
 a2179a <=( a424a ) or ( a425a );
 a2180a <=( a2179a ) or ( a2176a );
 a2183a <=( a422a ) or ( a423a );
 a2186a <=( a420a ) or ( a421a );
 a2187a <=( a2186a ) or ( a2183a );
 a2188a <=( a2187a ) or ( a2180a );
 a2191a <=( a418a ) or ( a419a );
 a2194a <=( a416a ) or ( a417a );
 a2195a <=( a2194a ) or ( a2191a );
 a2198a <=( a414a ) or ( a415a );
 a2201a <=( a412a ) or ( a413a );
 a2202a <=( a2201a ) or ( a2198a );
 a2203a <=( a2202a ) or ( a2195a );
 a2204a <=( a2203a ) or ( a2188a );
 a2205a <=( a2204a ) or ( a2173a );
 a2208a <=( a410a ) or ( a411a );
 a2211a <=( a408a ) or ( a409a );
 a2212a <=( a2211a ) or ( a2208a );
 a2215a <=( a406a ) or ( a407a );
 a2218a <=( a404a ) or ( a405a );
 a2219a <=( a2218a ) or ( a2215a );
 a2220a <=( a2219a ) or ( a2212a );
 a2223a <=( a402a ) or ( a403a );
 a2226a <=( a400a ) or ( a401a );
 a2227a <=( a2226a ) or ( a2223a );
 a2230a <=( a398a ) or ( a399a );
 a2233a <=( a396a ) or ( a397a );
 a2234a <=( a2233a ) or ( a2230a );
 a2235a <=( a2234a ) or ( a2227a );
 a2236a <=( a2235a ) or ( a2220a );
 a2239a <=( a394a ) or ( a395a );
 a2242a <=( a392a ) or ( a393a );
 a2243a <=( a2242a ) or ( a2239a );
 a2246a <=( a390a ) or ( a391a );
 a2249a <=( a388a ) or ( a389a );
 a2250a <=( a2249a ) or ( a2246a );
 a2251a <=( a2250a ) or ( a2243a );
 a2254a <=( a386a ) or ( a387a );
 a2257a <=( a384a ) or ( a385a );
 a2258a <=( a2257a ) or ( a2254a );
 a2261a <=( a382a ) or ( a383a );
 a2264a <=( a380a ) or ( a381a );
 a2265a <=( a2264a ) or ( a2261a );
 a2266a <=( a2265a ) or ( a2258a );
 a2267a <=( a2266a ) or ( a2251a );
 a2268a <=( a2267a ) or ( a2236a );
 a2269a <=( a2268a ) or ( a2205a );
 a2270a <=( a2269a ) or ( a2144a );
 a2274a <=( a377a ) or ( a378a );
 a2275a <=( a379a ) or ( a2274a );
 a2278a <=( a375a ) or ( a376a );
 a2281a <=( a373a ) or ( a374a );
 a2282a <=( a2281a ) or ( a2278a );
 a2283a <=( a2282a ) or ( a2275a );
 a2286a <=( a371a ) or ( a372a );
 a2289a <=( a369a ) or ( a370a );
 a2290a <=( a2289a ) or ( a2286a );
 a2293a <=( a367a ) or ( a368a );
 a2296a <=( a365a ) or ( a366a );
 a2297a <=( a2296a ) or ( a2293a );
 a2298a <=( a2297a ) or ( a2290a );
 a2299a <=( a2298a ) or ( a2283a );
 a2302a <=( a363a ) or ( a364a );
 a2305a <=( a361a ) or ( a362a );
 a2306a <=( a2305a ) or ( a2302a );
 a2309a <=( a359a ) or ( a360a );
 a2312a <=( a357a ) or ( a358a );
 a2313a <=( a2312a ) or ( a2309a );
 a2314a <=( a2313a ) or ( a2306a );
 a2317a <=( a355a ) or ( a356a );
 a2320a <=( a353a ) or ( a354a );
 a2321a <=( a2320a ) or ( a2317a );
 a2324a <=( a351a ) or ( a352a );
 a2327a <=( a349a ) or ( a350a );
 a2328a <=( a2327a ) or ( a2324a );
 a2329a <=( a2328a ) or ( a2321a );
 a2330a <=( a2329a ) or ( a2314a );
 a2331a <=( a2330a ) or ( a2299a );
 a2334a <=( a347a ) or ( a348a );
 a2337a <=( a345a ) or ( a346a );
 a2338a <=( a2337a ) or ( a2334a );
 a2341a <=( a343a ) or ( a344a );
 a2344a <=( a341a ) or ( a342a );
 a2345a <=( a2344a ) or ( a2341a );
 a2346a <=( a2345a ) or ( a2338a );
 a2349a <=( a339a ) or ( a340a );
 a2352a <=( a337a ) or ( a338a );
 a2353a <=( a2352a ) or ( a2349a );
 a2356a <=( a335a ) or ( a336a );
 a2359a <=( a333a ) or ( a334a );
 a2360a <=( a2359a ) or ( a2356a );
 a2361a <=( a2360a ) or ( a2353a );
 a2362a <=( a2361a ) or ( a2346a );
 a2365a <=( a331a ) or ( a332a );
 a2368a <=( a329a ) or ( a330a );
 a2369a <=( a2368a ) or ( a2365a );
 a2372a <=( a327a ) or ( a328a );
 a2375a <=( a325a ) or ( a326a );
 a2376a <=( a2375a ) or ( a2372a );
 a2377a <=( a2376a ) or ( a2369a );
 a2380a <=( a323a ) or ( a324a );
 a2383a <=( a321a ) or ( a322a );
 a2384a <=( a2383a ) or ( a2380a );
 a2387a <=( a319a ) or ( a320a );
 a2390a <=( a317a ) or ( a318a );
 a2391a <=( a2390a ) or ( a2387a );
 a2392a <=( a2391a ) or ( a2384a );
 a2393a <=( a2392a ) or ( a2377a );
 a2394a <=( a2393a ) or ( a2362a );
 a2395a <=( a2394a ) or ( a2331a );
 a2399a <=( a314a ) or ( a315a );
 a2400a <=( a316a ) or ( a2399a );
 a2403a <=( a312a ) or ( a313a );
 a2406a <=( a310a ) or ( a311a );
 a2407a <=( a2406a ) or ( a2403a );
 a2408a <=( a2407a ) or ( a2400a );
 a2411a <=( a308a ) or ( a309a );
 a2414a <=( a306a ) or ( a307a );
 a2415a <=( a2414a ) or ( a2411a );
 a2418a <=( a304a ) or ( a305a );
 a2421a <=( a302a ) or ( a303a );
 a2422a <=( a2421a ) or ( a2418a );
 a2423a <=( a2422a ) or ( a2415a );
 a2424a <=( a2423a ) or ( a2408a );
 a2427a <=( a300a ) or ( a301a );
 a2430a <=( a298a ) or ( a299a );
 a2431a <=( a2430a ) or ( a2427a );
 a2434a <=( a296a ) or ( a297a );
 a2437a <=( a294a ) or ( a295a );
 a2438a <=( a2437a ) or ( a2434a );
 a2439a <=( a2438a ) or ( a2431a );
 a2442a <=( a292a ) or ( a293a );
 a2445a <=( a290a ) or ( a291a );
 a2446a <=( a2445a ) or ( a2442a );
 a2449a <=( a288a ) or ( a289a );
 a2452a <=( a286a ) or ( a287a );
 a2453a <=( a2452a ) or ( a2449a );
 a2454a <=( a2453a ) or ( a2446a );
 a2455a <=( a2454a ) or ( a2439a );
 a2456a <=( a2455a ) or ( a2424a );
 a2459a <=( a284a ) or ( a285a );
 a2462a <=( a282a ) or ( a283a );
 a2463a <=( a2462a ) or ( a2459a );
 a2466a <=( a280a ) or ( a281a );
 a2469a <=( a278a ) or ( a279a );
 a2470a <=( a2469a ) or ( a2466a );
 a2471a <=( a2470a ) or ( a2463a );
 a2474a <=( a276a ) or ( a277a );
 a2477a <=( a274a ) or ( a275a );
 a2478a <=( a2477a ) or ( a2474a );
 a2481a <=( a272a ) or ( a273a );
 a2484a <=( a270a ) or ( a271a );
 a2485a <=( a2484a ) or ( a2481a );
 a2486a <=( a2485a ) or ( a2478a );
 a2487a <=( a2486a ) or ( a2471a );
 a2490a <=( a268a ) or ( a269a );
 a2493a <=( a266a ) or ( a267a );
 a2494a <=( a2493a ) or ( a2490a );
 a2497a <=( a264a ) or ( a265a );
 a2500a <=( a262a ) or ( a263a );
 a2501a <=( a2500a ) or ( a2497a );
 a2502a <=( a2501a ) or ( a2494a );
 a2505a <=( a260a ) or ( a261a );
 a2508a <=( a258a ) or ( a259a );
 a2509a <=( a2508a ) or ( a2505a );
 a2512a <=( a256a ) or ( a257a );
 a2515a <=( a254a ) or ( a255a );
 a2516a <=( a2515a ) or ( a2512a );
 a2517a <=( a2516a ) or ( a2509a );
 a2518a <=( a2517a ) or ( a2502a );
 a2519a <=( a2518a ) or ( a2487a );
 a2520a <=( a2519a ) or ( a2456a );
 a2521a <=( a2520a ) or ( a2395a );
 a2522a <=( a2521a ) or ( a2270a );
 a2526a <=( a251a ) or ( a252a );
 a2527a <=( a253a ) or ( a2526a );
 a2530a <=( a249a ) or ( a250a );
 a2533a <=( a247a ) or ( a248a );
 a2534a <=( a2533a ) or ( a2530a );
 a2535a <=( a2534a ) or ( a2527a );
 a2538a <=( a245a ) or ( a246a );
 a2541a <=( a243a ) or ( a244a );
 a2542a <=( a2541a ) or ( a2538a );
 a2545a <=( a241a ) or ( a242a );
 a2548a <=( a239a ) or ( a240a );
 a2549a <=( a2548a ) or ( a2545a );
 a2550a <=( a2549a ) or ( a2542a );
 a2551a <=( a2550a ) or ( a2535a );
 a2554a <=( a237a ) or ( a238a );
 a2557a <=( a235a ) or ( a236a );
 a2558a <=( a2557a ) or ( a2554a );
 a2561a <=( a233a ) or ( a234a );
 a2564a <=( a231a ) or ( a232a );
 a2565a <=( a2564a ) or ( a2561a );
 a2566a <=( a2565a ) or ( a2558a );
 a2569a <=( a229a ) or ( a230a );
 a2572a <=( a227a ) or ( a228a );
 a2573a <=( a2572a ) or ( a2569a );
 a2576a <=( a225a ) or ( a226a );
 a2579a <=( a223a ) or ( a224a );
 a2580a <=( a2579a ) or ( a2576a );
 a2581a <=( a2580a ) or ( a2573a );
 a2582a <=( a2581a ) or ( a2566a );
 a2583a <=( a2582a ) or ( a2551a );
 a2586a <=( a221a ) or ( a222a );
 a2589a <=( a219a ) or ( a220a );
 a2590a <=( a2589a ) or ( a2586a );
 a2593a <=( a217a ) or ( a218a );
 a2596a <=( a215a ) or ( a216a );
 a2597a <=( a2596a ) or ( a2593a );
 a2598a <=( a2597a ) or ( a2590a );
 a2601a <=( a213a ) or ( a214a );
 a2604a <=( a211a ) or ( a212a );
 a2605a <=( a2604a ) or ( a2601a );
 a2608a <=( a209a ) or ( a210a );
 a2611a <=( a207a ) or ( a208a );
 a2612a <=( a2611a ) or ( a2608a );
 a2613a <=( a2612a ) or ( a2605a );
 a2614a <=( a2613a ) or ( a2598a );
 a2617a <=( a205a ) or ( a206a );
 a2620a <=( a203a ) or ( a204a );
 a2621a <=( a2620a ) or ( a2617a );
 a2624a <=( a201a ) or ( a202a );
 a2627a <=( a199a ) or ( a200a );
 a2628a <=( a2627a ) or ( a2624a );
 a2629a <=( a2628a ) or ( a2621a );
 a2632a <=( a197a ) or ( a198a );
 a2635a <=( a195a ) or ( a196a );
 a2636a <=( a2635a ) or ( a2632a );
 a2639a <=( a193a ) or ( a194a );
 a2642a <=( a191a ) or ( a192a );
 a2643a <=( a2642a ) or ( a2639a );
 a2644a <=( a2643a ) or ( a2636a );
 a2645a <=( a2644a ) or ( a2629a );
 a2646a <=( a2645a ) or ( a2614a );
 a2647a <=( a2646a ) or ( a2583a );
 a2651a <=( a188a ) or ( a189a );
 a2652a <=( a190a ) or ( a2651a );
 a2655a <=( a186a ) or ( a187a );
 a2658a <=( a184a ) or ( a185a );
 a2659a <=( a2658a ) or ( a2655a );
 a2660a <=( a2659a ) or ( a2652a );
 a2663a <=( a182a ) or ( a183a );
 a2666a <=( a180a ) or ( a181a );
 a2667a <=( a2666a ) or ( a2663a );
 a2670a <=( a178a ) or ( a179a );
 a2673a <=( a176a ) or ( a177a );
 a2674a <=( a2673a ) or ( a2670a );
 a2675a <=( a2674a ) or ( a2667a );
 a2676a <=( a2675a ) or ( a2660a );
 a2679a <=( a174a ) or ( a175a );
 a2682a <=( a172a ) or ( a173a );
 a2683a <=( a2682a ) or ( a2679a );
 a2686a <=( a170a ) or ( a171a );
 a2689a <=( a168a ) or ( a169a );
 a2690a <=( a2689a ) or ( a2686a );
 a2691a <=( a2690a ) or ( a2683a );
 a2694a <=( a166a ) or ( a167a );
 a2697a <=( a164a ) or ( a165a );
 a2698a <=( a2697a ) or ( a2694a );
 a2701a <=( a162a ) or ( a163a );
 a2704a <=( a160a ) or ( a161a );
 a2705a <=( a2704a ) or ( a2701a );
 a2706a <=( a2705a ) or ( a2698a );
 a2707a <=( a2706a ) or ( a2691a );
 a2708a <=( a2707a ) or ( a2676a );
 a2711a <=( a158a ) or ( a159a );
 a2714a <=( a156a ) or ( a157a );
 a2715a <=( a2714a ) or ( a2711a );
 a2718a <=( a154a ) or ( a155a );
 a2721a <=( a152a ) or ( a153a );
 a2722a <=( a2721a ) or ( a2718a );
 a2723a <=( a2722a ) or ( a2715a );
 a2726a <=( a150a ) or ( a151a );
 a2729a <=( a148a ) or ( a149a );
 a2730a <=( a2729a ) or ( a2726a );
 a2733a <=( a146a ) or ( a147a );
 a2736a <=( a144a ) or ( a145a );
 a2737a <=( a2736a ) or ( a2733a );
 a2738a <=( a2737a ) or ( a2730a );
 a2739a <=( a2738a ) or ( a2723a );
 a2742a <=( a142a ) or ( a143a );
 a2745a <=( a140a ) or ( a141a );
 a2746a <=( a2745a ) or ( a2742a );
 a2749a <=( a138a ) or ( a139a );
 a2752a <=( a136a ) or ( a137a );
 a2753a <=( a2752a ) or ( a2749a );
 a2754a <=( a2753a ) or ( a2746a );
 a2757a <=( a134a ) or ( a135a );
 a2760a <=( a132a ) or ( a133a );
 a2761a <=( a2760a ) or ( a2757a );
 a2764a <=( a130a ) or ( a131a );
 a2767a <=( a128a ) or ( a129a );
 a2768a <=( a2767a ) or ( a2764a );
 a2769a <=( a2768a ) or ( a2761a );
 a2770a <=( a2769a ) or ( a2754a );
 a2771a <=( a2770a ) or ( a2739a );
 a2772a <=( a2771a ) or ( a2708a );
 a2773a <=( a2772a ) or ( a2647a );
 a2777a <=( a125a ) or ( a126a );
 a2778a <=( a127a ) or ( a2777a );
 a2781a <=( a123a ) or ( a124a );
 a2784a <=( a121a ) or ( a122a );
 a2785a <=( a2784a ) or ( a2781a );
 a2786a <=( a2785a ) or ( a2778a );
 a2789a <=( a119a ) or ( a120a );
 a2792a <=( a117a ) or ( a118a );
 a2793a <=( a2792a ) or ( a2789a );
 a2796a <=( a115a ) or ( a116a );
 a2799a <=( a113a ) or ( a114a );
 a2800a <=( a2799a ) or ( a2796a );
 a2801a <=( a2800a ) or ( a2793a );
 a2802a <=( a2801a ) or ( a2786a );
 a2805a <=( a111a ) or ( a112a );
 a2808a <=( a109a ) or ( a110a );
 a2809a <=( a2808a ) or ( a2805a );
 a2812a <=( a107a ) or ( a108a );
 a2815a <=( a105a ) or ( a106a );
 a2816a <=( a2815a ) or ( a2812a );
 a2817a <=( a2816a ) or ( a2809a );
 a2820a <=( a103a ) or ( a104a );
 a2823a <=( a101a ) or ( a102a );
 a2824a <=( a2823a ) or ( a2820a );
 a2827a <=( a99a ) or ( a100a );
 a2830a <=( a97a ) or ( a98a );
 a2831a <=( a2830a ) or ( a2827a );
 a2832a <=( a2831a ) or ( a2824a );
 a2833a <=( a2832a ) or ( a2817a );
 a2834a <=( a2833a ) or ( a2802a );
 a2837a <=( a95a ) or ( a96a );
 a2840a <=( a93a ) or ( a94a );
 a2841a <=( a2840a ) or ( a2837a );
 a2844a <=( a91a ) or ( a92a );
 a2847a <=( a89a ) or ( a90a );
 a2848a <=( a2847a ) or ( a2844a );
 a2849a <=( a2848a ) or ( a2841a );
 a2852a <=( a87a ) or ( a88a );
 a2855a <=( a85a ) or ( a86a );
 a2856a <=( a2855a ) or ( a2852a );
 a2859a <=( a83a ) or ( a84a );
 a2862a <=( a81a ) or ( a82a );
 a2863a <=( a2862a ) or ( a2859a );
 a2864a <=( a2863a ) or ( a2856a );
 a2865a <=( a2864a ) or ( a2849a );
 a2868a <=( a79a ) or ( a80a );
 a2871a <=( a77a ) or ( a78a );
 a2872a <=( a2871a ) or ( a2868a );
 a2875a <=( a75a ) or ( a76a );
 a2878a <=( a73a ) or ( a74a );
 a2879a <=( a2878a ) or ( a2875a );
 a2880a <=( a2879a ) or ( a2872a );
 a2883a <=( a71a ) or ( a72a );
 a2886a <=( a69a ) or ( a70a );
 a2887a <=( a2886a ) or ( a2883a );
 a2890a <=( a67a ) or ( a68a );
 a2893a <=( a65a ) or ( a66a );
 a2894a <=( a2893a ) or ( a2890a );
 a2895a <=( a2894a ) or ( a2887a );
 a2896a <=( a2895a ) or ( a2880a );
 a2897a <=( a2896a ) or ( a2865a );
 a2898a <=( a2897a ) or ( a2834a );
 a2901a <=( a63a ) or ( a64a );
 a2904a <=( a61a ) or ( a62a );
 a2905a <=( a2904a ) or ( a2901a );
 a2908a <=( a59a ) or ( a60a );
 a2911a <=( a57a ) or ( a58a );
 a2912a <=( a2911a ) or ( a2908a );
 a2913a <=( a2912a ) or ( a2905a );
 a2916a <=( a55a ) or ( a56a );
 a2919a <=( a53a ) or ( a54a );
 a2920a <=( a2919a ) or ( a2916a );
 a2923a <=( a51a ) or ( a52a );
 a2926a <=( a49a ) or ( a50a );
 a2927a <=( a2926a ) or ( a2923a );
 a2928a <=( a2927a ) or ( a2920a );
 a2929a <=( a2928a ) or ( a2913a );
 a2932a <=( a47a ) or ( a48a );
 a2935a <=( a45a ) or ( a46a );
 a2936a <=( a2935a ) or ( a2932a );
 a2939a <=( a43a ) or ( a44a );
 a2942a <=( a41a ) or ( a42a );
 a2943a <=( a2942a ) or ( a2939a );
 a2944a <=( a2943a ) or ( a2936a );
 a2947a <=( a39a ) or ( a40a );
 a2950a <=( a37a ) or ( a38a );
 a2951a <=( a2950a ) or ( a2947a );
 a2954a <=( a35a ) or ( a36a );
 a2957a <=( a33a ) or ( a34a );
 a2958a <=( a2957a ) or ( a2954a );
 a2959a <=( a2958a ) or ( a2951a );
 a2960a <=( a2959a ) or ( a2944a );
 a2961a <=( a2960a ) or ( a2929a );
 a2964a <=( a31a ) or ( a32a );
 a2967a <=( a29a ) or ( a30a );
 a2968a <=( a2967a ) or ( a2964a );
 a2971a <=( a27a ) or ( a28a );
 a2974a <=( a25a ) or ( a26a );
 a2975a <=( a2974a ) or ( a2971a );
 a2976a <=( a2975a ) or ( a2968a );
 a2979a <=( a23a ) or ( a24a );
 a2982a <=( a21a ) or ( a22a );
 a2983a <=( a2982a ) or ( a2979a );
 a2986a <=( a19a ) or ( a20a );
 a2989a <=( a17a ) or ( a18a );
 a2990a <=( a2989a ) or ( a2986a );
 a2991a <=( a2990a ) or ( a2983a );
 a2992a <=( a2991a ) or ( a2976a );
 a2995a <=( a15a ) or ( a16a );
 a2998a <=( a13a ) or ( a14a );
 a2999a <=( a2998a ) or ( a2995a );
 a3002a <=( a11a ) or ( a12a );
 a3005a <=( a9a ) or ( a10a );
 a3006a <=( a3005a ) or ( a3002a );
 a3007a <=( a3006a ) or ( a2999a );
 a3010a <=( a7a ) or ( a8a );
 a3013a <=( a5a ) or ( a6a );
 a3014a <=( a3013a ) or ( a3010a );
 a3017a <=( a3a ) or ( a4a );
 a3020a <=( a1a ) or ( a2a );
 a3021a <=( a3020a ) or ( a3017a );
 a3022a <=( a3021a ) or ( a3014a );
 a3023a <=( a3022a ) or ( a3007a );
 a3024a <=( a3023a ) or ( a2992a );
 a3025a <=( a3024a ) or ( a2961a );
 a3026a <=( a3025a ) or ( a2898a );
 a3027a <=( a3026a ) or ( a2773a );
 a3028a <=( a3027a ) or ( a2522a );
 a3036a <=( A234  and  A232 );
 a3040a <=( A234  and  A233 );
 a3044a <=( A235  and  A201 );
 a3048a <=( A235  and  A201 );
 a3052a <=( A235  and  A166 );
 a3056a <=( A235  and  A167 );
 a3060a <=( A234  and  A232 );
 a3064a <=( A234  and  A233 );
 a3067a <=( (not A232)  and  A202 );
 a3070a <=( A236  and  A233 );
 a3073a <=( A232  and  A202 );
 a3076a <=( A236  and  (not A233) );
 a3079a <=( A201  and  A199 );
 a3082a <=( A234  and  A232 );
 a3085a <=( A201  and  A199 );
 a3088a <=( A234  and  A233 );
 a3091a <=( A201  and  A200 );
 a3094a <=( A234  and  A232 );
 a3097a <=( A201  and  A200 );
 a3100a <=( A234  and  A233 );
 a3103a <=( A200  and  (not A199) );
 a3106a <=( A235  and  A203 );
 a3109a <=( (not A200)  and  A199 );
 a3112a <=( A235  and  A203 );
 a3115a <=( A166  and  A168 );
 a3118a <=( A234  and  A232 );
 a3121a <=( A166  and  A168 );
 a3124a <=( A234  and  A233 );
 a3127a <=( A167  and  A168 );
 a3130a <=( A234  and  A232 );
 a3133a <=( A167  and  A168 );
 a3136a <=( A234  and  A233 );
 a3139a <=( A167  and  A170 );
 a3142a <=( A235  and  (not A166) );
 a3145a <=( (not A167)  and  A170 );
 a3148a <=( A235  and  A166 );
 a3151a <=( (not A232)  and  A169 );
 a3154a <=( A236  and  A233 );
 a3157a <=( A232  and  A169 );
 a3160a <=( A236  and  (not A233) );
 a3163a <=( A201  and  A199 );
 a3167a <=( A236  and  A233 );
 a3168a <=( (not A232)  and  a3167a );
 a3171a <=( A201  and  A199 );
 a3175a <=( A236  and  (not A233) );
 a3176a <=( A232  and  a3175a );
 a3179a <=( A201  and  A200 );
 a3183a <=( A236  and  A233 );
 a3184a <=( (not A232)  and  a3183a );
 a3187a <=( A201  and  A200 );
 a3191a <=( A236  and  (not A233) );
 a3192a <=( A232  and  a3191a );
 a3195a <=( A200  and  (not A199) );
 a3199a <=( A234  and  A232 );
 a3200a <=( A203  and  a3199a );
 a3203a <=( A200  and  (not A199) );
 a3207a <=( A234  and  A233 );
 a3208a <=( A203  and  a3207a );
 a3211a <=( (not A200)  and  A199 );
 a3215a <=( A234  and  A232 );
 a3216a <=( A203  and  a3215a );
 a3219a <=( (not A200)  and  A199 );
 a3223a <=( A234  and  A233 );
 a3224a <=( A203  and  a3223a );
 a3227a <=( A166  and  A168 );
 a3231a <=( A236  and  A233 );
 a3232a <=( (not A232)  and  a3231a );
 a3235a <=( A166  and  A168 );
 a3239a <=( A236  and  (not A233) );
 a3240a <=( A232  and  a3239a );
 a3243a <=( A167  and  A168 );
 a3247a <=( A236  and  A233 );
 a3248a <=( (not A232)  and  a3247a );
 a3251a <=( A167  and  A168 );
 a3255a <=( A236  and  (not A233) );
 a3256a <=( A232  and  a3255a );
 a3259a <=( A167  and  A170 );
 a3263a <=( A234  and  A232 );
 a3264a <=( (not A166)  and  a3263a );
 a3267a <=( A167  and  A170 );
 a3271a <=( A234  and  A233 );
 a3272a <=( (not A166)  and  a3271a );
 a3275a <=( (not A167)  and  A170 );
 a3279a <=( A234  and  A232 );
 a3280a <=( A166  and  a3279a );
 a3283a <=( (not A167)  and  A170 );
 a3287a <=( A234  and  A233 );
 a3288a <=( A166  and  a3287a );
 a3292a <=( A203  and  A200 );
 a3293a <=( (not A199)  and  a3292a );
 a3297a <=( A236  and  A233 );
 a3298a <=( (not A232)  and  a3297a );
 a3302a <=( A203  and  A200 );
 a3303a <=( (not A199)  and  a3302a );
 a3307a <=( A236  and  (not A233) );
 a3308a <=( A232  and  a3307a );
 a3312a <=( A203  and  (not A200) );
 a3313a <=( A199  and  a3312a );
 a3317a <=( A236  and  A233 );
 a3318a <=( (not A232)  and  a3317a );
 a3322a <=( A203  and  (not A200) );
 a3323a <=( A199  and  a3322a );
 a3327a <=( A236  and  (not A233) );
 a3328a <=( A232  and  a3327a );
 a3332a <=( (not A166)  and  A167 );
 a3333a <=( A170  and  a3332a );
 a3337a <=( A236  and  A233 );
 a3338a <=( (not A232)  and  a3337a );
 a3342a <=( (not A166)  and  A167 );
 a3343a <=( A170  and  a3342a );
 a3347a <=( A236  and  (not A233) );
 a3348a <=( A232  and  a3347a );
 a3352a <=( A166  and  (not A167) );
 a3353a <=( A170  and  a3352a );
 a3357a <=( A236  and  A233 );
 a3358a <=( (not A232)  and  a3357a );
 a3362a <=( A166  and  (not A167) );
 a3363a <=( A170  and  a3362a );
 a3367a <=( A236  and  (not A233) );
 a3368a <=( A232  and  a3367a );
 a3372a <=( A268  and  A202 );
 a3373a <=( A169  and  a3372a );
 a3377a <=( (not A302)  and  (not A301) );
 a3378a <=( (not A300)  and  a3377a );
 a3382a <=( A268  and  A202 );
 a3383a <=( A169  and  a3382a );
 a3387a <=( (not A301)  and  (not A299) );
 a3388a <=( (not A298)  and  a3387a );
 a3392a <=( A202  and  A166 );
 a3393a <=( A168  and  a3392a );
 a3396a <=( (not A300)  and  A268 );
 a3399a <=( (not A302)  and  (not A301) );
 a3400a <=( a3399a  and  a3396a );
 a3404a <=( A202  and  A166 );
 a3405a <=( A168  and  a3404a );
 a3408a <=( (not A298)  and  A268 );
 a3411a <=( (not A301)  and  (not A299) );
 a3412a <=( a3411a  and  a3408a );
 a3416a <=( A202  and  A167 );
 a3417a <=( A168  and  a3416a );
 a3420a <=( (not A300)  and  A268 );
 a3423a <=( (not A302)  and  (not A301) );
 a3424a <=( a3423a  and  a3420a );
 a3428a <=( A202  and  A167 );
 a3429a <=( A168  and  a3428a );
 a3432a <=( (not A298)  and  A268 );
 a3435a <=( (not A301)  and  (not A299) );
 a3436a <=( a3435a  and  a3432a );
 a3440a <=( A268  and  A202 );
 a3441a <=( A169  and  a3440a );
 a3444a <=( A299  and  A298 );
 a3447a <=( (not A301)  and  (not A300) );
 a3448a <=( a3447a  and  a3444a );
 a3452a <=( A265  and  A202 );
 a3453a <=( A169  and  a3452a );
 a3456a <=( (not A300)  and  A267 );
 a3459a <=( (not A302)  and  (not A301) );
 a3460a <=( a3459a  and  a3456a );
 a3464a <=( A265  and  A202 );
 a3465a <=( A169  and  a3464a );
 a3468a <=( (not A298)  and  A267 );
 a3471a <=( (not A301)  and  (not A299) );
 a3472a <=( a3471a  and  a3468a );
 a3476a <=( A266  and  A202 );
 a3477a <=( A169  and  a3476a );
 a3480a <=( (not A300)  and  A267 );
 a3483a <=( (not A302)  and  (not A301) );
 a3484a <=( a3483a  and  a3480a );
 a3488a <=( A266  and  A202 );
 a3489a <=( A169  and  a3488a );
 a3492a <=( (not A298)  and  A267 );
 a3495a <=( (not A301)  and  (not A299) );
 a3496a <=( a3495a  and  a3492a );
 a3500a <=( A201  and  A199 );
 a3501a <=( A169  and  a3500a );
 a3504a <=( (not A300)  and  A268 );
 a3507a <=( (not A302)  and  (not A301) );
 a3508a <=( a3507a  and  a3504a );
 a3512a <=( A201  and  A199 );
 a3513a <=( A169  and  a3512a );
 a3516a <=( (not A298)  and  A268 );
 a3519a <=( (not A301)  and  (not A299) );
 a3520a <=( a3519a  and  a3516a );
 a3524a <=( A201  and  A200 );
 a3525a <=( A169  and  a3524a );
 a3528a <=( (not A300)  and  A268 );
 a3531a <=( (not A302)  and  (not A301) );
 a3532a <=( a3531a  and  a3528a );
 a3536a <=( A201  and  A200 );
 a3537a <=( A169  and  a3536a );
 a3540a <=( (not A298)  and  A268 );
 a3543a <=( (not A301)  and  (not A299) );
 a3544a <=( a3543a  and  a3540a );
 a3547a <=( A166  and  A168 );
 a3550a <=( A268  and  A202 );
 a3551a <=( a3550a  and  a3547a );
 a3554a <=( A299  and  A298 );
 a3557a <=( (not A301)  and  (not A300) );
 a3558a <=( a3557a  and  a3554a );
 a3561a <=( A166  and  A168 );
 a3564a <=( A265  and  A202 );
 a3565a <=( a3564a  and  a3561a );
 a3568a <=( (not A300)  and  A267 );
 a3571a <=( (not A302)  and  (not A301) );
 a3572a <=( a3571a  and  a3568a );
 a3575a <=( A166  and  A168 );
 a3578a <=( A265  and  A202 );
 a3579a <=( a3578a  and  a3575a );
 a3582a <=( (not A298)  and  A267 );
 a3585a <=( (not A301)  and  (not A299) );
 a3586a <=( a3585a  and  a3582a );
 a3589a <=( A166  and  A168 );
 a3592a <=( A266  and  A202 );
 a3593a <=( a3592a  and  a3589a );
 a3596a <=( (not A300)  and  A267 );
 a3599a <=( (not A302)  and  (not A301) );
 a3600a <=( a3599a  and  a3596a );
 a3603a <=( A166  and  A168 );
 a3606a <=( A266  and  A202 );
 a3607a <=( a3606a  and  a3603a );
 a3610a <=( (not A298)  and  A267 );
 a3613a <=( (not A301)  and  (not A299) );
 a3614a <=( a3613a  and  a3610a );
 a3617a <=( A166  and  A168 );
 a3620a <=( A201  and  A199 );
 a3621a <=( a3620a  and  a3617a );
 a3624a <=( (not A300)  and  A268 );
 a3627a <=( (not A302)  and  (not A301) );
 a3628a <=( a3627a  and  a3624a );
 a3631a <=( A166  and  A168 );
 a3634a <=( A201  and  A199 );
 a3635a <=( a3634a  and  a3631a );
 a3638a <=( (not A298)  and  A268 );
 a3641a <=( (not A301)  and  (not A299) );
 a3642a <=( a3641a  and  a3638a );
 a3645a <=( A166  and  A168 );
 a3648a <=( A201  and  A200 );
 a3649a <=( a3648a  and  a3645a );
 a3652a <=( (not A300)  and  A268 );
 a3655a <=( (not A302)  and  (not A301) );
 a3656a <=( a3655a  and  a3652a );
 a3659a <=( A166  and  A168 );
 a3662a <=( A201  and  A200 );
 a3663a <=( a3662a  and  a3659a );
 a3666a <=( (not A298)  and  A268 );
 a3669a <=( (not A301)  and  (not A299) );
 a3670a <=( a3669a  and  a3666a );
 a3673a <=( A167  and  A168 );
 a3676a <=( A268  and  A202 );
 a3677a <=( a3676a  and  a3673a );
 a3680a <=( A299  and  A298 );
 a3683a <=( (not A301)  and  (not A300) );
 a3684a <=( a3683a  and  a3680a );
 a3687a <=( A167  and  A168 );
 a3690a <=( A265  and  A202 );
 a3691a <=( a3690a  and  a3687a );
 a3694a <=( (not A300)  and  A267 );
 a3697a <=( (not A302)  and  (not A301) );
 a3698a <=( a3697a  and  a3694a );
 a3701a <=( A167  and  A168 );
 a3704a <=( A265  and  A202 );
 a3705a <=( a3704a  and  a3701a );
 a3708a <=( (not A298)  and  A267 );
 a3711a <=( (not A301)  and  (not A299) );
 a3712a <=( a3711a  and  a3708a );
 a3715a <=( A167  and  A168 );
 a3718a <=( A266  and  A202 );
 a3719a <=( a3718a  and  a3715a );
 a3722a <=( (not A300)  and  A267 );
 a3725a <=( (not A302)  and  (not A301) );
 a3726a <=( a3725a  and  a3722a );
 a3729a <=( A167  and  A168 );
 a3732a <=( A266  and  A202 );
 a3733a <=( a3732a  and  a3729a );
 a3736a <=( (not A298)  and  A267 );
 a3739a <=( (not A301)  and  (not A299) );
 a3740a <=( a3739a  and  a3736a );
 a3743a <=( A167  and  A168 );
 a3746a <=( A201  and  A199 );
 a3747a <=( a3746a  and  a3743a );
 a3750a <=( (not A300)  and  A268 );
 a3753a <=( (not A302)  and  (not A301) );
 a3754a <=( a3753a  and  a3750a );
 a3757a <=( A167  and  A168 );
 a3760a <=( A201  and  A199 );
 a3761a <=( a3760a  and  a3757a );
 a3764a <=( (not A298)  and  A268 );
 a3767a <=( (not A301)  and  (not A299) );
 a3768a <=( a3767a  and  a3764a );
 a3771a <=( A167  and  A168 );
 a3774a <=( A201  and  A200 );
 a3775a <=( a3774a  and  a3771a );
 a3778a <=( (not A300)  and  A268 );
 a3781a <=( (not A302)  and  (not A301) );
 a3782a <=( a3781a  and  a3778a );
 a3785a <=( A167  and  A168 );
 a3788a <=( A201  and  A200 );
 a3789a <=( a3788a  and  a3785a );
 a3792a <=( (not A298)  and  A268 );
 a3795a <=( (not A301)  and  (not A299) );
 a3796a <=( a3795a  and  a3792a );
 a3799a <=( A167  and  A170 );
 a3802a <=( A202  and  (not A166) );
 a3803a <=( a3802a  and  a3799a );
 a3806a <=( (not A300)  and  A268 );
 a3809a <=( (not A302)  and  (not A301) );
 a3810a <=( a3809a  and  a3806a );
 a3813a <=( A167  and  A170 );
 a3816a <=( A202  and  (not A166) );
 a3817a <=( a3816a  and  a3813a );
 a3820a <=( (not A298)  and  A268 );
 a3823a <=( (not A301)  and  (not A299) );
 a3824a <=( a3823a  and  a3820a );
 a3827a <=( (not A167)  and  A170 );
 a3830a <=( A202  and  A166 );
 a3831a <=( a3830a  and  a3827a );
 a3834a <=( (not A300)  and  A268 );
 a3837a <=( (not A302)  and  (not A301) );
 a3838a <=( a3837a  and  a3834a );
 a3841a <=( (not A167)  and  A170 );
 a3844a <=( A202  and  A166 );
 a3845a <=( a3844a  and  a3841a );
 a3848a <=( (not A298)  and  A268 );
 a3851a <=( (not A301)  and  (not A299) );
 a3852a <=( a3851a  and  a3848a );
 a3855a <=( A202  and  A169 );
 a3858a <=( A267  and  A265 );
 a3859a <=( a3858a  and  a3855a );
 a3862a <=( A299  and  A298 );
 a3865a <=( (not A301)  and  (not A300) );
 a3866a <=( a3865a  and  a3862a );
 a3869a <=( A202  and  A169 );
 a3872a <=( A267  and  A266 );
 a3873a <=( a3872a  and  a3869a );
 a3876a <=( A299  and  A298 );
 a3879a <=( (not A301)  and  (not A300) );
 a3880a <=( a3879a  and  a3876a );
 a3883a <=( A202  and  A169 );
 a3886a <=( A266  and  (not A265) );
 a3887a <=( a3886a  and  a3883a );
 a3890a <=( (not A300)  and  A269 );
 a3893a <=( (not A302)  and  (not A301) );
 a3894a <=( a3893a  and  a3890a );
 a3897a <=( A202  and  A169 );
 a3900a <=( A266  and  (not A265) );
 a3901a <=( a3900a  and  a3897a );
 a3904a <=( (not A298)  and  A269 );
 a3907a <=( (not A301)  and  (not A299) );
 a3908a <=( a3907a  and  a3904a );
 a3911a <=( A202  and  A169 );
 a3914a <=( (not A266)  and  A265 );
 a3915a <=( a3914a  and  a3911a );
 a3918a <=( (not A300)  and  A269 );
 a3921a <=( (not A302)  and  (not A301) );
 a3922a <=( a3921a  and  a3918a );
 a3925a <=( A202  and  A169 );
 a3928a <=( (not A266)  and  A265 );
 a3929a <=( a3928a  and  a3925a );
 a3932a <=( (not A298)  and  A269 );
 a3935a <=( (not A301)  and  (not A299) );
 a3936a <=( a3935a  and  a3932a );
 a3939a <=( (not A201)  and  A169 );
 a3942a <=( (not A203)  and  (not A202) );
 a3943a <=( a3942a  and  a3939a );
 a3946a <=( (not A268)  and  (not A267) );
 a3949a <=( A301  and  (not A269) );
 a3950a <=( a3949a  and  a3946a );
 a3953a <=( (not A201)  and  A169 );
 a3956a <=( (not A203)  and  (not A202) );
 a3957a <=( a3956a  and  a3953a );
 a3960a <=( (not A266)  and  (not A265) );
 a3963a <=( A301  and  (not A268) );
 a3964a <=( a3963a  and  a3960a );
 a3967a <=( A199  and  A169 );
 a3970a <=( A268  and  A201 );
 a3971a <=( a3970a  and  a3967a );
 a3974a <=( A299  and  A298 );
 a3977a <=( (not A301)  and  (not A300) );
 a3978a <=( a3977a  and  a3974a );
 a3981a <=( A199  and  A169 );
 a3984a <=( A265  and  A201 );
 a3985a <=( a3984a  and  a3981a );
 a3988a <=( (not A300)  and  A267 );
 a3991a <=( (not A302)  and  (not A301) );
 a3992a <=( a3991a  and  a3988a );
 a3995a <=( A199  and  A169 );
 a3998a <=( A265  and  A201 );
 a3999a <=( a3998a  and  a3995a );
 a4002a <=( (not A298)  and  A267 );
 a4005a <=( (not A301)  and  (not A299) );
 a4006a <=( a4005a  and  a4002a );
 a4009a <=( A199  and  A169 );
 a4012a <=( A266  and  A201 );
 a4013a <=( a4012a  and  a4009a );
 a4016a <=( (not A300)  and  A267 );
 a4019a <=( (not A302)  and  (not A301) );
 a4020a <=( a4019a  and  a4016a );
 a4023a <=( A199  and  A169 );
 a4026a <=( A266  and  A201 );
 a4027a <=( a4026a  and  a4023a );
 a4030a <=( (not A298)  and  A267 );
 a4033a <=( (not A301)  and  (not A299) );
 a4034a <=( a4033a  and  a4030a );
 a4037a <=( A200  and  A169 );
 a4040a <=( A268  and  A201 );
 a4041a <=( a4040a  and  a4037a );
 a4044a <=( A299  and  A298 );
 a4047a <=( (not A301)  and  (not A300) );
 a4048a <=( a4047a  and  a4044a );
 a4051a <=( A200  and  A169 );
 a4054a <=( A265  and  A201 );
 a4055a <=( a4054a  and  a4051a );
 a4058a <=( (not A300)  and  A267 );
 a4061a <=( (not A302)  and  (not A301) );
 a4062a <=( a4061a  and  a4058a );
 a4065a <=( A200  and  A169 );
 a4068a <=( A265  and  A201 );
 a4069a <=( a4068a  and  a4065a );
 a4072a <=( (not A298)  and  A267 );
 a4075a <=( (not A301)  and  (not A299) );
 a4076a <=( a4075a  and  a4072a );
 a4079a <=( A200  and  A169 );
 a4082a <=( A266  and  A201 );
 a4083a <=( a4082a  and  a4079a );
 a4086a <=( (not A300)  and  A267 );
 a4089a <=( (not A302)  and  (not A301) );
 a4090a <=( a4089a  and  a4086a );
 a4093a <=( A200  and  A169 );
 a4096a <=( A266  and  A201 );
 a4097a <=( a4096a  and  a4093a );
 a4100a <=( (not A298)  and  A267 );
 a4103a <=( (not A301)  and  (not A299) );
 a4104a <=( a4103a  and  a4100a );
 a4107a <=( (not A199)  and  A169 );
 a4110a <=( A203  and  A200 );
 a4111a <=( a4110a  and  a4107a );
 a4114a <=( (not A300)  and  A268 );
 a4117a <=( (not A302)  and  (not A301) );
 a4118a <=( a4117a  and  a4114a );
 a4121a <=( (not A199)  and  A169 );
 a4124a <=( A203  and  A200 );
 a4125a <=( a4124a  and  a4121a );
 a4128a <=( (not A298)  and  A268 );
 a4131a <=( (not A301)  and  (not A299) );
 a4132a <=( a4131a  and  a4128a );
 a4135a <=( A199  and  A169 );
 a4138a <=( A203  and  (not A200) );
 a4139a <=( a4138a  and  a4135a );
 a4142a <=( (not A300)  and  A268 );
 a4145a <=( (not A302)  and  (not A301) );
 a4146a <=( a4145a  and  a4142a );
 a4149a <=( A199  and  A169 );
 a4152a <=( A203  and  (not A200) );
 a4153a <=( a4152a  and  a4149a );
 a4156a <=( (not A298)  and  A268 );
 a4159a <=( (not A301)  and  (not A299) );
 a4160a <=( a4159a  and  a4156a );
 a4163a <=( (not A199)  and  A169 );
 a4166a <=( (not A202)  and  (not A200) );
 a4167a <=( a4166a  and  a4163a );
 a4170a <=( (not A268)  and  (not A267) );
 a4173a <=( A301  and  (not A269) );
 a4174a <=( a4173a  and  a4170a );
 a4177a <=( (not A199)  and  A169 );
 a4180a <=( (not A202)  and  (not A200) );
 a4181a <=( a4180a  and  a4177a );
 a4184a <=( (not A266)  and  (not A265) );
 a4187a <=( A301  and  (not A268) );
 a4188a <=( a4187a  and  a4184a );
 a4191a <=( (not A167)  and  (not A169) );
 a4194a <=( A202  and  (not A166) );
 a4195a <=( a4194a  and  a4191a );
 a4198a <=( (not A268)  and  (not A267) );
 a4201a <=( A301  and  (not A269) );
 a4202a <=( a4201a  and  a4198a );
 a4205a <=( (not A167)  and  (not A169) );
 a4208a <=( A202  and  (not A166) );
 a4209a <=( a4208a  and  a4205a );
 a4212a <=( (not A266)  and  (not A265) );
 a4215a <=( A301  and  (not A268) );
 a4216a <=( a4215a  and  a4212a );
 a4219a <=( (not A169)  and  (not A170) );
 a4222a <=( A202  and  (not A168) );
 a4223a <=( a4222a  and  a4219a );
 a4226a <=( (not A268)  and  (not A267) );
 a4229a <=( A301  and  (not A269) );
 a4230a <=( a4229a  and  a4226a );
 a4233a <=( (not A169)  and  (not A170) );
 a4236a <=( A202  and  (not A168) );
 a4237a <=( a4236a  and  a4233a );
 a4240a <=( (not A266)  and  (not A265) );
 a4243a <=( A301  and  (not A268) );
 a4244a <=( a4243a  and  a4240a );
 a4247a <=( A166  and  A168 );
 a4250a <=( A265  and  A202 );
 a4251a <=( a4250a  and  a4247a );
 a4254a <=( A298  and  A267 );
 a4258a <=( (not A301)  and  (not A300) );
 a4259a <=( A299  and  a4258a );
 a4260a <=( a4259a  and  a4254a );
 a4263a <=( A166  and  A168 );
 a4266a <=( A266  and  A202 );
 a4267a <=( a4266a  and  a4263a );
 a4270a <=( A298  and  A267 );
 a4274a <=( (not A301)  and  (not A300) );
 a4275a <=( A299  and  a4274a );
 a4276a <=( a4275a  and  a4270a );
 a4279a <=( A166  and  A168 );
 a4282a <=( (not A265)  and  A202 );
 a4283a <=( a4282a  and  a4279a );
 a4286a <=( A269  and  A266 );
 a4290a <=( (not A302)  and  (not A301) );
 a4291a <=( (not A300)  and  a4290a );
 a4292a <=( a4291a  and  a4286a );
 a4295a <=( A166  and  A168 );
 a4298a <=( (not A265)  and  A202 );
 a4299a <=( a4298a  and  a4295a );
 a4302a <=( A269  and  A266 );
 a4306a <=( (not A301)  and  (not A299) );
 a4307a <=( (not A298)  and  a4306a );
 a4308a <=( a4307a  and  a4302a );
 a4311a <=( A166  and  A168 );
 a4314a <=( A265  and  A202 );
 a4315a <=( a4314a  and  a4311a );
 a4318a <=( A269  and  (not A266) );
 a4322a <=( (not A302)  and  (not A301) );
 a4323a <=( (not A300)  and  a4322a );
 a4324a <=( a4323a  and  a4318a );
 a4327a <=( A166  and  A168 );
 a4330a <=( A265  and  A202 );
 a4331a <=( a4330a  and  a4327a );
 a4334a <=( A269  and  (not A266) );
 a4338a <=( (not A301)  and  (not A299) );
 a4339a <=( (not A298)  and  a4338a );
 a4340a <=( a4339a  and  a4334a );
 a4343a <=( A166  and  A168 );
 a4346a <=( (not A202)  and  (not A201) );
 a4347a <=( a4346a  and  a4343a );
 a4350a <=( (not A267)  and  (not A203) );
 a4354a <=( A301  and  (not A269) );
 a4355a <=( (not A268)  and  a4354a );
 a4356a <=( a4355a  and  a4350a );
 a4359a <=( A166  and  A168 );
 a4362a <=( (not A202)  and  (not A201) );
 a4363a <=( a4362a  and  a4359a );
 a4366a <=( (not A265)  and  (not A203) );
 a4370a <=( A301  and  (not A268) );
 a4371a <=( (not A266)  and  a4370a );
 a4372a <=( a4371a  and  a4366a );
 a4375a <=( A166  and  A168 );
 a4378a <=( A201  and  A199 );
 a4379a <=( a4378a  and  a4375a );
 a4382a <=( A298  and  A268 );
 a4386a <=( (not A301)  and  (not A300) );
 a4387a <=( A299  and  a4386a );
 a4388a <=( a4387a  and  a4382a );
 a4391a <=( A166  and  A168 );
 a4394a <=( A201  and  A199 );
 a4395a <=( a4394a  and  a4391a );
 a4398a <=( A267  and  A265 );
 a4402a <=( (not A302)  and  (not A301) );
 a4403a <=( (not A300)  and  a4402a );
 a4404a <=( a4403a  and  a4398a );
 a4407a <=( A166  and  A168 );
 a4410a <=( A201  and  A199 );
 a4411a <=( a4410a  and  a4407a );
 a4414a <=( A267  and  A265 );
 a4418a <=( (not A301)  and  (not A299) );
 a4419a <=( (not A298)  and  a4418a );
 a4420a <=( a4419a  and  a4414a );
 a4423a <=( A166  and  A168 );
 a4426a <=( A201  and  A199 );
 a4427a <=( a4426a  and  a4423a );
 a4430a <=( A267  and  A266 );
 a4434a <=( (not A302)  and  (not A301) );
 a4435a <=( (not A300)  and  a4434a );
 a4436a <=( a4435a  and  a4430a );
 a4439a <=( A166  and  A168 );
 a4442a <=( A201  and  A199 );
 a4443a <=( a4442a  and  a4439a );
 a4446a <=( A267  and  A266 );
 a4450a <=( (not A301)  and  (not A299) );
 a4451a <=( (not A298)  and  a4450a );
 a4452a <=( a4451a  and  a4446a );
 a4455a <=( A166  and  A168 );
 a4458a <=( A201  and  A200 );
 a4459a <=( a4458a  and  a4455a );
 a4462a <=( A298  and  A268 );
 a4466a <=( (not A301)  and  (not A300) );
 a4467a <=( A299  and  a4466a );
 a4468a <=( a4467a  and  a4462a );
 a4471a <=( A166  and  A168 );
 a4474a <=( A201  and  A200 );
 a4475a <=( a4474a  and  a4471a );
 a4478a <=( A267  and  A265 );
 a4482a <=( (not A302)  and  (not A301) );
 a4483a <=( (not A300)  and  a4482a );
 a4484a <=( a4483a  and  a4478a );
 a4487a <=( A166  and  A168 );
 a4490a <=( A201  and  A200 );
 a4491a <=( a4490a  and  a4487a );
 a4494a <=( A267  and  A265 );
 a4498a <=( (not A301)  and  (not A299) );
 a4499a <=( (not A298)  and  a4498a );
 a4500a <=( a4499a  and  a4494a );
 a4503a <=( A166  and  A168 );
 a4506a <=( A201  and  A200 );
 a4507a <=( a4506a  and  a4503a );
 a4510a <=( A267  and  A266 );
 a4514a <=( (not A302)  and  (not A301) );
 a4515a <=( (not A300)  and  a4514a );
 a4516a <=( a4515a  and  a4510a );
 a4519a <=( A166  and  A168 );
 a4522a <=( A201  and  A200 );
 a4523a <=( a4522a  and  a4519a );
 a4526a <=( A267  and  A266 );
 a4530a <=( (not A301)  and  (not A299) );
 a4531a <=( (not A298)  and  a4530a );
 a4532a <=( a4531a  and  a4526a );
 a4535a <=( A166  and  A168 );
 a4538a <=( A200  and  (not A199) );
 a4539a <=( a4538a  and  a4535a );
 a4542a <=( A268  and  A203 );
 a4546a <=( (not A302)  and  (not A301) );
 a4547a <=( (not A300)  and  a4546a );
 a4548a <=( a4547a  and  a4542a );
 a4551a <=( A166  and  A168 );
 a4554a <=( A200  and  (not A199) );
 a4555a <=( a4554a  and  a4551a );
 a4558a <=( A268  and  A203 );
 a4562a <=( (not A301)  and  (not A299) );
 a4563a <=( (not A298)  and  a4562a );
 a4564a <=( a4563a  and  a4558a );
 a4567a <=( A166  and  A168 );
 a4570a <=( (not A200)  and  A199 );
 a4571a <=( a4570a  and  a4567a );
 a4574a <=( A268  and  A203 );
 a4578a <=( (not A302)  and  (not A301) );
 a4579a <=( (not A300)  and  a4578a );
 a4580a <=( a4579a  and  a4574a );
 a4583a <=( A166  and  A168 );
 a4586a <=( (not A200)  and  A199 );
 a4587a <=( a4586a  and  a4583a );
 a4590a <=( A268  and  A203 );
 a4594a <=( (not A301)  and  (not A299) );
 a4595a <=( (not A298)  and  a4594a );
 a4596a <=( a4595a  and  a4590a );
 a4599a <=( A166  and  A168 );
 a4602a <=( (not A200)  and  (not A199) );
 a4603a <=( a4602a  and  a4599a );
 a4606a <=( (not A267)  and  (not A202) );
 a4610a <=( A301  and  (not A269) );
 a4611a <=( (not A268)  and  a4610a );
 a4612a <=( a4611a  and  a4606a );
 a4615a <=( A166  and  A168 );
 a4618a <=( (not A200)  and  (not A199) );
 a4619a <=( a4618a  and  a4615a );
 a4622a <=( (not A265)  and  (not A202) );
 a4626a <=( A301  and  (not A268) );
 a4627a <=( (not A266)  and  a4626a );
 a4628a <=( a4627a  and  a4622a );
 a4631a <=( A167  and  A168 );
 a4634a <=( A265  and  A202 );
 a4635a <=( a4634a  and  a4631a );
 a4638a <=( A298  and  A267 );
 a4642a <=( (not A301)  and  (not A300) );
 a4643a <=( A299  and  a4642a );
 a4644a <=( a4643a  and  a4638a );
 a4647a <=( A167  and  A168 );
 a4650a <=( A266  and  A202 );
 a4651a <=( a4650a  and  a4647a );
 a4654a <=( A298  and  A267 );
 a4658a <=( (not A301)  and  (not A300) );
 a4659a <=( A299  and  a4658a );
 a4660a <=( a4659a  and  a4654a );
 a4663a <=( A167  and  A168 );
 a4666a <=( (not A265)  and  A202 );
 a4667a <=( a4666a  and  a4663a );
 a4670a <=( A269  and  A266 );
 a4674a <=( (not A302)  and  (not A301) );
 a4675a <=( (not A300)  and  a4674a );
 a4676a <=( a4675a  and  a4670a );
 a4679a <=( A167  and  A168 );
 a4682a <=( (not A265)  and  A202 );
 a4683a <=( a4682a  and  a4679a );
 a4686a <=( A269  and  A266 );
 a4690a <=( (not A301)  and  (not A299) );
 a4691a <=( (not A298)  and  a4690a );
 a4692a <=( a4691a  and  a4686a );
 a4695a <=( A167  and  A168 );
 a4698a <=( A265  and  A202 );
 a4699a <=( a4698a  and  a4695a );
 a4702a <=( A269  and  (not A266) );
 a4706a <=( (not A302)  and  (not A301) );
 a4707a <=( (not A300)  and  a4706a );
 a4708a <=( a4707a  and  a4702a );
 a4711a <=( A167  and  A168 );
 a4714a <=( A265  and  A202 );
 a4715a <=( a4714a  and  a4711a );
 a4718a <=( A269  and  (not A266) );
 a4722a <=( (not A301)  and  (not A299) );
 a4723a <=( (not A298)  and  a4722a );
 a4724a <=( a4723a  and  a4718a );
 a4727a <=( A167  and  A168 );
 a4730a <=( (not A202)  and  (not A201) );
 a4731a <=( a4730a  and  a4727a );
 a4734a <=( (not A267)  and  (not A203) );
 a4738a <=( A301  and  (not A269) );
 a4739a <=( (not A268)  and  a4738a );
 a4740a <=( a4739a  and  a4734a );
 a4743a <=( A167  and  A168 );
 a4746a <=( (not A202)  and  (not A201) );
 a4747a <=( a4746a  and  a4743a );
 a4750a <=( (not A265)  and  (not A203) );
 a4754a <=( A301  and  (not A268) );
 a4755a <=( (not A266)  and  a4754a );
 a4756a <=( a4755a  and  a4750a );
 a4759a <=( A167  and  A168 );
 a4762a <=( A201  and  A199 );
 a4763a <=( a4762a  and  a4759a );
 a4766a <=( A298  and  A268 );
 a4770a <=( (not A301)  and  (not A300) );
 a4771a <=( A299  and  a4770a );
 a4772a <=( a4771a  and  a4766a );
 a4775a <=( A167  and  A168 );
 a4778a <=( A201  and  A199 );
 a4779a <=( a4778a  and  a4775a );
 a4782a <=( A267  and  A265 );
 a4786a <=( (not A302)  and  (not A301) );
 a4787a <=( (not A300)  and  a4786a );
 a4788a <=( a4787a  and  a4782a );
 a4791a <=( A167  and  A168 );
 a4794a <=( A201  and  A199 );
 a4795a <=( a4794a  and  a4791a );
 a4798a <=( A267  and  A265 );
 a4802a <=( (not A301)  and  (not A299) );
 a4803a <=( (not A298)  and  a4802a );
 a4804a <=( a4803a  and  a4798a );
 a4807a <=( A167  and  A168 );
 a4810a <=( A201  and  A199 );
 a4811a <=( a4810a  and  a4807a );
 a4814a <=( A267  and  A266 );
 a4818a <=( (not A302)  and  (not A301) );
 a4819a <=( (not A300)  and  a4818a );
 a4820a <=( a4819a  and  a4814a );
 a4823a <=( A167  and  A168 );
 a4826a <=( A201  and  A199 );
 a4827a <=( a4826a  and  a4823a );
 a4830a <=( A267  and  A266 );
 a4834a <=( (not A301)  and  (not A299) );
 a4835a <=( (not A298)  and  a4834a );
 a4836a <=( a4835a  and  a4830a );
 a4839a <=( A167  and  A168 );
 a4842a <=( A201  and  A200 );
 a4843a <=( a4842a  and  a4839a );
 a4846a <=( A298  and  A268 );
 a4850a <=( (not A301)  and  (not A300) );
 a4851a <=( A299  and  a4850a );
 a4852a <=( a4851a  and  a4846a );
 a4855a <=( A167  and  A168 );
 a4858a <=( A201  and  A200 );
 a4859a <=( a4858a  and  a4855a );
 a4862a <=( A267  and  A265 );
 a4866a <=( (not A302)  and  (not A301) );
 a4867a <=( (not A300)  and  a4866a );
 a4868a <=( a4867a  and  a4862a );
 a4871a <=( A167  and  A168 );
 a4874a <=( A201  and  A200 );
 a4875a <=( a4874a  and  a4871a );
 a4878a <=( A267  and  A265 );
 a4882a <=( (not A301)  and  (not A299) );
 a4883a <=( (not A298)  and  a4882a );
 a4884a <=( a4883a  and  a4878a );
 a4887a <=( A167  and  A168 );
 a4890a <=( A201  and  A200 );
 a4891a <=( a4890a  and  a4887a );
 a4894a <=( A267  and  A266 );
 a4898a <=( (not A302)  and  (not A301) );
 a4899a <=( (not A300)  and  a4898a );
 a4900a <=( a4899a  and  a4894a );
 a4903a <=( A167  and  A168 );
 a4906a <=( A201  and  A200 );
 a4907a <=( a4906a  and  a4903a );
 a4910a <=( A267  and  A266 );
 a4914a <=( (not A301)  and  (not A299) );
 a4915a <=( (not A298)  and  a4914a );
 a4916a <=( a4915a  and  a4910a );
 a4919a <=( A167  and  A168 );
 a4922a <=( A200  and  (not A199) );
 a4923a <=( a4922a  and  a4919a );
 a4926a <=( A268  and  A203 );
 a4930a <=( (not A302)  and  (not A301) );
 a4931a <=( (not A300)  and  a4930a );
 a4932a <=( a4931a  and  a4926a );
 a4935a <=( A167  and  A168 );
 a4938a <=( A200  and  (not A199) );
 a4939a <=( a4938a  and  a4935a );
 a4942a <=( A268  and  A203 );
 a4946a <=( (not A301)  and  (not A299) );
 a4947a <=( (not A298)  and  a4946a );
 a4948a <=( a4947a  and  a4942a );
 a4951a <=( A167  and  A168 );
 a4954a <=( (not A200)  and  A199 );
 a4955a <=( a4954a  and  a4951a );
 a4958a <=( A268  and  A203 );
 a4962a <=( (not A302)  and  (not A301) );
 a4963a <=( (not A300)  and  a4962a );
 a4964a <=( a4963a  and  a4958a );
 a4967a <=( A167  and  A168 );
 a4970a <=( (not A200)  and  A199 );
 a4971a <=( a4970a  and  a4967a );
 a4974a <=( A268  and  A203 );
 a4978a <=( (not A301)  and  (not A299) );
 a4979a <=( (not A298)  and  a4978a );
 a4980a <=( a4979a  and  a4974a );
 a4983a <=( A167  and  A168 );
 a4986a <=( (not A200)  and  (not A199) );
 a4987a <=( a4986a  and  a4983a );
 a4990a <=( (not A267)  and  (not A202) );
 a4994a <=( A301  and  (not A269) );
 a4995a <=( (not A268)  and  a4994a );
 a4996a <=( a4995a  and  a4990a );
 a4999a <=( A167  and  A168 );
 a5002a <=( (not A200)  and  (not A199) );
 a5003a <=( a5002a  and  a4999a );
 a5006a <=( (not A265)  and  (not A202) );
 a5010a <=( A301  and  (not A268) );
 a5011a <=( (not A266)  and  a5010a );
 a5012a <=( a5011a  and  a5006a );
 a5015a <=( A167  and  A170 );
 a5018a <=( A202  and  (not A166) );
 a5019a <=( a5018a  and  a5015a );
 a5022a <=( A298  and  A268 );
 a5026a <=( (not A301)  and  (not A300) );
 a5027a <=( A299  and  a5026a );
 a5028a <=( a5027a  and  a5022a );
 a5031a <=( A167  and  A170 );
 a5034a <=( A202  and  (not A166) );
 a5035a <=( a5034a  and  a5031a );
 a5038a <=( A267  and  A265 );
 a5042a <=( (not A302)  and  (not A301) );
 a5043a <=( (not A300)  and  a5042a );
 a5044a <=( a5043a  and  a5038a );
 a5047a <=( A167  and  A170 );
 a5050a <=( A202  and  (not A166) );
 a5051a <=( a5050a  and  a5047a );
 a5054a <=( A267  and  A265 );
 a5058a <=( (not A301)  and  (not A299) );
 a5059a <=( (not A298)  and  a5058a );
 a5060a <=( a5059a  and  a5054a );
 a5063a <=( A167  and  A170 );
 a5066a <=( A202  and  (not A166) );
 a5067a <=( a5066a  and  a5063a );
 a5070a <=( A267  and  A266 );
 a5074a <=( (not A302)  and  (not A301) );
 a5075a <=( (not A300)  and  a5074a );
 a5076a <=( a5075a  and  a5070a );
 a5079a <=( A167  and  A170 );
 a5082a <=( A202  and  (not A166) );
 a5083a <=( a5082a  and  a5079a );
 a5086a <=( A267  and  A266 );
 a5090a <=( (not A301)  and  (not A299) );
 a5091a <=( (not A298)  and  a5090a );
 a5092a <=( a5091a  and  a5086a );
 a5095a <=( A167  and  A170 );
 a5098a <=( A199  and  (not A166) );
 a5099a <=( a5098a  and  a5095a );
 a5102a <=( A268  and  A201 );
 a5106a <=( (not A302)  and  (not A301) );
 a5107a <=( (not A300)  and  a5106a );
 a5108a <=( a5107a  and  a5102a );
 a5111a <=( A167  and  A170 );
 a5114a <=( A199  and  (not A166) );
 a5115a <=( a5114a  and  a5111a );
 a5118a <=( A268  and  A201 );
 a5122a <=( (not A301)  and  (not A299) );
 a5123a <=( (not A298)  and  a5122a );
 a5124a <=( a5123a  and  a5118a );
 a5127a <=( A167  and  A170 );
 a5130a <=( A200  and  (not A166) );
 a5131a <=( a5130a  and  a5127a );
 a5134a <=( A268  and  A201 );
 a5138a <=( (not A302)  and  (not A301) );
 a5139a <=( (not A300)  and  a5138a );
 a5140a <=( a5139a  and  a5134a );
 a5143a <=( A167  and  A170 );
 a5146a <=( A200  and  (not A166) );
 a5147a <=( a5146a  and  a5143a );
 a5150a <=( A268  and  A201 );
 a5154a <=( (not A301)  and  (not A299) );
 a5155a <=( (not A298)  and  a5154a );
 a5156a <=( a5155a  and  a5150a );
 a5159a <=( (not A167)  and  A170 );
 a5162a <=( A202  and  A166 );
 a5163a <=( a5162a  and  a5159a );
 a5166a <=( A298  and  A268 );
 a5170a <=( (not A301)  and  (not A300) );
 a5171a <=( A299  and  a5170a );
 a5172a <=( a5171a  and  a5166a );
 a5175a <=( (not A167)  and  A170 );
 a5178a <=( A202  and  A166 );
 a5179a <=( a5178a  and  a5175a );
 a5182a <=( A267  and  A265 );
 a5186a <=( (not A302)  and  (not A301) );
 a5187a <=( (not A300)  and  a5186a );
 a5188a <=( a5187a  and  a5182a );
 a5191a <=( (not A167)  and  A170 );
 a5194a <=( A202  and  A166 );
 a5195a <=( a5194a  and  a5191a );
 a5198a <=( A267  and  A265 );
 a5202a <=( (not A301)  and  (not A299) );
 a5203a <=( (not A298)  and  a5202a );
 a5204a <=( a5203a  and  a5198a );
 a5207a <=( (not A167)  and  A170 );
 a5210a <=( A202  and  A166 );
 a5211a <=( a5210a  and  a5207a );
 a5214a <=( A267  and  A266 );
 a5218a <=( (not A302)  and  (not A301) );
 a5219a <=( (not A300)  and  a5218a );
 a5220a <=( a5219a  and  a5214a );
 a5223a <=( (not A167)  and  A170 );
 a5226a <=( A202  and  A166 );
 a5227a <=( a5226a  and  a5223a );
 a5230a <=( A267  and  A266 );
 a5234a <=( (not A301)  and  (not A299) );
 a5235a <=( (not A298)  and  a5234a );
 a5236a <=( a5235a  and  a5230a );
 a5239a <=( (not A167)  and  A170 );
 a5242a <=( A199  and  A166 );
 a5243a <=( a5242a  and  a5239a );
 a5246a <=( A268  and  A201 );
 a5250a <=( (not A302)  and  (not A301) );
 a5251a <=( (not A300)  and  a5250a );
 a5252a <=( a5251a  and  a5246a );
 a5255a <=( (not A167)  and  A170 );
 a5258a <=( A199  and  A166 );
 a5259a <=( a5258a  and  a5255a );
 a5262a <=( A268  and  A201 );
 a5266a <=( (not A301)  and  (not A299) );
 a5267a <=( (not A298)  and  a5266a );
 a5268a <=( a5267a  and  a5262a );
 a5271a <=( (not A167)  and  A170 );
 a5274a <=( A200  and  A166 );
 a5275a <=( a5274a  and  a5271a );
 a5278a <=( A268  and  A201 );
 a5282a <=( (not A302)  and  (not A301) );
 a5283a <=( (not A300)  and  a5282a );
 a5284a <=( a5283a  and  a5278a );
 a5287a <=( (not A167)  and  A170 );
 a5290a <=( A200  and  A166 );
 a5291a <=( a5290a  and  a5287a );
 a5294a <=( A268  and  A201 );
 a5298a <=( (not A301)  and  (not A299) );
 a5299a <=( (not A298)  and  a5298a );
 a5300a <=( a5299a  and  a5294a );
 a5303a <=( A202  and  A169 );
 a5306a <=( A266  and  (not A265) );
 a5307a <=( a5306a  and  a5303a );
 a5310a <=( A298  and  A269 );
 a5314a <=( (not A301)  and  (not A300) );
 a5315a <=( A299  and  a5314a );
 a5316a <=( a5315a  and  a5310a );
 a5319a <=( A202  and  A169 );
 a5322a <=( (not A266)  and  A265 );
 a5323a <=( a5322a  and  a5319a );
 a5326a <=( A298  and  A269 );
 a5330a <=( (not A301)  and  (not A300) );
 a5331a <=( A299  and  a5330a );
 a5332a <=( a5331a  and  a5326a );
 a5335a <=( (not A201)  and  A169 );
 a5338a <=( (not A203)  and  (not A202) );
 a5339a <=( a5338a  and  a5335a );
 a5342a <=( (not A268)  and  (not A267) );
 a5346a <=( A300  and  A299 );
 a5347a <=( (not A269)  and  a5346a );
 a5348a <=( a5347a  and  a5342a );
 a5351a <=( (not A201)  and  A169 );
 a5354a <=( (not A203)  and  (not A202) );
 a5355a <=( a5354a  and  a5351a );
 a5358a <=( (not A268)  and  (not A267) );
 a5362a <=( A300  and  A298 );
 a5363a <=( (not A269)  and  a5362a );
 a5364a <=( a5363a  and  a5358a );
 a5367a <=( (not A201)  and  A169 );
 a5370a <=( (not A203)  and  (not A202) );
 a5371a <=( a5370a  and  a5367a );
 a5374a <=( A266  and  A265 );
 a5378a <=( A301  and  (not A268) );
 a5379a <=( (not A267)  and  a5378a );
 a5380a <=( a5379a  and  a5374a );
 a5383a <=( (not A201)  and  A169 );
 a5386a <=( (not A203)  and  (not A202) );
 a5387a <=( a5386a  and  a5383a );
 a5390a <=( (not A266)  and  (not A265) );
 a5394a <=( A300  and  A299 );
 a5395a <=( (not A268)  and  a5394a );
 a5396a <=( a5395a  and  a5390a );
 a5399a <=( (not A201)  and  A169 );
 a5402a <=( (not A203)  and  (not A202) );
 a5403a <=( a5402a  and  a5399a );
 a5406a <=( (not A266)  and  (not A265) );
 a5410a <=( A300  and  A298 );
 a5411a <=( (not A268)  and  a5410a );
 a5412a <=( a5411a  and  a5406a );
 a5415a <=( A199  and  A169 );
 a5418a <=( A265  and  A201 );
 a5419a <=( a5418a  and  a5415a );
 a5422a <=( A298  and  A267 );
 a5426a <=( (not A301)  and  (not A300) );
 a5427a <=( A299  and  a5426a );
 a5428a <=( a5427a  and  a5422a );
 a5431a <=( A199  and  A169 );
 a5434a <=( A266  and  A201 );
 a5435a <=( a5434a  and  a5431a );
 a5438a <=( A298  and  A267 );
 a5442a <=( (not A301)  and  (not A300) );
 a5443a <=( A299  and  a5442a );
 a5444a <=( a5443a  and  a5438a );
 a5447a <=( A199  and  A169 );
 a5450a <=( (not A265)  and  A201 );
 a5451a <=( a5450a  and  a5447a );
 a5454a <=( A269  and  A266 );
 a5458a <=( (not A302)  and  (not A301) );
 a5459a <=( (not A300)  and  a5458a );
 a5460a <=( a5459a  and  a5454a );
 a5463a <=( A199  and  A169 );
 a5466a <=( (not A265)  and  A201 );
 a5467a <=( a5466a  and  a5463a );
 a5470a <=( A269  and  A266 );
 a5474a <=( (not A301)  and  (not A299) );
 a5475a <=( (not A298)  and  a5474a );
 a5476a <=( a5475a  and  a5470a );
 a5479a <=( A199  and  A169 );
 a5482a <=( A265  and  A201 );
 a5483a <=( a5482a  and  a5479a );
 a5486a <=( A269  and  (not A266) );
 a5490a <=( (not A302)  and  (not A301) );
 a5491a <=( (not A300)  and  a5490a );
 a5492a <=( a5491a  and  a5486a );
 a5495a <=( A199  and  A169 );
 a5498a <=( A265  and  A201 );
 a5499a <=( a5498a  and  a5495a );
 a5502a <=( A269  and  (not A266) );
 a5506a <=( (not A301)  and  (not A299) );
 a5507a <=( (not A298)  and  a5506a );
 a5508a <=( a5507a  and  a5502a );
 a5511a <=( A200  and  A169 );
 a5514a <=( A265  and  A201 );
 a5515a <=( a5514a  and  a5511a );
 a5518a <=( A298  and  A267 );
 a5522a <=( (not A301)  and  (not A300) );
 a5523a <=( A299  and  a5522a );
 a5524a <=( a5523a  and  a5518a );
 a5527a <=( A200  and  A169 );
 a5530a <=( A266  and  A201 );
 a5531a <=( a5530a  and  a5527a );
 a5534a <=( A298  and  A267 );
 a5538a <=( (not A301)  and  (not A300) );
 a5539a <=( A299  and  a5538a );
 a5540a <=( a5539a  and  a5534a );
 a5543a <=( A200  and  A169 );
 a5546a <=( (not A265)  and  A201 );
 a5547a <=( a5546a  and  a5543a );
 a5550a <=( A269  and  A266 );
 a5554a <=( (not A302)  and  (not A301) );
 a5555a <=( (not A300)  and  a5554a );
 a5556a <=( a5555a  and  a5550a );
 a5559a <=( A200  and  A169 );
 a5562a <=( (not A265)  and  A201 );
 a5563a <=( a5562a  and  a5559a );
 a5566a <=( A269  and  A266 );
 a5570a <=( (not A301)  and  (not A299) );
 a5571a <=( (not A298)  and  a5570a );
 a5572a <=( a5571a  and  a5566a );
 a5575a <=( A200  and  A169 );
 a5578a <=( A265  and  A201 );
 a5579a <=( a5578a  and  a5575a );
 a5582a <=( A269  and  (not A266) );
 a5586a <=( (not A302)  and  (not A301) );
 a5587a <=( (not A300)  and  a5586a );
 a5588a <=( a5587a  and  a5582a );
 a5591a <=( A200  and  A169 );
 a5594a <=( A265  and  A201 );
 a5595a <=( a5594a  and  a5591a );
 a5598a <=( A269  and  (not A266) );
 a5602a <=( (not A301)  and  (not A299) );
 a5603a <=( (not A298)  and  a5602a );
 a5604a <=( a5603a  and  a5598a );
 a5607a <=( A199  and  A169 );
 a5610a <=( (not A201)  and  A200 );
 a5611a <=( a5610a  and  a5607a );
 a5614a <=( (not A267)  and  (not A202) );
 a5618a <=( A301  and  (not A269) );
 a5619a <=( (not A268)  and  a5618a );
 a5620a <=( a5619a  and  a5614a );
 a5623a <=( A199  and  A169 );
 a5626a <=( (not A201)  and  A200 );
 a5627a <=( a5626a  and  a5623a );
 a5630a <=( (not A265)  and  (not A202) );
 a5634a <=( A301  and  (not A268) );
 a5635a <=( (not A266)  and  a5634a );
 a5636a <=( a5635a  and  a5630a );
 a5639a <=( (not A199)  and  A169 );
 a5642a <=( A203  and  A200 );
 a5643a <=( a5642a  and  a5639a );
 a5646a <=( A298  and  A268 );
 a5650a <=( (not A301)  and  (not A300) );
 a5651a <=( A299  and  a5650a );
 a5652a <=( a5651a  and  a5646a );
 a5655a <=( (not A199)  and  A169 );
 a5658a <=( A203  and  A200 );
 a5659a <=( a5658a  and  a5655a );
 a5662a <=( A267  and  A265 );
 a5666a <=( (not A302)  and  (not A301) );
 a5667a <=( (not A300)  and  a5666a );
 a5668a <=( a5667a  and  a5662a );
 a5671a <=( (not A199)  and  A169 );
 a5674a <=( A203  and  A200 );
 a5675a <=( a5674a  and  a5671a );
 a5678a <=( A267  and  A265 );
 a5682a <=( (not A301)  and  (not A299) );
 a5683a <=( (not A298)  and  a5682a );
 a5684a <=( a5683a  and  a5678a );
 a5687a <=( (not A199)  and  A169 );
 a5690a <=( A203  and  A200 );
 a5691a <=( a5690a  and  a5687a );
 a5694a <=( A267  and  A266 );
 a5698a <=( (not A302)  and  (not A301) );
 a5699a <=( (not A300)  and  a5698a );
 a5700a <=( a5699a  and  a5694a );
 a5703a <=( (not A199)  and  A169 );
 a5706a <=( A203  and  A200 );
 a5707a <=( a5706a  and  a5703a );
 a5710a <=( A267  and  A266 );
 a5714a <=( (not A301)  and  (not A299) );
 a5715a <=( (not A298)  and  a5714a );
 a5716a <=( a5715a  and  a5710a );
 a5719a <=( A199  and  A169 );
 a5722a <=( A203  and  (not A200) );
 a5723a <=( a5722a  and  a5719a );
 a5726a <=( A298  and  A268 );
 a5730a <=( (not A301)  and  (not A300) );
 a5731a <=( A299  and  a5730a );
 a5732a <=( a5731a  and  a5726a );
 a5735a <=( A199  and  A169 );
 a5738a <=( A203  and  (not A200) );
 a5739a <=( a5738a  and  a5735a );
 a5742a <=( A267  and  A265 );
 a5746a <=( (not A302)  and  (not A301) );
 a5747a <=( (not A300)  and  a5746a );
 a5748a <=( a5747a  and  a5742a );
 a5751a <=( A199  and  A169 );
 a5754a <=( A203  and  (not A200) );
 a5755a <=( a5754a  and  a5751a );
 a5758a <=( A267  and  A265 );
 a5762a <=( (not A301)  and  (not A299) );
 a5763a <=( (not A298)  and  a5762a );
 a5764a <=( a5763a  and  a5758a );
 a5767a <=( A199  and  A169 );
 a5770a <=( A203  and  (not A200) );
 a5771a <=( a5770a  and  a5767a );
 a5774a <=( A267  and  A266 );
 a5778a <=( (not A302)  and  (not A301) );
 a5779a <=( (not A300)  and  a5778a );
 a5780a <=( a5779a  and  a5774a );
 a5783a <=( A199  and  A169 );
 a5786a <=( A203  and  (not A200) );
 a5787a <=( a5786a  and  a5783a );
 a5790a <=( A267  and  A266 );
 a5794a <=( (not A301)  and  (not A299) );
 a5795a <=( (not A298)  and  a5794a );
 a5796a <=( a5795a  and  a5790a );
 a5799a <=( (not A199)  and  A169 );
 a5802a <=( (not A202)  and  (not A200) );
 a5803a <=( a5802a  and  a5799a );
 a5806a <=( (not A268)  and  (not A267) );
 a5810a <=( A300  and  A299 );
 a5811a <=( (not A269)  and  a5810a );
 a5812a <=( a5811a  and  a5806a );
 a5815a <=( (not A199)  and  A169 );
 a5818a <=( (not A202)  and  (not A200) );
 a5819a <=( a5818a  and  a5815a );
 a5822a <=( (not A268)  and  (not A267) );
 a5826a <=( A300  and  A298 );
 a5827a <=( (not A269)  and  a5826a );
 a5828a <=( a5827a  and  a5822a );
 a5831a <=( (not A199)  and  A169 );
 a5834a <=( (not A202)  and  (not A200) );
 a5835a <=( a5834a  and  a5831a );
 a5838a <=( A266  and  A265 );
 a5842a <=( A301  and  (not A268) );
 a5843a <=( (not A267)  and  a5842a );
 a5844a <=( a5843a  and  a5838a );
 a5847a <=( (not A199)  and  A169 );
 a5850a <=( (not A202)  and  (not A200) );
 a5851a <=( a5850a  and  a5847a );
 a5854a <=( (not A266)  and  (not A265) );
 a5858a <=( A300  and  A299 );
 a5859a <=( (not A268)  and  a5858a );
 a5860a <=( a5859a  and  a5854a );
 a5863a <=( (not A199)  and  A169 );
 a5866a <=( (not A202)  and  (not A200) );
 a5867a <=( a5866a  and  a5863a );
 a5870a <=( (not A266)  and  (not A265) );
 a5874a <=( A300  and  A298 );
 a5875a <=( (not A268)  and  a5874a );
 a5876a <=( a5875a  and  a5870a );
 a5879a <=( (not A167)  and  (not A169) );
 a5882a <=( A202  and  (not A166) );
 a5883a <=( a5882a  and  a5879a );
 a5886a <=( (not A268)  and  (not A267) );
 a5890a <=( A300  and  A299 );
 a5891a <=( (not A269)  and  a5890a );
 a5892a <=( a5891a  and  a5886a );
 a5895a <=( (not A167)  and  (not A169) );
 a5898a <=( A202  and  (not A166) );
 a5899a <=( a5898a  and  a5895a );
 a5902a <=( (not A268)  and  (not A267) );
 a5906a <=( A300  and  A298 );
 a5907a <=( (not A269)  and  a5906a );
 a5908a <=( a5907a  and  a5902a );
 a5911a <=( (not A167)  and  (not A169) );
 a5914a <=( A202  and  (not A166) );
 a5915a <=( a5914a  and  a5911a );
 a5918a <=( A266  and  A265 );
 a5922a <=( A301  and  (not A268) );
 a5923a <=( (not A267)  and  a5922a );
 a5924a <=( a5923a  and  a5918a );
 a5927a <=( (not A167)  and  (not A169) );
 a5930a <=( A202  and  (not A166) );
 a5931a <=( a5930a  and  a5927a );
 a5934a <=( (not A266)  and  (not A265) );
 a5938a <=( A300  and  A299 );
 a5939a <=( (not A268)  and  a5938a );
 a5940a <=( a5939a  and  a5934a );
 a5943a <=( (not A167)  and  (not A169) );
 a5946a <=( A202  and  (not A166) );
 a5947a <=( a5946a  and  a5943a );
 a5950a <=( (not A266)  and  (not A265) );
 a5954a <=( A300  and  A298 );
 a5955a <=( (not A268)  and  a5954a );
 a5956a <=( a5955a  and  a5950a );
 a5959a <=( (not A167)  and  (not A169) );
 a5962a <=( A199  and  (not A166) );
 a5963a <=( a5962a  and  a5959a );
 a5966a <=( (not A267)  and  A201 );
 a5970a <=( A301  and  (not A269) );
 a5971a <=( (not A268)  and  a5970a );
 a5972a <=( a5971a  and  a5966a );
 a5975a <=( (not A167)  and  (not A169) );
 a5978a <=( A199  and  (not A166) );
 a5979a <=( a5978a  and  a5975a );
 a5982a <=( (not A265)  and  A201 );
 a5986a <=( A301  and  (not A268) );
 a5987a <=( (not A266)  and  a5986a );
 a5988a <=( a5987a  and  a5982a );
 a5991a <=( (not A167)  and  (not A169) );
 a5994a <=( A200  and  (not A166) );
 a5995a <=( a5994a  and  a5991a );
 a5998a <=( (not A267)  and  A201 );
 a6002a <=( A301  and  (not A269) );
 a6003a <=( (not A268)  and  a6002a );
 a6004a <=( a6003a  and  a5998a );
 a6007a <=( (not A167)  and  (not A169) );
 a6010a <=( A200  and  (not A166) );
 a6011a <=( a6010a  and  a6007a );
 a6014a <=( (not A265)  and  A201 );
 a6018a <=( A301  and  (not A268) );
 a6019a <=( (not A266)  and  a6018a );
 a6020a <=( a6019a  and  a6014a );
 a6023a <=( (not A168)  and  (not A169) );
 a6026a <=( A166  and  A167 );
 a6027a <=( a6026a  and  a6023a );
 a6030a <=( (not A267)  and  A202 );
 a6034a <=( A301  and  (not A269) );
 a6035a <=( (not A268)  and  a6034a );
 a6036a <=( a6035a  and  a6030a );
 a6039a <=( (not A168)  and  (not A169) );
 a6042a <=( A166  and  A167 );
 a6043a <=( a6042a  and  a6039a );
 a6046a <=( (not A265)  and  A202 );
 a6050a <=( A301  and  (not A268) );
 a6051a <=( (not A266)  and  a6050a );
 a6052a <=( a6051a  and  a6046a );
 a6055a <=( (not A169)  and  (not A170) );
 a6058a <=( A202  and  (not A168) );
 a6059a <=( a6058a  and  a6055a );
 a6062a <=( (not A268)  and  (not A267) );
 a6066a <=( A300  and  A299 );
 a6067a <=( (not A269)  and  a6066a );
 a6068a <=( a6067a  and  a6062a );
 a6071a <=( (not A169)  and  (not A170) );
 a6074a <=( A202  and  (not A168) );
 a6075a <=( a6074a  and  a6071a );
 a6078a <=( (not A268)  and  (not A267) );
 a6082a <=( A300  and  A298 );
 a6083a <=( (not A269)  and  a6082a );
 a6084a <=( a6083a  and  a6078a );
 a6087a <=( (not A169)  and  (not A170) );
 a6090a <=( A202  and  (not A168) );
 a6091a <=( a6090a  and  a6087a );
 a6094a <=( A266  and  A265 );
 a6098a <=( A301  and  (not A268) );
 a6099a <=( (not A267)  and  a6098a );
 a6100a <=( a6099a  and  a6094a );
 a6103a <=( (not A169)  and  (not A170) );
 a6106a <=( A202  and  (not A168) );
 a6107a <=( a6106a  and  a6103a );
 a6110a <=( (not A266)  and  (not A265) );
 a6114a <=( A300  and  A299 );
 a6115a <=( (not A268)  and  a6114a );
 a6116a <=( a6115a  and  a6110a );
 a6119a <=( (not A169)  and  (not A170) );
 a6122a <=( A202  and  (not A168) );
 a6123a <=( a6122a  and  a6119a );
 a6126a <=( (not A266)  and  (not A265) );
 a6130a <=( A300  and  A298 );
 a6131a <=( (not A268)  and  a6130a );
 a6132a <=( a6131a  and  a6126a );
 a6135a <=( (not A169)  and  (not A170) );
 a6138a <=( A199  and  (not A168) );
 a6139a <=( a6138a  and  a6135a );
 a6142a <=( (not A267)  and  A201 );
 a6146a <=( A301  and  (not A269) );
 a6147a <=( (not A268)  and  a6146a );
 a6148a <=( a6147a  and  a6142a );
 a6151a <=( (not A169)  and  (not A170) );
 a6154a <=( A199  and  (not A168) );
 a6155a <=( a6154a  and  a6151a );
 a6158a <=( (not A265)  and  A201 );
 a6162a <=( A301  and  (not A268) );
 a6163a <=( (not A266)  and  a6162a );
 a6164a <=( a6163a  and  a6158a );
 a6167a <=( (not A169)  and  (not A170) );
 a6170a <=( A200  and  (not A168) );
 a6171a <=( a6170a  and  a6167a );
 a6174a <=( (not A267)  and  A201 );
 a6178a <=( A301  and  (not A269) );
 a6179a <=( (not A268)  and  a6178a );
 a6180a <=( a6179a  and  a6174a );
 a6183a <=( (not A169)  and  (not A170) );
 a6186a <=( A200  and  (not A168) );
 a6187a <=( a6186a  and  a6183a );
 a6190a <=( (not A265)  and  A201 );
 a6194a <=( A301  and  (not A268) );
 a6195a <=( (not A266)  and  a6194a );
 a6196a <=( a6195a  and  a6190a );
 a6199a <=( A166  and  A168 );
 a6203a <=( A266  and  (not A265) );
 a6204a <=( A202  and  a6203a );
 a6205a <=( a6204a  and  a6199a );
 a6208a <=( A298  and  A269 );
 a6212a <=( (not A301)  and  (not A300) );
 a6213a <=( A299  and  a6212a );
 a6214a <=( a6213a  and  a6208a );
 a6217a <=( A166  and  A168 );
 a6221a <=( (not A266)  and  A265 );
 a6222a <=( A202  and  a6221a );
 a6223a <=( a6222a  and  a6217a );
 a6226a <=( A298  and  A269 );
 a6230a <=( (not A301)  and  (not A300) );
 a6231a <=( A299  and  a6230a );
 a6232a <=( a6231a  and  a6226a );
 a6235a <=( A166  and  A168 );
 a6239a <=( (not A203)  and  (not A202) );
 a6240a <=( (not A201)  and  a6239a );
 a6241a <=( a6240a  and  a6235a );
 a6244a <=( (not A268)  and  (not A267) );
 a6248a <=( A300  and  A299 );
 a6249a <=( (not A269)  and  a6248a );
 a6250a <=( a6249a  and  a6244a );
 a6253a <=( A166  and  A168 );
 a6257a <=( (not A203)  and  (not A202) );
 a6258a <=( (not A201)  and  a6257a );
 a6259a <=( a6258a  and  a6253a );
 a6262a <=( (not A268)  and  (not A267) );
 a6266a <=( A300  and  A298 );
 a6267a <=( (not A269)  and  a6266a );
 a6268a <=( a6267a  and  a6262a );
 a6271a <=( A166  and  A168 );
 a6275a <=( (not A203)  and  (not A202) );
 a6276a <=( (not A201)  and  a6275a );
 a6277a <=( a6276a  and  a6271a );
 a6280a <=( A266  and  A265 );
 a6284a <=( A301  and  (not A268) );
 a6285a <=( (not A267)  and  a6284a );
 a6286a <=( a6285a  and  a6280a );
 a6289a <=( A166  and  A168 );
 a6293a <=( (not A203)  and  (not A202) );
 a6294a <=( (not A201)  and  a6293a );
 a6295a <=( a6294a  and  a6289a );
 a6298a <=( (not A266)  and  (not A265) );
 a6302a <=( A300  and  A299 );
 a6303a <=( (not A268)  and  a6302a );
 a6304a <=( a6303a  and  a6298a );
 a6307a <=( A166  and  A168 );
 a6311a <=( (not A203)  and  (not A202) );
 a6312a <=( (not A201)  and  a6311a );
 a6313a <=( a6312a  and  a6307a );
 a6316a <=( (not A266)  and  (not A265) );
 a6320a <=( A300  and  A298 );
 a6321a <=( (not A268)  and  a6320a );
 a6322a <=( a6321a  and  a6316a );
 a6325a <=( A166  and  A168 );
 a6329a <=( A265  and  A201 );
 a6330a <=( A199  and  a6329a );
 a6331a <=( a6330a  and  a6325a );
 a6334a <=( A298  and  A267 );
 a6338a <=( (not A301)  and  (not A300) );
 a6339a <=( A299  and  a6338a );
 a6340a <=( a6339a  and  a6334a );
 a6343a <=( A166  and  A168 );
 a6347a <=( A266  and  A201 );
 a6348a <=( A199  and  a6347a );
 a6349a <=( a6348a  and  a6343a );
 a6352a <=( A298  and  A267 );
 a6356a <=( (not A301)  and  (not A300) );
 a6357a <=( A299  and  a6356a );
 a6358a <=( a6357a  and  a6352a );
 a6361a <=( A166  and  A168 );
 a6365a <=( (not A265)  and  A201 );
 a6366a <=( A199  and  a6365a );
 a6367a <=( a6366a  and  a6361a );
 a6370a <=( A269  and  A266 );
 a6374a <=( (not A302)  and  (not A301) );
 a6375a <=( (not A300)  and  a6374a );
 a6376a <=( a6375a  and  a6370a );
 a6379a <=( A166  and  A168 );
 a6383a <=( (not A265)  and  A201 );
 a6384a <=( A199  and  a6383a );
 a6385a <=( a6384a  and  a6379a );
 a6388a <=( A269  and  A266 );
 a6392a <=( (not A301)  and  (not A299) );
 a6393a <=( (not A298)  and  a6392a );
 a6394a <=( a6393a  and  a6388a );
 a6397a <=( A166  and  A168 );
 a6401a <=( A265  and  A201 );
 a6402a <=( A199  and  a6401a );
 a6403a <=( a6402a  and  a6397a );
 a6406a <=( A269  and  (not A266) );
 a6410a <=( (not A302)  and  (not A301) );
 a6411a <=( (not A300)  and  a6410a );
 a6412a <=( a6411a  and  a6406a );
 a6415a <=( A166  and  A168 );
 a6419a <=( A265  and  A201 );
 a6420a <=( A199  and  a6419a );
 a6421a <=( a6420a  and  a6415a );
 a6424a <=( A269  and  (not A266) );
 a6428a <=( (not A301)  and  (not A299) );
 a6429a <=( (not A298)  and  a6428a );
 a6430a <=( a6429a  and  a6424a );
 a6433a <=( A166  and  A168 );
 a6437a <=( A265  and  A201 );
 a6438a <=( A200  and  a6437a );
 a6439a <=( a6438a  and  a6433a );
 a6442a <=( A298  and  A267 );
 a6446a <=( (not A301)  and  (not A300) );
 a6447a <=( A299  and  a6446a );
 a6448a <=( a6447a  and  a6442a );
 a6451a <=( A166  and  A168 );
 a6455a <=( A266  and  A201 );
 a6456a <=( A200  and  a6455a );
 a6457a <=( a6456a  and  a6451a );
 a6460a <=( A298  and  A267 );
 a6464a <=( (not A301)  and  (not A300) );
 a6465a <=( A299  and  a6464a );
 a6466a <=( a6465a  and  a6460a );
 a6469a <=( A166  and  A168 );
 a6473a <=( (not A265)  and  A201 );
 a6474a <=( A200  and  a6473a );
 a6475a <=( a6474a  and  a6469a );
 a6478a <=( A269  and  A266 );
 a6482a <=( (not A302)  and  (not A301) );
 a6483a <=( (not A300)  and  a6482a );
 a6484a <=( a6483a  and  a6478a );
 a6487a <=( A166  and  A168 );
 a6491a <=( (not A265)  and  A201 );
 a6492a <=( A200  and  a6491a );
 a6493a <=( a6492a  and  a6487a );
 a6496a <=( A269  and  A266 );
 a6500a <=( (not A301)  and  (not A299) );
 a6501a <=( (not A298)  and  a6500a );
 a6502a <=( a6501a  and  a6496a );
 a6505a <=( A166  and  A168 );
 a6509a <=( A265  and  A201 );
 a6510a <=( A200  and  a6509a );
 a6511a <=( a6510a  and  a6505a );
 a6514a <=( A269  and  (not A266) );
 a6518a <=( (not A302)  and  (not A301) );
 a6519a <=( (not A300)  and  a6518a );
 a6520a <=( a6519a  and  a6514a );
 a6523a <=( A166  and  A168 );
 a6527a <=( A265  and  A201 );
 a6528a <=( A200  and  a6527a );
 a6529a <=( a6528a  and  a6523a );
 a6532a <=( A269  and  (not A266) );
 a6536a <=( (not A301)  and  (not A299) );
 a6537a <=( (not A298)  and  a6536a );
 a6538a <=( a6537a  and  a6532a );
 a6541a <=( A166  and  A168 );
 a6545a <=( (not A201)  and  A200 );
 a6546a <=( A199  and  a6545a );
 a6547a <=( a6546a  and  a6541a );
 a6550a <=( (not A267)  and  (not A202) );
 a6554a <=( A301  and  (not A269) );
 a6555a <=( (not A268)  and  a6554a );
 a6556a <=( a6555a  and  a6550a );
 a6559a <=( A166  and  A168 );
 a6563a <=( (not A201)  and  A200 );
 a6564a <=( A199  and  a6563a );
 a6565a <=( a6564a  and  a6559a );
 a6568a <=( (not A265)  and  (not A202) );
 a6572a <=( A301  and  (not A268) );
 a6573a <=( (not A266)  and  a6572a );
 a6574a <=( a6573a  and  a6568a );
 a6577a <=( A166  and  A168 );
 a6581a <=( A203  and  A200 );
 a6582a <=( (not A199)  and  a6581a );
 a6583a <=( a6582a  and  a6577a );
 a6586a <=( A298  and  A268 );
 a6590a <=( (not A301)  and  (not A300) );
 a6591a <=( A299  and  a6590a );
 a6592a <=( a6591a  and  a6586a );
 a6595a <=( A166  and  A168 );
 a6599a <=( A203  and  A200 );
 a6600a <=( (not A199)  and  a6599a );
 a6601a <=( a6600a  and  a6595a );
 a6604a <=( A267  and  A265 );
 a6608a <=( (not A302)  and  (not A301) );
 a6609a <=( (not A300)  and  a6608a );
 a6610a <=( a6609a  and  a6604a );
 a6613a <=( A166  and  A168 );
 a6617a <=( A203  and  A200 );
 a6618a <=( (not A199)  and  a6617a );
 a6619a <=( a6618a  and  a6613a );
 a6622a <=( A267  and  A265 );
 a6626a <=( (not A301)  and  (not A299) );
 a6627a <=( (not A298)  and  a6626a );
 a6628a <=( a6627a  and  a6622a );
 a6631a <=( A166  and  A168 );
 a6635a <=( A203  and  A200 );
 a6636a <=( (not A199)  and  a6635a );
 a6637a <=( a6636a  and  a6631a );
 a6640a <=( A267  and  A266 );
 a6644a <=( (not A302)  and  (not A301) );
 a6645a <=( (not A300)  and  a6644a );
 a6646a <=( a6645a  and  a6640a );
 a6649a <=( A166  and  A168 );
 a6653a <=( A203  and  A200 );
 a6654a <=( (not A199)  and  a6653a );
 a6655a <=( a6654a  and  a6649a );
 a6658a <=( A267  and  A266 );
 a6662a <=( (not A301)  and  (not A299) );
 a6663a <=( (not A298)  and  a6662a );
 a6664a <=( a6663a  and  a6658a );
 a6667a <=( A166  and  A168 );
 a6671a <=( A203  and  (not A200) );
 a6672a <=( A199  and  a6671a );
 a6673a <=( a6672a  and  a6667a );
 a6676a <=( A298  and  A268 );
 a6680a <=( (not A301)  and  (not A300) );
 a6681a <=( A299  and  a6680a );
 a6682a <=( a6681a  and  a6676a );
 a6685a <=( A166  and  A168 );
 a6689a <=( A203  and  (not A200) );
 a6690a <=( A199  and  a6689a );
 a6691a <=( a6690a  and  a6685a );
 a6694a <=( A267  and  A265 );
 a6698a <=( (not A302)  and  (not A301) );
 a6699a <=( (not A300)  and  a6698a );
 a6700a <=( a6699a  and  a6694a );
 a6703a <=( A166  and  A168 );
 a6707a <=( A203  and  (not A200) );
 a6708a <=( A199  and  a6707a );
 a6709a <=( a6708a  and  a6703a );
 a6712a <=( A267  and  A265 );
 a6716a <=( (not A301)  and  (not A299) );
 a6717a <=( (not A298)  and  a6716a );
 a6718a <=( a6717a  and  a6712a );
 a6721a <=( A166  and  A168 );
 a6725a <=( A203  and  (not A200) );
 a6726a <=( A199  and  a6725a );
 a6727a <=( a6726a  and  a6721a );
 a6730a <=( A267  and  A266 );
 a6734a <=( (not A302)  and  (not A301) );
 a6735a <=( (not A300)  and  a6734a );
 a6736a <=( a6735a  and  a6730a );
 a6739a <=( A166  and  A168 );
 a6743a <=( A203  and  (not A200) );
 a6744a <=( A199  and  a6743a );
 a6745a <=( a6744a  and  a6739a );
 a6748a <=( A267  and  A266 );
 a6752a <=( (not A301)  and  (not A299) );
 a6753a <=( (not A298)  and  a6752a );
 a6754a <=( a6753a  and  a6748a );
 a6757a <=( A166  and  A168 );
 a6761a <=( (not A202)  and  (not A200) );
 a6762a <=( (not A199)  and  a6761a );
 a6763a <=( a6762a  and  a6757a );
 a6766a <=( (not A268)  and  (not A267) );
 a6770a <=( A300  and  A299 );
 a6771a <=( (not A269)  and  a6770a );
 a6772a <=( a6771a  and  a6766a );
 a6775a <=( A166  and  A168 );
 a6779a <=( (not A202)  and  (not A200) );
 a6780a <=( (not A199)  and  a6779a );
 a6781a <=( a6780a  and  a6775a );
 a6784a <=( (not A268)  and  (not A267) );
 a6788a <=( A300  and  A298 );
 a6789a <=( (not A269)  and  a6788a );
 a6790a <=( a6789a  and  a6784a );
 a6793a <=( A166  and  A168 );
 a6797a <=( (not A202)  and  (not A200) );
 a6798a <=( (not A199)  and  a6797a );
 a6799a <=( a6798a  and  a6793a );
 a6802a <=( A266  and  A265 );
 a6806a <=( A301  and  (not A268) );
 a6807a <=( (not A267)  and  a6806a );
 a6808a <=( a6807a  and  a6802a );
 a6811a <=( A166  and  A168 );
 a6815a <=( (not A202)  and  (not A200) );
 a6816a <=( (not A199)  and  a6815a );
 a6817a <=( a6816a  and  a6811a );
 a6820a <=( (not A266)  and  (not A265) );
 a6824a <=( A300  and  A299 );
 a6825a <=( (not A268)  and  a6824a );
 a6826a <=( a6825a  and  a6820a );
 a6829a <=( A166  and  A168 );
 a6833a <=( (not A202)  and  (not A200) );
 a6834a <=( (not A199)  and  a6833a );
 a6835a <=( a6834a  and  a6829a );
 a6838a <=( (not A266)  and  (not A265) );
 a6842a <=( A300  and  A298 );
 a6843a <=( (not A268)  and  a6842a );
 a6844a <=( a6843a  and  a6838a );
 a6847a <=( A167  and  A168 );
 a6851a <=( A266  and  (not A265) );
 a6852a <=( A202  and  a6851a );
 a6853a <=( a6852a  and  a6847a );
 a6856a <=( A298  and  A269 );
 a6860a <=( (not A301)  and  (not A300) );
 a6861a <=( A299  and  a6860a );
 a6862a <=( a6861a  and  a6856a );
 a6865a <=( A167  and  A168 );
 a6869a <=( (not A266)  and  A265 );
 a6870a <=( A202  and  a6869a );
 a6871a <=( a6870a  and  a6865a );
 a6874a <=( A298  and  A269 );
 a6878a <=( (not A301)  and  (not A300) );
 a6879a <=( A299  and  a6878a );
 a6880a <=( a6879a  and  a6874a );
 a6883a <=( A167  and  A168 );
 a6887a <=( (not A203)  and  (not A202) );
 a6888a <=( (not A201)  and  a6887a );
 a6889a <=( a6888a  and  a6883a );
 a6892a <=( (not A268)  and  (not A267) );
 a6896a <=( A300  and  A299 );
 a6897a <=( (not A269)  and  a6896a );
 a6898a <=( a6897a  and  a6892a );
 a6901a <=( A167  and  A168 );
 a6905a <=( (not A203)  and  (not A202) );
 a6906a <=( (not A201)  and  a6905a );
 a6907a <=( a6906a  and  a6901a );
 a6910a <=( (not A268)  and  (not A267) );
 a6914a <=( A300  and  A298 );
 a6915a <=( (not A269)  and  a6914a );
 a6916a <=( a6915a  and  a6910a );
 a6919a <=( A167  and  A168 );
 a6923a <=( (not A203)  and  (not A202) );
 a6924a <=( (not A201)  and  a6923a );
 a6925a <=( a6924a  and  a6919a );
 a6928a <=( A266  and  A265 );
 a6932a <=( A301  and  (not A268) );
 a6933a <=( (not A267)  and  a6932a );
 a6934a <=( a6933a  and  a6928a );
 a6937a <=( A167  and  A168 );
 a6941a <=( (not A203)  and  (not A202) );
 a6942a <=( (not A201)  and  a6941a );
 a6943a <=( a6942a  and  a6937a );
 a6946a <=( (not A266)  and  (not A265) );
 a6950a <=( A300  and  A299 );
 a6951a <=( (not A268)  and  a6950a );
 a6952a <=( a6951a  and  a6946a );
 a6955a <=( A167  and  A168 );
 a6959a <=( (not A203)  and  (not A202) );
 a6960a <=( (not A201)  and  a6959a );
 a6961a <=( a6960a  and  a6955a );
 a6964a <=( (not A266)  and  (not A265) );
 a6968a <=( A300  and  A298 );
 a6969a <=( (not A268)  and  a6968a );
 a6970a <=( a6969a  and  a6964a );
 a6973a <=( A167  and  A168 );
 a6977a <=( A265  and  A201 );
 a6978a <=( A199  and  a6977a );
 a6979a <=( a6978a  and  a6973a );
 a6982a <=( A298  and  A267 );
 a6986a <=( (not A301)  and  (not A300) );
 a6987a <=( A299  and  a6986a );
 a6988a <=( a6987a  and  a6982a );
 a6991a <=( A167  and  A168 );
 a6995a <=( A266  and  A201 );
 a6996a <=( A199  and  a6995a );
 a6997a <=( a6996a  and  a6991a );
 a7000a <=( A298  and  A267 );
 a7004a <=( (not A301)  and  (not A300) );
 a7005a <=( A299  and  a7004a );
 a7006a <=( a7005a  and  a7000a );
 a7009a <=( A167  and  A168 );
 a7013a <=( (not A265)  and  A201 );
 a7014a <=( A199  and  a7013a );
 a7015a <=( a7014a  and  a7009a );
 a7018a <=( A269  and  A266 );
 a7022a <=( (not A302)  and  (not A301) );
 a7023a <=( (not A300)  and  a7022a );
 a7024a <=( a7023a  and  a7018a );
 a7027a <=( A167  and  A168 );
 a7031a <=( (not A265)  and  A201 );
 a7032a <=( A199  and  a7031a );
 a7033a <=( a7032a  and  a7027a );
 a7036a <=( A269  and  A266 );
 a7040a <=( (not A301)  and  (not A299) );
 a7041a <=( (not A298)  and  a7040a );
 a7042a <=( a7041a  and  a7036a );
 a7045a <=( A167  and  A168 );
 a7049a <=( A265  and  A201 );
 a7050a <=( A199  and  a7049a );
 a7051a <=( a7050a  and  a7045a );
 a7054a <=( A269  and  (not A266) );
 a7058a <=( (not A302)  and  (not A301) );
 a7059a <=( (not A300)  and  a7058a );
 a7060a <=( a7059a  and  a7054a );
 a7063a <=( A167  and  A168 );
 a7067a <=( A265  and  A201 );
 a7068a <=( A199  and  a7067a );
 a7069a <=( a7068a  and  a7063a );
 a7072a <=( A269  and  (not A266) );
 a7076a <=( (not A301)  and  (not A299) );
 a7077a <=( (not A298)  and  a7076a );
 a7078a <=( a7077a  and  a7072a );
 a7081a <=( A167  and  A168 );
 a7085a <=( A265  and  A201 );
 a7086a <=( A200  and  a7085a );
 a7087a <=( a7086a  and  a7081a );
 a7090a <=( A298  and  A267 );
 a7094a <=( (not A301)  and  (not A300) );
 a7095a <=( A299  and  a7094a );
 a7096a <=( a7095a  and  a7090a );
 a7099a <=( A167  and  A168 );
 a7103a <=( A266  and  A201 );
 a7104a <=( A200  and  a7103a );
 a7105a <=( a7104a  and  a7099a );
 a7108a <=( A298  and  A267 );
 a7112a <=( (not A301)  and  (not A300) );
 a7113a <=( A299  and  a7112a );
 a7114a <=( a7113a  and  a7108a );
 a7117a <=( A167  and  A168 );
 a7121a <=( (not A265)  and  A201 );
 a7122a <=( A200  and  a7121a );
 a7123a <=( a7122a  and  a7117a );
 a7126a <=( A269  and  A266 );
 a7130a <=( (not A302)  and  (not A301) );
 a7131a <=( (not A300)  and  a7130a );
 a7132a <=( a7131a  and  a7126a );
 a7135a <=( A167  and  A168 );
 a7139a <=( (not A265)  and  A201 );
 a7140a <=( A200  and  a7139a );
 a7141a <=( a7140a  and  a7135a );
 a7144a <=( A269  and  A266 );
 a7148a <=( (not A301)  and  (not A299) );
 a7149a <=( (not A298)  and  a7148a );
 a7150a <=( a7149a  and  a7144a );
 a7153a <=( A167  and  A168 );
 a7157a <=( A265  and  A201 );
 a7158a <=( A200  and  a7157a );
 a7159a <=( a7158a  and  a7153a );
 a7162a <=( A269  and  (not A266) );
 a7166a <=( (not A302)  and  (not A301) );
 a7167a <=( (not A300)  and  a7166a );
 a7168a <=( a7167a  and  a7162a );
 a7171a <=( A167  and  A168 );
 a7175a <=( A265  and  A201 );
 a7176a <=( A200  and  a7175a );
 a7177a <=( a7176a  and  a7171a );
 a7180a <=( A269  and  (not A266) );
 a7184a <=( (not A301)  and  (not A299) );
 a7185a <=( (not A298)  and  a7184a );
 a7186a <=( a7185a  and  a7180a );
 a7189a <=( A167  and  A168 );
 a7193a <=( (not A201)  and  A200 );
 a7194a <=( A199  and  a7193a );
 a7195a <=( a7194a  and  a7189a );
 a7198a <=( (not A267)  and  (not A202) );
 a7202a <=( A301  and  (not A269) );
 a7203a <=( (not A268)  and  a7202a );
 a7204a <=( a7203a  and  a7198a );
 a7207a <=( A167  and  A168 );
 a7211a <=( (not A201)  and  A200 );
 a7212a <=( A199  and  a7211a );
 a7213a <=( a7212a  and  a7207a );
 a7216a <=( (not A265)  and  (not A202) );
 a7220a <=( A301  and  (not A268) );
 a7221a <=( (not A266)  and  a7220a );
 a7222a <=( a7221a  and  a7216a );
 a7225a <=( A167  and  A168 );
 a7229a <=( A203  and  A200 );
 a7230a <=( (not A199)  and  a7229a );
 a7231a <=( a7230a  and  a7225a );
 a7234a <=( A298  and  A268 );
 a7238a <=( (not A301)  and  (not A300) );
 a7239a <=( A299  and  a7238a );
 a7240a <=( a7239a  and  a7234a );
 a7243a <=( A167  and  A168 );
 a7247a <=( A203  and  A200 );
 a7248a <=( (not A199)  and  a7247a );
 a7249a <=( a7248a  and  a7243a );
 a7252a <=( A267  and  A265 );
 a7256a <=( (not A302)  and  (not A301) );
 a7257a <=( (not A300)  and  a7256a );
 a7258a <=( a7257a  and  a7252a );
 a7261a <=( A167  and  A168 );
 a7265a <=( A203  and  A200 );
 a7266a <=( (not A199)  and  a7265a );
 a7267a <=( a7266a  and  a7261a );
 a7270a <=( A267  and  A265 );
 a7274a <=( (not A301)  and  (not A299) );
 a7275a <=( (not A298)  and  a7274a );
 a7276a <=( a7275a  and  a7270a );
 a7279a <=( A167  and  A168 );
 a7283a <=( A203  and  A200 );
 a7284a <=( (not A199)  and  a7283a );
 a7285a <=( a7284a  and  a7279a );
 a7288a <=( A267  and  A266 );
 a7292a <=( (not A302)  and  (not A301) );
 a7293a <=( (not A300)  and  a7292a );
 a7294a <=( a7293a  and  a7288a );
 a7297a <=( A167  and  A168 );
 a7301a <=( A203  and  A200 );
 a7302a <=( (not A199)  and  a7301a );
 a7303a <=( a7302a  and  a7297a );
 a7306a <=( A267  and  A266 );
 a7310a <=( (not A301)  and  (not A299) );
 a7311a <=( (not A298)  and  a7310a );
 a7312a <=( a7311a  and  a7306a );
 a7315a <=( A167  and  A168 );
 a7319a <=( A203  and  (not A200) );
 a7320a <=( A199  and  a7319a );
 a7321a <=( a7320a  and  a7315a );
 a7324a <=( A298  and  A268 );
 a7328a <=( (not A301)  and  (not A300) );
 a7329a <=( A299  and  a7328a );
 a7330a <=( a7329a  and  a7324a );
 a7333a <=( A167  and  A168 );
 a7337a <=( A203  and  (not A200) );
 a7338a <=( A199  and  a7337a );
 a7339a <=( a7338a  and  a7333a );
 a7342a <=( A267  and  A265 );
 a7346a <=( (not A302)  and  (not A301) );
 a7347a <=( (not A300)  and  a7346a );
 a7348a <=( a7347a  and  a7342a );
 a7351a <=( A167  and  A168 );
 a7355a <=( A203  and  (not A200) );
 a7356a <=( A199  and  a7355a );
 a7357a <=( a7356a  and  a7351a );
 a7360a <=( A267  and  A265 );
 a7364a <=( (not A301)  and  (not A299) );
 a7365a <=( (not A298)  and  a7364a );
 a7366a <=( a7365a  and  a7360a );
 a7369a <=( A167  and  A168 );
 a7373a <=( A203  and  (not A200) );
 a7374a <=( A199  and  a7373a );
 a7375a <=( a7374a  and  a7369a );
 a7378a <=( A267  and  A266 );
 a7382a <=( (not A302)  and  (not A301) );
 a7383a <=( (not A300)  and  a7382a );
 a7384a <=( a7383a  and  a7378a );
 a7387a <=( A167  and  A168 );
 a7391a <=( A203  and  (not A200) );
 a7392a <=( A199  and  a7391a );
 a7393a <=( a7392a  and  a7387a );
 a7396a <=( A267  and  A266 );
 a7400a <=( (not A301)  and  (not A299) );
 a7401a <=( (not A298)  and  a7400a );
 a7402a <=( a7401a  and  a7396a );
 a7405a <=( A167  and  A168 );
 a7409a <=( (not A202)  and  (not A200) );
 a7410a <=( (not A199)  and  a7409a );
 a7411a <=( a7410a  and  a7405a );
 a7414a <=( (not A268)  and  (not A267) );
 a7418a <=( A300  and  A299 );
 a7419a <=( (not A269)  and  a7418a );
 a7420a <=( a7419a  and  a7414a );
 a7423a <=( A167  and  A168 );
 a7427a <=( (not A202)  and  (not A200) );
 a7428a <=( (not A199)  and  a7427a );
 a7429a <=( a7428a  and  a7423a );
 a7432a <=( (not A268)  and  (not A267) );
 a7436a <=( A300  and  A298 );
 a7437a <=( (not A269)  and  a7436a );
 a7438a <=( a7437a  and  a7432a );
 a7441a <=( A167  and  A168 );
 a7445a <=( (not A202)  and  (not A200) );
 a7446a <=( (not A199)  and  a7445a );
 a7447a <=( a7446a  and  a7441a );
 a7450a <=( A266  and  A265 );
 a7454a <=( A301  and  (not A268) );
 a7455a <=( (not A267)  and  a7454a );
 a7456a <=( a7455a  and  a7450a );
 a7459a <=( A167  and  A168 );
 a7463a <=( (not A202)  and  (not A200) );
 a7464a <=( (not A199)  and  a7463a );
 a7465a <=( a7464a  and  a7459a );
 a7468a <=( (not A266)  and  (not A265) );
 a7472a <=( A300  and  A299 );
 a7473a <=( (not A268)  and  a7472a );
 a7474a <=( a7473a  and  a7468a );
 a7477a <=( A167  and  A168 );
 a7481a <=( (not A202)  and  (not A200) );
 a7482a <=( (not A199)  and  a7481a );
 a7483a <=( a7482a  and  a7477a );
 a7486a <=( (not A266)  and  (not A265) );
 a7490a <=( A300  and  A298 );
 a7491a <=( (not A268)  and  a7490a );
 a7492a <=( a7491a  and  a7486a );
 a7495a <=( A167  and  A170 );
 a7499a <=( A265  and  A202 );
 a7500a <=( (not A166)  and  a7499a );
 a7501a <=( a7500a  and  a7495a );
 a7504a <=( A298  and  A267 );
 a7508a <=( (not A301)  and  (not A300) );
 a7509a <=( A299  and  a7508a );
 a7510a <=( a7509a  and  a7504a );
 a7513a <=( A167  and  A170 );
 a7517a <=( A266  and  A202 );
 a7518a <=( (not A166)  and  a7517a );
 a7519a <=( a7518a  and  a7513a );
 a7522a <=( A298  and  A267 );
 a7526a <=( (not A301)  and  (not A300) );
 a7527a <=( A299  and  a7526a );
 a7528a <=( a7527a  and  a7522a );
 a7531a <=( A167  and  A170 );
 a7535a <=( (not A265)  and  A202 );
 a7536a <=( (not A166)  and  a7535a );
 a7537a <=( a7536a  and  a7531a );
 a7540a <=( A269  and  A266 );
 a7544a <=( (not A302)  and  (not A301) );
 a7545a <=( (not A300)  and  a7544a );
 a7546a <=( a7545a  and  a7540a );
 a7549a <=( A167  and  A170 );
 a7553a <=( (not A265)  and  A202 );
 a7554a <=( (not A166)  and  a7553a );
 a7555a <=( a7554a  and  a7549a );
 a7558a <=( A269  and  A266 );
 a7562a <=( (not A301)  and  (not A299) );
 a7563a <=( (not A298)  and  a7562a );
 a7564a <=( a7563a  and  a7558a );
 a7567a <=( A167  and  A170 );
 a7571a <=( A265  and  A202 );
 a7572a <=( (not A166)  and  a7571a );
 a7573a <=( a7572a  and  a7567a );
 a7576a <=( A269  and  (not A266) );
 a7580a <=( (not A302)  and  (not A301) );
 a7581a <=( (not A300)  and  a7580a );
 a7582a <=( a7581a  and  a7576a );
 a7585a <=( A167  and  A170 );
 a7589a <=( A265  and  A202 );
 a7590a <=( (not A166)  and  a7589a );
 a7591a <=( a7590a  and  a7585a );
 a7594a <=( A269  and  (not A266) );
 a7598a <=( (not A301)  and  (not A299) );
 a7599a <=( (not A298)  and  a7598a );
 a7600a <=( a7599a  and  a7594a );
 a7603a <=( A167  and  A170 );
 a7607a <=( (not A202)  and  (not A201) );
 a7608a <=( (not A166)  and  a7607a );
 a7609a <=( a7608a  and  a7603a );
 a7612a <=( (not A267)  and  (not A203) );
 a7616a <=( A301  and  (not A269) );
 a7617a <=( (not A268)  and  a7616a );
 a7618a <=( a7617a  and  a7612a );
 a7621a <=( A167  and  A170 );
 a7625a <=( (not A202)  and  (not A201) );
 a7626a <=( (not A166)  and  a7625a );
 a7627a <=( a7626a  and  a7621a );
 a7630a <=( (not A265)  and  (not A203) );
 a7634a <=( A301  and  (not A268) );
 a7635a <=( (not A266)  and  a7634a );
 a7636a <=( a7635a  and  a7630a );
 a7639a <=( A167  and  A170 );
 a7643a <=( A201  and  A199 );
 a7644a <=( (not A166)  and  a7643a );
 a7645a <=( a7644a  and  a7639a );
 a7648a <=( A298  and  A268 );
 a7652a <=( (not A301)  and  (not A300) );
 a7653a <=( A299  and  a7652a );
 a7654a <=( a7653a  and  a7648a );
 a7657a <=( A167  and  A170 );
 a7661a <=( A201  and  A199 );
 a7662a <=( (not A166)  and  a7661a );
 a7663a <=( a7662a  and  a7657a );
 a7666a <=( A267  and  A265 );
 a7670a <=( (not A302)  and  (not A301) );
 a7671a <=( (not A300)  and  a7670a );
 a7672a <=( a7671a  and  a7666a );
 a7675a <=( A167  and  A170 );
 a7679a <=( A201  and  A199 );
 a7680a <=( (not A166)  and  a7679a );
 a7681a <=( a7680a  and  a7675a );
 a7684a <=( A267  and  A265 );
 a7688a <=( (not A301)  and  (not A299) );
 a7689a <=( (not A298)  and  a7688a );
 a7690a <=( a7689a  and  a7684a );
 a7693a <=( A167  and  A170 );
 a7697a <=( A201  and  A199 );
 a7698a <=( (not A166)  and  a7697a );
 a7699a <=( a7698a  and  a7693a );
 a7702a <=( A267  and  A266 );
 a7706a <=( (not A302)  and  (not A301) );
 a7707a <=( (not A300)  and  a7706a );
 a7708a <=( a7707a  and  a7702a );
 a7711a <=( A167  and  A170 );
 a7715a <=( A201  and  A199 );
 a7716a <=( (not A166)  and  a7715a );
 a7717a <=( a7716a  and  a7711a );
 a7720a <=( A267  and  A266 );
 a7724a <=( (not A301)  and  (not A299) );
 a7725a <=( (not A298)  and  a7724a );
 a7726a <=( a7725a  and  a7720a );
 a7729a <=( A167  and  A170 );
 a7733a <=( A201  and  A200 );
 a7734a <=( (not A166)  and  a7733a );
 a7735a <=( a7734a  and  a7729a );
 a7738a <=( A298  and  A268 );
 a7742a <=( (not A301)  and  (not A300) );
 a7743a <=( A299  and  a7742a );
 a7744a <=( a7743a  and  a7738a );
 a7747a <=( A167  and  A170 );
 a7751a <=( A201  and  A200 );
 a7752a <=( (not A166)  and  a7751a );
 a7753a <=( a7752a  and  a7747a );
 a7756a <=( A267  and  A265 );
 a7760a <=( (not A302)  and  (not A301) );
 a7761a <=( (not A300)  and  a7760a );
 a7762a <=( a7761a  and  a7756a );
 a7765a <=( A167  and  A170 );
 a7769a <=( A201  and  A200 );
 a7770a <=( (not A166)  and  a7769a );
 a7771a <=( a7770a  and  a7765a );
 a7774a <=( A267  and  A265 );
 a7778a <=( (not A301)  and  (not A299) );
 a7779a <=( (not A298)  and  a7778a );
 a7780a <=( a7779a  and  a7774a );
 a7783a <=( A167  and  A170 );
 a7787a <=( A201  and  A200 );
 a7788a <=( (not A166)  and  a7787a );
 a7789a <=( a7788a  and  a7783a );
 a7792a <=( A267  and  A266 );
 a7796a <=( (not A302)  and  (not A301) );
 a7797a <=( (not A300)  and  a7796a );
 a7798a <=( a7797a  and  a7792a );
 a7801a <=( A167  and  A170 );
 a7805a <=( A201  and  A200 );
 a7806a <=( (not A166)  and  a7805a );
 a7807a <=( a7806a  and  a7801a );
 a7810a <=( A267  and  A266 );
 a7814a <=( (not A301)  and  (not A299) );
 a7815a <=( (not A298)  and  a7814a );
 a7816a <=( a7815a  and  a7810a );
 a7819a <=( A167  and  A170 );
 a7823a <=( A200  and  (not A199) );
 a7824a <=( (not A166)  and  a7823a );
 a7825a <=( a7824a  and  a7819a );
 a7828a <=( A268  and  A203 );
 a7832a <=( (not A302)  and  (not A301) );
 a7833a <=( (not A300)  and  a7832a );
 a7834a <=( a7833a  and  a7828a );
 a7837a <=( A167  and  A170 );
 a7841a <=( A200  and  (not A199) );
 a7842a <=( (not A166)  and  a7841a );
 a7843a <=( a7842a  and  a7837a );
 a7846a <=( A268  and  A203 );
 a7850a <=( (not A301)  and  (not A299) );
 a7851a <=( (not A298)  and  a7850a );
 a7852a <=( a7851a  and  a7846a );
 a7855a <=( A167  and  A170 );
 a7859a <=( (not A200)  and  A199 );
 a7860a <=( (not A166)  and  a7859a );
 a7861a <=( a7860a  and  a7855a );
 a7864a <=( A268  and  A203 );
 a7868a <=( (not A302)  and  (not A301) );
 a7869a <=( (not A300)  and  a7868a );
 a7870a <=( a7869a  and  a7864a );
 a7873a <=( A167  and  A170 );
 a7877a <=( (not A200)  and  A199 );
 a7878a <=( (not A166)  and  a7877a );
 a7879a <=( a7878a  and  a7873a );
 a7882a <=( A268  and  A203 );
 a7886a <=( (not A301)  and  (not A299) );
 a7887a <=( (not A298)  and  a7886a );
 a7888a <=( a7887a  and  a7882a );
 a7891a <=( A167  and  A170 );
 a7895a <=( (not A200)  and  (not A199) );
 a7896a <=( (not A166)  and  a7895a );
 a7897a <=( a7896a  and  a7891a );
 a7900a <=( (not A267)  and  (not A202) );
 a7904a <=( A301  and  (not A269) );
 a7905a <=( (not A268)  and  a7904a );
 a7906a <=( a7905a  and  a7900a );
 a7909a <=( A167  and  A170 );
 a7913a <=( (not A200)  and  (not A199) );
 a7914a <=( (not A166)  and  a7913a );
 a7915a <=( a7914a  and  a7909a );
 a7918a <=( (not A265)  and  (not A202) );
 a7922a <=( A301  and  (not A268) );
 a7923a <=( (not A266)  and  a7922a );
 a7924a <=( a7923a  and  a7918a );
 a7927a <=( (not A167)  and  A170 );
 a7931a <=( A265  and  A202 );
 a7932a <=( A166  and  a7931a );
 a7933a <=( a7932a  and  a7927a );
 a7936a <=( A298  and  A267 );
 a7940a <=( (not A301)  and  (not A300) );
 a7941a <=( A299  and  a7940a );
 a7942a <=( a7941a  and  a7936a );
 a7945a <=( (not A167)  and  A170 );
 a7949a <=( A266  and  A202 );
 a7950a <=( A166  and  a7949a );
 a7951a <=( a7950a  and  a7945a );
 a7954a <=( A298  and  A267 );
 a7958a <=( (not A301)  and  (not A300) );
 a7959a <=( A299  and  a7958a );
 a7960a <=( a7959a  and  a7954a );
 a7963a <=( (not A167)  and  A170 );
 a7967a <=( (not A265)  and  A202 );
 a7968a <=( A166  and  a7967a );
 a7969a <=( a7968a  and  a7963a );
 a7972a <=( A269  and  A266 );
 a7976a <=( (not A302)  and  (not A301) );
 a7977a <=( (not A300)  and  a7976a );
 a7978a <=( a7977a  and  a7972a );
 a7981a <=( (not A167)  and  A170 );
 a7985a <=( (not A265)  and  A202 );
 a7986a <=( A166  and  a7985a );
 a7987a <=( a7986a  and  a7981a );
 a7990a <=( A269  and  A266 );
 a7994a <=( (not A301)  and  (not A299) );
 a7995a <=( (not A298)  and  a7994a );
 a7996a <=( a7995a  and  a7990a );
 a7999a <=( (not A167)  and  A170 );
 a8003a <=( A265  and  A202 );
 a8004a <=( A166  and  a8003a );
 a8005a <=( a8004a  and  a7999a );
 a8008a <=( A269  and  (not A266) );
 a8012a <=( (not A302)  and  (not A301) );
 a8013a <=( (not A300)  and  a8012a );
 a8014a <=( a8013a  and  a8008a );
 a8017a <=( (not A167)  and  A170 );
 a8021a <=( A265  and  A202 );
 a8022a <=( A166  and  a8021a );
 a8023a <=( a8022a  and  a8017a );
 a8026a <=( A269  and  (not A266) );
 a8030a <=( (not A301)  and  (not A299) );
 a8031a <=( (not A298)  and  a8030a );
 a8032a <=( a8031a  and  a8026a );
 a8035a <=( (not A167)  and  A170 );
 a8039a <=( (not A202)  and  (not A201) );
 a8040a <=( A166  and  a8039a );
 a8041a <=( a8040a  and  a8035a );
 a8044a <=( (not A267)  and  (not A203) );
 a8048a <=( A301  and  (not A269) );
 a8049a <=( (not A268)  and  a8048a );
 a8050a <=( a8049a  and  a8044a );
 a8053a <=( (not A167)  and  A170 );
 a8057a <=( (not A202)  and  (not A201) );
 a8058a <=( A166  and  a8057a );
 a8059a <=( a8058a  and  a8053a );
 a8062a <=( (not A265)  and  (not A203) );
 a8066a <=( A301  and  (not A268) );
 a8067a <=( (not A266)  and  a8066a );
 a8068a <=( a8067a  and  a8062a );
 a8071a <=( (not A167)  and  A170 );
 a8075a <=( A201  and  A199 );
 a8076a <=( A166  and  a8075a );
 a8077a <=( a8076a  and  a8071a );
 a8080a <=( A298  and  A268 );
 a8084a <=( (not A301)  and  (not A300) );
 a8085a <=( A299  and  a8084a );
 a8086a <=( a8085a  and  a8080a );
 a8089a <=( (not A167)  and  A170 );
 a8093a <=( A201  and  A199 );
 a8094a <=( A166  and  a8093a );
 a8095a <=( a8094a  and  a8089a );
 a8098a <=( A267  and  A265 );
 a8102a <=( (not A302)  and  (not A301) );
 a8103a <=( (not A300)  and  a8102a );
 a8104a <=( a8103a  and  a8098a );
 a8107a <=( (not A167)  and  A170 );
 a8111a <=( A201  and  A199 );
 a8112a <=( A166  and  a8111a );
 a8113a <=( a8112a  and  a8107a );
 a8116a <=( A267  and  A265 );
 a8120a <=( (not A301)  and  (not A299) );
 a8121a <=( (not A298)  and  a8120a );
 a8122a <=( a8121a  and  a8116a );
 a8125a <=( (not A167)  and  A170 );
 a8129a <=( A201  and  A199 );
 a8130a <=( A166  and  a8129a );
 a8131a <=( a8130a  and  a8125a );
 a8134a <=( A267  and  A266 );
 a8138a <=( (not A302)  and  (not A301) );
 a8139a <=( (not A300)  and  a8138a );
 a8140a <=( a8139a  and  a8134a );
 a8143a <=( (not A167)  and  A170 );
 a8147a <=( A201  and  A199 );
 a8148a <=( A166  and  a8147a );
 a8149a <=( a8148a  and  a8143a );
 a8152a <=( A267  and  A266 );
 a8156a <=( (not A301)  and  (not A299) );
 a8157a <=( (not A298)  and  a8156a );
 a8158a <=( a8157a  and  a8152a );
 a8161a <=( (not A167)  and  A170 );
 a8165a <=( A201  and  A200 );
 a8166a <=( A166  and  a8165a );
 a8167a <=( a8166a  and  a8161a );
 a8170a <=( A298  and  A268 );
 a8174a <=( (not A301)  and  (not A300) );
 a8175a <=( A299  and  a8174a );
 a8176a <=( a8175a  and  a8170a );
 a8179a <=( (not A167)  and  A170 );
 a8183a <=( A201  and  A200 );
 a8184a <=( A166  and  a8183a );
 a8185a <=( a8184a  and  a8179a );
 a8188a <=( A267  and  A265 );
 a8192a <=( (not A302)  and  (not A301) );
 a8193a <=( (not A300)  and  a8192a );
 a8194a <=( a8193a  and  a8188a );
 a8197a <=( (not A167)  and  A170 );
 a8201a <=( A201  and  A200 );
 a8202a <=( A166  and  a8201a );
 a8203a <=( a8202a  and  a8197a );
 a8206a <=( A267  and  A265 );
 a8210a <=( (not A301)  and  (not A299) );
 a8211a <=( (not A298)  and  a8210a );
 a8212a <=( a8211a  and  a8206a );
 a8215a <=( (not A167)  and  A170 );
 a8219a <=( A201  and  A200 );
 a8220a <=( A166  and  a8219a );
 a8221a <=( a8220a  and  a8215a );
 a8224a <=( A267  and  A266 );
 a8228a <=( (not A302)  and  (not A301) );
 a8229a <=( (not A300)  and  a8228a );
 a8230a <=( a8229a  and  a8224a );
 a8233a <=( (not A167)  and  A170 );
 a8237a <=( A201  and  A200 );
 a8238a <=( A166  and  a8237a );
 a8239a <=( a8238a  and  a8233a );
 a8242a <=( A267  and  A266 );
 a8246a <=( (not A301)  and  (not A299) );
 a8247a <=( (not A298)  and  a8246a );
 a8248a <=( a8247a  and  a8242a );
 a8251a <=( (not A167)  and  A170 );
 a8255a <=( A200  and  (not A199) );
 a8256a <=( A166  and  a8255a );
 a8257a <=( a8256a  and  a8251a );
 a8260a <=( A268  and  A203 );
 a8264a <=( (not A302)  and  (not A301) );
 a8265a <=( (not A300)  and  a8264a );
 a8266a <=( a8265a  and  a8260a );
 a8269a <=( (not A167)  and  A170 );
 a8273a <=( A200  and  (not A199) );
 a8274a <=( A166  and  a8273a );
 a8275a <=( a8274a  and  a8269a );
 a8278a <=( A268  and  A203 );
 a8282a <=( (not A301)  and  (not A299) );
 a8283a <=( (not A298)  and  a8282a );
 a8284a <=( a8283a  and  a8278a );
 a8287a <=( (not A167)  and  A170 );
 a8291a <=( (not A200)  and  A199 );
 a8292a <=( A166  and  a8291a );
 a8293a <=( a8292a  and  a8287a );
 a8296a <=( A268  and  A203 );
 a8300a <=( (not A302)  and  (not A301) );
 a8301a <=( (not A300)  and  a8300a );
 a8302a <=( a8301a  and  a8296a );
 a8305a <=( (not A167)  and  A170 );
 a8309a <=( (not A200)  and  A199 );
 a8310a <=( A166  and  a8309a );
 a8311a <=( a8310a  and  a8305a );
 a8314a <=( A268  and  A203 );
 a8318a <=( (not A301)  and  (not A299) );
 a8319a <=( (not A298)  and  a8318a );
 a8320a <=( a8319a  and  a8314a );
 a8323a <=( (not A167)  and  A170 );
 a8327a <=( (not A200)  and  (not A199) );
 a8328a <=( A166  and  a8327a );
 a8329a <=( a8328a  and  a8323a );
 a8332a <=( (not A267)  and  (not A202) );
 a8336a <=( A301  and  (not A269) );
 a8337a <=( (not A268)  and  a8336a );
 a8338a <=( a8337a  and  a8332a );
 a8341a <=( (not A167)  and  A170 );
 a8345a <=( (not A200)  and  (not A199) );
 a8346a <=( A166  and  a8345a );
 a8347a <=( a8346a  and  a8341a );
 a8350a <=( (not A265)  and  (not A202) );
 a8354a <=( A301  and  (not A268) );
 a8355a <=( (not A266)  and  a8354a );
 a8356a <=( a8355a  and  a8350a );
 a8359a <=( (not A201)  and  A169 );
 a8363a <=( (not A267)  and  (not A203) );
 a8364a <=( (not A202)  and  a8363a );
 a8365a <=( a8364a  and  a8359a );
 a8368a <=( (not A269)  and  (not A268) );
 a8372a <=( A302  and  (not A299) );
 a8373a <=( A298  and  a8372a );
 a8374a <=( a8373a  and  a8368a );
 a8377a <=( (not A201)  and  A169 );
 a8381a <=( (not A267)  and  (not A203) );
 a8382a <=( (not A202)  and  a8381a );
 a8383a <=( a8382a  and  a8377a );
 a8386a <=( (not A269)  and  (not A268) );
 a8390a <=( A302  and  A299 );
 a8391a <=( (not A298)  and  a8390a );
 a8392a <=( a8391a  and  a8386a );
 a8395a <=( (not A201)  and  A169 );
 a8399a <=( A265  and  (not A203) );
 a8400a <=( (not A202)  and  a8399a );
 a8401a <=( a8400a  and  a8395a );
 a8404a <=( (not A267)  and  A266 );
 a8408a <=( A300  and  A299 );
 a8409a <=( (not A268)  and  a8408a );
 a8410a <=( a8409a  and  a8404a );
 a8413a <=( (not A201)  and  A169 );
 a8417a <=( A265  and  (not A203) );
 a8418a <=( (not A202)  and  a8417a );
 a8419a <=( a8418a  and  a8413a );
 a8422a <=( (not A267)  and  A266 );
 a8426a <=( A300  and  A298 );
 a8427a <=( (not A268)  and  a8426a );
 a8428a <=( a8427a  and  a8422a );
 a8431a <=( (not A201)  and  A169 );
 a8435a <=( (not A265)  and  (not A203) );
 a8436a <=( (not A202)  and  a8435a );
 a8437a <=( a8436a  and  a8431a );
 a8440a <=( (not A268)  and  (not A266) );
 a8444a <=( A302  and  (not A299) );
 a8445a <=( A298  and  a8444a );
 a8446a <=( a8445a  and  a8440a );
 a8449a <=( (not A201)  and  A169 );
 a8453a <=( (not A265)  and  (not A203) );
 a8454a <=( (not A202)  and  a8453a );
 a8455a <=( a8454a  and  a8449a );
 a8458a <=( (not A268)  and  (not A266) );
 a8462a <=( A302  and  A299 );
 a8463a <=( (not A298)  and  a8462a );
 a8464a <=( a8463a  and  a8458a );
 a8467a <=( A199  and  A169 );
 a8471a <=( A266  and  (not A265) );
 a8472a <=( A201  and  a8471a );
 a8473a <=( a8472a  and  a8467a );
 a8476a <=( A298  and  A269 );
 a8480a <=( (not A301)  and  (not A300) );
 a8481a <=( A299  and  a8480a );
 a8482a <=( a8481a  and  a8476a );
 a8485a <=( A199  and  A169 );
 a8489a <=( (not A266)  and  A265 );
 a8490a <=( A201  and  a8489a );
 a8491a <=( a8490a  and  a8485a );
 a8494a <=( A298  and  A269 );
 a8498a <=( (not A301)  and  (not A300) );
 a8499a <=( A299  and  a8498a );
 a8500a <=( a8499a  and  a8494a );
 a8503a <=( A200  and  A169 );
 a8507a <=( A266  and  (not A265) );
 a8508a <=( A201  and  a8507a );
 a8509a <=( a8508a  and  a8503a );
 a8512a <=( A298  and  A269 );
 a8516a <=( (not A301)  and  (not A300) );
 a8517a <=( A299  and  a8516a );
 a8518a <=( a8517a  and  a8512a );
 a8521a <=( A200  and  A169 );
 a8525a <=( (not A266)  and  A265 );
 a8526a <=( A201  and  a8525a );
 a8527a <=( a8526a  and  a8521a );
 a8530a <=( A298  and  A269 );
 a8534a <=( (not A301)  and  (not A300) );
 a8535a <=( A299  and  a8534a );
 a8536a <=( a8535a  and  a8530a );
 a8539a <=( A199  and  A169 );
 a8543a <=( (not A202)  and  (not A201) );
 a8544a <=( A200  and  a8543a );
 a8545a <=( a8544a  and  a8539a );
 a8548a <=( (not A268)  and  (not A267) );
 a8552a <=( A300  and  A299 );
 a8553a <=( (not A269)  and  a8552a );
 a8554a <=( a8553a  and  a8548a );
 a8557a <=( A199  and  A169 );
 a8561a <=( (not A202)  and  (not A201) );
 a8562a <=( A200  and  a8561a );
 a8563a <=( a8562a  and  a8557a );
 a8566a <=( (not A268)  and  (not A267) );
 a8570a <=( A300  and  A298 );
 a8571a <=( (not A269)  and  a8570a );
 a8572a <=( a8571a  and  a8566a );
 a8575a <=( A199  and  A169 );
 a8579a <=( (not A202)  and  (not A201) );
 a8580a <=( A200  and  a8579a );
 a8581a <=( a8580a  and  a8575a );
 a8584a <=( A266  and  A265 );
 a8588a <=( A301  and  (not A268) );
 a8589a <=( (not A267)  and  a8588a );
 a8590a <=( a8589a  and  a8584a );
 a8593a <=( A199  and  A169 );
 a8597a <=( (not A202)  and  (not A201) );
 a8598a <=( A200  and  a8597a );
 a8599a <=( a8598a  and  a8593a );
 a8602a <=( (not A266)  and  (not A265) );
 a8606a <=( A300  and  A299 );
 a8607a <=( (not A268)  and  a8606a );
 a8608a <=( a8607a  and  a8602a );
 a8611a <=( A199  and  A169 );
 a8615a <=( (not A202)  and  (not A201) );
 a8616a <=( A200  and  a8615a );
 a8617a <=( a8616a  and  a8611a );
 a8620a <=( (not A266)  and  (not A265) );
 a8624a <=( A300  and  A298 );
 a8625a <=( (not A268)  and  a8624a );
 a8626a <=( a8625a  and  a8620a );
 a8629a <=( (not A199)  and  A169 );
 a8633a <=( A265  and  A203 );
 a8634a <=( A200  and  a8633a );
 a8635a <=( a8634a  and  a8629a );
 a8638a <=( A298  and  A267 );
 a8642a <=( (not A301)  and  (not A300) );
 a8643a <=( A299  and  a8642a );
 a8644a <=( a8643a  and  a8638a );
 a8647a <=( (not A199)  and  A169 );
 a8651a <=( A266  and  A203 );
 a8652a <=( A200  and  a8651a );
 a8653a <=( a8652a  and  a8647a );
 a8656a <=( A298  and  A267 );
 a8660a <=( (not A301)  and  (not A300) );
 a8661a <=( A299  and  a8660a );
 a8662a <=( a8661a  and  a8656a );
 a8665a <=( (not A199)  and  A169 );
 a8669a <=( (not A265)  and  A203 );
 a8670a <=( A200  and  a8669a );
 a8671a <=( a8670a  and  a8665a );
 a8674a <=( A269  and  A266 );
 a8678a <=( (not A302)  and  (not A301) );
 a8679a <=( (not A300)  and  a8678a );
 a8680a <=( a8679a  and  a8674a );
 a8683a <=( (not A199)  and  A169 );
 a8687a <=( (not A265)  and  A203 );
 a8688a <=( A200  and  a8687a );
 a8689a <=( a8688a  and  a8683a );
 a8692a <=( A269  and  A266 );
 a8696a <=( (not A301)  and  (not A299) );
 a8697a <=( (not A298)  and  a8696a );
 a8698a <=( a8697a  and  a8692a );
 a8701a <=( (not A199)  and  A169 );
 a8705a <=( A265  and  A203 );
 a8706a <=( A200  and  a8705a );
 a8707a <=( a8706a  and  a8701a );
 a8710a <=( A269  and  (not A266) );
 a8714a <=( (not A302)  and  (not A301) );
 a8715a <=( (not A300)  and  a8714a );
 a8716a <=( a8715a  and  a8710a );
 a8719a <=( (not A199)  and  A169 );
 a8723a <=( A265  and  A203 );
 a8724a <=( A200  and  a8723a );
 a8725a <=( a8724a  and  a8719a );
 a8728a <=( A269  and  (not A266) );
 a8732a <=( (not A301)  and  (not A299) );
 a8733a <=( (not A298)  and  a8732a );
 a8734a <=( a8733a  and  a8728a );
 a8737a <=( A199  and  A169 );
 a8741a <=( A265  and  A203 );
 a8742a <=( (not A200)  and  a8741a );
 a8743a <=( a8742a  and  a8737a );
 a8746a <=( A298  and  A267 );
 a8750a <=( (not A301)  and  (not A300) );
 a8751a <=( A299  and  a8750a );
 a8752a <=( a8751a  and  a8746a );
 a8755a <=( A199  and  A169 );
 a8759a <=( A266  and  A203 );
 a8760a <=( (not A200)  and  a8759a );
 a8761a <=( a8760a  and  a8755a );
 a8764a <=( A298  and  A267 );
 a8768a <=( (not A301)  and  (not A300) );
 a8769a <=( A299  and  a8768a );
 a8770a <=( a8769a  and  a8764a );
 a8773a <=( A199  and  A169 );
 a8777a <=( (not A265)  and  A203 );
 a8778a <=( (not A200)  and  a8777a );
 a8779a <=( a8778a  and  a8773a );
 a8782a <=( A269  and  A266 );
 a8786a <=( (not A302)  and  (not A301) );
 a8787a <=( (not A300)  and  a8786a );
 a8788a <=( a8787a  and  a8782a );
 a8791a <=( A199  and  A169 );
 a8795a <=( (not A265)  and  A203 );
 a8796a <=( (not A200)  and  a8795a );
 a8797a <=( a8796a  and  a8791a );
 a8800a <=( A269  and  A266 );
 a8804a <=( (not A301)  and  (not A299) );
 a8805a <=( (not A298)  and  a8804a );
 a8806a <=( a8805a  and  a8800a );
 a8809a <=( A199  and  A169 );
 a8813a <=( A265  and  A203 );
 a8814a <=( (not A200)  and  a8813a );
 a8815a <=( a8814a  and  a8809a );
 a8818a <=( A269  and  (not A266) );
 a8822a <=( (not A302)  and  (not A301) );
 a8823a <=( (not A300)  and  a8822a );
 a8824a <=( a8823a  and  a8818a );
 a8827a <=( A199  and  A169 );
 a8831a <=( A265  and  A203 );
 a8832a <=( (not A200)  and  a8831a );
 a8833a <=( a8832a  and  a8827a );
 a8836a <=( A269  and  (not A266) );
 a8840a <=( (not A301)  and  (not A299) );
 a8841a <=( (not A298)  and  a8840a );
 a8842a <=( a8841a  and  a8836a );
 a8845a <=( (not A199)  and  A169 );
 a8849a <=( (not A267)  and  (not A202) );
 a8850a <=( (not A200)  and  a8849a );
 a8851a <=( a8850a  and  a8845a );
 a8854a <=( (not A269)  and  (not A268) );
 a8858a <=( A302  and  (not A299) );
 a8859a <=( A298  and  a8858a );
 a8860a <=( a8859a  and  a8854a );
 a8863a <=( (not A199)  and  A169 );
 a8867a <=( (not A267)  and  (not A202) );
 a8868a <=( (not A200)  and  a8867a );
 a8869a <=( a8868a  and  a8863a );
 a8872a <=( (not A269)  and  (not A268) );
 a8876a <=( A302  and  A299 );
 a8877a <=( (not A298)  and  a8876a );
 a8878a <=( a8877a  and  a8872a );
 a8881a <=( (not A199)  and  A169 );
 a8885a <=( A265  and  (not A202) );
 a8886a <=( (not A200)  and  a8885a );
 a8887a <=( a8886a  and  a8881a );
 a8890a <=( (not A267)  and  A266 );
 a8894a <=( A300  and  A299 );
 a8895a <=( (not A268)  and  a8894a );
 a8896a <=( a8895a  and  a8890a );
 a8899a <=( (not A199)  and  A169 );
 a8903a <=( A265  and  (not A202) );
 a8904a <=( (not A200)  and  a8903a );
 a8905a <=( a8904a  and  a8899a );
 a8908a <=( (not A267)  and  A266 );
 a8912a <=( A300  and  A298 );
 a8913a <=( (not A268)  and  a8912a );
 a8914a <=( a8913a  and  a8908a );
 a8917a <=( (not A199)  and  A169 );
 a8921a <=( (not A265)  and  (not A202) );
 a8922a <=( (not A200)  and  a8921a );
 a8923a <=( a8922a  and  a8917a );
 a8926a <=( (not A268)  and  (not A266) );
 a8930a <=( A302  and  (not A299) );
 a8931a <=( A298  and  a8930a );
 a8932a <=( a8931a  and  a8926a );
 a8935a <=( (not A199)  and  A169 );
 a8939a <=( (not A265)  and  (not A202) );
 a8940a <=( (not A200)  and  a8939a );
 a8941a <=( a8940a  and  a8935a );
 a8944a <=( (not A268)  and  (not A266) );
 a8948a <=( A302  and  A299 );
 a8949a <=( (not A298)  and  a8948a );
 a8950a <=( a8949a  and  a8944a );
 a8953a <=( (not A167)  and  (not A169) );
 a8957a <=( (not A267)  and  A202 );
 a8958a <=( (not A166)  and  a8957a );
 a8959a <=( a8958a  and  a8953a );
 a8962a <=( (not A269)  and  (not A268) );
 a8966a <=( A302  and  (not A299) );
 a8967a <=( A298  and  a8966a );
 a8968a <=( a8967a  and  a8962a );
 a8971a <=( (not A167)  and  (not A169) );
 a8975a <=( (not A267)  and  A202 );
 a8976a <=( (not A166)  and  a8975a );
 a8977a <=( a8976a  and  a8971a );
 a8980a <=( (not A269)  and  (not A268) );
 a8984a <=( A302  and  A299 );
 a8985a <=( (not A298)  and  a8984a );
 a8986a <=( a8985a  and  a8980a );
 a8989a <=( (not A167)  and  (not A169) );
 a8993a <=( A265  and  A202 );
 a8994a <=( (not A166)  and  a8993a );
 a8995a <=( a8994a  and  a8989a );
 a8998a <=( (not A267)  and  A266 );
 a9002a <=( A300  and  A299 );
 a9003a <=( (not A268)  and  a9002a );
 a9004a <=( a9003a  and  a8998a );
 a9007a <=( (not A167)  and  (not A169) );
 a9011a <=( A265  and  A202 );
 a9012a <=( (not A166)  and  a9011a );
 a9013a <=( a9012a  and  a9007a );
 a9016a <=( (not A267)  and  A266 );
 a9020a <=( A300  and  A298 );
 a9021a <=( (not A268)  and  a9020a );
 a9022a <=( a9021a  and  a9016a );
 a9025a <=( (not A167)  and  (not A169) );
 a9029a <=( (not A265)  and  A202 );
 a9030a <=( (not A166)  and  a9029a );
 a9031a <=( a9030a  and  a9025a );
 a9034a <=( (not A268)  and  (not A266) );
 a9038a <=( A302  and  (not A299) );
 a9039a <=( A298  and  a9038a );
 a9040a <=( a9039a  and  a9034a );
 a9043a <=( (not A167)  and  (not A169) );
 a9047a <=( (not A265)  and  A202 );
 a9048a <=( (not A166)  and  a9047a );
 a9049a <=( a9048a  and  a9043a );
 a9052a <=( (not A268)  and  (not A266) );
 a9056a <=( A302  and  A299 );
 a9057a <=( (not A298)  and  a9056a );
 a9058a <=( a9057a  and  a9052a );
 a9061a <=( (not A167)  and  (not A169) );
 a9065a <=( (not A202)  and  (not A201) );
 a9066a <=( (not A166)  and  a9065a );
 a9067a <=( a9066a  and  a9061a );
 a9070a <=( A268  and  (not A203) );
 a9074a <=( (not A302)  and  (not A301) );
 a9075a <=( (not A300)  and  a9074a );
 a9076a <=( a9075a  and  a9070a );
 a9079a <=( (not A167)  and  (not A169) );
 a9083a <=( (not A202)  and  (not A201) );
 a9084a <=( (not A166)  and  a9083a );
 a9085a <=( a9084a  and  a9079a );
 a9088a <=( A268  and  (not A203) );
 a9092a <=( (not A301)  and  (not A299) );
 a9093a <=( (not A298)  and  a9092a );
 a9094a <=( a9093a  and  a9088a );
 a9097a <=( (not A167)  and  (not A169) );
 a9101a <=( A201  and  A199 );
 a9102a <=( (not A166)  and  a9101a );
 a9103a <=( a9102a  and  a9097a );
 a9106a <=( (not A268)  and  (not A267) );
 a9110a <=( A300  and  A299 );
 a9111a <=( (not A269)  and  a9110a );
 a9112a <=( a9111a  and  a9106a );
 a9115a <=( (not A167)  and  (not A169) );
 a9119a <=( A201  and  A199 );
 a9120a <=( (not A166)  and  a9119a );
 a9121a <=( a9120a  and  a9115a );
 a9124a <=( (not A268)  and  (not A267) );
 a9128a <=( A300  and  A298 );
 a9129a <=( (not A269)  and  a9128a );
 a9130a <=( a9129a  and  a9124a );
 a9133a <=( (not A167)  and  (not A169) );
 a9137a <=( A201  and  A199 );
 a9138a <=( (not A166)  and  a9137a );
 a9139a <=( a9138a  and  a9133a );
 a9142a <=( A266  and  A265 );
 a9146a <=( A301  and  (not A268) );
 a9147a <=( (not A267)  and  a9146a );
 a9148a <=( a9147a  and  a9142a );
 a9151a <=( (not A167)  and  (not A169) );
 a9155a <=( A201  and  A199 );
 a9156a <=( (not A166)  and  a9155a );
 a9157a <=( a9156a  and  a9151a );
 a9160a <=( (not A266)  and  (not A265) );
 a9164a <=( A300  and  A299 );
 a9165a <=( (not A268)  and  a9164a );
 a9166a <=( a9165a  and  a9160a );
 a9169a <=( (not A167)  and  (not A169) );
 a9173a <=( A201  and  A199 );
 a9174a <=( (not A166)  and  a9173a );
 a9175a <=( a9174a  and  a9169a );
 a9178a <=( (not A266)  and  (not A265) );
 a9182a <=( A300  and  A298 );
 a9183a <=( (not A268)  and  a9182a );
 a9184a <=( a9183a  and  a9178a );
 a9187a <=( (not A167)  and  (not A169) );
 a9191a <=( A201  and  A200 );
 a9192a <=( (not A166)  and  a9191a );
 a9193a <=( a9192a  and  a9187a );
 a9196a <=( (not A268)  and  (not A267) );
 a9200a <=( A300  and  A299 );
 a9201a <=( (not A269)  and  a9200a );
 a9202a <=( a9201a  and  a9196a );
 a9205a <=( (not A167)  and  (not A169) );
 a9209a <=( A201  and  A200 );
 a9210a <=( (not A166)  and  a9209a );
 a9211a <=( a9210a  and  a9205a );
 a9214a <=( (not A268)  and  (not A267) );
 a9218a <=( A300  and  A298 );
 a9219a <=( (not A269)  and  a9218a );
 a9220a <=( a9219a  and  a9214a );
 a9223a <=( (not A167)  and  (not A169) );
 a9227a <=( A201  and  A200 );
 a9228a <=( (not A166)  and  a9227a );
 a9229a <=( a9228a  and  a9223a );
 a9232a <=( A266  and  A265 );
 a9236a <=( A301  and  (not A268) );
 a9237a <=( (not A267)  and  a9236a );
 a9238a <=( a9237a  and  a9232a );
 a9241a <=( (not A167)  and  (not A169) );
 a9245a <=( A201  and  A200 );
 a9246a <=( (not A166)  and  a9245a );
 a9247a <=( a9246a  and  a9241a );
 a9250a <=( (not A266)  and  (not A265) );
 a9254a <=( A300  and  A299 );
 a9255a <=( (not A268)  and  a9254a );
 a9256a <=( a9255a  and  a9250a );
 a9259a <=( (not A167)  and  (not A169) );
 a9263a <=( A201  and  A200 );
 a9264a <=( (not A166)  and  a9263a );
 a9265a <=( a9264a  and  a9259a );
 a9268a <=( (not A266)  and  (not A265) );
 a9272a <=( A300  and  A298 );
 a9273a <=( (not A268)  and  a9272a );
 a9274a <=( a9273a  and  a9268a );
 a9277a <=( (not A167)  and  (not A169) );
 a9281a <=( A200  and  (not A199) );
 a9282a <=( (not A166)  and  a9281a );
 a9283a <=( a9282a  and  a9277a );
 a9286a <=( (not A267)  and  A203 );
 a9290a <=( A301  and  (not A269) );
 a9291a <=( (not A268)  and  a9290a );
 a9292a <=( a9291a  and  a9286a );
 a9295a <=( (not A167)  and  (not A169) );
 a9299a <=( A200  and  (not A199) );
 a9300a <=( (not A166)  and  a9299a );
 a9301a <=( a9300a  and  a9295a );
 a9304a <=( (not A265)  and  A203 );
 a9308a <=( A301  and  (not A268) );
 a9309a <=( (not A266)  and  a9308a );
 a9310a <=( a9309a  and  a9304a );
 a9313a <=( (not A167)  and  (not A169) );
 a9317a <=( (not A200)  and  A199 );
 a9318a <=( (not A166)  and  a9317a );
 a9319a <=( a9318a  and  a9313a );
 a9322a <=( (not A267)  and  A203 );
 a9326a <=( A301  and  (not A269) );
 a9327a <=( (not A268)  and  a9326a );
 a9328a <=( a9327a  and  a9322a );
 a9331a <=( (not A167)  and  (not A169) );
 a9335a <=( (not A200)  and  A199 );
 a9336a <=( (not A166)  and  a9335a );
 a9337a <=( a9336a  and  a9331a );
 a9340a <=( (not A265)  and  A203 );
 a9344a <=( A301  and  (not A268) );
 a9345a <=( (not A266)  and  a9344a );
 a9346a <=( a9345a  and  a9340a );
 a9349a <=( (not A167)  and  (not A169) );
 a9353a <=( (not A200)  and  (not A199) );
 a9354a <=( (not A166)  and  a9353a );
 a9355a <=( a9354a  and  a9349a );
 a9358a <=( A268  and  (not A202) );
 a9362a <=( (not A302)  and  (not A301) );
 a9363a <=( (not A300)  and  a9362a );
 a9364a <=( a9363a  and  a9358a );
 a9367a <=( (not A167)  and  (not A169) );
 a9371a <=( (not A200)  and  (not A199) );
 a9372a <=( (not A166)  and  a9371a );
 a9373a <=( a9372a  and  a9367a );
 a9376a <=( A268  and  (not A202) );
 a9380a <=( (not A301)  and  (not A299) );
 a9381a <=( (not A298)  and  a9380a );
 a9382a <=( a9381a  and  a9376a );
 a9385a <=( (not A168)  and  (not A169) );
 a9389a <=( A202  and  A166 );
 a9390a <=( A167  and  a9389a );
 a9391a <=( a9390a  and  a9385a );
 a9394a <=( (not A268)  and  (not A267) );
 a9398a <=( A300  and  A299 );
 a9399a <=( (not A269)  and  a9398a );
 a9400a <=( a9399a  and  a9394a );
 a9403a <=( (not A168)  and  (not A169) );
 a9407a <=( A202  and  A166 );
 a9408a <=( A167  and  a9407a );
 a9409a <=( a9408a  and  a9403a );
 a9412a <=( (not A268)  and  (not A267) );
 a9416a <=( A300  and  A298 );
 a9417a <=( (not A269)  and  a9416a );
 a9418a <=( a9417a  and  a9412a );
 a9421a <=( (not A168)  and  (not A169) );
 a9425a <=( A202  and  A166 );
 a9426a <=( A167  and  a9425a );
 a9427a <=( a9426a  and  a9421a );
 a9430a <=( A266  and  A265 );
 a9434a <=( A301  and  (not A268) );
 a9435a <=( (not A267)  and  a9434a );
 a9436a <=( a9435a  and  a9430a );
 a9439a <=( (not A168)  and  (not A169) );
 a9443a <=( A202  and  A166 );
 a9444a <=( A167  and  a9443a );
 a9445a <=( a9444a  and  a9439a );
 a9448a <=( (not A266)  and  (not A265) );
 a9452a <=( A300  and  A299 );
 a9453a <=( (not A268)  and  a9452a );
 a9454a <=( a9453a  and  a9448a );
 a9457a <=( (not A168)  and  (not A169) );
 a9461a <=( A202  and  A166 );
 a9462a <=( A167  and  a9461a );
 a9463a <=( a9462a  and  a9457a );
 a9466a <=( (not A266)  and  (not A265) );
 a9470a <=( A300  and  A298 );
 a9471a <=( (not A268)  and  a9470a );
 a9472a <=( a9471a  and  a9466a );
 a9475a <=( (not A168)  and  (not A169) );
 a9479a <=( A199  and  A166 );
 a9480a <=( A167  and  a9479a );
 a9481a <=( a9480a  and  a9475a );
 a9484a <=( (not A267)  and  A201 );
 a9488a <=( A301  and  (not A269) );
 a9489a <=( (not A268)  and  a9488a );
 a9490a <=( a9489a  and  a9484a );
 a9493a <=( (not A168)  and  (not A169) );
 a9497a <=( A199  and  A166 );
 a9498a <=( A167  and  a9497a );
 a9499a <=( a9498a  and  a9493a );
 a9502a <=( (not A265)  and  A201 );
 a9506a <=( A301  and  (not A268) );
 a9507a <=( (not A266)  and  a9506a );
 a9508a <=( a9507a  and  a9502a );
 a9511a <=( (not A168)  and  (not A169) );
 a9515a <=( A200  and  A166 );
 a9516a <=( A167  and  a9515a );
 a9517a <=( a9516a  and  a9511a );
 a9520a <=( (not A267)  and  A201 );
 a9524a <=( A301  and  (not A269) );
 a9525a <=( (not A268)  and  a9524a );
 a9526a <=( a9525a  and  a9520a );
 a9529a <=( (not A168)  and  (not A169) );
 a9533a <=( A200  and  A166 );
 a9534a <=( A167  and  a9533a );
 a9535a <=( a9534a  and  a9529a );
 a9538a <=( (not A265)  and  A201 );
 a9542a <=( A301  and  (not A268) );
 a9543a <=( (not A266)  and  a9542a );
 a9544a <=( a9543a  and  a9538a );
 a9547a <=( (not A169)  and  (not A170) );
 a9551a <=( (not A267)  and  A202 );
 a9552a <=( (not A168)  and  a9551a );
 a9553a <=( a9552a  and  a9547a );
 a9556a <=( (not A269)  and  (not A268) );
 a9560a <=( A302  and  (not A299) );
 a9561a <=( A298  and  a9560a );
 a9562a <=( a9561a  and  a9556a );
 a9565a <=( (not A169)  and  (not A170) );
 a9569a <=( (not A267)  and  A202 );
 a9570a <=( (not A168)  and  a9569a );
 a9571a <=( a9570a  and  a9565a );
 a9574a <=( (not A269)  and  (not A268) );
 a9578a <=( A302  and  A299 );
 a9579a <=( (not A298)  and  a9578a );
 a9580a <=( a9579a  and  a9574a );
 a9583a <=( (not A169)  and  (not A170) );
 a9587a <=( A265  and  A202 );
 a9588a <=( (not A168)  and  a9587a );
 a9589a <=( a9588a  and  a9583a );
 a9592a <=( (not A267)  and  A266 );
 a9596a <=( A300  and  A299 );
 a9597a <=( (not A268)  and  a9596a );
 a9598a <=( a9597a  and  a9592a );
 a9601a <=( (not A169)  and  (not A170) );
 a9605a <=( A265  and  A202 );
 a9606a <=( (not A168)  and  a9605a );
 a9607a <=( a9606a  and  a9601a );
 a9610a <=( (not A267)  and  A266 );
 a9614a <=( A300  and  A298 );
 a9615a <=( (not A268)  and  a9614a );
 a9616a <=( a9615a  and  a9610a );
 a9619a <=( (not A169)  and  (not A170) );
 a9623a <=( (not A265)  and  A202 );
 a9624a <=( (not A168)  and  a9623a );
 a9625a <=( a9624a  and  a9619a );
 a9628a <=( (not A268)  and  (not A266) );
 a9632a <=( A302  and  (not A299) );
 a9633a <=( A298  and  a9632a );
 a9634a <=( a9633a  and  a9628a );
 a9637a <=( (not A169)  and  (not A170) );
 a9641a <=( (not A265)  and  A202 );
 a9642a <=( (not A168)  and  a9641a );
 a9643a <=( a9642a  and  a9637a );
 a9646a <=( (not A268)  and  (not A266) );
 a9650a <=( A302  and  A299 );
 a9651a <=( (not A298)  and  a9650a );
 a9652a <=( a9651a  and  a9646a );
 a9655a <=( (not A169)  and  (not A170) );
 a9659a <=( (not A202)  and  (not A201) );
 a9660a <=( (not A168)  and  a9659a );
 a9661a <=( a9660a  and  a9655a );
 a9664a <=( A268  and  (not A203) );
 a9668a <=( (not A302)  and  (not A301) );
 a9669a <=( (not A300)  and  a9668a );
 a9670a <=( a9669a  and  a9664a );
 a9673a <=( (not A169)  and  (not A170) );
 a9677a <=( (not A202)  and  (not A201) );
 a9678a <=( (not A168)  and  a9677a );
 a9679a <=( a9678a  and  a9673a );
 a9682a <=( A268  and  (not A203) );
 a9686a <=( (not A301)  and  (not A299) );
 a9687a <=( (not A298)  and  a9686a );
 a9688a <=( a9687a  and  a9682a );
 a9691a <=( (not A169)  and  (not A170) );
 a9695a <=( A201  and  A199 );
 a9696a <=( (not A168)  and  a9695a );
 a9697a <=( a9696a  and  a9691a );
 a9700a <=( (not A268)  and  (not A267) );
 a9704a <=( A300  and  A299 );
 a9705a <=( (not A269)  and  a9704a );
 a9706a <=( a9705a  and  a9700a );
 a9709a <=( (not A169)  and  (not A170) );
 a9713a <=( A201  and  A199 );
 a9714a <=( (not A168)  and  a9713a );
 a9715a <=( a9714a  and  a9709a );
 a9718a <=( (not A268)  and  (not A267) );
 a9722a <=( A300  and  A298 );
 a9723a <=( (not A269)  and  a9722a );
 a9724a <=( a9723a  and  a9718a );
 a9727a <=( (not A169)  and  (not A170) );
 a9731a <=( A201  and  A199 );
 a9732a <=( (not A168)  and  a9731a );
 a9733a <=( a9732a  and  a9727a );
 a9736a <=( A266  and  A265 );
 a9740a <=( A301  and  (not A268) );
 a9741a <=( (not A267)  and  a9740a );
 a9742a <=( a9741a  and  a9736a );
 a9745a <=( (not A169)  and  (not A170) );
 a9749a <=( A201  and  A199 );
 a9750a <=( (not A168)  and  a9749a );
 a9751a <=( a9750a  and  a9745a );
 a9754a <=( (not A266)  and  (not A265) );
 a9758a <=( A300  and  A299 );
 a9759a <=( (not A268)  and  a9758a );
 a9760a <=( a9759a  and  a9754a );
 a9763a <=( (not A169)  and  (not A170) );
 a9767a <=( A201  and  A199 );
 a9768a <=( (not A168)  and  a9767a );
 a9769a <=( a9768a  and  a9763a );
 a9772a <=( (not A266)  and  (not A265) );
 a9776a <=( A300  and  A298 );
 a9777a <=( (not A268)  and  a9776a );
 a9778a <=( a9777a  and  a9772a );
 a9781a <=( (not A169)  and  (not A170) );
 a9785a <=( A201  and  A200 );
 a9786a <=( (not A168)  and  a9785a );
 a9787a <=( a9786a  and  a9781a );
 a9790a <=( (not A268)  and  (not A267) );
 a9794a <=( A300  and  A299 );
 a9795a <=( (not A269)  and  a9794a );
 a9796a <=( a9795a  and  a9790a );
 a9799a <=( (not A169)  and  (not A170) );
 a9803a <=( A201  and  A200 );
 a9804a <=( (not A168)  and  a9803a );
 a9805a <=( a9804a  and  a9799a );
 a9808a <=( (not A268)  and  (not A267) );
 a9812a <=( A300  and  A298 );
 a9813a <=( (not A269)  and  a9812a );
 a9814a <=( a9813a  and  a9808a );
 a9817a <=( (not A169)  and  (not A170) );
 a9821a <=( A201  and  A200 );
 a9822a <=( (not A168)  and  a9821a );
 a9823a <=( a9822a  and  a9817a );
 a9826a <=( A266  and  A265 );
 a9830a <=( A301  and  (not A268) );
 a9831a <=( (not A267)  and  a9830a );
 a9832a <=( a9831a  and  a9826a );
 a9835a <=( (not A169)  and  (not A170) );
 a9839a <=( A201  and  A200 );
 a9840a <=( (not A168)  and  a9839a );
 a9841a <=( a9840a  and  a9835a );
 a9844a <=( (not A266)  and  (not A265) );
 a9848a <=( A300  and  A299 );
 a9849a <=( (not A268)  and  a9848a );
 a9850a <=( a9849a  and  a9844a );
 a9853a <=( (not A169)  and  (not A170) );
 a9857a <=( A201  and  A200 );
 a9858a <=( (not A168)  and  a9857a );
 a9859a <=( a9858a  and  a9853a );
 a9862a <=( (not A266)  and  (not A265) );
 a9866a <=( A300  and  A298 );
 a9867a <=( (not A268)  and  a9866a );
 a9868a <=( a9867a  and  a9862a );
 a9871a <=( (not A169)  and  (not A170) );
 a9875a <=( A200  and  (not A199) );
 a9876a <=( (not A168)  and  a9875a );
 a9877a <=( a9876a  and  a9871a );
 a9880a <=( (not A267)  and  A203 );
 a9884a <=( A301  and  (not A269) );
 a9885a <=( (not A268)  and  a9884a );
 a9886a <=( a9885a  and  a9880a );
 a9889a <=( (not A169)  and  (not A170) );
 a9893a <=( A200  and  (not A199) );
 a9894a <=( (not A168)  and  a9893a );
 a9895a <=( a9894a  and  a9889a );
 a9898a <=( (not A265)  and  A203 );
 a9902a <=( A301  and  (not A268) );
 a9903a <=( (not A266)  and  a9902a );
 a9904a <=( a9903a  and  a9898a );
 a9907a <=( (not A169)  and  (not A170) );
 a9911a <=( (not A200)  and  A199 );
 a9912a <=( (not A168)  and  a9911a );
 a9913a <=( a9912a  and  a9907a );
 a9916a <=( (not A267)  and  A203 );
 a9920a <=( A301  and  (not A269) );
 a9921a <=( (not A268)  and  a9920a );
 a9922a <=( a9921a  and  a9916a );
 a9925a <=( (not A169)  and  (not A170) );
 a9929a <=( (not A200)  and  A199 );
 a9930a <=( (not A168)  and  a9929a );
 a9931a <=( a9930a  and  a9925a );
 a9934a <=( (not A265)  and  A203 );
 a9938a <=( A301  and  (not A268) );
 a9939a <=( (not A266)  and  a9938a );
 a9940a <=( a9939a  and  a9934a );
 a9943a <=( (not A169)  and  (not A170) );
 a9947a <=( (not A200)  and  (not A199) );
 a9948a <=( (not A168)  and  a9947a );
 a9949a <=( a9948a  and  a9943a );
 a9952a <=( A268  and  (not A202) );
 a9956a <=( (not A302)  and  (not A301) );
 a9957a <=( (not A300)  and  a9956a );
 a9958a <=( a9957a  and  a9952a );
 a9961a <=( (not A169)  and  (not A170) );
 a9965a <=( (not A200)  and  (not A199) );
 a9966a <=( (not A168)  and  a9965a );
 a9967a <=( a9966a  and  a9961a );
 a9970a <=( A268  and  (not A202) );
 a9974a <=( (not A301)  and  (not A299) );
 a9975a <=( (not A298)  and  a9974a );
 a9976a <=( a9975a  and  a9970a );
 a9979a <=( A166  and  A168 );
 a9983a <=( (not A203)  and  (not A202) );
 a9984a <=( (not A201)  and  a9983a );
 a9985a <=( a9984a  and  a9979a );
 a9989a <=( (not A269)  and  (not A268) );
 a9990a <=( (not A267)  and  a9989a );
 a9994a <=( A302  and  (not A299) );
 a9995a <=( A298  and  a9994a );
 a9996a <=( a9995a  and  a9990a );
 a9999a <=( A166  and  A168 );
 a10003a <=( (not A203)  and  (not A202) );
 a10004a <=( (not A201)  and  a10003a );
 a10005a <=( a10004a  and  a9999a );
 a10009a <=( (not A269)  and  (not A268) );
 a10010a <=( (not A267)  and  a10009a );
 a10014a <=( A302  and  A299 );
 a10015a <=( (not A298)  and  a10014a );
 a10016a <=( a10015a  and  a10010a );
 a10019a <=( A166  and  A168 );
 a10023a <=( (not A203)  and  (not A202) );
 a10024a <=( (not A201)  and  a10023a );
 a10025a <=( a10024a  and  a10019a );
 a10029a <=( (not A267)  and  A266 );
 a10030a <=( A265  and  a10029a );
 a10034a <=( A300  and  A299 );
 a10035a <=( (not A268)  and  a10034a );
 a10036a <=( a10035a  and  a10030a );
 a10039a <=( A166  and  A168 );
 a10043a <=( (not A203)  and  (not A202) );
 a10044a <=( (not A201)  and  a10043a );
 a10045a <=( a10044a  and  a10039a );
 a10049a <=( (not A267)  and  A266 );
 a10050a <=( A265  and  a10049a );
 a10054a <=( A300  and  A298 );
 a10055a <=( (not A268)  and  a10054a );
 a10056a <=( a10055a  and  a10050a );
 a10059a <=( A166  and  A168 );
 a10063a <=( (not A203)  and  (not A202) );
 a10064a <=( (not A201)  and  a10063a );
 a10065a <=( a10064a  and  a10059a );
 a10069a <=( (not A268)  and  (not A266) );
 a10070a <=( (not A265)  and  a10069a );
 a10074a <=( A302  and  (not A299) );
 a10075a <=( A298  and  a10074a );
 a10076a <=( a10075a  and  a10070a );
 a10079a <=( A166  and  A168 );
 a10083a <=( (not A203)  and  (not A202) );
 a10084a <=( (not A201)  and  a10083a );
 a10085a <=( a10084a  and  a10079a );
 a10089a <=( (not A268)  and  (not A266) );
 a10090a <=( (not A265)  and  a10089a );
 a10094a <=( A302  and  A299 );
 a10095a <=( (not A298)  and  a10094a );
 a10096a <=( a10095a  and  a10090a );
 a10099a <=( A166  and  A168 );
 a10103a <=( (not A265)  and  A201 );
 a10104a <=( A199  and  a10103a );
 a10105a <=( a10104a  and  a10099a );
 a10109a <=( A298  and  A269 );
 a10110a <=( A266  and  a10109a );
 a10114a <=( (not A301)  and  (not A300) );
 a10115a <=( A299  and  a10114a );
 a10116a <=( a10115a  and  a10110a );
 a10119a <=( A166  and  A168 );
 a10123a <=( A265  and  A201 );
 a10124a <=( A199  and  a10123a );
 a10125a <=( a10124a  and  a10119a );
 a10129a <=( A298  and  A269 );
 a10130a <=( (not A266)  and  a10129a );
 a10134a <=( (not A301)  and  (not A300) );
 a10135a <=( A299  and  a10134a );
 a10136a <=( a10135a  and  a10130a );
 a10139a <=( A166  and  A168 );
 a10143a <=( (not A265)  and  A201 );
 a10144a <=( A200  and  a10143a );
 a10145a <=( a10144a  and  a10139a );
 a10149a <=( A298  and  A269 );
 a10150a <=( A266  and  a10149a );
 a10154a <=( (not A301)  and  (not A300) );
 a10155a <=( A299  and  a10154a );
 a10156a <=( a10155a  and  a10150a );
 a10159a <=( A166  and  A168 );
 a10163a <=( A265  and  A201 );
 a10164a <=( A200  and  a10163a );
 a10165a <=( a10164a  and  a10159a );
 a10169a <=( A298  and  A269 );
 a10170a <=( (not A266)  and  a10169a );
 a10174a <=( (not A301)  and  (not A300) );
 a10175a <=( A299  and  a10174a );
 a10176a <=( a10175a  and  a10170a );
 a10179a <=( A166  and  A168 );
 a10183a <=( (not A201)  and  A200 );
 a10184a <=( A199  and  a10183a );
 a10185a <=( a10184a  and  a10179a );
 a10189a <=( (not A268)  and  (not A267) );
 a10190a <=( (not A202)  and  a10189a );
 a10194a <=( A300  and  A299 );
 a10195a <=( (not A269)  and  a10194a );
 a10196a <=( a10195a  and  a10190a );
 a10199a <=( A166  and  A168 );
 a10203a <=( (not A201)  and  A200 );
 a10204a <=( A199  and  a10203a );
 a10205a <=( a10204a  and  a10199a );
 a10209a <=( (not A268)  and  (not A267) );
 a10210a <=( (not A202)  and  a10209a );
 a10214a <=( A300  and  A298 );
 a10215a <=( (not A269)  and  a10214a );
 a10216a <=( a10215a  and  a10210a );
 a10219a <=( A166  and  A168 );
 a10223a <=( (not A201)  and  A200 );
 a10224a <=( A199  and  a10223a );
 a10225a <=( a10224a  and  a10219a );
 a10229a <=( A266  and  A265 );
 a10230a <=( (not A202)  and  a10229a );
 a10234a <=( A301  and  (not A268) );
 a10235a <=( (not A267)  and  a10234a );
 a10236a <=( a10235a  and  a10230a );
 a10239a <=( A166  and  A168 );
 a10243a <=( (not A201)  and  A200 );
 a10244a <=( A199  and  a10243a );
 a10245a <=( a10244a  and  a10239a );
 a10249a <=( (not A266)  and  (not A265) );
 a10250a <=( (not A202)  and  a10249a );
 a10254a <=( A300  and  A299 );
 a10255a <=( (not A268)  and  a10254a );
 a10256a <=( a10255a  and  a10250a );
 a10259a <=( A166  and  A168 );
 a10263a <=( (not A201)  and  A200 );
 a10264a <=( A199  and  a10263a );
 a10265a <=( a10264a  and  a10259a );
 a10269a <=( (not A266)  and  (not A265) );
 a10270a <=( (not A202)  and  a10269a );
 a10274a <=( A300  and  A298 );
 a10275a <=( (not A268)  and  a10274a );
 a10276a <=( a10275a  and  a10270a );
 a10279a <=( A166  and  A168 );
 a10283a <=( A203  and  A200 );
 a10284a <=( (not A199)  and  a10283a );
 a10285a <=( a10284a  and  a10279a );
 a10289a <=( A298  and  A267 );
 a10290a <=( A265  and  a10289a );
 a10294a <=( (not A301)  and  (not A300) );
 a10295a <=( A299  and  a10294a );
 a10296a <=( a10295a  and  a10290a );
 a10299a <=( A166  and  A168 );
 a10303a <=( A203  and  A200 );
 a10304a <=( (not A199)  and  a10303a );
 a10305a <=( a10304a  and  a10299a );
 a10309a <=( A298  and  A267 );
 a10310a <=( A266  and  a10309a );
 a10314a <=( (not A301)  and  (not A300) );
 a10315a <=( A299  and  a10314a );
 a10316a <=( a10315a  and  a10310a );
 a10319a <=( A166  and  A168 );
 a10323a <=( A203  and  A200 );
 a10324a <=( (not A199)  and  a10323a );
 a10325a <=( a10324a  and  a10319a );
 a10329a <=( A269  and  A266 );
 a10330a <=( (not A265)  and  a10329a );
 a10334a <=( (not A302)  and  (not A301) );
 a10335a <=( (not A300)  and  a10334a );
 a10336a <=( a10335a  and  a10330a );
 a10339a <=( A166  and  A168 );
 a10343a <=( A203  and  A200 );
 a10344a <=( (not A199)  and  a10343a );
 a10345a <=( a10344a  and  a10339a );
 a10349a <=( A269  and  A266 );
 a10350a <=( (not A265)  and  a10349a );
 a10354a <=( (not A301)  and  (not A299) );
 a10355a <=( (not A298)  and  a10354a );
 a10356a <=( a10355a  and  a10350a );
 a10359a <=( A166  and  A168 );
 a10363a <=( A203  and  A200 );
 a10364a <=( (not A199)  and  a10363a );
 a10365a <=( a10364a  and  a10359a );
 a10369a <=( A269  and  (not A266) );
 a10370a <=( A265  and  a10369a );
 a10374a <=( (not A302)  and  (not A301) );
 a10375a <=( (not A300)  and  a10374a );
 a10376a <=( a10375a  and  a10370a );
 a10379a <=( A166  and  A168 );
 a10383a <=( A203  and  A200 );
 a10384a <=( (not A199)  and  a10383a );
 a10385a <=( a10384a  and  a10379a );
 a10389a <=( A269  and  (not A266) );
 a10390a <=( A265  and  a10389a );
 a10394a <=( (not A301)  and  (not A299) );
 a10395a <=( (not A298)  and  a10394a );
 a10396a <=( a10395a  and  a10390a );
 a10399a <=( A166  and  A168 );
 a10403a <=( A203  and  (not A200) );
 a10404a <=( A199  and  a10403a );
 a10405a <=( a10404a  and  a10399a );
 a10409a <=( A298  and  A267 );
 a10410a <=( A265  and  a10409a );
 a10414a <=( (not A301)  and  (not A300) );
 a10415a <=( A299  and  a10414a );
 a10416a <=( a10415a  and  a10410a );
 a10419a <=( A166  and  A168 );
 a10423a <=( A203  and  (not A200) );
 a10424a <=( A199  and  a10423a );
 a10425a <=( a10424a  and  a10419a );
 a10429a <=( A298  and  A267 );
 a10430a <=( A266  and  a10429a );
 a10434a <=( (not A301)  and  (not A300) );
 a10435a <=( A299  and  a10434a );
 a10436a <=( a10435a  and  a10430a );
 a10439a <=( A166  and  A168 );
 a10443a <=( A203  and  (not A200) );
 a10444a <=( A199  and  a10443a );
 a10445a <=( a10444a  and  a10439a );
 a10449a <=( A269  and  A266 );
 a10450a <=( (not A265)  and  a10449a );
 a10454a <=( (not A302)  and  (not A301) );
 a10455a <=( (not A300)  and  a10454a );
 a10456a <=( a10455a  and  a10450a );
 a10459a <=( A166  and  A168 );
 a10463a <=( A203  and  (not A200) );
 a10464a <=( A199  and  a10463a );
 a10465a <=( a10464a  and  a10459a );
 a10469a <=( A269  and  A266 );
 a10470a <=( (not A265)  and  a10469a );
 a10474a <=( (not A301)  and  (not A299) );
 a10475a <=( (not A298)  and  a10474a );
 a10476a <=( a10475a  and  a10470a );
 a10479a <=( A166  and  A168 );
 a10483a <=( A203  and  (not A200) );
 a10484a <=( A199  and  a10483a );
 a10485a <=( a10484a  and  a10479a );
 a10489a <=( A269  and  (not A266) );
 a10490a <=( A265  and  a10489a );
 a10494a <=( (not A302)  and  (not A301) );
 a10495a <=( (not A300)  and  a10494a );
 a10496a <=( a10495a  and  a10490a );
 a10499a <=( A166  and  A168 );
 a10503a <=( A203  and  (not A200) );
 a10504a <=( A199  and  a10503a );
 a10505a <=( a10504a  and  a10499a );
 a10509a <=( A269  and  (not A266) );
 a10510a <=( A265  and  a10509a );
 a10514a <=( (not A301)  and  (not A299) );
 a10515a <=( (not A298)  and  a10514a );
 a10516a <=( a10515a  and  a10510a );
 a10519a <=( A166  and  A168 );
 a10523a <=( (not A202)  and  (not A200) );
 a10524a <=( (not A199)  and  a10523a );
 a10525a <=( a10524a  and  a10519a );
 a10529a <=( (not A269)  and  (not A268) );
 a10530a <=( (not A267)  and  a10529a );
 a10534a <=( A302  and  (not A299) );
 a10535a <=( A298  and  a10534a );
 a10536a <=( a10535a  and  a10530a );
 a10539a <=( A166  and  A168 );
 a10543a <=( (not A202)  and  (not A200) );
 a10544a <=( (not A199)  and  a10543a );
 a10545a <=( a10544a  and  a10539a );
 a10549a <=( (not A269)  and  (not A268) );
 a10550a <=( (not A267)  and  a10549a );
 a10554a <=( A302  and  A299 );
 a10555a <=( (not A298)  and  a10554a );
 a10556a <=( a10555a  and  a10550a );
 a10559a <=( A166  and  A168 );
 a10563a <=( (not A202)  and  (not A200) );
 a10564a <=( (not A199)  and  a10563a );
 a10565a <=( a10564a  and  a10559a );
 a10569a <=( (not A267)  and  A266 );
 a10570a <=( A265  and  a10569a );
 a10574a <=( A300  and  A299 );
 a10575a <=( (not A268)  and  a10574a );
 a10576a <=( a10575a  and  a10570a );
 a10579a <=( A166  and  A168 );
 a10583a <=( (not A202)  and  (not A200) );
 a10584a <=( (not A199)  and  a10583a );
 a10585a <=( a10584a  and  a10579a );
 a10589a <=( (not A267)  and  A266 );
 a10590a <=( A265  and  a10589a );
 a10594a <=( A300  and  A298 );
 a10595a <=( (not A268)  and  a10594a );
 a10596a <=( a10595a  and  a10590a );
 a10599a <=( A166  and  A168 );
 a10603a <=( (not A202)  and  (not A200) );
 a10604a <=( (not A199)  and  a10603a );
 a10605a <=( a10604a  and  a10599a );
 a10609a <=( (not A268)  and  (not A266) );
 a10610a <=( (not A265)  and  a10609a );
 a10614a <=( A302  and  (not A299) );
 a10615a <=( A298  and  a10614a );
 a10616a <=( a10615a  and  a10610a );
 a10619a <=( A166  and  A168 );
 a10623a <=( (not A202)  and  (not A200) );
 a10624a <=( (not A199)  and  a10623a );
 a10625a <=( a10624a  and  a10619a );
 a10629a <=( (not A268)  and  (not A266) );
 a10630a <=( (not A265)  and  a10629a );
 a10634a <=( A302  and  A299 );
 a10635a <=( (not A298)  and  a10634a );
 a10636a <=( a10635a  and  a10630a );
 a10639a <=( A167  and  A168 );
 a10643a <=( (not A203)  and  (not A202) );
 a10644a <=( (not A201)  and  a10643a );
 a10645a <=( a10644a  and  a10639a );
 a10649a <=( (not A269)  and  (not A268) );
 a10650a <=( (not A267)  and  a10649a );
 a10654a <=( A302  and  (not A299) );
 a10655a <=( A298  and  a10654a );
 a10656a <=( a10655a  and  a10650a );
 a10659a <=( A167  and  A168 );
 a10663a <=( (not A203)  and  (not A202) );
 a10664a <=( (not A201)  and  a10663a );
 a10665a <=( a10664a  and  a10659a );
 a10669a <=( (not A269)  and  (not A268) );
 a10670a <=( (not A267)  and  a10669a );
 a10674a <=( A302  and  A299 );
 a10675a <=( (not A298)  and  a10674a );
 a10676a <=( a10675a  and  a10670a );
 a10679a <=( A167  and  A168 );
 a10683a <=( (not A203)  and  (not A202) );
 a10684a <=( (not A201)  and  a10683a );
 a10685a <=( a10684a  and  a10679a );
 a10689a <=( (not A267)  and  A266 );
 a10690a <=( A265  and  a10689a );
 a10694a <=( A300  and  A299 );
 a10695a <=( (not A268)  and  a10694a );
 a10696a <=( a10695a  and  a10690a );
 a10699a <=( A167  and  A168 );
 a10703a <=( (not A203)  and  (not A202) );
 a10704a <=( (not A201)  and  a10703a );
 a10705a <=( a10704a  and  a10699a );
 a10709a <=( (not A267)  and  A266 );
 a10710a <=( A265  and  a10709a );
 a10714a <=( A300  and  A298 );
 a10715a <=( (not A268)  and  a10714a );
 a10716a <=( a10715a  and  a10710a );
 a10719a <=( A167  and  A168 );
 a10723a <=( (not A203)  and  (not A202) );
 a10724a <=( (not A201)  and  a10723a );
 a10725a <=( a10724a  and  a10719a );
 a10729a <=( (not A268)  and  (not A266) );
 a10730a <=( (not A265)  and  a10729a );
 a10734a <=( A302  and  (not A299) );
 a10735a <=( A298  and  a10734a );
 a10736a <=( a10735a  and  a10730a );
 a10739a <=( A167  and  A168 );
 a10743a <=( (not A203)  and  (not A202) );
 a10744a <=( (not A201)  and  a10743a );
 a10745a <=( a10744a  and  a10739a );
 a10749a <=( (not A268)  and  (not A266) );
 a10750a <=( (not A265)  and  a10749a );
 a10754a <=( A302  and  A299 );
 a10755a <=( (not A298)  and  a10754a );
 a10756a <=( a10755a  and  a10750a );
 a10759a <=( A167  and  A168 );
 a10763a <=( (not A265)  and  A201 );
 a10764a <=( A199  and  a10763a );
 a10765a <=( a10764a  and  a10759a );
 a10769a <=( A298  and  A269 );
 a10770a <=( A266  and  a10769a );
 a10774a <=( (not A301)  and  (not A300) );
 a10775a <=( A299  and  a10774a );
 a10776a <=( a10775a  and  a10770a );
 a10779a <=( A167  and  A168 );
 a10783a <=( A265  and  A201 );
 a10784a <=( A199  and  a10783a );
 a10785a <=( a10784a  and  a10779a );
 a10789a <=( A298  and  A269 );
 a10790a <=( (not A266)  and  a10789a );
 a10794a <=( (not A301)  and  (not A300) );
 a10795a <=( A299  and  a10794a );
 a10796a <=( a10795a  and  a10790a );
 a10799a <=( A167  and  A168 );
 a10803a <=( (not A265)  and  A201 );
 a10804a <=( A200  and  a10803a );
 a10805a <=( a10804a  and  a10799a );
 a10809a <=( A298  and  A269 );
 a10810a <=( A266  and  a10809a );
 a10814a <=( (not A301)  and  (not A300) );
 a10815a <=( A299  and  a10814a );
 a10816a <=( a10815a  and  a10810a );
 a10819a <=( A167  and  A168 );
 a10823a <=( A265  and  A201 );
 a10824a <=( A200  and  a10823a );
 a10825a <=( a10824a  and  a10819a );
 a10829a <=( A298  and  A269 );
 a10830a <=( (not A266)  and  a10829a );
 a10834a <=( (not A301)  and  (not A300) );
 a10835a <=( A299  and  a10834a );
 a10836a <=( a10835a  and  a10830a );
 a10839a <=( A167  and  A168 );
 a10843a <=( (not A201)  and  A200 );
 a10844a <=( A199  and  a10843a );
 a10845a <=( a10844a  and  a10839a );
 a10849a <=( (not A268)  and  (not A267) );
 a10850a <=( (not A202)  and  a10849a );
 a10854a <=( A300  and  A299 );
 a10855a <=( (not A269)  and  a10854a );
 a10856a <=( a10855a  and  a10850a );
 a10859a <=( A167  and  A168 );
 a10863a <=( (not A201)  and  A200 );
 a10864a <=( A199  and  a10863a );
 a10865a <=( a10864a  and  a10859a );
 a10869a <=( (not A268)  and  (not A267) );
 a10870a <=( (not A202)  and  a10869a );
 a10874a <=( A300  and  A298 );
 a10875a <=( (not A269)  and  a10874a );
 a10876a <=( a10875a  and  a10870a );
 a10879a <=( A167  and  A168 );
 a10883a <=( (not A201)  and  A200 );
 a10884a <=( A199  and  a10883a );
 a10885a <=( a10884a  and  a10879a );
 a10889a <=( A266  and  A265 );
 a10890a <=( (not A202)  and  a10889a );
 a10894a <=( A301  and  (not A268) );
 a10895a <=( (not A267)  and  a10894a );
 a10896a <=( a10895a  and  a10890a );
 a10899a <=( A167  and  A168 );
 a10903a <=( (not A201)  and  A200 );
 a10904a <=( A199  and  a10903a );
 a10905a <=( a10904a  and  a10899a );
 a10909a <=( (not A266)  and  (not A265) );
 a10910a <=( (not A202)  and  a10909a );
 a10914a <=( A300  and  A299 );
 a10915a <=( (not A268)  and  a10914a );
 a10916a <=( a10915a  and  a10910a );
 a10919a <=( A167  and  A168 );
 a10923a <=( (not A201)  and  A200 );
 a10924a <=( A199  and  a10923a );
 a10925a <=( a10924a  and  a10919a );
 a10929a <=( (not A266)  and  (not A265) );
 a10930a <=( (not A202)  and  a10929a );
 a10934a <=( A300  and  A298 );
 a10935a <=( (not A268)  and  a10934a );
 a10936a <=( a10935a  and  a10930a );
 a10939a <=( A167  and  A168 );
 a10943a <=( A203  and  A200 );
 a10944a <=( (not A199)  and  a10943a );
 a10945a <=( a10944a  and  a10939a );
 a10949a <=( A298  and  A267 );
 a10950a <=( A265  and  a10949a );
 a10954a <=( (not A301)  and  (not A300) );
 a10955a <=( A299  and  a10954a );
 a10956a <=( a10955a  and  a10950a );
 a10959a <=( A167  and  A168 );
 a10963a <=( A203  and  A200 );
 a10964a <=( (not A199)  and  a10963a );
 a10965a <=( a10964a  and  a10959a );
 a10969a <=( A298  and  A267 );
 a10970a <=( A266  and  a10969a );
 a10974a <=( (not A301)  and  (not A300) );
 a10975a <=( A299  and  a10974a );
 a10976a <=( a10975a  and  a10970a );
 a10979a <=( A167  and  A168 );
 a10983a <=( A203  and  A200 );
 a10984a <=( (not A199)  and  a10983a );
 a10985a <=( a10984a  and  a10979a );
 a10989a <=( A269  and  A266 );
 a10990a <=( (not A265)  and  a10989a );
 a10994a <=( (not A302)  and  (not A301) );
 a10995a <=( (not A300)  and  a10994a );
 a10996a <=( a10995a  and  a10990a );
 a10999a <=( A167  and  A168 );
 a11003a <=( A203  and  A200 );
 a11004a <=( (not A199)  and  a11003a );
 a11005a <=( a11004a  and  a10999a );
 a11009a <=( A269  and  A266 );
 a11010a <=( (not A265)  and  a11009a );
 a11014a <=( (not A301)  and  (not A299) );
 a11015a <=( (not A298)  and  a11014a );
 a11016a <=( a11015a  and  a11010a );
 a11019a <=( A167  and  A168 );
 a11023a <=( A203  and  A200 );
 a11024a <=( (not A199)  and  a11023a );
 a11025a <=( a11024a  and  a11019a );
 a11029a <=( A269  and  (not A266) );
 a11030a <=( A265  and  a11029a );
 a11034a <=( (not A302)  and  (not A301) );
 a11035a <=( (not A300)  and  a11034a );
 a11036a <=( a11035a  and  a11030a );
 a11039a <=( A167  and  A168 );
 a11043a <=( A203  and  A200 );
 a11044a <=( (not A199)  and  a11043a );
 a11045a <=( a11044a  and  a11039a );
 a11049a <=( A269  and  (not A266) );
 a11050a <=( A265  and  a11049a );
 a11054a <=( (not A301)  and  (not A299) );
 a11055a <=( (not A298)  and  a11054a );
 a11056a <=( a11055a  and  a11050a );
 a11059a <=( A167  and  A168 );
 a11063a <=( A203  and  (not A200) );
 a11064a <=( A199  and  a11063a );
 a11065a <=( a11064a  and  a11059a );
 a11069a <=( A298  and  A267 );
 a11070a <=( A265  and  a11069a );
 a11074a <=( (not A301)  and  (not A300) );
 a11075a <=( A299  and  a11074a );
 a11076a <=( a11075a  and  a11070a );
 a11079a <=( A167  and  A168 );
 a11083a <=( A203  and  (not A200) );
 a11084a <=( A199  and  a11083a );
 a11085a <=( a11084a  and  a11079a );
 a11089a <=( A298  and  A267 );
 a11090a <=( A266  and  a11089a );
 a11094a <=( (not A301)  and  (not A300) );
 a11095a <=( A299  and  a11094a );
 a11096a <=( a11095a  and  a11090a );
 a11099a <=( A167  and  A168 );
 a11103a <=( A203  and  (not A200) );
 a11104a <=( A199  and  a11103a );
 a11105a <=( a11104a  and  a11099a );
 a11109a <=( A269  and  A266 );
 a11110a <=( (not A265)  and  a11109a );
 a11114a <=( (not A302)  and  (not A301) );
 a11115a <=( (not A300)  and  a11114a );
 a11116a <=( a11115a  and  a11110a );
 a11119a <=( A167  and  A168 );
 a11123a <=( A203  and  (not A200) );
 a11124a <=( A199  and  a11123a );
 a11125a <=( a11124a  and  a11119a );
 a11129a <=( A269  and  A266 );
 a11130a <=( (not A265)  and  a11129a );
 a11134a <=( (not A301)  and  (not A299) );
 a11135a <=( (not A298)  and  a11134a );
 a11136a <=( a11135a  and  a11130a );
 a11139a <=( A167  and  A168 );
 a11143a <=( A203  and  (not A200) );
 a11144a <=( A199  and  a11143a );
 a11145a <=( a11144a  and  a11139a );
 a11149a <=( A269  and  (not A266) );
 a11150a <=( A265  and  a11149a );
 a11154a <=( (not A302)  and  (not A301) );
 a11155a <=( (not A300)  and  a11154a );
 a11156a <=( a11155a  and  a11150a );
 a11159a <=( A167  and  A168 );
 a11163a <=( A203  and  (not A200) );
 a11164a <=( A199  and  a11163a );
 a11165a <=( a11164a  and  a11159a );
 a11169a <=( A269  and  (not A266) );
 a11170a <=( A265  and  a11169a );
 a11174a <=( (not A301)  and  (not A299) );
 a11175a <=( (not A298)  and  a11174a );
 a11176a <=( a11175a  and  a11170a );
 a11179a <=( A167  and  A168 );
 a11183a <=( (not A202)  and  (not A200) );
 a11184a <=( (not A199)  and  a11183a );
 a11185a <=( a11184a  and  a11179a );
 a11189a <=( (not A269)  and  (not A268) );
 a11190a <=( (not A267)  and  a11189a );
 a11194a <=( A302  and  (not A299) );
 a11195a <=( A298  and  a11194a );
 a11196a <=( a11195a  and  a11190a );
 a11199a <=( A167  and  A168 );
 a11203a <=( (not A202)  and  (not A200) );
 a11204a <=( (not A199)  and  a11203a );
 a11205a <=( a11204a  and  a11199a );
 a11209a <=( (not A269)  and  (not A268) );
 a11210a <=( (not A267)  and  a11209a );
 a11214a <=( A302  and  A299 );
 a11215a <=( (not A298)  and  a11214a );
 a11216a <=( a11215a  and  a11210a );
 a11219a <=( A167  and  A168 );
 a11223a <=( (not A202)  and  (not A200) );
 a11224a <=( (not A199)  and  a11223a );
 a11225a <=( a11224a  and  a11219a );
 a11229a <=( (not A267)  and  A266 );
 a11230a <=( A265  and  a11229a );
 a11234a <=( A300  and  A299 );
 a11235a <=( (not A268)  and  a11234a );
 a11236a <=( a11235a  and  a11230a );
 a11239a <=( A167  and  A168 );
 a11243a <=( (not A202)  and  (not A200) );
 a11244a <=( (not A199)  and  a11243a );
 a11245a <=( a11244a  and  a11239a );
 a11249a <=( (not A267)  and  A266 );
 a11250a <=( A265  and  a11249a );
 a11254a <=( A300  and  A298 );
 a11255a <=( (not A268)  and  a11254a );
 a11256a <=( a11255a  and  a11250a );
 a11259a <=( A167  and  A168 );
 a11263a <=( (not A202)  and  (not A200) );
 a11264a <=( (not A199)  and  a11263a );
 a11265a <=( a11264a  and  a11259a );
 a11269a <=( (not A268)  and  (not A266) );
 a11270a <=( (not A265)  and  a11269a );
 a11274a <=( A302  and  (not A299) );
 a11275a <=( A298  and  a11274a );
 a11276a <=( a11275a  and  a11270a );
 a11279a <=( A167  and  A168 );
 a11283a <=( (not A202)  and  (not A200) );
 a11284a <=( (not A199)  and  a11283a );
 a11285a <=( a11284a  and  a11279a );
 a11289a <=( (not A268)  and  (not A266) );
 a11290a <=( (not A265)  and  a11289a );
 a11294a <=( A302  and  A299 );
 a11295a <=( (not A298)  and  a11294a );
 a11296a <=( a11295a  and  a11290a );
 a11299a <=( A167  and  A170 );
 a11303a <=( (not A265)  and  A202 );
 a11304a <=( (not A166)  and  a11303a );
 a11305a <=( a11304a  and  a11299a );
 a11309a <=( A298  and  A269 );
 a11310a <=( A266  and  a11309a );
 a11314a <=( (not A301)  and  (not A300) );
 a11315a <=( A299  and  a11314a );
 a11316a <=( a11315a  and  a11310a );
 a11319a <=( A167  and  A170 );
 a11323a <=( A265  and  A202 );
 a11324a <=( (not A166)  and  a11323a );
 a11325a <=( a11324a  and  a11319a );
 a11329a <=( A298  and  A269 );
 a11330a <=( (not A266)  and  a11329a );
 a11334a <=( (not A301)  and  (not A300) );
 a11335a <=( A299  and  a11334a );
 a11336a <=( a11335a  and  a11330a );
 a11339a <=( A167  and  A170 );
 a11343a <=( (not A202)  and  (not A201) );
 a11344a <=( (not A166)  and  a11343a );
 a11345a <=( a11344a  and  a11339a );
 a11349a <=( (not A268)  and  (not A267) );
 a11350a <=( (not A203)  and  a11349a );
 a11354a <=( A300  and  A299 );
 a11355a <=( (not A269)  and  a11354a );
 a11356a <=( a11355a  and  a11350a );
 a11359a <=( A167  and  A170 );
 a11363a <=( (not A202)  and  (not A201) );
 a11364a <=( (not A166)  and  a11363a );
 a11365a <=( a11364a  and  a11359a );
 a11369a <=( (not A268)  and  (not A267) );
 a11370a <=( (not A203)  and  a11369a );
 a11374a <=( A300  and  A298 );
 a11375a <=( (not A269)  and  a11374a );
 a11376a <=( a11375a  and  a11370a );
 a11379a <=( A167  and  A170 );
 a11383a <=( (not A202)  and  (not A201) );
 a11384a <=( (not A166)  and  a11383a );
 a11385a <=( a11384a  and  a11379a );
 a11389a <=( A266  and  A265 );
 a11390a <=( (not A203)  and  a11389a );
 a11394a <=( A301  and  (not A268) );
 a11395a <=( (not A267)  and  a11394a );
 a11396a <=( a11395a  and  a11390a );
 a11399a <=( A167  and  A170 );
 a11403a <=( (not A202)  and  (not A201) );
 a11404a <=( (not A166)  and  a11403a );
 a11405a <=( a11404a  and  a11399a );
 a11409a <=( (not A266)  and  (not A265) );
 a11410a <=( (not A203)  and  a11409a );
 a11414a <=( A300  and  A299 );
 a11415a <=( (not A268)  and  a11414a );
 a11416a <=( a11415a  and  a11410a );
 a11419a <=( A167  and  A170 );
 a11423a <=( (not A202)  and  (not A201) );
 a11424a <=( (not A166)  and  a11423a );
 a11425a <=( a11424a  and  a11419a );
 a11429a <=( (not A266)  and  (not A265) );
 a11430a <=( (not A203)  and  a11429a );
 a11434a <=( A300  and  A298 );
 a11435a <=( (not A268)  and  a11434a );
 a11436a <=( a11435a  and  a11430a );
 a11439a <=( A167  and  A170 );
 a11443a <=( A201  and  A199 );
 a11444a <=( (not A166)  and  a11443a );
 a11445a <=( a11444a  and  a11439a );
 a11449a <=( A298  and  A267 );
 a11450a <=( A265  and  a11449a );
 a11454a <=( (not A301)  and  (not A300) );
 a11455a <=( A299  and  a11454a );
 a11456a <=( a11455a  and  a11450a );
 a11459a <=( A167  and  A170 );
 a11463a <=( A201  and  A199 );
 a11464a <=( (not A166)  and  a11463a );
 a11465a <=( a11464a  and  a11459a );
 a11469a <=( A298  and  A267 );
 a11470a <=( A266  and  a11469a );
 a11474a <=( (not A301)  and  (not A300) );
 a11475a <=( A299  and  a11474a );
 a11476a <=( a11475a  and  a11470a );
 a11479a <=( A167  and  A170 );
 a11483a <=( A201  and  A199 );
 a11484a <=( (not A166)  and  a11483a );
 a11485a <=( a11484a  and  a11479a );
 a11489a <=( A269  and  A266 );
 a11490a <=( (not A265)  and  a11489a );
 a11494a <=( (not A302)  and  (not A301) );
 a11495a <=( (not A300)  and  a11494a );
 a11496a <=( a11495a  and  a11490a );
 a11499a <=( A167  and  A170 );
 a11503a <=( A201  and  A199 );
 a11504a <=( (not A166)  and  a11503a );
 a11505a <=( a11504a  and  a11499a );
 a11509a <=( A269  and  A266 );
 a11510a <=( (not A265)  and  a11509a );
 a11514a <=( (not A301)  and  (not A299) );
 a11515a <=( (not A298)  and  a11514a );
 a11516a <=( a11515a  and  a11510a );
 a11519a <=( A167  and  A170 );
 a11523a <=( A201  and  A199 );
 a11524a <=( (not A166)  and  a11523a );
 a11525a <=( a11524a  and  a11519a );
 a11529a <=( A269  and  (not A266) );
 a11530a <=( A265  and  a11529a );
 a11534a <=( (not A302)  and  (not A301) );
 a11535a <=( (not A300)  and  a11534a );
 a11536a <=( a11535a  and  a11530a );
 a11539a <=( A167  and  A170 );
 a11543a <=( A201  and  A199 );
 a11544a <=( (not A166)  and  a11543a );
 a11545a <=( a11544a  and  a11539a );
 a11549a <=( A269  and  (not A266) );
 a11550a <=( A265  and  a11549a );
 a11554a <=( (not A301)  and  (not A299) );
 a11555a <=( (not A298)  and  a11554a );
 a11556a <=( a11555a  and  a11550a );
 a11559a <=( A167  and  A170 );
 a11563a <=( A201  and  A200 );
 a11564a <=( (not A166)  and  a11563a );
 a11565a <=( a11564a  and  a11559a );
 a11569a <=( A298  and  A267 );
 a11570a <=( A265  and  a11569a );
 a11574a <=( (not A301)  and  (not A300) );
 a11575a <=( A299  and  a11574a );
 a11576a <=( a11575a  and  a11570a );
 a11579a <=( A167  and  A170 );
 a11583a <=( A201  and  A200 );
 a11584a <=( (not A166)  and  a11583a );
 a11585a <=( a11584a  and  a11579a );
 a11589a <=( A298  and  A267 );
 a11590a <=( A266  and  a11589a );
 a11594a <=( (not A301)  and  (not A300) );
 a11595a <=( A299  and  a11594a );
 a11596a <=( a11595a  and  a11590a );
 a11599a <=( A167  and  A170 );
 a11603a <=( A201  and  A200 );
 a11604a <=( (not A166)  and  a11603a );
 a11605a <=( a11604a  and  a11599a );
 a11609a <=( A269  and  A266 );
 a11610a <=( (not A265)  and  a11609a );
 a11614a <=( (not A302)  and  (not A301) );
 a11615a <=( (not A300)  and  a11614a );
 a11616a <=( a11615a  and  a11610a );
 a11619a <=( A167  and  A170 );
 a11623a <=( A201  and  A200 );
 a11624a <=( (not A166)  and  a11623a );
 a11625a <=( a11624a  and  a11619a );
 a11629a <=( A269  and  A266 );
 a11630a <=( (not A265)  and  a11629a );
 a11634a <=( (not A301)  and  (not A299) );
 a11635a <=( (not A298)  and  a11634a );
 a11636a <=( a11635a  and  a11630a );
 a11639a <=( A167  and  A170 );
 a11643a <=( A201  and  A200 );
 a11644a <=( (not A166)  and  a11643a );
 a11645a <=( a11644a  and  a11639a );
 a11649a <=( A269  and  (not A266) );
 a11650a <=( A265  and  a11649a );
 a11654a <=( (not A302)  and  (not A301) );
 a11655a <=( (not A300)  and  a11654a );
 a11656a <=( a11655a  and  a11650a );
 a11659a <=( A167  and  A170 );
 a11663a <=( A201  and  A200 );
 a11664a <=( (not A166)  and  a11663a );
 a11665a <=( a11664a  and  a11659a );
 a11669a <=( A269  and  (not A266) );
 a11670a <=( A265  and  a11669a );
 a11674a <=( (not A301)  and  (not A299) );
 a11675a <=( (not A298)  and  a11674a );
 a11676a <=( a11675a  and  a11670a );
 a11679a <=( A167  and  A170 );
 a11683a <=( A200  and  A199 );
 a11684a <=( (not A166)  and  a11683a );
 a11685a <=( a11684a  and  a11679a );
 a11689a <=( (not A267)  and  (not A202) );
 a11690a <=( (not A201)  and  a11689a );
 a11694a <=( A301  and  (not A269) );
 a11695a <=( (not A268)  and  a11694a );
 a11696a <=( a11695a  and  a11690a );
 a11699a <=( A167  and  A170 );
 a11703a <=( A200  and  A199 );
 a11704a <=( (not A166)  and  a11703a );
 a11705a <=( a11704a  and  a11699a );
 a11709a <=( (not A265)  and  (not A202) );
 a11710a <=( (not A201)  and  a11709a );
 a11714a <=( A301  and  (not A268) );
 a11715a <=( (not A266)  and  a11714a );
 a11716a <=( a11715a  and  a11710a );
 a11719a <=( A167  and  A170 );
 a11723a <=( A200  and  (not A199) );
 a11724a <=( (not A166)  and  a11723a );
 a11725a <=( a11724a  and  a11719a );
 a11729a <=( A298  and  A268 );
 a11730a <=( A203  and  a11729a );
 a11734a <=( (not A301)  and  (not A300) );
 a11735a <=( A299  and  a11734a );
 a11736a <=( a11735a  and  a11730a );
 a11739a <=( A167  and  A170 );
 a11743a <=( A200  and  (not A199) );
 a11744a <=( (not A166)  and  a11743a );
 a11745a <=( a11744a  and  a11739a );
 a11749a <=( A267  and  A265 );
 a11750a <=( A203  and  a11749a );
 a11754a <=( (not A302)  and  (not A301) );
 a11755a <=( (not A300)  and  a11754a );
 a11756a <=( a11755a  and  a11750a );
 a11759a <=( A167  and  A170 );
 a11763a <=( A200  and  (not A199) );
 a11764a <=( (not A166)  and  a11763a );
 a11765a <=( a11764a  and  a11759a );
 a11769a <=( A267  and  A265 );
 a11770a <=( A203  and  a11769a );
 a11774a <=( (not A301)  and  (not A299) );
 a11775a <=( (not A298)  and  a11774a );
 a11776a <=( a11775a  and  a11770a );
 a11779a <=( A167  and  A170 );
 a11783a <=( A200  and  (not A199) );
 a11784a <=( (not A166)  and  a11783a );
 a11785a <=( a11784a  and  a11779a );
 a11789a <=( A267  and  A266 );
 a11790a <=( A203  and  a11789a );
 a11794a <=( (not A302)  and  (not A301) );
 a11795a <=( (not A300)  and  a11794a );
 a11796a <=( a11795a  and  a11790a );
 a11799a <=( A167  and  A170 );
 a11803a <=( A200  and  (not A199) );
 a11804a <=( (not A166)  and  a11803a );
 a11805a <=( a11804a  and  a11799a );
 a11809a <=( A267  and  A266 );
 a11810a <=( A203  and  a11809a );
 a11814a <=( (not A301)  and  (not A299) );
 a11815a <=( (not A298)  and  a11814a );
 a11816a <=( a11815a  and  a11810a );
 a11819a <=( A167  and  A170 );
 a11823a <=( (not A200)  and  A199 );
 a11824a <=( (not A166)  and  a11823a );
 a11825a <=( a11824a  and  a11819a );
 a11829a <=( A298  and  A268 );
 a11830a <=( A203  and  a11829a );
 a11834a <=( (not A301)  and  (not A300) );
 a11835a <=( A299  and  a11834a );
 a11836a <=( a11835a  and  a11830a );
 a11839a <=( A167  and  A170 );
 a11843a <=( (not A200)  and  A199 );
 a11844a <=( (not A166)  and  a11843a );
 a11845a <=( a11844a  and  a11839a );
 a11849a <=( A267  and  A265 );
 a11850a <=( A203  and  a11849a );
 a11854a <=( (not A302)  and  (not A301) );
 a11855a <=( (not A300)  and  a11854a );
 a11856a <=( a11855a  and  a11850a );
 a11859a <=( A167  and  A170 );
 a11863a <=( (not A200)  and  A199 );
 a11864a <=( (not A166)  and  a11863a );
 a11865a <=( a11864a  and  a11859a );
 a11869a <=( A267  and  A265 );
 a11870a <=( A203  and  a11869a );
 a11874a <=( (not A301)  and  (not A299) );
 a11875a <=( (not A298)  and  a11874a );
 a11876a <=( a11875a  and  a11870a );
 a11879a <=( A167  and  A170 );
 a11883a <=( (not A200)  and  A199 );
 a11884a <=( (not A166)  and  a11883a );
 a11885a <=( a11884a  and  a11879a );
 a11889a <=( A267  and  A266 );
 a11890a <=( A203  and  a11889a );
 a11894a <=( (not A302)  and  (not A301) );
 a11895a <=( (not A300)  and  a11894a );
 a11896a <=( a11895a  and  a11890a );
 a11899a <=( A167  and  A170 );
 a11903a <=( (not A200)  and  A199 );
 a11904a <=( (not A166)  and  a11903a );
 a11905a <=( a11904a  and  a11899a );
 a11909a <=( A267  and  A266 );
 a11910a <=( A203  and  a11909a );
 a11914a <=( (not A301)  and  (not A299) );
 a11915a <=( (not A298)  and  a11914a );
 a11916a <=( a11915a  and  a11910a );
 a11919a <=( A167  and  A170 );
 a11923a <=( (not A200)  and  (not A199) );
 a11924a <=( (not A166)  and  a11923a );
 a11925a <=( a11924a  and  a11919a );
 a11929a <=( (not A268)  and  (not A267) );
 a11930a <=( (not A202)  and  a11929a );
 a11934a <=( A300  and  A299 );
 a11935a <=( (not A269)  and  a11934a );
 a11936a <=( a11935a  and  a11930a );
 a11939a <=( A167  and  A170 );
 a11943a <=( (not A200)  and  (not A199) );
 a11944a <=( (not A166)  and  a11943a );
 a11945a <=( a11944a  and  a11939a );
 a11949a <=( (not A268)  and  (not A267) );
 a11950a <=( (not A202)  and  a11949a );
 a11954a <=( A300  and  A298 );
 a11955a <=( (not A269)  and  a11954a );
 a11956a <=( a11955a  and  a11950a );
 a11959a <=( A167  and  A170 );
 a11963a <=( (not A200)  and  (not A199) );
 a11964a <=( (not A166)  and  a11963a );
 a11965a <=( a11964a  and  a11959a );
 a11969a <=( A266  and  A265 );
 a11970a <=( (not A202)  and  a11969a );
 a11974a <=( A301  and  (not A268) );
 a11975a <=( (not A267)  and  a11974a );
 a11976a <=( a11975a  and  a11970a );
 a11979a <=( A167  and  A170 );
 a11983a <=( (not A200)  and  (not A199) );
 a11984a <=( (not A166)  and  a11983a );
 a11985a <=( a11984a  and  a11979a );
 a11989a <=( (not A266)  and  (not A265) );
 a11990a <=( (not A202)  and  a11989a );
 a11994a <=( A300  and  A299 );
 a11995a <=( (not A268)  and  a11994a );
 a11996a <=( a11995a  and  a11990a );
 a11999a <=( A167  and  A170 );
 a12003a <=( (not A200)  and  (not A199) );
 a12004a <=( (not A166)  and  a12003a );
 a12005a <=( a12004a  and  a11999a );
 a12009a <=( (not A266)  and  (not A265) );
 a12010a <=( (not A202)  and  a12009a );
 a12014a <=( A300  and  A298 );
 a12015a <=( (not A268)  and  a12014a );
 a12016a <=( a12015a  and  a12010a );
 a12019a <=( (not A167)  and  A170 );
 a12023a <=( (not A265)  and  A202 );
 a12024a <=( A166  and  a12023a );
 a12025a <=( a12024a  and  a12019a );
 a12029a <=( A298  and  A269 );
 a12030a <=( A266  and  a12029a );
 a12034a <=( (not A301)  and  (not A300) );
 a12035a <=( A299  and  a12034a );
 a12036a <=( a12035a  and  a12030a );
 a12039a <=( (not A167)  and  A170 );
 a12043a <=( A265  and  A202 );
 a12044a <=( A166  and  a12043a );
 a12045a <=( a12044a  and  a12039a );
 a12049a <=( A298  and  A269 );
 a12050a <=( (not A266)  and  a12049a );
 a12054a <=( (not A301)  and  (not A300) );
 a12055a <=( A299  and  a12054a );
 a12056a <=( a12055a  and  a12050a );
 a12059a <=( (not A167)  and  A170 );
 a12063a <=( (not A202)  and  (not A201) );
 a12064a <=( A166  and  a12063a );
 a12065a <=( a12064a  and  a12059a );
 a12069a <=( (not A268)  and  (not A267) );
 a12070a <=( (not A203)  and  a12069a );
 a12074a <=( A300  and  A299 );
 a12075a <=( (not A269)  and  a12074a );
 a12076a <=( a12075a  and  a12070a );
 a12079a <=( (not A167)  and  A170 );
 a12083a <=( (not A202)  and  (not A201) );
 a12084a <=( A166  and  a12083a );
 a12085a <=( a12084a  and  a12079a );
 a12089a <=( (not A268)  and  (not A267) );
 a12090a <=( (not A203)  and  a12089a );
 a12094a <=( A300  and  A298 );
 a12095a <=( (not A269)  and  a12094a );
 a12096a <=( a12095a  and  a12090a );
 a12099a <=( (not A167)  and  A170 );
 a12103a <=( (not A202)  and  (not A201) );
 a12104a <=( A166  and  a12103a );
 a12105a <=( a12104a  and  a12099a );
 a12109a <=( A266  and  A265 );
 a12110a <=( (not A203)  and  a12109a );
 a12114a <=( A301  and  (not A268) );
 a12115a <=( (not A267)  and  a12114a );
 a12116a <=( a12115a  and  a12110a );
 a12119a <=( (not A167)  and  A170 );
 a12123a <=( (not A202)  and  (not A201) );
 a12124a <=( A166  and  a12123a );
 a12125a <=( a12124a  and  a12119a );
 a12129a <=( (not A266)  and  (not A265) );
 a12130a <=( (not A203)  and  a12129a );
 a12134a <=( A300  and  A299 );
 a12135a <=( (not A268)  and  a12134a );
 a12136a <=( a12135a  and  a12130a );
 a12139a <=( (not A167)  and  A170 );
 a12143a <=( (not A202)  and  (not A201) );
 a12144a <=( A166  and  a12143a );
 a12145a <=( a12144a  and  a12139a );
 a12149a <=( (not A266)  and  (not A265) );
 a12150a <=( (not A203)  and  a12149a );
 a12154a <=( A300  and  A298 );
 a12155a <=( (not A268)  and  a12154a );
 a12156a <=( a12155a  and  a12150a );
 a12159a <=( (not A167)  and  A170 );
 a12163a <=( A201  and  A199 );
 a12164a <=( A166  and  a12163a );
 a12165a <=( a12164a  and  a12159a );
 a12169a <=( A298  and  A267 );
 a12170a <=( A265  and  a12169a );
 a12174a <=( (not A301)  and  (not A300) );
 a12175a <=( A299  and  a12174a );
 a12176a <=( a12175a  and  a12170a );
 a12179a <=( (not A167)  and  A170 );
 a12183a <=( A201  and  A199 );
 a12184a <=( A166  and  a12183a );
 a12185a <=( a12184a  and  a12179a );
 a12189a <=( A298  and  A267 );
 a12190a <=( A266  and  a12189a );
 a12194a <=( (not A301)  and  (not A300) );
 a12195a <=( A299  and  a12194a );
 a12196a <=( a12195a  and  a12190a );
 a12199a <=( (not A167)  and  A170 );
 a12203a <=( A201  and  A199 );
 a12204a <=( A166  and  a12203a );
 a12205a <=( a12204a  and  a12199a );
 a12209a <=( A269  and  A266 );
 a12210a <=( (not A265)  and  a12209a );
 a12214a <=( (not A302)  and  (not A301) );
 a12215a <=( (not A300)  and  a12214a );
 a12216a <=( a12215a  and  a12210a );
 a12219a <=( (not A167)  and  A170 );
 a12223a <=( A201  and  A199 );
 a12224a <=( A166  and  a12223a );
 a12225a <=( a12224a  and  a12219a );
 a12229a <=( A269  and  A266 );
 a12230a <=( (not A265)  and  a12229a );
 a12234a <=( (not A301)  and  (not A299) );
 a12235a <=( (not A298)  and  a12234a );
 a12236a <=( a12235a  and  a12230a );
 a12239a <=( (not A167)  and  A170 );
 a12243a <=( A201  and  A199 );
 a12244a <=( A166  and  a12243a );
 a12245a <=( a12244a  and  a12239a );
 a12249a <=( A269  and  (not A266) );
 a12250a <=( A265  and  a12249a );
 a12254a <=( (not A302)  and  (not A301) );
 a12255a <=( (not A300)  and  a12254a );
 a12256a <=( a12255a  and  a12250a );
 a12259a <=( (not A167)  and  A170 );
 a12263a <=( A201  and  A199 );
 a12264a <=( A166  and  a12263a );
 a12265a <=( a12264a  and  a12259a );
 a12269a <=( A269  and  (not A266) );
 a12270a <=( A265  and  a12269a );
 a12274a <=( (not A301)  and  (not A299) );
 a12275a <=( (not A298)  and  a12274a );
 a12276a <=( a12275a  and  a12270a );
 a12279a <=( (not A167)  and  A170 );
 a12283a <=( A201  and  A200 );
 a12284a <=( A166  and  a12283a );
 a12285a <=( a12284a  and  a12279a );
 a12289a <=( A298  and  A267 );
 a12290a <=( A265  and  a12289a );
 a12294a <=( (not A301)  and  (not A300) );
 a12295a <=( A299  and  a12294a );
 a12296a <=( a12295a  and  a12290a );
 a12299a <=( (not A167)  and  A170 );
 a12303a <=( A201  and  A200 );
 a12304a <=( A166  and  a12303a );
 a12305a <=( a12304a  and  a12299a );
 a12309a <=( A298  and  A267 );
 a12310a <=( A266  and  a12309a );
 a12314a <=( (not A301)  and  (not A300) );
 a12315a <=( A299  and  a12314a );
 a12316a <=( a12315a  and  a12310a );
 a12319a <=( (not A167)  and  A170 );
 a12323a <=( A201  and  A200 );
 a12324a <=( A166  and  a12323a );
 a12325a <=( a12324a  and  a12319a );
 a12329a <=( A269  and  A266 );
 a12330a <=( (not A265)  and  a12329a );
 a12334a <=( (not A302)  and  (not A301) );
 a12335a <=( (not A300)  and  a12334a );
 a12336a <=( a12335a  and  a12330a );
 a12339a <=( (not A167)  and  A170 );
 a12343a <=( A201  and  A200 );
 a12344a <=( A166  and  a12343a );
 a12345a <=( a12344a  and  a12339a );
 a12349a <=( A269  and  A266 );
 a12350a <=( (not A265)  and  a12349a );
 a12354a <=( (not A301)  and  (not A299) );
 a12355a <=( (not A298)  and  a12354a );
 a12356a <=( a12355a  and  a12350a );
 a12359a <=( (not A167)  and  A170 );
 a12363a <=( A201  and  A200 );
 a12364a <=( A166  and  a12363a );
 a12365a <=( a12364a  and  a12359a );
 a12369a <=( A269  and  (not A266) );
 a12370a <=( A265  and  a12369a );
 a12374a <=( (not A302)  and  (not A301) );
 a12375a <=( (not A300)  and  a12374a );
 a12376a <=( a12375a  and  a12370a );
 a12379a <=( (not A167)  and  A170 );
 a12383a <=( A201  and  A200 );
 a12384a <=( A166  and  a12383a );
 a12385a <=( a12384a  and  a12379a );
 a12389a <=( A269  and  (not A266) );
 a12390a <=( A265  and  a12389a );
 a12394a <=( (not A301)  and  (not A299) );
 a12395a <=( (not A298)  and  a12394a );
 a12396a <=( a12395a  and  a12390a );
 a12399a <=( (not A167)  and  A170 );
 a12403a <=( A200  and  A199 );
 a12404a <=( A166  and  a12403a );
 a12405a <=( a12404a  and  a12399a );
 a12409a <=( (not A267)  and  (not A202) );
 a12410a <=( (not A201)  and  a12409a );
 a12414a <=( A301  and  (not A269) );
 a12415a <=( (not A268)  and  a12414a );
 a12416a <=( a12415a  and  a12410a );
 a12419a <=( (not A167)  and  A170 );
 a12423a <=( A200  and  A199 );
 a12424a <=( A166  and  a12423a );
 a12425a <=( a12424a  and  a12419a );
 a12429a <=( (not A265)  and  (not A202) );
 a12430a <=( (not A201)  and  a12429a );
 a12434a <=( A301  and  (not A268) );
 a12435a <=( (not A266)  and  a12434a );
 a12436a <=( a12435a  and  a12430a );
 a12439a <=( (not A167)  and  A170 );
 a12443a <=( A200  and  (not A199) );
 a12444a <=( A166  and  a12443a );
 a12445a <=( a12444a  and  a12439a );
 a12449a <=( A298  and  A268 );
 a12450a <=( A203  and  a12449a );
 a12454a <=( (not A301)  and  (not A300) );
 a12455a <=( A299  and  a12454a );
 a12456a <=( a12455a  and  a12450a );
 a12459a <=( (not A167)  and  A170 );
 a12463a <=( A200  and  (not A199) );
 a12464a <=( A166  and  a12463a );
 a12465a <=( a12464a  and  a12459a );
 a12469a <=( A267  and  A265 );
 a12470a <=( A203  and  a12469a );
 a12474a <=( (not A302)  and  (not A301) );
 a12475a <=( (not A300)  and  a12474a );
 a12476a <=( a12475a  and  a12470a );
 a12479a <=( (not A167)  and  A170 );
 a12483a <=( A200  and  (not A199) );
 a12484a <=( A166  and  a12483a );
 a12485a <=( a12484a  and  a12479a );
 a12489a <=( A267  and  A265 );
 a12490a <=( A203  and  a12489a );
 a12494a <=( (not A301)  and  (not A299) );
 a12495a <=( (not A298)  and  a12494a );
 a12496a <=( a12495a  and  a12490a );
 a12499a <=( (not A167)  and  A170 );
 a12503a <=( A200  and  (not A199) );
 a12504a <=( A166  and  a12503a );
 a12505a <=( a12504a  and  a12499a );
 a12509a <=( A267  and  A266 );
 a12510a <=( A203  and  a12509a );
 a12514a <=( (not A302)  and  (not A301) );
 a12515a <=( (not A300)  and  a12514a );
 a12516a <=( a12515a  and  a12510a );
 a12519a <=( (not A167)  and  A170 );
 a12523a <=( A200  and  (not A199) );
 a12524a <=( A166  and  a12523a );
 a12525a <=( a12524a  and  a12519a );
 a12529a <=( A267  and  A266 );
 a12530a <=( A203  and  a12529a );
 a12534a <=( (not A301)  and  (not A299) );
 a12535a <=( (not A298)  and  a12534a );
 a12536a <=( a12535a  and  a12530a );
 a12539a <=( (not A167)  and  A170 );
 a12543a <=( (not A200)  and  A199 );
 a12544a <=( A166  and  a12543a );
 a12545a <=( a12544a  and  a12539a );
 a12549a <=( A298  and  A268 );
 a12550a <=( A203  and  a12549a );
 a12554a <=( (not A301)  and  (not A300) );
 a12555a <=( A299  and  a12554a );
 a12556a <=( a12555a  and  a12550a );
 a12559a <=( (not A167)  and  A170 );
 a12563a <=( (not A200)  and  A199 );
 a12564a <=( A166  and  a12563a );
 a12565a <=( a12564a  and  a12559a );
 a12569a <=( A267  and  A265 );
 a12570a <=( A203  and  a12569a );
 a12574a <=( (not A302)  and  (not A301) );
 a12575a <=( (not A300)  and  a12574a );
 a12576a <=( a12575a  and  a12570a );
 a12579a <=( (not A167)  and  A170 );
 a12583a <=( (not A200)  and  A199 );
 a12584a <=( A166  and  a12583a );
 a12585a <=( a12584a  and  a12579a );
 a12589a <=( A267  and  A265 );
 a12590a <=( A203  and  a12589a );
 a12594a <=( (not A301)  and  (not A299) );
 a12595a <=( (not A298)  and  a12594a );
 a12596a <=( a12595a  and  a12590a );
 a12599a <=( (not A167)  and  A170 );
 a12603a <=( (not A200)  and  A199 );
 a12604a <=( A166  and  a12603a );
 a12605a <=( a12604a  and  a12599a );
 a12609a <=( A267  and  A266 );
 a12610a <=( A203  and  a12609a );
 a12614a <=( (not A302)  and  (not A301) );
 a12615a <=( (not A300)  and  a12614a );
 a12616a <=( a12615a  and  a12610a );
 a12619a <=( (not A167)  and  A170 );
 a12623a <=( (not A200)  and  A199 );
 a12624a <=( A166  and  a12623a );
 a12625a <=( a12624a  and  a12619a );
 a12629a <=( A267  and  A266 );
 a12630a <=( A203  and  a12629a );
 a12634a <=( (not A301)  and  (not A299) );
 a12635a <=( (not A298)  and  a12634a );
 a12636a <=( a12635a  and  a12630a );
 a12639a <=( (not A167)  and  A170 );
 a12643a <=( (not A200)  and  (not A199) );
 a12644a <=( A166  and  a12643a );
 a12645a <=( a12644a  and  a12639a );
 a12649a <=( (not A268)  and  (not A267) );
 a12650a <=( (not A202)  and  a12649a );
 a12654a <=( A300  and  A299 );
 a12655a <=( (not A269)  and  a12654a );
 a12656a <=( a12655a  and  a12650a );
 a12659a <=( (not A167)  and  A170 );
 a12663a <=( (not A200)  and  (not A199) );
 a12664a <=( A166  and  a12663a );
 a12665a <=( a12664a  and  a12659a );
 a12669a <=( (not A268)  and  (not A267) );
 a12670a <=( (not A202)  and  a12669a );
 a12674a <=( A300  and  A298 );
 a12675a <=( (not A269)  and  a12674a );
 a12676a <=( a12675a  and  a12670a );
 a12679a <=( (not A167)  and  A170 );
 a12683a <=( (not A200)  and  (not A199) );
 a12684a <=( A166  and  a12683a );
 a12685a <=( a12684a  and  a12679a );
 a12689a <=( A266  and  A265 );
 a12690a <=( (not A202)  and  a12689a );
 a12694a <=( A301  and  (not A268) );
 a12695a <=( (not A267)  and  a12694a );
 a12696a <=( a12695a  and  a12690a );
 a12699a <=( (not A167)  and  A170 );
 a12703a <=( (not A200)  and  (not A199) );
 a12704a <=( A166  and  a12703a );
 a12705a <=( a12704a  and  a12699a );
 a12709a <=( (not A266)  and  (not A265) );
 a12710a <=( (not A202)  and  a12709a );
 a12714a <=( A300  and  A299 );
 a12715a <=( (not A268)  and  a12714a );
 a12716a <=( a12715a  and  a12710a );
 a12719a <=( (not A167)  and  A170 );
 a12723a <=( (not A200)  and  (not A199) );
 a12724a <=( A166  and  a12723a );
 a12725a <=( a12724a  and  a12719a );
 a12729a <=( (not A266)  and  (not A265) );
 a12730a <=( (not A202)  and  a12729a );
 a12734a <=( A300  and  A298 );
 a12735a <=( (not A268)  and  a12734a );
 a12736a <=( a12735a  and  a12730a );
 a12739a <=( (not A201)  and  A169 );
 a12743a <=( A265  and  (not A203) );
 a12744a <=( (not A202)  and  a12743a );
 a12745a <=( a12744a  and  a12739a );
 a12749a <=( (not A268)  and  (not A267) );
 a12750a <=( A266  and  a12749a );
 a12754a <=( A302  and  (not A299) );
 a12755a <=( A298  and  a12754a );
 a12756a <=( a12755a  and  a12750a );
 a12759a <=( (not A201)  and  A169 );
 a12763a <=( A265  and  (not A203) );
 a12764a <=( (not A202)  and  a12763a );
 a12765a <=( a12764a  and  a12759a );
 a12769a <=( (not A268)  and  (not A267) );
 a12770a <=( A266  and  a12769a );
 a12774a <=( A302  and  A299 );
 a12775a <=( (not A298)  and  a12774a );
 a12776a <=( a12775a  and  a12770a );
 a12779a <=( A199  and  A169 );
 a12783a <=( (not A202)  and  (not A201) );
 a12784a <=( A200  and  a12783a );
 a12785a <=( a12784a  and  a12779a );
 a12789a <=( (not A269)  and  (not A268) );
 a12790a <=( (not A267)  and  a12789a );
 a12794a <=( A302  and  (not A299) );
 a12795a <=( A298  and  a12794a );
 a12796a <=( a12795a  and  a12790a );
 a12799a <=( A199  and  A169 );
 a12803a <=( (not A202)  and  (not A201) );
 a12804a <=( A200  and  a12803a );
 a12805a <=( a12804a  and  a12799a );
 a12809a <=( (not A269)  and  (not A268) );
 a12810a <=( (not A267)  and  a12809a );
 a12814a <=( A302  and  A299 );
 a12815a <=( (not A298)  and  a12814a );
 a12816a <=( a12815a  and  a12810a );
 a12819a <=( A199  and  A169 );
 a12823a <=( (not A202)  and  (not A201) );
 a12824a <=( A200  and  a12823a );
 a12825a <=( a12824a  and  a12819a );
 a12829a <=( (not A267)  and  A266 );
 a12830a <=( A265  and  a12829a );
 a12834a <=( A300  and  A299 );
 a12835a <=( (not A268)  and  a12834a );
 a12836a <=( a12835a  and  a12830a );
 a12839a <=( A199  and  A169 );
 a12843a <=( (not A202)  and  (not A201) );
 a12844a <=( A200  and  a12843a );
 a12845a <=( a12844a  and  a12839a );
 a12849a <=( (not A267)  and  A266 );
 a12850a <=( A265  and  a12849a );
 a12854a <=( A300  and  A298 );
 a12855a <=( (not A268)  and  a12854a );
 a12856a <=( a12855a  and  a12850a );
 a12859a <=( A199  and  A169 );
 a12863a <=( (not A202)  and  (not A201) );
 a12864a <=( A200  and  a12863a );
 a12865a <=( a12864a  and  a12859a );
 a12869a <=( (not A268)  and  (not A266) );
 a12870a <=( (not A265)  and  a12869a );
 a12874a <=( A302  and  (not A299) );
 a12875a <=( A298  and  a12874a );
 a12876a <=( a12875a  and  a12870a );
 a12879a <=( A199  and  A169 );
 a12883a <=( (not A202)  and  (not A201) );
 a12884a <=( A200  and  a12883a );
 a12885a <=( a12884a  and  a12879a );
 a12889a <=( (not A268)  and  (not A266) );
 a12890a <=( (not A265)  and  a12889a );
 a12894a <=( A302  and  A299 );
 a12895a <=( (not A298)  and  a12894a );
 a12896a <=( a12895a  and  a12890a );
 a12899a <=( (not A199)  and  A169 );
 a12903a <=( (not A265)  and  A203 );
 a12904a <=( A200  and  a12903a );
 a12905a <=( a12904a  and  a12899a );
 a12909a <=( A298  and  A269 );
 a12910a <=( A266  and  a12909a );
 a12914a <=( (not A301)  and  (not A300) );
 a12915a <=( A299  and  a12914a );
 a12916a <=( a12915a  and  a12910a );
 a12919a <=( (not A199)  and  A169 );
 a12923a <=( A265  and  A203 );
 a12924a <=( A200  and  a12923a );
 a12925a <=( a12924a  and  a12919a );
 a12929a <=( A298  and  A269 );
 a12930a <=( (not A266)  and  a12929a );
 a12934a <=( (not A301)  and  (not A300) );
 a12935a <=( A299  and  a12934a );
 a12936a <=( a12935a  and  a12930a );
 a12939a <=( A199  and  A169 );
 a12943a <=( (not A265)  and  A203 );
 a12944a <=( (not A200)  and  a12943a );
 a12945a <=( a12944a  and  a12939a );
 a12949a <=( A298  and  A269 );
 a12950a <=( A266  and  a12949a );
 a12954a <=( (not A301)  and  (not A300) );
 a12955a <=( A299  and  a12954a );
 a12956a <=( a12955a  and  a12950a );
 a12959a <=( A199  and  A169 );
 a12963a <=( A265  and  A203 );
 a12964a <=( (not A200)  and  a12963a );
 a12965a <=( a12964a  and  a12959a );
 a12969a <=( A298  and  A269 );
 a12970a <=( (not A266)  and  a12969a );
 a12974a <=( (not A301)  and  (not A300) );
 a12975a <=( A299  and  a12974a );
 a12976a <=( a12975a  and  a12970a );
 a12979a <=( (not A199)  and  A169 );
 a12983a <=( A265  and  (not A202) );
 a12984a <=( (not A200)  and  a12983a );
 a12985a <=( a12984a  and  a12979a );
 a12989a <=( (not A268)  and  (not A267) );
 a12990a <=( A266  and  a12989a );
 a12994a <=( A302  and  (not A299) );
 a12995a <=( A298  and  a12994a );
 a12996a <=( a12995a  and  a12990a );
 a12999a <=( (not A199)  and  A169 );
 a13003a <=( A265  and  (not A202) );
 a13004a <=( (not A200)  and  a13003a );
 a13005a <=( a13004a  and  a12999a );
 a13009a <=( (not A268)  and  (not A267) );
 a13010a <=( A266  and  a13009a );
 a13014a <=( A302  and  A299 );
 a13015a <=( (not A298)  and  a13014a );
 a13016a <=( a13015a  and  a13010a );
 a13019a <=( (not A167)  and  (not A169) );
 a13023a <=( A265  and  A202 );
 a13024a <=( (not A166)  and  a13023a );
 a13025a <=( a13024a  and  a13019a );
 a13029a <=( (not A268)  and  (not A267) );
 a13030a <=( A266  and  a13029a );
 a13034a <=( A302  and  (not A299) );
 a13035a <=( A298  and  a13034a );
 a13036a <=( a13035a  and  a13030a );
 a13039a <=( (not A167)  and  (not A169) );
 a13043a <=( A265  and  A202 );
 a13044a <=( (not A166)  and  a13043a );
 a13045a <=( a13044a  and  a13039a );
 a13049a <=( (not A268)  and  (not A267) );
 a13050a <=( A266  and  a13049a );
 a13054a <=( A302  and  A299 );
 a13055a <=( (not A298)  and  a13054a );
 a13056a <=( a13055a  and  a13050a );
 a13059a <=( (not A167)  and  (not A169) );
 a13063a <=( (not A202)  and  (not A201) );
 a13064a <=( (not A166)  and  a13063a );
 a13065a <=( a13064a  and  a13059a );
 a13069a <=( A298  and  A268 );
 a13070a <=( (not A203)  and  a13069a );
 a13074a <=( (not A301)  and  (not A300) );
 a13075a <=( A299  and  a13074a );
 a13076a <=( a13075a  and  a13070a );
 a13079a <=( (not A167)  and  (not A169) );
 a13083a <=( (not A202)  and  (not A201) );
 a13084a <=( (not A166)  and  a13083a );
 a13085a <=( a13084a  and  a13079a );
 a13089a <=( A267  and  A265 );
 a13090a <=( (not A203)  and  a13089a );
 a13094a <=( (not A302)  and  (not A301) );
 a13095a <=( (not A300)  and  a13094a );
 a13096a <=( a13095a  and  a13090a );
 a13099a <=( (not A167)  and  (not A169) );
 a13103a <=( (not A202)  and  (not A201) );
 a13104a <=( (not A166)  and  a13103a );
 a13105a <=( a13104a  and  a13099a );
 a13109a <=( A267  and  A265 );
 a13110a <=( (not A203)  and  a13109a );
 a13114a <=( (not A301)  and  (not A299) );
 a13115a <=( (not A298)  and  a13114a );
 a13116a <=( a13115a  and  a13110a );
 a13119a <=( (not A167)  and  (not A169) );
 a13123a <=( (not A202)  and  (not A201) );
 a13124a <=( (not A166)  and  a13123a );
 a13125a <=( a13124a  and  a13119a );
 a13129a <=( A267  and  A266 );
 a13130a <=( (not A203)  and  a13129a );
 a13134a <=( (not A302)  and  (not A301) );
 a13135a <=( (not A300)  and  a13134a );
 a13136a <=( a13135a  and  a13130a );
 a13139a <=( (not A167)  and  (not A169) );
 a13143a <=( (not A202)  and  (not A201) );
 a13144a <=( (not A166)  and  a13143a );
 a13145a <=( a13144a  and  a13139a );
 a13149a <=( A267  and  A266 );
 a13150a <=( (not A203)  and  a13149a );
 a13154a <=( (not A301)  and  (not A299) );
 a13155a <=( (not A298)  and  a13154a );
 a13156a <=( a13155a  and  a13150a );
 a13159a <=( (not A167)  and  (not A169) );
 a13163a <=( A201  and  A199 );
 a13164a <=( (not A166)  and  a13163a );
 a13165a <=( a13164a  and  a13159a );
 a13169a <=( (not A269)  and  (not A268) );
 a13170a <=( (not A267)  and  a13169a );
 a13174a <=( A302  and  (not A299) );
 a13175a <=( A298  and  a13174a );
 a13176a <=( a13175a  and  a13170a );
 a13179a <=( (not A167)  and  (not A169) );
 a13183a <=( A201  and  A199 );
 a13184a <=( (not A166)  and  a13183a );
 a13185a <=( a13184a  and  a13179a );
 a13189a <=( (not A269)  and  (not A268) );
 a13190a <=( (not A267)  and  a13189a );
 a13194a <=( A302  and  A299 );
 a13195a <=( (not A298)  and  a13194a );
 a13196a <=( a13195a  and  a13190a );
 a13199a <=( (not A167)  and  (not A169) );
 a13203a <=( A201  and  A199 );
 a13204a <=( (not A166)  and  a13203a );
 a13205a <=( a13204a  and  a13199a );
 a13209a <=( (not A267)  and  A266 );
 a13210a <=( A265  and  a13209a );
 a13214a <=( A300  and  A299 );
 a13215a <=( (not A268)  and  a13214a );
 a13216a <=( a13215a  and  a13210a );
 a13219a <=( (not A167)  and  (not A169) );
 a13223a <=( A201  and  A199 );
 a13224a <=( (not A166)  and  a13223a );
 a13225a <=( a13224a  and  a13219a );
 a13229a <=( (not A267)  and  A266 );
 a13230a <=( A265  and  a13229a );
 a13234a <=( A300  and  A298 );
 a13235a <=( (not A268)  and  a13234a );
 a13236a <=( a13235a  and  a13230a );
 a13239a <=( (not A167)  and  (not A169) );
 a13243a <=( A201  and  A199 );
 a13244a <=( (not A166)  and  a13243a );
 a13245a <=( a13244a  and  a13239a );
 a13249a <=( (not A268)  and  (not A266) );
 a13250a <=( (not A265)  and  a13249a );
 a13254a <=( A302  and  (not A299) );
 a13255a <=( A298  and  a13254a );
 a13256a <=( a13255a  and  a13250a );
 a13259a <=( (not A167)  and  (not A169) );
 a13263a <=( A201  and  A199 );
 a13264a <=( (not A166)  and  a13263a );
 a13265a <=( a13264a  and  a13259a );
 a13269a <=( (not A268)  and  (not A266) );
 a13270a <=( (not A265)  and  a13269a );
 a13274a <=( A302  and  A299 );
 a13275a <=( (not A298)  and  a13274a );
 a13276a <=( a13275a  and  a13270a );
 a13279a <=( (not A167)  and  (not A169) );
 a13283a <=( A201  and  A200 );
 a13284a <=( (not A166)  and  a13283a );
 a13285a <=( a13284a  and  a13279a );
 a13289a <=( (not A269)  and  (not A268) );
 a13290a <=( (not A267)  and  a13289a );
 a13294a <=( A302  and  (not A299) );
 a13295a <=( A298  and  a13294a );
 a13296a <=( a13295a  and  a13290a );
 a13299a <=( (not A167)  and  (not A169) );
 a13303a <=( A201  and  A200 );
 a13304a <=( (not A166)  and  a13303a );
 a13305a <=( a13304a  and  a13299a );
 a13309a <=( (not A269)  and  (not A268) );
 a13310a <=( (not A267)  and  a13309a );
 a13314a <=( A302  and  A299 );
 a13315a <=( (not A298)  and  a13314a );
 a13316a <=( a13315a  and  a13310a );
 a13319a <=( (not A167)  and  (not A169) );
 a13323a <=( A201  and  A200 );
 a13324a <=( (not A166)  and  a13323a );
 a13325a <=( a13324a  and  a13319a );
 a13329a <=( (not A267)  and  A266 );
 a13330a <=( A265  and  a13329a );
 a13334a <=( A300  and  A299 );
 a13335a <=( (not A268)  and  a13334a );
 a13336a <=( a13335a  and  a13330a );
 a13339a <=( (not A167)  and  (not A169) );
 a13343a <=( A201  and  A200 );
 a13344a <=( (not A166)  and  a13343a );
 a13345a <=( a13344a  and  a13339a );
 a13349a <=( (not A267)  and  A266 );
 a13350a <=( A265  and  a13349a );
 a13354a <=( A300  and  A298 );
 a13355a <=( (not A268)  and  a13354a );
 a13356a <=( a13355a  and  a13350a );
 a13359a <=( (not A167)  and  (not A169) );
 a13363a <=( A201  and  A200 );
 a13364a <=( (not A166)  and  a13363a );
 a13365a <=( a13364a  and  a13359a );
 a13369a <=( (not A268)  and  (not A266) );
 a13370a <=( (not A265)  and  a13369a );
 a13374a <=( A302  and  (not A299) );
 a13375a <=( A298  and  a13374a );
 a13376a <=( a13375a  and  a13370a );
 a13379a <=( (not A167)  and  (not A169) );
 a13383a <=( A201  and  A200 );
 a13384a <=( (not A166)  and  a13383a );
 a13385a <=( a13384a  and  a13379a );
 a13389a <=( (not A268)  and  (not A266) );
 a13390a <=( (not A265)  and  a13389a );
 a13394a <=( A302  and  A299 );
 a13395a <=( (not A298)  and  a13394a );
 a13396a <=( a13395a  and  a13390a );
 a13399a <=( (not A167)  and  (not A169) );
 a13403a <=( A200  and  A199 );
 a13404a <=( (not A166)  and  a13403a );
 a13405a <=( a13404a  and  a13399a );
 a13409a <=( A268  and  (not A202) );
 a13410a <=( (not A201)  and  a13409a );
 a13414a <=( (not A302)  and  (not A301) );
 a13415a <=( (not A300)  and  a13414a );
 a13416a <=( a13415a  and  a13410a );
 a13419a <=( (not A167)  and  (not A169) );
 a13423a <=( A200  and  A199 );
 a13424a <=( (not A166)  and  a13423a );
 a13425a <=( a13424a  and  a13419a );
 a13429a <=( A268  and  (not A202) );
 a13430a <=( (not A201)  and  a13429a );
 a13434a <=( (not A301)  and  (not A299) );
 a13435a <=( (not A298)  and  a13434a );
 a13436a <=( a13435a  and  a13430a );
 a13439a <=( (not A167)  and  (not A169) );
 a13443a <=( A200  and  (not A199) );
 a13444a <=( (not A166)  and  a13443a );
 a13445a <=( a13444a  and  a13439a );
 a13449a <=( (not A268)  and  (not A267) );
 a13450a <=( A203  and  a13449a );
 a13454a <=( A300  and  A299 );
 a13455a <=( (not A269)  and  a13454a );
 a13456a <=( a13455a  and  a13450a );
 a13459a <=( (not A167)  and  (not A169) );
 a13463a <=( A200  and  (not A199) );
 a13464a <=( (not A166)  and  a13463a );
 a13465a <=( a13464a  and  a13459a );
 a13469a <=( (not A268)  and  (not A267) );
 a13470a <=( A203  and  a13469a );
 a13474a <=( A300  and  A298 );
 a13475a <=( (not A269)  and  a13474a );
 a13476a <=( a13475a  and  a13470a );
 a13479a <=( (not A167)  and  (not A169) );
 a13483a <=( A200  and  (not A199) );
 a13484a <=( (not A166)  and  a13483a );
 a13485a <=( a13484a  and  a13479a );
 a13489a <=( A266  and  A265 );
 a13490a <=( A203  and  a13489a );
 a13494a <=( A301  and  (not A268) );
 a13495a <=( (not A267)  and  a13494a );
 a13496a <=( a13495a  and  a13490a );
 a13499a <=( (not A167)  and  (not A169) );
 a13503a <=( A200  and  (not A199) );
 a13504a <=( (not A166)  and  a13503a );
 a13505a <=( a13504a  and  a13499a );
 a13509a <=( (not A266)  and  (not A265) );
 a13510a <=( A203  and  a13509a );
 a13514a <=( A300  and  A299 );
 a13515a <=( (not A268)  and  a13514a );
 a13516a <=( a13515a  and  a13510a );
 a13519a <=( (not A167)  and  (not A169) );
 a13523a <=( A200  and  (not A199) );
 a13524a <=( (not A166)  and  a13523a );
 a13525a <=( a13524a  and  a13519a );
 a13529a <=( (not A266)  and  (not A265) );
 a13530a <=( A203  and  a13529a );
 a13534a <=( A300  and  A298 );
 a13535a <=( (not A268)  and  a13534a );
 a13536a <=( a13535a  and  a13530a );
 a13539a <=( (not A167)  and  (not A169) );
 a13543a <=( (not A200)  and  A199 );
 a13544a <=( (not A166)  and  a13543a );
 a13545a <=( a13544a  and  a13539a );
 a13549a <=( (not A268)  and  (not A267) );
 a13550a <=( A203  and  a13549a );
 a13554a <=( A300  and  A299 );
 a13555a <=( (not A269)  and  a13554a );
 a13556a <=( a13555a  and  a13550a );
 a13559a <=( (not A167)  and  (not A169) );
 a13563a <=( (not A200)  and  A199 );
 a13564a <=( (not A166)  and  a13563a );
 a13565a <=( a13564a  and  a13559a );
 a13569a <=( (not A268)  and  (not A267) );
 a13570a <=( A203  and  a13569a );
 a13574a <=( A300  and  A298 );
 a13575a <=( (not A269)  and  a13574a );
 a13576a <=( a13575a  and  a13570a );
 a13579a <=( (not A167)  and  (not A169) );
 a13583a <=( (not A200)  and  A199 );
 a13584a <=( (not A166)  and  a13583a );
 a13585a <=( a13584a  and  a13579a );
 a13589a <=( A266  and  A265 );
 a13590a <=( A203  and  a13589a );
 a13594a <=( A301  and  (not A268) );
 a13595a <=( (not A267)  and  a13594a );
 a13596a <=( a13595a  and  a13590a );
 a13599a <=( (not A167)  and  (not A169) );
 a13603a <=( (not A200)  and  A199 );
 a13604a <=( (not A166)  and  a13603a );
 a13605a <=( a13604a  and  a13599a );
 a13609a <=( (not A266)  and  (not A265) );
 a13610a <=( A203  and  a13609a );
 a13614a <=( A300  and  A299 );
 a13615a <=( (not A268)  and  a13614a );
 a13616a <=( a13615a  and  a13610a );
 a13619a <=( (not A167)  and  (not A169) );
 a13623a <=( (not A200)  and  A199 );
 a13624a <=( (not A166)  and  a13623a );
 a13625a <=( a13624a  and  a13619a );
 a13629a <=( (not A266)  and  (not A265) );
 a13630a <=( A203  and  a13629a );
 a13634a <=( A300  and  A298 );
 a13635a <=( (not A268)  and  a13634a );
 a13636a <=( a13635a  and  a13630a );
 a13639a <=( (not A167)  and  (not A169) );
 a13643a <=( (not A200)  and  (not A199) );
 a13644a <=( (not A166)  and  a13643a );
 a13645a <=( a13644a  and  a13639a );
 a13649a <=( A298  and  A268 );
 a13650a <=( (not A202)  and  a13649a );
 a13654a <=( (not A301)  and  (not A300) );
 a13655a <=( A299  and  a13654a );
 a13656a <=( a13655a  and  a13650a );
 a13659a <=( (not A167)  and  (not A169) );
 a13663a <=( (not A200)  and  (not A199) );
 a13664a <=( (not A166)  and  a13663a );
 a13665a <=( a13664a  and  a13659a );
 a13669a <=( A267  and  A265 );
 a13670a <=( (not A202)  and  a13669a );
 a13674a <=( (not A302)  and  (not A301) );
 a13675a <=( (not A300)  and  a13674a );
 a13676a <=( a13675a  and  a13670a );
 a13679a <=( (not A167)  and  (not A169) );
 a13683a <=( (not A200)  and  (not A199) );
 a13684a <=( (not A166)  and  a13683a );
 a13685a <=( a13684a  and  a13679a );
 a13689a <=( A267  and  A265 );
 a13690a <=( (not A202)  and  a13689a );
 a13694a <=( (not A301)  and  (not A299) );
 a13695a <=( (not A298)  and  a13694a );
 a13696a <=( a13695a  and  a13690a );
 a13699a <=( (not A167)  and  (not A169) );
 a13703a <=( (not A200)  and  (not A199) );
 a13704a <=( (not A166)  and  a13703a );
 a13705a <=( a13704a  and  a13699a );
 a13709a <=( A267  and  A266 );
 a13710a <=( (not A202)  and  a13709a );
 a13714a <=( (not A302)  and  (not A301) );
 a13715a <=( (not A300)  and  a13714a );
 a13716a <=( a13715a  and  a13710a );
 a13719a <=( (not A167)  and  (not A169) );
 a13723a <=( (not A200)  and  (not A199) );
 a13724a <=( (not A166)  and  a13723a );
 a13725a <=( a13724a  and  a13719a );
 a13729a <=( A267  and  A266 );
 a13730a <=( (not A202)  and  a13729a );
 a13734a <=( (not A301)  and  (not A299) );
 a13735a <=( (not A298)  and  a13734a );
 a13736a <=( a13735a  and  a13730a );
 a13739a <=( (not A168)  and  (not A169) );
 a13743a <=( A202  and  A166 );
 a13744a <=( A167  and  a13743a );
 a13745a <=( a13744a  and  a13739a );
 a13749a <=( (not A269)  and  (not A268) );
 a13750a <=( (not A267)  and  a13749a );
 a13754a <=( A302  and  (not A299) );
 a13755a <=( A298  and  a13754a );
 a13756a <=( a13755a  and  a13750a );
 a13759a <=( (not A168)  and  (not A169) );
 a13763a <=( A202  and  A166 );
 a13764a <=( A167  and  a13763a );
 a13765a <=( a13764a  and  a13759a );
 a13769a <=( (not A269)  and  (not A268) );
 a13770a <=( (not A267)  and  a13769a );
 a13774a <=( A302  and  A299 );
 a13775a <=( (not A298)  and  a13774a );
 a13776a <=( a13775a  and  a13770a );
 a13779a <=( (not A168)  and  (not A169) );
 a13783a <=( A202  and  A166 );
 a13784a <=( A167  and  a13783a );
 a13785a <=( a13784a  and  a13779a );
 a13789a <=( (not A267)  and  A266 );
 a13790a <=( A265  and  a13789a );
 a13794a <=( A300  and  A299 );
 a13795a <=( (not A268)  and  a13794a );
 a13796a <=( a13795a  and  a13790a );
 a13799a <=( (not A168)  and  (not A169) );
 a13803a <=( A202  and  A166 );
 a13804a <=( A167  and  a13803a );
 a13805a <=( a13804a  and  a13799a );
 a13809a <=( (not A267)  and  A266 );
 a13810a <=( A265  and  a13809a );
 a13814a <=( A300  and  A298 );
 a13815a <=( (not A268)  and  a13814a );
 a13816a <=( a13815a  and  a13810a );
 a13819a <=( (not A168)  and  (not A169) );
 a13823a <=( A202  and  A166 );
 a13824a <=( A167  and  a13823a );
 a13825a <=( a13824a  and  a13819a );
 a13829a <=( (not A268)  and  (not A266) );
 a13830a <=( (not A265)  and  a13829a );
 a13834a <=( A302  and  (not A299) );
 a13835a <=( A298  and  a13834a );
 a13836a <=( a13835a  and  a13830a );
 a13839a <=( (not A168)  and  (not A169) );
 a13843a <=( A202  and  A166 );
 a13844a <=( A167  and  a13843a );
 a13845a <=( a13844a  and  a13839a );
 a13849a <=( (not A268)  and  (not A266) );
 a13850a <=( (not A265)  and  a13849a );
 a13854a <=( A302  and  A299 );
 a13855a <=( (not A298)  and  a13854a );
 a13856a <=( a13855a  and  a13850a );
 a13859a <=( (not A168)  and  (not A169) );
 a13863a <=( (not A201)  and  A166 );
 a13864a <=( A167  and  a13863a );
 a13865a <=( a13864a  and  a13859a );
 a13869a <=( A268  and  (not A203) );
 a13870a <=( (not A202)  and  a13869a );
 a13874a <=( (not A302)  and  (not A301) );
 a13875a <=( (not A300)  and  a13874a );
 a13876a <=( a13875a  and  a13870a );
 a13879a <=( (not A168)  and  (not A169) );
 a13883a <=( (not A201)  and  A166 );
 a13884a <=( A167  and  a13883a );
 a13885a <=( a13884a  and  a13879a );
 a13889a <=( A268  and  (not A203) );
 a13890a <=( (not A202)  and  a13889a );
 a13894a <=( (not A301)  and  (not A299) );
 a13895a <=( (not A298)  and  a13894a );
 a13896a <=( a13895a  and  a13890a );
 a13899a <=( (not A168)  and  (not A169) );
 a13903a <=( A199  and  A166 );
 a13904a <=( A167  and  a13903a );
 a13905a <=( a13904a  and  a13899a );
 a13909a <=( (not A268)  and  (not A267) );
 a13910a <=( A201  and  a13909a );
 a13914a <=( A300  and  A299 );
 a13915a <=( (not A269)  and  a13914a );
 a13916a <=( a13915a  and  a13910a );
 a13919a <=( (not A168)  and  (not A169) );
 a13923a <=( A199  and  A166 );
 a13924a <=( A167  and  a13923a );
 a13925a <=( a13924a  and  a13919a );
 a13929a <=( (not A268)  and  (not A267) );
 a13930a <=( A201  and  a13929a );
 a13934a <=( A300  and  A298 );
 a13935a <=( (not A269)  and  a13934a );
 a13936a <=( a13935a  and  a13930a );
 a13939a <=( (not A168)  and  (not A169) );
 a13943a <=( A199  and  A166 );
 a13944a <=( A167  and  a13943a );
 a13945a <=( a13944a  and  a13939a );
 a13949a <=( A266  and  A265 );
 a13950a <=( A201  and  a13949a );
 a13954a <=( A301  and  (not A268) );
 a13955a <=( (not A267)  and  a13954a );
 a13956a <=( a13955a  and  a13950a );
 a13959a <=( (not A168)  and  (not A169) );
 a13963a <=( A199  and  A166 );
 a13964a <=( A167  and  a13963a );
 a13965a <=( a13964a  and  a13959a );
 a13969a <=( (not A266)  and  (not A265) );
 a13970a <=( A201  and  a13969a );
 a13974a <=( A300  and  A299 );
 a13975a <=( (not A268)  and  a13974a );
 a13976a <=( a13975a  and  a13970a );
 a13979a <=( (not A168)  and  (not A169) );
 a13983a <=( A199  and  A166 );
 a13984a <=( A167  and  a13983a );
 a13985a <=( a13984a  and  a13979a );
 a13989a <=( (not A266)  and  (not A265) );
 a13990a <=( A201  and  a13989a );
 a13994a <=( A300  and  A298 );
 a13995a <=( (not A268)  and  a13994a );
 a13996a <=( a13995a  and  a13990a );
 a13999a <=( (not A168)  and  (not A169) );
 a14003a <=( A200  and  A166 );
 a14004a <=( A167  and  a14003a );
 a14005a <=( a14004a  and  a13999a );
 a14009a <=( (not A268)  and  (not A267) );
 a14010a <=( A201  and  a14009a );
 a14014a <=( A300  and  A299 );
 a14015a <=( (not A269)  and  a14014a );
 a14016a <=( a14015a  and  a14010a );
 a14019a <=( (not A168)  and  (not A169) );
 a14023a <=( A200  and  A166 );
 a14024a <=( A167  and  a14023a );
 a14025a <=( a14024a  and  a14019a );
 a14029a <=( (not A268)  and  (not A267) );
 a14030a <=( A201  and  a14029a );
 a14034a <=( A300  and  A298 );
 a14035a <=( (not A269)  and  a14034a );
 a14036a <=( a14035a  and  a14030a );
 a14039a <=( (not A168)  and  (not A169) );
 a14043a <=( A200  and  A166 );
 a14044a <=( A167  and  a14043a );
 a14045a <=( a14044a  and  a14039a );
 a14049a <=( A266  and  A265 );
 a14050a <=( A201  and  a14049a );
 a14054a <=( A301  and  (not A268) );
 a14055a <=( (not A267)  and  a14054a );
 a14056a <=( a14055a  and  a14050a );
 a14059a <=( (not A168)  and  (not A169) );
 a14063a <=( A200  and  A166 );
 a14064a <=( A167  and  a14063a );
 a14065a <=( a14064a  and  a14059a );
 a14069a <=( (not A266)  and  (not A265) );
 a14070a <=( A201  and  a14069a );
 a14074a <=( A300  and  A299 );
 a14075a <=( (not A268)  and  a14074a );
 a14076a <=( a14075a  and  a14070a );
 a14079a <=( (not A168)  and  (not A169) );
 a14083a <=( A200  and  A166 );
 a14084a <=( A167  and  a14083a );
 a14085a <=( a14084a  and  a14079a );
 a14089a <=( (not A266)  and  (not A265) );
 a14090a <=( A201  and  a14089a );
 a14094a <=( A300  and  A298 );
 a14095a <=( (not A268)  and  a14094a );
 a14096a <=( a14095a  and  a14090a );
 a14099a <=( (not A168)  and  (not A169) );
 a14103a <=( (not A199)  and  A166 );
 a14104a <=( A167  and  a14103a );
 a14105a <=( a14104a  and  a14099a );
 a14109a <=( (not A267)  and  A203 );
 a14110a <=( A200  and  a14109a );
 a14114a <=( A301  and  (not A269) );
 a14115a <=( (not A268)  and  a14114a );
 a14116a <=( a14115a  and  a14110a );
 a14119a <=( (not A168)  and  (not A169) );
 a14123a <=( (not A199)  and  A166 );
 a14124a <=( A167  and  a14123a );
 a14125a <=( a14124a  and  a14119a );
 a14129a <=( (not A265)  and  A203 );
 a14130a <=( A200  and  a14129a );
 a14134a <=( A301  and  (not A268) );
 a14135a <=( (not A266)  and  a14134a );
 a14136a <=( a14135a  and  a14130a );
 a14139a <=( (not A168)  and  (not A169) );
 a14143a <=( A199  and  A166 );
 a14144a <=( A167  and  a14143a );
 a14145a <=( a14144a  and  a14139a );
 a14149a <=( (not A267)  and  A203 );
 a14150a <=( (not A200)  and  a14149a );
 a14154a <=( A301  and  (not A269) );
 a14155a <=( (not A268)  and  a14154a );
 a14156a <=( a14155a  and  a14150a );
 a14159a <=( (not A168)  and  (not A169) );
 a14163a <=( A199  and  A166 );
 a14164a <=( A167  and  a14163a );
 a14165a <=( a14164a  and  a14159a );
 a14169a <=( (not A265)  and  A203 );
 a14170a <=( (not A200)  and  a14169a );
 a14174a <=( A301  and  (not A268) );
 a14175a <=( (not A266)  and  a14174a );
 a14176a <=( a14175a  and  a14170a );
 a14179a <=( (not A168)  and  (not A169) );
 a14183a <=( (not A199)  and  A166 );
 a14184a <=( A167  and  a14183a );
 a14185a <=( a14184a  and  a14179a );
 a14189a <=( A268  and  (not A202) );
 a14190a <=( (not A200)  and  a14189a );
 a14194a <=( (not A302)  and  (not A301) );
 a14195a <=( (not A300)  and  a14194a );
 a14196a <=( a14195a  and  a14190a );
 a14199a <=( (not A168)  and  (not A169) );
 a14203a <=( (not A199)  and  A166 );
 a14204a <=( A167  and  a14203a );
 a14205a <=( a14204a  and  a14199a );
 a14209a <=( A268  and  (not A202) );
 a14210a <=( (not A200)  and  a14209a );
 a14214a <=( (not A301)  and  (not A299) );
 a14215a <=( (not A298)  and  a14214a );
 a14216a <=( a14215a  and  a14210a );
 a14219a <=( (not A169)  and  (not A170) );
 a14223a <=( A265  and  A202 );
 a14224a <=( (not A168)  and  a14223a );
 a14225a <=( a14224a  and  a14219a );
 a14229a <=( (not A268)  and  (not A267) );
 a14230a <=( A266  and  a14229a );
 a14234a <=( A302  and  (not A299) );
 a14235a <=( A298  and  a14234a );
 a14236a <=( a14235a  and  a14230a );
 a14239a <=( (not A169)  and  (not A170) );
 a14243a <=( A265  and  A202 );
 a14244a <=( (not A168)  and  a14243a );
 a14245a <=( a14244a  and  a14239a );
 a14249a <=( (not A268)  and  (not A267) );
 a14250a <=( A266  and  a14249a );
 a14254a <=( A302  and  A299 );
 a14255a <=( (not A298)  and  a14254a );
 a14256a <=( a14255a  and  a14250a );
 a14259a <=( (not A169)  and  (not A170) );
 a14263a <=( (not A202)  and  (not A201) );
 a14264a <=( (not A168)  and  a14263a );
 a14265a <=( a14264a  and  a14259a );
 a14269a <=( A298  and  A268 );
 a14270a <=( (not A203)  and  a14269a );
 a14274a <=( (not A301)  and  (not A300) );
 a14275a <=( A299  and  a14274a );
 a14276a <=( a14275a  and  a14270a );
 a14279a <=( (not A169)  and  (not A170) );
 a14283a <=( (not A202)  and  (not A201) );
 a14284a <=( (not A168)  and  a14283a );
 a14285a <=( a14284a  and  a14279a );
 a14289a <=( A267  and  A265 );
 a14290a <=( (not A203)  and  a14289a );
 a14294a <=( (not A302)  and  (not A301) );
 a14295a <=( (not A300)  and  a14294a );
 a14296a <=( a14295a  and  a14290a );
 a14299a <=( (not A169)  and  (not A170) );
 a14303a <=( (not A202)  and  (not A201) );
 a14304a <=( (not A168)  and  a14303a );
 a14305a <=( a14304a  and  a14299a );
 a14309a <=( A267  and  A265 );
 a14310a <=( (not A203)  and  a14309a );
 a14314a <=( (not A301)  and  (not A299) );
 a14315a <=( (not A298)  and  a14314a );
 a14316a <=( a14315a  and  a14310a );
 a14319a <=( (not A169)  and  (not A170) );
 a14323a <=( (not A202)  and  (not A201) );
 a14324a <=( (not A168)  and  a14323a );
 a14325a <=( a14324a  and  a14319a );
 a14329a <=( A267  and  A266 );
 a14330a <=( (not A203)  and  a14329a );
 a14334a <=( (not A302)  and  (not A301) );
 a14335a <=( (not A300)  and  a14334a );
 a14336a <=( a14335a  and  a14330a );
 a14339a <=( (not A169)  and  (not A170) );
 a14343a <=( (not A202)  and  (not A201) );
 a14344a <=( (not A168)  and  a14343a );
 a14345a <=( a14344a  and  a14339a );
 a14349a <=( A267  and  A266 );
 a14350a <=( (not A203)  and  a14349a );
 a14354a <=( (not A301)  and  (not A299) );
 a14355a <=( (not A298)  and  a14354a );
 a14356a <=( a14355a  and  a14350a );
 a14359a <=( (not A169)  and  (not A170) );
 a14363a <=( A201  and  A199 );
 a14364a <=( (not A168)  and  a14363a );
 a14365a <=( a14364a  and  a14359a );
 a14369a <=( (not A269)  and  (not A268) );
 a14370a <=( (not A267)  and  a14369a );
 a14374a <=( A302  and  (not A299) );
 a14375a <=( A298  and  a14374a );
 a14376a <=( a14375a  and  a14370a );
 a14379a <=( (not A169)  and  (not A170) );
 a14383a <=( A201  and  A199 );
 a14384a <=( (not A168)  and  a14383a );
 a14385a <=( a14384a  and  a14379a );
 a14389a <=( (not A269)  and  (not A268) );
 a14390a <=( (not A267)  and  a14389a );
 a14394a <=( A302  and  A299 );
 a14395a <=( (not A298)  and  a14394a );
 a14396a <=( a14395a  and  a14390a );
 a14399a <=( (not A169)  and  (not A170) );
 a14403a <=( A201  and  A199 );
 a14404a <=( (not A168)  and  a14403a );
 a14405a <=( a14404a  and  a14399a );
 a14409a <=( (not A267)  and  A266 );
 a14410a <=( A265  and  a14409a );
 a14414a <=( A300  and  A299 );
 a14415a <=( (not A268)  and  a14414a );
 a14416a <=( a14415a  and  a14410a );
 a14419a <=( (not A169)  and  (not A170) );
 a14423a <=( A201  and  A199 );
 a14424a <=( (not A168)  and  a14423a );
 a14425a <=( a14424a  and  a14419a );
 a14429a <=( (not A267)  and  A266 );
 a14430a <=( A265  and  a14429a );
 a14434a <=( A300  and  A298 );
 a14435a <=( (not A268)  and  a14434a );
 a14436a <=( a14435a  and  a14430a );
 a14439a <=( (not A169)  and  (not A170) );
 a14443a <=( A201  and  A199 );
 a14444a <=( (not A168)  and  a14443a );
 a14445a <=( a14444a  and  a14439a );
 a14449a <=( (not A268)  and  (not A266) );
 a14450a <=( (not A265)  and  a14449a );
 a14454a <=( A302  and  (not A299) );
 a14455a <=( A298  and  a14454a );
 a14456a <=( a14455a  and  a14450a );
 a14459a <=( (not A169)  and  (not A170) );
 a14463a <=( A201  and  A199 );
 a14464a <=( (not A168)  and  a14463a );
 a14465a <=( a14464a  and  a14459a );
 a14469a <=( (not A268)  and  (not A266) );
 a14470a <=( (not A265)  and  a14469a );
 a14474a <=( A302  and  A299 );
 a14475a <=( (not A298)  and  a14474a );
 a14476a <=( a14475a  and  a14470a );
 a14479a <=( (not A169)  and  (not A170) );
 a14483a <=( A201  and  A200 );
 a14484a <=( (not A168)  and  a14483a );
 a14485a <=( a14484a  and  a14479a );
 a14489a <=( (not A269)  and  (not A268) );
 a14490a <=( (not A267)  and  a14489a );
 a14494a <=( A302  and  (not A299) );
 a14495a <=( A298  and  a14494a );
 a14496a <=( a14495a  and  a14490a );
 a14499a <=( (not A169)  and  (not A170) );
 a14503a <=( A201  and  A200 );
 a14504a <=( (not A168)  and  a14503a );
 a14505a <=( a14504a  and  a14499a );
 a14509a <=( (not A269)  and  (not A268) );
 a14510a <=( (not A267)  and  a14509a );
 a14514a <=( A302  and  A299 );
 a14515a <=( (not A298)  and  a14514a );
 a14516a <=( a14515a  and  a14510a );
 a14519a <=( (not A169)  and  (not A170) );
 a14523a <=( A201  and  A200 );
 a14524a <=( (not A168)  and  a14523a );
 a14525a <=( a14524a  and  a14519a );
 a14529a <=( (not A267)  and  A266 );
 a14530a <=( A265  and  a14529a );
 a14534a <=( A300  and  A299 );
 a14535a <=( (not A268)  and  a14534a );
 a14536a <=( a14535a  and  a14530a );
 a14539a <=( (not A169)  and  (not A170) );
 a14543a <=( A201  and  A200 );
 a14544a <=( (not A168)  and  a14543a );
 a14545a <=( a14544a  and  a14539a );
 a14549a <=( (not A267)  and  A266 );
 a14550a <=( A265  and  a14549a );
 a14554a <=( A300  and  A298 );
 a14555a <=( (not A268)  and  a14554a );
 a14556a <=( a14555a  and  a14550a );
 a14559a <=( (not A169)  and  (not A170) );
 a14563a <=( A201  and  A200 );
 a14564a <=( (not A168)  and  a14563a );
 a14565a <=( a14564a  and  a14559a );
 a14569a <=( (not A268)  and  (not A266) );
 a14570a <=( (not A265)  and  a14569a );
 a14574a <=( A302  and  (not A299) );
 a14575a <=( A298  and  a14574a );
 a14576a <=( a14575a  and  a14570a );
 a14579a <=( (not A169)  and  (not A170) );
 a14583a <=( A201  and  A200 );
 a14584a <=( (not A168)  and  a14583a );
 a14585a <=( a14584a  and  a14579a );
 a14589a <=( (not A268)  and  (not A266) );
 a14590a <=( (not A265)  and  a14589a );
 a14594a <=( A302  and  A299 );
 a14595a <=( (not A298)  and  a14594a );
 a14596a <=( a14595a  and  a14590a );
 a14599a <=( (not A169)  and  (not A170) );
 a14603a <=( A200  and  A199 );
 a14604a <=( (not A168)  and  a14603a );
 a14605a <=( a14604a  and  a14599a );
 a14609a <=( A268  and  (not A202) );
 a14610a <=( (not A201)  and  a14609a );
 a14614a <=( (not A302)  and  (not A301) );
 a14615a <=( (not A300)  and  a14614a );
 a14616a <=( a14615a  and  a14610a );
 a14619a <=( (not A169)  and  (not A170) );
 a14623a <=( A200  and  A199 );
 a14624a <=( (not A168)  and  a14623a );
 a14625a <=( a14624a  and  a14619a );
 a14629a <=( A268  and  (not A202) );
 a14630a <=( (not A201)  and  a14629a );
 a14634a <=( (not A301)  and  (not A299) );
 a14635a <=( (not A298)  and  a14634a );
 a14636a <=( a14635a  and  a14630a );
 a14639a <=( (not A169)  and  (not A170) );
 a14643a <=( A200  and  (not A199) );
 a14644a <=( (not A168)  and  a14643a );
 a14645a <=( a14644a  and  a14639a );
 a14649a <=( (not A268)  and  (not A267) );
 a14650a <=( A203  and  a14649a );
 a14654a <=( A300  and  A299 );
 a14655a <=( (not A269)  and  a14654a );
 a14656a <=( a14655a  and  a14650a );
 a14659a <=( (not A169)  and  (not A170) );
 a14663a <=( A200  and  (not A199) );
 a14664a <=( (not A168)  and  a14663a );
 a14665a <=( a14664a  and  a14659a );
 a14669a <=( (not A268)  and  (not A267) );
 a14670a <=( A203  and  a14669a );
 a14674a <=( A300  and  A298 );
 a14675a <=( (not A269)  and  a14674a );
 a14676a <=( a14675a  and  a14670a );
 a14679a <=( (not A169)  and  (not A170) );
 a14683a <=( A200  and  (not A199) );
 a14684a <=( (not A168)  and  a14683a );
 a14685a <=( a14684a  and  a14679a );
 a14689a <=( A266  and  A265 );
 a14690a <=( A203  and  a14689a );
 a14694a <=( A301  and  (not A268) );
 a14695a <=( (not A267)  and  a14694a );
 a14696a <=( a14695a  and  a14690a );
 a14699a <=( (not A169)  and  (not A170) );
 a14703a <=( A200  and  (not A199) );
 a14704a <=( (not A168)  and  a14703a );
 a14705a <=( a14704a  and  a14699a );
 a14709a <=( (not A266)  and  (not A265) );
 a14710a <=( A203  and  a14709a );
 a14714a <=( A300  and  A299 );
 a14715a <=( (not A268)  and  a14714a );
 a14716a <=( a14715a  and  a14710a );
 a14719a <=( (not A169)  and  (not A170) );
 a14723a <=( A200  and  (not A199) );
 a14724a <=( (not A168)  and  a14723a );
 a14725a <=( a14724a  and  a14719a );
 a14729a <=( (not A266)  and  (not A265) );
 a14730a <=( A203  and  a14729a );
 a14734a <=( A300  and  A298 );
 a14735a <=( (not A268)  and  a14734a );
 a14736a <=( a14735a  and  a14730a );
 a14739a <=( (not A169)  and  (not A170) );
 a14743a <=( (not A200)  and  A199 );
 a14744a <=( (not A168)  and  a14743a );
 a14745a <=( a14744a  and  a14739a );
 a14749a <=( (not A268)  and  (not A267) );
 a14750a <=( A203  and  a14749a );
 a14754a <=( A300  and  A299 );
 a14755a <=( (not A269)  and  a14754a );
 a14756a <=( a14755a  and  a14750a );
 a14759a <=( (not A169)  and  (not A170) );
 a14763a <=( (not A200)  and  A199 );
 a14764a <=( (not A168)  and  a14763a );
 a14765a <=( a14764a  and  a14759a );
 a14769a <=( (not A268)  and  (not A267) );
 a14770a <=( A203  and  a14769a );
 a14774a <=( A300  and  A298 );
 a14775a <=( (not A269)  and  a14774a );
 a14776a <=( a14775a  and  a14770a );
 a14779a <=( (not A169)  and  (not A170) );
 a14783a <=( (not A200)  and  A199 );
 a14784a <=( (not A168)  and  a14783a );
 a14785a <=( a14784a  and  a14779a );
 a14789a <=( A266  and  A265 );
 a14790a <=( A203  and  a14789a );
 a14794a <=( A301  and  (not A268) );
 a14795a <=( (not A267)  and  a14794a );
 a14796a <=( a14795a  and  a14790a );
 a14799a <=( (not A169)  and  (not A170) );
 a14803a <=( (not A200)  and  A199 );
 a14804a <=( (not A168)  and  a14803a );
 a14805a <=( a14804a  and  a14799a );
 a14809a <=( (not A266)  and  (not A265) );
 a14810a <=( A203  and  a14809a );
 a14814a <=( A300  and  A299 );
 a14815a <=( (not A268)  and  a14814a );
 a14816a <=( a14815a  and  a14810a );
 a14819a <=( (not A169)  and  (not A170) );
 a14823a <=( (not A200)  and  A199 );
 a14824a <=( (not A168)  and  a14823a );
 a14825a <=( a14824a  and  a14819a );
 a14829a <=( (not A266)  and  (not A265) );
 a14830a <=( A203  and  a14829a );
 a14834a <=( A300  and  A298 );
 a14835a <=( (not A268)  and  a14834a );
 a14836a <=( a14835a  and  a14830a );
 a14839a <=( (not A169)  and  (not A170) );
 a14843a <=( (not A200)  and  (not A199) );
 a14844a <=( (not A168)  and  a14843a );
 a14845a <=( a14844a  and  a14839a );
 a14849a <=( A298  and  A268 );
 a14850a <=( (not A202)  and  a14849a );
 a14854a <=( (not A301)  and  (not A300) );
 a14855a <=( A299  and  a14854a );
 a14856a <=( a14855a  and  a14850a );
 a14859a <=( (not A169)  and  (not A170) );
 a14863a <=( (not A200)  and  (not A199) );
 a14864a <=( (not A168)  and  a14863a );
 a14865a <=( a14864a  and  a14859a );
 a14869a <=( A267  and  A265 );
 a14870a <=( (not A202)  and  a14869a );
 a14874a <=( (not A302)  and  (not A301) );
 a14875a <=( (not A300)  and  a14874a );
 a14876a <=( a14875a  and  a14870a );
 a14879a <=( (not A169)  and  (not A170) );
 a14883a <=( (not A200)  and  (not A199) );
 a14884a <=( (not A168)  and  a14883a );
 a14885a <=( a14884a  and  a14879a );
 a14889a <=( A267  and  A265 );
 a14890a <=( (not A202)  and  a14889a );
 a14894a <=( (not A301)  and  (not A299) );
 a14895a <=( (not A298)  and  a14894a );
 a14896a <=( a14895a  and  a14890a );
 a14899a <=( (not A169)  and  (not A170) );
 a14903a <=( (not A200)  and  (not A199) );
 a14904a <=( (not A168)  and  a14903a );
 a14905a <=( a14904a  and  a14899a );
 a14909a <=( A267  and  A266 );
 a14910a <=( (not A202)  and  a14909a );
 a14914a <=( (not A302)  and  (not A301) );
 a14915a <=( (not A300)  and  a14914a );
 a14916a <=( a14915a  and  a14910a );
 a14919a <=( (not A169)  and  (not A170) );
 a14923a <=( (not A200)  and  (not A199) );
 a14924a <=( (not A168)  and  a14923a );
 a14925a <=( a14924a  and  a14919a );
 a14929a <=( A267  and  A266 );
 a14930a <=( (not A202)  and  a14929a );
 a14934a <=( (not A301)  and  (not A299) );
 a14935a <=( (not A298)  and  a14934a );
 a14936a <=( a14935a  and  a14930a );
 a14940a <=( (not A201)  and  A166 );
 a14941a <=( A168  and  a14940a );
 a14945a <=( A265  and  (not A203) );
 a14946a <=( (not A202)  and  a14945a );
 a14947a <=( a14946a  and  a14941a );
 a14951a <=( (not A268)  and  (not A267) );
 a14952a <=( A266  and  a14951a );
 a14956a <=( A302  and  (not A299) );
 a14957a <=( A298  and  a14956a );
 a14958a <=( a14957a  and  a14952a );
 a14962a <=( (not A201)  and  A166 );
 a14963a <=( A168  and  a14962a );
 a14967a <=( A265  and  (not A203) );
 a14968a <=( (not A202)  and  a14967a );
 a14969a <=( a14968a  and  a14963a );
 a14973a <=( (not A268)  and  (not A267) );
 a14974a <=( A266  and  a14973a );
 a14978a <=( A302  and  A299 );
 a14979a <=( (not A298)  and  a14978a );
 a14980a <=( a14979a  and  a14974a );
 a14984a <=( A199  and  A166 );
 a14985a <=( A168  and  a14984a );
 a14989a <=( (not A202)  and  (not A201) );
 a14990a <=( A200  and  a14989a );
 a14991a <=( a14990a  and  a14985a );
 a14995a <=( (not A269)  and  (not A268) );
 a14996a <=( (not A267)  and  a14995a );
 a15000a <=( A302  and  (not A299) );
 a15001a <=( A298  and  a15000a );
 a15002a <=( a15001a  and  a14996a );
 a15006a <=( A199  and  A166 );
 a15007a <=( A168  and  a15006a );
 a15011a <=( (not A202)  and  (not A201) );
 a15012a <=( A200  and  a15011a );
 a15013a <=( a15012a  and  a15007a );
 a15017a <=( (not A269)  and  (not A268) );
 a15018a <=( (not A267)  and  a15017a );
 a15022a <=( A302  and  A299 );
 a15023a <=( (not A298)  and  a15022a );
 a15024a <=( a15023a  and  a15018a );
 a15028a <=( A199  and  A166 );
 a15029a <=( A168  and  a15028a );
 a15033a <=( (not A202)  and  (not A201) );
 a15034a <=( A200  and  a15033a );
 a15035a <=( a15034a  and  a15029a );
 a15039a <=( (not A267)  and  A266 );
 a15040a <=( A265  and  a15039a );
 a15044a <=( A300  and  A299 );
 a15045a <=( (not A268)  and  a15044a );
 a15046a <=( a15045a  and  a15040a );
 a15050a <=( A199  and  A166 );
 a15051a <=( A168  and  a15050a );
 a15055a <=( (not A202)  and  (not A201) );
 a15056a <=( A200  and  a15055a );
 a15057a <=( a15056a  and  a15051a );
 a15061a <=( (not A267)  and  A266 );
 a15062a <=( A265  and  a15061a );
 a15066a <=( A300  and  A298 );
 a15067a <=( (not A268)  and  a15066a );
 a15068a <=( a15067a  and  a15062a );
 a15072a <=( A199  and  A166 );
 a15073a <=( A168  and  a15072a );
 a15077a <=( (not A202)  and  (not A201) );
 a15078a <=( A200  and  a15077a );
 a15079a <=( a15078a  and  a15073a );
 a15083a <=( (not A268)  and  (not A266) );
 a15084a <=( (not A265)  and  a15083a );
 a15088a <=( A302  and  (not A299) );
 a15089a <=( A298  and  a15088a );
 a15090a <=( a15089a  and  a15084a );
 a15094a <=( A199  and  A166 );
 a15095a <=( A168  and  a15094a );
 a15099a <=( (not A202)  and  (not A201) );
 a15100a <=( A200  and  a15099a );
 a15101a <=( a15100a  and  a15095a );
 a15105a <=( (not A268)  and  (not A266) );
 a15106a <=( (not A265)  and  a15105a );
 a15110a <=( A302  and  A299 );
 a15111a <=( (not A298)  and  a15110a );
 a15112a <=( a15111a  and  a15106a );
 a15116a <=( (not A199)  and  A166 );
 a15117a <=( A168  and  a15116a );
 a15121a <=( (not A265)  and  A203 );
 a15122a <=( A200  and  a15121a );
 a15123a <=( a15122a  and  a15117a );
 a15127a <=( A298  and  A269 );
 a15128a <=( A266  and  a15127a );
 a15132a <=( (not A301)  and  (not A300) );
 a15133a <=( A299  and  a15132a );
 a15134a <=( a15133a  and  a15128a );
 a15138a <=( (not A199)  and  A166 );
 a15139a <=( A168  and  a15138a );
 a15143a <=( A265  and  A203 );
 a15144a <=( A200  and  a15143a );
 a15145a <=( a15144a  and  a15139a );
 a15149a <=( A298  and  A269 );
 a15150a <=( (not A266)  and  a15149a );
 a15154a <=( (not A301)  and  (not A300) );
 a15155a <=( A299  and  a15154a );
 a15156a <=( a15155a  and  a15150a );
 a15160a <=( A199  and  A166 );
 a15161a <=( A168  and  a15160a );
 a15165a <=( (not A265)  and  A203 );
 a15166a <=( (not A200)  and  a15165a );
 a15167a <=( a15166a  and  a15161a );
 a15171a <=( A298  and  A269 );
 a15172a <=( A266  and  a15171a );
 a15176a <=( (not A301)  and  (not A300) );
 a15177a <=( A299  and  a15176a );
 a15178a <=( a15177a  and  a15172a );
 a15182a <=( A199  and  A166 );
 a15183a <=( A168  and  a15182a );
 a15187a <=( A265  and  A203 );
 a15188a <=( (not A200)  and  a15187a );
 a15189a <=( a15188a  and  a15183a );
 a15193a <=( A298  and  A269 );
 a15194a <=( (not A266)  and  a15193a );
 a15198a <=( (not A301)  and  (not A300) );
 a15199a <=( A299  and  a15198a );
 a15200a <=( a15199a  and  a15194a );
 a15204a <=( (not A199)  and  A166 );
 a15205a <=( A168  and  a15204a );
 a15209a <=( A265  and  (not A202) );
 a15210a <=( (not A200)  and  a15209a );
 a15211a <=( a15210a  and  a15205a );
 a15215a <=( (not A268)  and  (not A267) );
 a15216a <=( A266  and  a15215a );
 a15220a <=( A302  and  (not A299) );
 a15221a <=( A298  and  a15220a );
 a15222a <=( a15221a  and  a15216a );
 a15226a <=( (not A199)  and  A166 );
 a15227a <=( A168  and  a15226a );
 a15231a <=( A265  and  (not A202) );
 a15232a <=( (not A200)  and  a15231a );
 a15233a <=( a15232a  and  a15227a );
 a15237a <=( (not A268)  and  (not A267) );
 a15238a <=( A266  and  a15237a );
 a15242a <=( A302  and  A299 );
 a15243a <=( (not A298)  and  a15242a );
 a15244a <=( a15243a  and  a15238a );
 a15248a <=( (not A201)  and  A167 );
 a15249a <=( A168  and  a15248a );
 a15253a <=( A265  and  (not A203) );
 a15254a <=( (not A202)  and  a15253a );
 a15255a <=( a15254a  and  a15249a );
 a15259a <=( (not A268)  and  (not A267) );
 a15260a <=( A266  and  a15259a );
 a15264a <=( A302  and  (not A299) );
 a15265a <=( A298  and  a15264a );
 a15266a <=( a15265a  and  a15260a );
 a15270a <=( (not A201)  and  A167 );
 a15271a <=( A168  and  a15270a );
 a15275a <=( A265  and  (not A203) );
 a15276a <=( (not A202)  and  a15275a );
 a15277a <=( a15276a  and  a15271a );
 a15281a <=( (not A268)  and  (not A267) );
 a15282a <=( A266  and  a15281a );
 a15286a <=( A302  and  A299 );
 a15287a <=( (not A298)  and  a15286a );
 a15288a <=( a15287a  and  a15282a );
 a15292a <=( A199  and  A167 );
 a15293a <=( A168  and  a15292a );
 a15297a <=( (not A202)  and  (not A201) );
 a15298a <=( A200  and  a15297a );
 a15299a <=( a15298a  and  a15293a );
 a15303a <=( (not A269)  and  (not A268) );
 a15304a <=( (not A267)  and  a15303a );
 a15308a <=( A302  and  (not A299) );
 a15309a <=( A298  and  a15308a );
 a15310a <=( a15309a  and  a15304a );
 a15314a <=( A199  and  A167 );
 a15315a <=( A168  and  a15314a );
 a15319a <=( (not A202)  and  (not A201) );
 a15320a <=( A200  and  a15319a );
 a15321a <=( a15320a  and  a15315a );
 a15325a <=( (not A269)  and  (not A268) );
 a15326a <=( (not A267)  and  a15325a );
 a15330a <=( A302  and  A299 );
 a15331a <=( (not A298)  and  a15330a );
 a15332a <=( a15331a  and  a15326a );
 a15336a <=( A199  and  A167 );
 a15337a <=( A168  and  a15336a );
 a15341a <=( (not A202)  and  (not A201) );
 a15342a <=( A200  and  a15341a );
 a15343a <=( a15342a  and  a15337a );
 a15347a <=( (not A267)  and  A266 );
 a15348a <=( A265  and  a15347a );
 a15352a <=( A300  and  A299 );
 a15353a <=( (not A268)  and  a15352a );
 a15354a <=( a15353a  and  a15348a );
 a15358a <=( A199  and  A167 );
 a15359a <=( A168  and  a15358a );
 a15363a <=( (not A202)  and  (not A201) );
 a15364a <=( A200  and  a15363a );
 a15365a <=( a15364a  and  a15359a );
 a15369a <=( (not A267)  and  A266 );
 a15370a <=( A265  and  a15369a );
 a15374a <=( A300  and  A298 );
 a15375a <=( (not A268)  and  a15374a );
 a15376a <=( a15375a  and  a15370a );
 a15380a <=( A199  and  A167 );
 a15381a <=( A168  and  a15380a );
 a15385a <=( (not A202)  and  (not A201) );
 a15386a <=( A200  and  a15385a );
 a15387a <=( a15386a  and  a15381a );
 a15391a <=( (not A268)  and  (not A266) );
 a15392a <=( (not A265)  and  a15391a );
 a15396a <=( A302  and  (not A299) );
 a15397a <=( A298  and  a15396a );
 a15398a <=( a15397a  and  a15392a );
 a15402a <=( A199  and  A167 );
 a15403a <=( A168  and  a15402a );
 a15407a <=( (not A202)  and  (not A201) );
 a15408a <=( A200  and  a15407a );
 a15409a <=( a15408a  and  a15403a );
 a15413a <=( (not A268)  and  (not A266) );
 a15414a <=( (not A265)  and  a15413a );
 a15418a <=( A302  and  A299 );
 a15419a <=( (not A298)  and  a15418a );
 a15420a <=( a15419a  and  a15414a );
 a15424a <=( (not A199)  and  A167 );
 a15425a <=( A168  and  a15424a );
 a15429a <=( (not A265)  and  A203 );
 a15430a <=( A200  and  a15429a );
 a15431a <=( a15430a  and  a15425a );
 a15435a <=( A298  and  A269 );
 a15436a <=( A266  and  a15435a );
 a15440a <=( (not A301)  and  (not A300) );
 a15441a <=( A299  and  a15440a );
 a15442a <=( a15441a  and  a15436a );
 a15446a <=( (not A199)  and  A167 );
 a15447a <=( A168  and  a15446a );
 a15451a <=( A265  and  A203 );
 a15452a <=( A200  and  a15451a );
 a15453a <=( a15452a  and  a15447a );
 a15457a <=( A298  and  A269 );
 a15458a <=( (not A266)  and  a15457a );
 a15462a <=( (not A301)  and  (not A300) );
 a15463a <=( A299  and  a15462a );
 a15464a <=( a15463a  and  a15458a );
 a15468a <=( A199  and  A167 );
 a15469a <=( A168  and  a15468a );
 a15473a <=( (not A265)  and  A203 );
 a15474a <=( (not A200)  and  a15473a );
 a15475a <=( a15474a  and  a15469a );
 a15479a <=( A298  and  A269 );
 a15480a <=( A266  and  a15479a );
 a15484a <=( (not A301)  and  (not A300) );
 a15485a <=( A299  and  a15484a );
 a15486a <=( a15485a  and  a15480a );
 a15490a <=( A199  and  A167 );
 a15491a <=( A168  and  a15490a );
 a15495a <=( A265  and  A203 );
 a15496a <=( (not A200)  and  a15495a );
 a15497a <=( a15496a  and  a15491a );
 a15501a <=( A298  and  A269 );
 a15502a <=( (not A266)  and  a15501a );
 a15506a <=( (not A301)  and  (not A300) );
 a15507a <=( A299  and  a15506a );
 a15508a <=( a15507a  and  a15502a );
 a15512a <=( (not A199)  and  A167 );
 a15513a <=( A168  and  a15512a );
 a15517a <=( A265  and  (not A202) );
 a15518a <=( (not A200)  and  a15517a );
 a15519a <=( a15518a  and  a15513a );
 a15523a <=( (not A268)  and  (not A267) );
 a15524a <=( A266  and  a15523a );
 a15528a <=( A302  and  (not A299) );
 a15529a <=( A298  and  a15528a );
 a15530a <=( a15529a  and  a15524a );
 a15534a <=( (not A199)  and  A167 );
 a15535a <=( A168  and  a15534a );
 a15539a <=( A265  and  (not A202) );
 a15540a <=( (not A200)  and  a15539a );
 a15541a <=( a15540a  and  a15535a );
 a15545a <=( (not A268)  and  (not A267) );
 a15546a <=( A266  and  a15545a );
 a15550a <=( A302  and  A299 );
 a15551a <=( (not A298)  and  a15550a );
 a15552a <=( a15551a  and  a15546a );
 a15556a <=( (not A166)  and  A167 );
 a15557a <=( A170  and  a15556a );
 a15561a <=( (not A203)  and  (not A202) );
 a15562a <=( (not A201)  and  a15561a );
 a15563a <=( a15562a  and  a15557a );
 a15567a <=( (not A269)  and  (not A268) );
 a15568a <=( (not A267)  and  a15567a );
 a15572a <=( A302  and  (not A299) );
 a15573a <=( A298  and  a15572a );
 a15574a <=( a15573a  and  a15568a );
 a15578a <=( (not A166)  and  A167 );
 a15579a <=( A170  and  a15578a );
 a15583a <=( (not A203)  and  (not A202) );
 a15584a <=( (not A201)  and  a15583a );
 a15585a <=( a15584a  and  a15579a );
 a15589a <=( (not A269)  and  (not A268) );
 a15590a <=( (not A267)  and  a15589a );
 a15594a <=( A302  and  A299 );
 a15595a <=( (not A298)  and  a15594a );
 a15596a <=( a15595a  and  a15590a );
 a15600a <=( (not A166)  and  A167 );
 a15601a <=( A170  and  a15600a );
 a15605a <=( (not A203)  and  (not A202) );
 a15606a <=( (not A201)  and  a15605a );
 a15607a <=( a15606a  and  a15601a );
 a15611a <=( (not A267)  and  A266 );
 a15612a <=( A265  and  a15611a );
 a15616a <=( A300  and  A299 );
 a15617a <=( (not A268)  and  a15616a );
 a15618a <=( a15617a  and  a15612a );
 a15622a <=( (not A166)  and  A167 );
 a15623a <=( A170  and  a15622a );
 a15627a <=( (not A203)  and  (not A202) );
 a15628a <=( (not A201)  and  a15627a );
 a15629a <=( a15628a  and  a15623a );
 a15633a <=( (not A267)  and  A266 );
 a15634a <=( A265  and  a15633a );
 a15638a <=( A300  and  A298 );
 a15639a <=( (not A268)  and  a15638a );
 a15640a <=( a15639a  and  a15634a );
 a15644a <=( (not A166)  and  A167 );
 a15645a <=( A170  and  a15644a );
 a15649a <=( (not A203)  and  (not A202) );
 a15650a <=( (not A201)  and  a15649a );
 a15651a <=( a15650a  and  a15645a );
 a15655a <=( (not A268)  and  (not A266) );
 a15656a <=( (not A265)  and  a15655a );
 a15660a <=( A302  and  (not A299) );
 a15661a <=( A298  and  a15660a );
 a15662a <=( a15661a  and  a15656a );
 a15666a <=( (not A166)  and  A167 );
 a15667a <=( A170  and  a15666a );
 a15671a <=( (not A203)  and  (not A202) );
 a15672a <=( (not A201)  and  a15671a );
 a15673a <=( a15672a  and  a15667a );
 a15677a <=( (not A268)  and  (not A266) );
 a15678a <=( (not A265)  and  a15677a );
 a15682a <=( A302  and  A299 );
 a15683a <=( (not A298)  and  a15682a );
 a15684a <=( a15683a  and  a15678a );
 a15688a <=( (not A166)  and  A167 );
 a15689a <=( A170  and  a15688a );
 a15693a <=( (not A265)  and  A201 );
 a15694a <=( A199  and  a15693a );
 a15695a <=( a15694a  and  a15689a );
 a15699a <=( A298  and  A269 );
 a15700a <=( A266  and  a15699a );
 a15704a <=( (not A301)  and  (not A300) );
 a15705a <=( A299  and  a15704a );
 a15706a <=( a15705a  and  a15700a );
 a15710a <=( (not A166)  and  A167 );
 a15711a <=( A170  and  a15710a );
 a15715a <=( A265  and  A201 );
 a15716a <=( A199  and  a15715a );
 a15717a <=( a15716a  and  a15711a );
 a15721a <=( A298  and  A269 );
 a15722a <=( (not A266)  and  a15721a );
 a15726a <=( (not A301)  and  (not A300) );
 a15727a <=( A299  and  a15726a );
 a15728a <=( a15727a  and  a15722a );
 a15732a <=( (not A166)  and  A167 );
 a15733a <=( A170  and  a15732a );
 a15737a <=( (not A265)  and  A201 );
 a15738a <=( A200  and  a15737a );
 a15739a <=( a15738a  and  a15733a );
 a15743a <=( A298  and  A269 );
 a15744a <=( A266  and  a15743a );
 a15748a <=( (not A301)  and  (not A300) );
 a15749a <=( A299  and  a15748a );
 a15750a <=( a15749a  and  a15744a );
 a15754a <=( (not A166)  and  A167 );
 a15755a <=( A170  and  a15754a );
 a15759a <=( A265  and  A201 );
 a15760a <=( A200  and  a15759a );
 a15761a <=( a15760a  and  a15755a );
 a15765a <=( A298  and  A269 );
 a15766a <=( (not A266)  and  a15765a );
 a15770a <=( (not A301)  and  (not A300) );
 a15771a <=( A299  and  a15770a );
 a15772a <=( a15771a  and  a15766a );
 a15776a <=( (not A166)  and  A167 );
 a15777a <=( A170  and  a15776a );
 a15781a <=( (not A201)  and  A200 );
 a15782a <=( A199  and  a15781a );
 a15783a <=( a15782a  and  a15777a );
 a15787a <=( (not A268)  and  (not A267) );
 a15788a <=( (not A202)  and  a15787a );
 a15792a <=( A300  and  A299 );
 a15793a <=( (not A269)  and  a15792a );
 a15794a <=( a15793a  and  a15788a );
 a15798a <=( (not A166)  and  A167 );
 a15799a <=( A170  and  a15798a );
 a15803a <=( (not A201)  and  A200 );
 a15804a <=( A199  and  a15803a );
 a15805a <=( a15804a  and  a15799a );
 a15809a <=( (not A268)  and  (not A267) );
 a15810a <=( (not A202)  and  a15809a );
 a15814a <=( A300  and  A298 );
 a15815a <=( (not A269)  and  a15814a );
 a15816a <=( a15815a  and  a15810a );
 a15820a <=( (not A166)  and  A167 );
 a15821a <=( A170  and  a15820a );
 a15825a <=( (not A201)  and  A200 );
 a15826a <=( A199  and  a15825a );
 a15827a <=( a15826a  and  a15821a );
 a15831a <=( A266  and  A265 );
 a15832a <=( (not A202)  and  a15831a );
 a15836a <=( A301  and  (not A268) );
 a15837a <=( (not A267)  and  a15836a );
 a15838a <=( a15837a  and  a15832a );
 a15842a <=( (not A166)  and  A167 );
 a15843a <=( A170  and  a15842a );
 a15847a <=( (not A201)  and  A200 );
 a15848a <=( A199  and  a15847a );
 a15849a <=( a15848a  and  a15843a );
 a15853a <=( (not A266)  and  (not A265) );
 a15854a <=( (not A202)  and  a15853a );
 a15858a <=( A300  and  A299 );
 a15859a <=( (not A268)  and  a15858a );
 a15860a <=( a15859a  and  a15854a );
 a15864a <=( (not A166)  and  A167 );
 a15865a <=( A170  and  a15864a );
 a15869a <=( (not A201)  and  A200 );
 a15870a <=( A199  and  a15869a );
 a15871a <=( a15870a  and  a15865a );
 a15875a <=( (not A266)  and  (not A265) );
 a15876a <=( (not A202)  and  a15875a );
 a15880a <=( A300  and  A298 );
 a15881a <=( (not A268)  and  a15880a );
 a15882a <=( a15881a  and  a15876a );
 a15886a <=( (not A166)  and  A167 );
 a15887a <=( A170  and  a15886a );
 a15891a <=( A203  and  A200 );
 a15892a <=( (not A199)  and  a15891a );
 a15893a <=( a15892a  and  a15887a );
 a15897a <=( A298  and  A267 );
 a15898a <=( A265  and  a15897a );
 a15902a <=( (not A301)  and  (not A300) );
 a15903a <=( A299  and  a15902a );
 a15904a <=( a15903a  and  a15898a );
 a15908a <=( (not A166)  and  A167 );
 a15909a <=( A170  and  a15908a );
 a15913a <=( A203  and  A200 );
 a15914a <=( (not A199)  and  a15913a );
 a15915a <=( a15914a  and  a15909a );
 a15919a <=( A298  and  A267 );
 a15920a <=( A266  and  a15919a );
 a15924a <=( (not A301)  and  (not A300) );
 a15925a <=( A299  and  a15924a );
 a15926a <=( a15925a  and  a15920a );
 a15930a <=( (not A166)  and  A167 );
 a15931a <=( A170  and  a15930a );
 a15935a <=( A203  and  A200 );
 a15936a <=( (not A199)  and  a15935a );
 a15937a <=( a15936a  and  a15931a );
 a15941a <=( A269  and  A266 );
 a15942a <=( (not A265)  and  a15941a );
 a15946a <=( (not A302)  and  (not A301) );
 a15947a <=( (not A300)  and  a15946a );
 a15948a <=( a15947a  and  a15942a );
 a15952a <=( (not A166)  and  A167 );
 a15953a <=( A170  and  a15952a );
 a15957a <=( A203  and  A200 );
 a15958a <=( (not A199)  and  a15957a );
 a15959a <=( a15958a  and  a15953a );
 a15963a <=( A269  and  A266 );
 a15964a <=( (not A265)  and  a15963a );
 a15968a <=( (not A301)  and  (not A299) );
 a15969a <=( (not A298)  and  a15968a );
 a15970a <=( a15969a  and  a15964a );
 a15974a <=( (not A166)  and  A167 );
 a15975a <=( A170  and  a15974a );
 a15979a <=( A203  and  A200 );
 a15980a <=( (not A199)  and  a15979a );
 a15981a <=( a15980a  and  a15975a );
 a15985a <=( A269  and  (not A266) );
 a15986a <=( A265  and  a15985a );
 a15990a <=( (not A302)  and  (not A301) );
 a15991a <=( (not A300)  and  a15990a );
 a15992a <=( a15991a  and  a15986a );
 a15996a <=( (not A166)  and  A167 );
 a15997a <=( A170  and  a15996a );
 a16001a <=( A203  and  A200 );
 a16002a <=( (not A199)  and  a16001a );
 a16003a <=( a16002a  and  a15997a );
 a16007a <=( A269  and  (not A266) );
 a16008a <=( A265  and  a16007a );
 a16012a <=( (not A301)  and  (not A299) );
 a16013a <=( (not A298)  and  a16012a );
 a16014a <=( a16013a  and  a16008a );
 a16018a <=( (not A166)  and  A167 );
 a16019a <=( A170  and  a16018a );
 a16023a <=( A203  and  (not A200) );
 a16024a <=( A199  and  a16023a );
 a16025a <=( a16024a  and  a16019a );
 a16029a <=( A298  and  A267 );
 a16030a <=( A265  and  a16029a );
 a16034a <=( (not A301)  and  (not A300) );
 a16035a <=( A299  and  a16034a );
 a16036a <=( a16035a  and  a16030a );
 a16040a <=( (not A166)  and  A167 );
 a16041a <=( A170  and  a16040a );
 a16045a <=( A203  and  (not A200) );
 a16046a <=( A199  and  a16045a );
 a16047a <=( a16046a  and  a16041a );
 a16051a <=( A298  and  A267 );
 a16052a <=( A266  and  a16051a );
 a16056a <=( (not A301)  and  (not A300) );
 a16057a <=( A299  and  a16056a );
 a16058a <=( a16057a  and  a16052a );
 a16062a <=( (not A166)  and  A167 );
 a16063a <=( A170  and  a16062a );
 a16067a <=( A203  and  (not A200) );
 a16068a <=( A199  and  a16067a );
 a16069a <=( a16068a  and  a16063a );
 a16073a <=( A269  and  A266 );
 a16074a <=( (not A265)  and  a16073a );
 a16078a <=( (not A302)  and  (not A301) );
 a16079a <=( (not A300)  and  a16078a );
 a16080a <=( a16079a  and  a16074a );
 a16084a <=( (not A166)  and  A167 );
 a16085a <=( A170  and  a16084a );
 a16089a <=( A203  and  (not A200) );
 a16090a <=( A199  and  a16089a );
 a16091a <=( a16090a  and  a16085a );
 a16095a <=( A269  and  A266 );
 a16096a <=( (not A265)  and  a16095a );
 a16100a <=( (not A301)  and  (not A299) );
 a16101a <=( (not A298)  and  a16100a );
 a16102a <=( a16101a  and  a16096a );
 a16106a <=( (not A166)  and  A167 );
 a16107a <=( A170  and  a16106a );
 a16111a <=( A203  and  (not A200) );
 a16112a <=( A199  and  a16111a );
 a16113a <=( a16112a  and  a16107a );
 a16117a <=( A269  and  (not A266) );
 a16118a <=( A265  and  a16117a );
 a16122a <=( (not A302)  and  (not A301) );
 a16123a <=( (not A300)  and  a16122a );
 a16124a <=( a16123a  and  a16118a );
 a16128a <=( (not A166)  and  A167 );
 a16129a <=( A170  and  a16128a );
 a16133a <=( A203  and  (not A200) );
 a16134a <=( A199  and  a16133a );
 a16135a <=( a16134a  and  a16129a );
 a16139a <=( A269  and  (not A266) );
 a16140a <=( A265  and  a16139a );
 a16144a <=( (not A301)  and  (not A299) );
 a16145a <=( (not A298)  and  a16144a );
 a16146a <=( a16145a  and  a16140a );
 a16150a <=( (not A166)  and  A167 );
 a16151a <=( A170  and  a16150a );
 a16155a <=( (not A202)  and  (not A200) );
 a16156a <=( (not A199)  and  a16155a );
 a16157a <=( a16156a  and  a16151a );
 a16161a <=( (not A269)  and  (not A268) );
 a16162a <=( (not A267)  and  a16161a );
 a16166a <=( A302  and  (not A299) );
 a16167a <=( A298  and  a16166a );
 a16168a <=( a16167a  and  a16162a );
 a16172a <=( (not A166)  and  A167 );
 a16173a <=( A170  and  a16172a );
 a16177a <=( (not A202)  and  (not A200) );
 a16178a <=( (not A199)  and  a16177a );
 a16179a <=( a16178a  and  a16173a );
 a16183a <=( (not A269)  and  (not A268) );
 a16184a <=( (not A267)  and  a16183a );
 a16188a <=( A302  and  A299 );
 a16189a <=( (not A298)  and  a16188a );
 a16190a <=( a16189a  and  a16184a );
 a16194a <=( (not A166)  and  A167 );
 a16195a <=( A170  and  a16194a );
 a16199a <=( (not A202)  and  (not A200) );
 a16200a <=( (not A199)  and  a16199a );
 a16201a <=( a16200a  and  a16195a );
 a16205a <=( (not A267)  and  A266 );
 a16206a <=( A265  and  a16205a );
 a16210a <=( A300  and  A299 );
 a16211a <=( (not A268)  and  a16210a );
 a16212a <=( a16211a  and  a16206a );
 a16216a <=( (not A166)  and  A167 );
 a16217a <=( A170  and  a16216a );
 a16221a <=( (not A202)  and  (not A200) );
 a16222a <=( (not A199)  and  a16221a );
 a16223a <=( a16222a  and  a16217a );
 a16227a <=( (not A267)  and  A266 );
 a16228a <=( A265  and  a16227a );
 a16232a <=( A300  and  A298 );
 a16233a <=( (not A268)  and  a16232a );
 a16234a <=( a16233a  and  a16228a );
 a16238a <=( (not A166)  and  A167 );
 a16239a <=( A170  and  a16238a );
 a16243a <=( (not A202)  and  (not A200) );
 a16244a <=( (not A199)  and  a16243a );
 a16245a <=( a16244a  and  a16239a );
 a16249a <=( (not A268)  and  (not A266) );
 a16250a <=( (not A265)  and  a16249a );
 a16254a <=( A302  and  (not A299) );
 a16255a <=( A298  and  a16254a );
 a16256a <=( a16255a  and  a16250a );
 a16260a <=( (not A166)  and  A167 );
 a16261a <=( A170  and  a16260a );
 a16265a <=( (not A202)  and  (not A200) );
 a16266a <=( (not A199)  and  a16265a );
 a16267a <=( a16266a  and  a16261a );
 a16271a <=( (not A268)  and  (not A266) );
 a16272a <=( (not A265)  and  a16271a );
 a16276a <=( A302  and  A299 );
 a16277a <=( (not A298)  and  a16276a );
 a16278a <=( a16277a  and  a16272a );
 a16282a <=( A166  and  (not A167) );
 a16283a <=( A170  and  a16282a );
 a16287a <=( (not A203)  and  (not A202) );
 a16288a <=( (not A201)  and  a16287a );
 a16289a <=( a16288a  and  a16283a );
 a16293a <=( (not A269)  and  (not A268) );
 a16294a <=( (not A267)  and  a16293a );
 a16298a <=( A302  and  (not A299) );
 a16299a <=( A298  and  a16298a );
 a16300a <=( a16299a  and  a16294a );
 a16304a <=( A166  and  (not A167) );
 a16305a <=( A170  and  a16304a );
 a16309a <=( (not A203)  and  (not A202) );
 a16310a <=( (not A201)  and  a16309a );
 a16311a <=( a16310a  and  a16305a );
 a16315a <=( (not A269)  and  (not A268) );
 a16316a <=( (not A267)  and  a16315a );
 a16320a <=( A302  and  A299 );
 a16321a <=( (not A298)  and  a16320a );
 a16322a <=( a16321a  and  a16316a );
 a16326a <=( A166  and  (not A167) );
 a16327a <=( A170  and  a16326a );
 a16331a <=( (not A203)  and  (not A202) );
 a16332a <=( (not A201)  and  a16331a );
 a16333a <=( a16332a  and  a16327a );
 a16337a <=( (not A267)  and  A266 );
 a16338a <=( A265  and  a16337a );
 a16342a <=( A300  and  A299 );
 a16343a <=( (not A268)  and  a16342a );
 a16344a <=( a16343a  and  a16338a );
 a16348a <=( A166  and  (not A167) );
 a16349a <=( A170  and  a16348a );
 a16353a <=( (not A203)  and  (not A202) );
 a16354a <=( (not A201)  and  a16353a );
 a16355a <=( a16354a  and  a16349a );
 a16359a <=( (not A267)  and  A266 );
 a16360a <=( A265  and  a16359a );
 a16364a <=( A300  and  A298 );
 a16365a <=( (not A268)  and  a16364a );
 a16366a <=( a16365a  and  a16360a );
 a16370a <=( A166  and  (not A167) );
 a16371a <=( A170  and  a16370a );
 a16375a <=( (not A203)  and  (not A202) );
 a16376a <=( (not A201)  and  a16375a );
 a16377a <=( a16376a  and  a16371a );
 a16381a <=( (not A268)  and  (not A266) );
 a16382a <=( (not A265)  and  a16381a );
 a16386a <=( A302  and  (not A299) );
 a16387a <=( A298  and  a16386a );
 a16388a <=( a16387a  and  a16382a );
 a16392a <=( A166  and  (not A167) );
 a16393a <=( A170  and  a16392a );
 a16397a <=( (not A203)  and  (not A202) );
 a16398a <=( (not A201)  and  a16397a );
 a16399a <=( a16398a  and  a16393a );
 a16403a <=( (not A268)  and  (not A266) );
 a16404a <=( (not A265)  and  a16403a );
 a16408a <=( A302  and  A299 );
 a16409a <=( (not A298)  and  a16408a );
 a16410a <=( a16409a  and  a16404a );
 a16414a <=( A166  and  (not A167) );
 a16415a <=( A170  and  a16414a );
 a16419a <=( (not A265)  and  A201 );
 a16420a <=( A199  and  a16419a );
 a16421a <=( a16420a  and  a16415a );
 a16425a <=( A298  and  A269 );
 a16426a <=( A266  and  a16425a );
 a16430a <=( (not A301)  and  (not A300) );
 a16431a <=( A299  and  a16430a );
 a16432a <=( a16431a  and  a16426a );
 a16436a <=( A166  and  (not A167) );
 a16437a <=( A170  and  a16436a );
 a16441a <=( A265  and  A201 );
 a16442a <=( A199  and  a16441a );
 a16443a <=( a16442a  and  a16437a );
 a16447a <=( A298  and  A269 );
 a16448a <=( (not A266)  and  a16447a );
 a16452a <=( (not A301)  and  (not A300) );
 a16453a <=( A299  and  a16452a );
 a16454a <=( a16453a  and  a16448a );
 a16458a <=( A166  and  (not A167) );
 a16459a <=( A170  and  a16458a );
 a16463a <=( (not A265)  and  A201 );
 a16464a <=( A200  and  a16463a );
 a16465a <=( a16464a  and  a16459a );
 a16469a <=( A298  and  A269 );
 a16470a <=( A266  and  a16469a );
 a16474a <=( (not A301)  and  (not A300) );
 a16475a <=( A299  and  a16474a );
 a16476a <=( a16475a  and  a16470a );
 a16480a <=( A166  and  (not A167) );
 a16481a <=( A170  and  a16480a );
 a16485a <=( A265  and  A201 );
 a16486a <=( A200  and  a16485a );
 a16487a <=( a16486a  and  a16481a );
 a16491a <=( A298  and  A269 );
 a16492a <=( (not A266)  and  a16491a );
 a16496a <=( (not A301)  and  (not A300) );
 a16497a <=( A299  and  a16496a );
 a16498a <=( a16497a  and  a16492a );
 a16502a <=( A166  and  (not A167) );
 a16503a <=( A170  and  a16502a );
 a16507a <=( (not A201)  and  A200 );
 a16508a <=( A199  and  a16507a );
 a16509a <=( a16508a  and  a16503a );
 a16513a <=( (not A268)  and  (not A267) );
 a16514a <=( (not A202)  and  a16513a );
 a16518a <=( A300  and  A299 );
 a16519a <=( (not A269)  and  a16518a );
 a16520a <=( a16519a  and  a16514a );
 a16524a <=( A166  and  (not A167) );
 a16525a <=( A170  and  a16524a );
 a16529a <=( (not A201)  and  A200 );
 a16530a <=( A199  and  a16529a );
 a16531a <=( a16530a  and  a16525a );
 a16535a <=( (not A268)  and  (not A267) );
 a16536a <=( (not A202)  and  a16535a );
 a16540a <=( A300  and  A298 );
 a16541a <=( (not A269)  and  a16540a );
 a16542a <=( a16541a  and  a16536a );
 a16546a <=( A166  and  (not A167) );
 a16547a <=( A170  and  a16546a );
 a16551a <=( (not A201)  and  A200 );
 a16552a <=( A199  and  a16551a );
 a16553a <=( a16552a  and  a16547a );
 a16557a <=( A266  and  A265 );
 a16558a <=( (not A202)  and  a16557a );
 a16562a <=( A301  and  (not A268) );
 a16563a <=( (not A267)  and  a16562a );
 a16564a <=( a16563a  and  a16558a );
 a16568a <=( A166  and  (not A167) );
 a16569a <=( A170  and  a16568a );
 a16573a <=( (not A201)  and  A200 );
 a16574a <=( A199  and  a16573a );
 a16575a <=( a16574a  and  a16569a );
 a16579a <=( (not A266)  and  (not A265) );
 a16580a <=( (not A202)  and  a16579a );
 a16584a <=( A300  and  A299 );
 a16585a <=( (not A268)  and  a16584a );
 a16586a <=( a16585a  and  a16580a );
 a16590a <=( A166  and  (not A167) );
 a16591a <=( A170  and  a16590a );
 a16595a <=( (not A201)  and  A200 );
 a16596a <=( A199  and  a16595a );
 a16597a <=( a16596a  and  a16591a );
 a16601a <=( (not A266)  and  (not A265) );
 a16602a <=( (not A202)  and  a16601a );
 a16606a <=( A300  and  A298 );
 a16607a <=( (not A268)  and  a16606a );
 a16608a <=( a16607a  and  a16602a );
 a16612a <=( A166  and  (not A167) );
 a16613a <=( A170  and  a16612a );
 a16617a <=( A203  and  A200 );
 a16618a <=( (not A199)  and  a16617a );
 a16619a <=( a16618a  and  a16613a );
 a16623a <=( A298  and  A267 );
 a16624a <=( A265  and  a16623a );
 a16628a <=( (not A301)  and  (not A300) );
 a16629a <=( A299  and  a16628a );
 a16630a <=( a16629a  and  a16624a );
 a16634a <=( A166  and  (not A167) );
 a16635a <=( A170  and  a16634a );
 a16639a <=( A203  and  A200 );
 a16640a <=( (not A199)  and  a16639a );
 a16641a <=( a16640a  and  a16635a );
 a16645a <=( A298  and  A267 );
 a16646a <=( A266  and  a16645a );
 a16650a <=( (not A301)  and  (not A300) );
 a16651a <=( A299  and  a16650a );
 a16652a <=( a16651a  and  a16646a );
 a16656a <=( A166  and  (not A167) );
 a16657a <=( A170  and  a16656a );
 a16661a <=( A203  and  A200 );
 a16662a <=( (not A199)  and  a16661a );
 a16663a <=( a16662a  and  a16657a );
 a16667a <=( A269  and  A266 );
 a16668a <=( (not A265)  and  a16667a );
 a16672a <=( (not A302)  and  (not A301) );
 a16673a <=( (not A300)  and  a16672a );
 a16674a <=( a16673a  and  a16668a );
 a16678a <=( A166  and  (not A167) );
 a16679a <=( A170  and  a16678a );
 a16683a <=( A203  and  A200 );
 a16684a <=( (not A199)  and  a16683a );
 a16685a <=( a16684a  and  a16679a );
 a16689a <=( A269  and  A266 );
 a16690a <=( (not A265)  and  a16689a );
 a16694a <=( (not A301)  and  (not A299) );
 a16695a <=( (not A298)  and  a16694a );
 a16696a <=( a16695a  and  a16690a );
 a16700a <=( A166  and  (not A167) );
 a16701a <=( A170  and  a16700a );
 a16705a <=( A203  and  A200 );
 a16706a <=( (not A199)  and  a16705a );
 a16707a <=( a16706a  and  a16701a );
 a16711a <=( A269  and  (not A266) );
 a16712a <=( A265  and  a16711a );
 a16716a <=( (not A302)  and  (not A301) );
 a16717a <=( (not A300)  and  a16716a );
 a16718a <=( a16717a  and  a16712a );
 a16722a <=( A166  and  (not A167) );
 a16723a <=( A170  and  a16722a );
 a16727a <=( A203  and  A200 );
 a16728a <=( (not A199)  and  a16727a );
 a16729a <=( a16728a  and  a16723a );
 a16733a <=( A269  and  (not A266) );
 a16734a <=( A265  and  a16733a );
 a16738a <=( (not A301)  and  (not A299) );
 a16739a <=( (not A298)  and  a16738a );
 a16740a <=( a16739a  and  a16734a );
 a16744a <=( A166  and  (not A167) );
 a16745a <=( A170  and  a16744a );
 a16749a <=( A203  and  (not A200) );
 a16750a <=( A199  and  a16749a );
 a16751a <=( a16750a  and  a16745a );
 a16755a <=( A298  and  A267 );
 a16756a <=( A265  and  a16755a );
 a16760a <=( (not A301)  and  (not A300) );
 a16761a <=( A299  and  a16760a );
 a16762a <=( a16761a  and  a16756a );
 a16766a <=( A166  and  (not A167) );
 a16767a <=( A170  and  a16766a );
 a16771a <=( A203  and  (not A200) );
 a16772a <=( A199  and  a16771a );
 a16773a <=( a16772a  and  a16767a );
 a16777a <=( A298  and  A267 );
 a16778a <=( A266  and  a16777a );
 a16782a <=( (not A301)  and  (not A300) );
 a16783a <=( A299  and  a16782a );
 a16784a <=( a16783a  and  a16778a );
 a16788a <=( A166  and  (not A167) );
 a16789a <=( A170  and  a16788a );
 a16793a <=( A203  and  (not A200) );
 a16794a <=( A199  and  a16793a );
 a16795a <=( a16794a  and  a16789a );
 a16799a <=( A269  and  A266 );
 a16800a <=( (not A265)  and  a16799a );
 a16804a <=( (not A302)  and  (not A301) );
 a16805a <=( (not A300)  and  a16804a );
 a16806a <=( a16805a  and  a16800a );
 a16810a <=( A166  and  (not A167) );
 a16811a <=( A170  and  a16810a );
 a16815a <=( A203  and  (not A200) );
 a16816a <=( A199  and  a16815a );
 a16817a <=( a16816a  and  a16811a );
 a16821a <=( A269  and  A266 );
 a16822a <=( (not A265)  and  a16821a );
 a16826a <=( (not A301)  and  (not A299) );
 a16827a <=( (not A298)  and  a16826a );
 a16828a <=( a16827a  and  a16822a );
 a16832a <=( A166  and  (not A167) );
 a16833a <=( A170  and  a16832a );
 a16837a <=( A203  and  (not A200) );
 a16838a <=( A199  and  a16837a );
 a16839a <=( a16838a  and  a16833a );
 a16843a <=( A269  and  (not A266) );
 a16844a <=( A265  and  a16843a );
 a16848a <=( (not A302)  and  (not A301) );
 a16849a <=( (not A300)  and  a16848a );
 a16850a <=( a16849a  and  a16844a );
 a16854a <=( A166  and  (not A167) );
 a16855a <=( A170  and  a16854a );
 a16859a <=( A203  and  (not A200) );
 a16860a <=( A199  and  a16859a );
 a16861a <=( a16860a  and  a16855a );
 a16865a <=( A269  and  (not A266) );
 a16866a <=( A265  and  a16865a );
 a16870a <=( (not A301)  and  (not A299) );
 a16871a <=( (not A298)  and  a16870a );
 a16872a <=( a16871a  and  a16866a );
 a16876a <=( A166  and  (not A167) );
 a16877a <=( A170  and  a16876a );
 a16881a <=( (not A202)  and  (not A200) );
 a16882a <=( (not A199)  and  a16881a );
 a16883a <=( a16882a  and  a16877a );
 a16887a <=( (not A269)  and  (not A268) );
 a16888a <=( (not A267)  and  a16887a );
 a16892a <=( A302  and  (not A299) );
 a16893a <=( A298  and  a16892a );
 a16894a <=( a16893a  and  a16888a );
 a16898a <=( A166  and  (not A167) );
 a16899a <=( A170  and  a16898a );
 a16903a <=( (not A202)  and  (not A200) );
 a16904a <=( (not A199)  and  a16903a );
 a16905a <=( a16904a  and  a16899a );
 a16909a <=( (not A269)  and  (not A268) );
 a16910a <=( (not A267)  and  a16909a );
 a16914a <=( A302  and  A299 );
 a16915a <=( (not A298)  and  a16914a );
 a16916a <=( a16915a  and  a16910a );
 a16920a <=( A166  and  (not A167) );
 a16921a <=( A170  and  a16920a );
 a16925a <=( (not A202)  and  (not A200) );
 a16926a <=( (not A199)  and  a16925a );
 a16927a <=( a16926a  and  a16921a );
 a16931a <=( (not A267)  and  A266 );
 a16932a <=( A265  and  a16931a );
 a16936a <=( A300  and  A299 );
 a16937a <=( (not A268)  and  a16936a );
 a16938a <=( a16937a  and  a16932a );
 a16942a <=( A166  and  (not A167) );
 a16943a <=( A170  and  a16942a );
 a16947a <=( (not A202)  and  (not A200) );
 a16948a <=( (not A199)  and  a16947a );
 a16949a <=( a16948a  and  a16943a );
 a16953a <=( (not A267)  and  A266 );
 a16954a <=( A265  and  a16953a );
 a16958a <=( A300  and  A298 );
 a16959a <=( (not A268)  and  a16958a );
 a16960a <=( a16959a  and  a16954a );
 a16964a <=( A166  and  (not A167) );
 a16965a <=( A170  and  a16964a );
 a16969a <=( (not A202)  and  (not A200) );
 a16970a <=( (not A199)  and  a16969a );
 a16971a <=( a16970a  and  a16965a );
 a16975a <=( (not A268)  and  (not A266) );
 a16976a <=( (not A265)  and  a16975a );
 a16980a <=( A302  and  (not A299) );
 a16981a <=( A298  and  a16980a );
 a16982a <=( a16981a  and  a16976a );
 a16986a <=( A166  and  (not A167) );
 a16987a <=( A170  and  a16986a );
 a16991a <=( (not A202)  and  (not A200) );
 a16992a <=( (not A199)  and  a16991a );
 a16993a <=( a16992a  and  a16987a );
 a16997a <=( (not A268)  and  (not A266) );
 a16998a <=( (not A265)  and  a16997a );
 a17002a <=( A302  and  A299 );
 a17003a <=( (not A298)  and  a17002a );
 a17004a <=( a17003a  and  a16998a );
 a17008a <=( A200  and  A199 );
 a17009a <=( A169  and  a17008a );
 a17013a <=( A265  and  (not A202) );
 a17014a <=( (not A201)  and  a17013a );
 a17015a <=( a17014a  and  a17009a );
 a17019a <=( (not A268)  and  (not A267) );
 a17020a <=( A266  and  a17019a );
 a17024a <=( A302  and  (not A299) );
 a17025a <=( A298  and  a17024a );
 a17026a <=( a17025a  and  a17020a );
 a17030a <=( A200  and  A199 );
 a17031a <=( A169  and  a17030a );
 a17035a <=( A265  and  (not A202) );
 a17036a <=( (not A201)  and  a17035a );
 a17037a <=( a17036a  and  a17031a );
 a17041a <=( (not A268)  and  (not A267) );
 a17042a <=( A266  and  a17041a );
 a17046a <=( A302  and  A299 );
 a17047a <=( (not A298)  and  a17046a );
 a17048a <=( a17047a  and  a17042a );
 a17052a <=( (not A166)  and  (not A167) );
 a17053a <=( (not A169)  and  a17052a );
 a17057a <=( (not A203)  and  (not A202) );
 a17058a <=( (not A201)  and  a17057a );
 a17059a <=( a17058a  and  a17053a );
 a17063a <=( A298  and  A267 );
 a17064a <=( A265  and  a17063a );
 a17068a <=( (not A301)  and  (not A300) );
 a17069a <=( A299  and  a17068a );
 a17070a <=( a17069a  and  a17064a );
 a17074a <=( (not A166)  and  (not A167) );
 a17075a <=( (not A169)  and  a17074a );
 a17079a <=( (not A203)  and  (not A202) );
 a17080a <=( (not A201)  and  a17079a );
 a17081a <=( a17080a  and  a17075a );
 a17085a <=( A298  and  A267 );
 a17086a <=( A266  and  a17085a );
 a17090a <=( (not A301)  and  (not A300) );
 a17091a <=( A299  and  a17090a );
 a17092a <=( a17091a  and  a17086a );
 a17096a <=( (not A166)  and  (not A167) );
 a17097a <=( (not A169)  and  a17096a );
 a17101a <=( (not A203)  and  (not A202) );
 a17102a <=( (not A201)  and  a17101a );
 a17103a <=( a17102a  and  a17097a );
 a17107a <=( A269  and  A266 );
 a17108a <=( (not A265)  and  a17107a );
 a17112a <=( (not A302)  and  (not A301) );
 a17113a <=( (not A300)  and  a17112a );
 a17114a <=( a17113a  and  a17108a );
 a17118a <=( (not A166)  and  (not A167) );
 a17119a <=( (not A169)  and  a17118a );
 a17123a <=( (not A203)  and  (not A202) );
 a17124a <=( (not A201)  and  a17123a );
 a17125a <=( a17124a  and  a17119a );
 a17129a <=( A269  and  A266 );
 a17130a <=( (not A265)  and  a17129a );
 a17134a <=( (not A301)  and  (not A299) );
 a17135a <=( (not A298)  and  a17134a );
 a17136a <=( a17135a  and  a17130a );
 a17140a <=( (not A166)  and  (not A167) );
 a17141a <=( (not A169)  and  a17140a );
 a17145a <=( (not A203)  and  (not A202) );
 a17146a <=( (not A201)  and  a17145a );
 a17147a <=( a17146a  and  a17141a );
 a17151a <=( A269  and  (not A266) );
 a17152a <=( A265  and  a17151a );
 a17156a <=( (not A302)  and  (not A301) );
 a17157a <=( (not A300)  and  a17156a );
 a17158a <=( a17157a  and  a17152a );
 a17162a <=( (not A166)  and  (not A167) );
 a17163a <=( (not A169)  and  a17162a );
 a17167a <=( (not A203)  and  (not A202) );
 a17168a <=( (not A201)  and  a17167a );
 a17169a <=( a17168a  and  a17163a );
 a17173a <=( A269  and  (not A266) );
 a17174a <=( A265  and  a17173a );
 a17178a <=( (not A301)  and  (not A299) );
 a17179a <=( (not A298)  and  a17178a );
 a17180a <=( a17179a  and  a17174a );
 a17184a <=( (not A166)  and  (not A167) );
 a17185a <=( (not A169)  and  a17184a );
 a17189a <=( A265  and  A201 );
 a17190a <=( A199  and  a17189a );
 a17191a <=( a17190a  and  a17185a );
 a17195a <=( (not A268)  and  (not A267) );
 a17196a <=( A266  and  a17195a );
 a17200a <=( A302  and  (not A299) );
 a17201a <=( A298  and  a17200a );
 a17202a <=( a17201a  and  a17196a );
 a17206a <=( (not A166)  and  (not A167) );
 a17207a <=( (not A169)  and  a17206a );
 a17211a <=( A265  and  A201 );
 a17212a <=( A199  and  a17211a );
 a17213a <=( a17212a  and  a17207a );
 a17217a <=( (not A268)  and  (not A267) );
 a17218a <=( A266  and  a17217a );
 a17222a <=( A302  and  A299 );
 a17223a <=( (not A298)  and  a17222a );
 a17224a <=( a17223a  and  a17218a );
 a17228a <=( (not A166)  and  (not A167) );
 a17229a <=( (not A169)  and  a17228a );
 a17233a <=( A265  and  A201 );
 a17234a <=( A200  and  a17233a );
 a17235a <=( a17234a  and  a17229a );
 a17239a <=( (not A268)  and  (not A267) );
 a17240a <=( A266  and  a17239a );
 a17244a <=( A302  and  (not A299) );
 a17245a <=( A298  and  a17244a );
 a17246a <=( a17245a  and  a17240a );
 a17250a <=( (not A166)  and  (not A167) );
 a17251a <=( (not A169)  and  a17250a );
 a17255a <=( A265  and  A201 );
 a17256a <=( A200  and  a17255a );
 a17257a <=( a17256a  and  a17251a );
 a17261a <=( (not A268)  and  (not A267) );
 a17262a <=( A266  and  a17261a );
 a17266a <=( A302  and  A299 );
 a17267a <=( (not A298)  and  a17266a );
 a17268a <=( a17267a  and  a17262a );
 a17272a <=( (not A166)  and  (not A167) );
 a17273a <=( (not A169)  and  a17272a );
 a17277a <=( (not A201)  and  A200 );
 a17278a <=( A199  and  a17277a );
 a17279a <=( a17278a  and  a17273a );
 a17283a <=( A298  and  A268 );
 a17284a <=( (not A202)  and  a17283a );
 a17288a <=( (not A301)  and  (not A300) );
 a17289a <=( A299  and  a17288a );
 a17290a <=( a17289a  and  a17284a );
 a17294a <=( (not A166)  and  (not A167) );
 a17295a <=( (not A169)  and  a17294a );
 a17299a <=( (not A201)  and  A200 );
 a17300a <=( A199  and  a17299a );
 a17301a <=( a17300a  and  a17295a );
 a17305a <=( A267  and  A265 );
 a17306a <=( (not A202)  and  a17305a );
 a17310a <=( (not A302)  and  (not A301) );
 a17311a <=( (not A300)  and  a17310a );
 a17312a <=( a17311a  and  a17306a );
 a17316a <=( (not A166)  and  (not A167) );
 a17317a <=( (not A169)  and  a17316a );
 a17321a <=( (not A201)  and  A200 );
 a17322a <=( A199  and  a17321a );
 a17323a <=( a17322a  and  a17317a );
 a17327a <=( A267  and  A265 );
 a17328a <=( (not A202)  and  a17327a );
 a17332a <=( (not A301)  and  (not A299) );
 a17333a <=( (not A298)  and  a17332a );
 a17334a <=( a17333a  and  a17328a );
 a17338a <=( (not A166)  and  (not A167) );
 a17339a <=( (not A169)  and  a17338a );
 a17343a <=( (not A201)  and  A200 );
 a17344a <=( A199  and  a17343a );
 a17345a <=( a17344a  and  a17339a );
 a17349a <=( A267  and  A266 );
 a17350a <=( (not A202)  and  a17349a );
 a17354a <=( (not A302)  and  (not A301) );
 a17355a <=( (not A300)  and  a17354a );
 a17356a <=( a17355a  and  a17350a );
 a17360a <=( (not A166)  and  (not A167) );
 a17361a <=( (not A169)  and  a17360a );
 a17365a <=( (not A201)  and  A200 );
 a17366a <=( A199  and  a17365a );
 a17367a <=( a17366a  and  a17361a );
 a17371a <=( A267  and  A266 );
 a17372a <=( (not A202)  and  a17371a );
 a17376a <=( (not A301)  and  (not A299) );
 a17377a <=( (not A298)  and  a17376a );
 a17378a <=( a17377a  and  a17372a );
 a17382a <=( (not A166)  and  (not A167) );
 a17383a <=( (not A169)  and  a17382a );
 a17387a <=( A203  and  A200 );
 a17388a <=( (not A199)  and  a17387a );
 a17389a <=( a17388a  and  a17383a );
 a17393a <=( (not A269)  and  (not A268) );
 a17394a <=( (not A267)  and  a17393a );
 a17398a <=( A302  and  (not A299) );
 a17399a <=( A298  and  a17398a );
 a17400a <=( a17399a  and  a17394a );
 a17404a <=( (not A166)  and  (not A167) );
 a17405a <=( (not A169)  and  a17404a );
 a17409a <=( A203  and  A200 );
 a17410a <=( (not A199)  and  a17409a );
 a17411a <=( a17410a  and  a17405a );
 a17415a <=( (not A269)  and  (not A268) );
 a17416a <=( (not A267)  and  a17415a );
 a17420a <=( A302  and  A299 );
 a17421a <=( (not A298)  and  a17420a );
 a17422a <=( a17421a  and  a17416a );
 a17426a <=( (not A166)  and  (not A167) );
 a17427a <=( (not A169)  and  a17426a );
 a17431a <=( A203  and  A200 );
 a17432a <=( (not A199)  and  a17431a );
 a17433a <=( a17432a  and  a17427a );
 a17437a <=( (not A267)  and  A266 );
 a17438a <=( A265  and  a17437a );
 a17442a <=( A300  and  A299 );
 a17443a <=( (not A268)  and  a17442a );
 a17444a <=( a17443a  and  a17438a );
 a17448a <=( (not A166)  and  (not A167) );
 a17449a <=( (not A169)  and  a17448a );
 a17453a <=( A203  and  A200 );
 a17454a <=( (not A199)  and  a17453a );
 a17455a <=( a17454a  and  a17449a );
 a17459a <=( (not A267)  and  A266 );
 a17460a <=( A265  and  a17459a );
 a17464a <=( A300  and  A298 );
 a17465a <=( (not A268)  and  a17464a );
 a17466a <=( a17465a  and  a17460a );
 a17470a <=( (not A166)  and  (not A167) );
 a17471a <=( (not A169)  and  a17470a );
 a17475a <=( A203  and  A200 );
 a17476a <=( (not A199)  and  a17475a );
 a17477a <=( a17476a  and  a17471a );
 a17481a <=( (not A268)  and  (not A266) );
 a17482a <=( (not A265)  and  a17481a );
 a17486a <=( A302  and  (not A299) );
 a17487a <=( A298  and  a17486a );
 a17488a <=( a17487a  and  a17482a );
 a17492a <=( (not A166)  and  (not A167) );
 a17493a <=( (not A169)  and  a17492a );
 a17497a <=( A203  and  A200 );
 a17498a <=( (not A199)  and  a17497a );
 a17499a <=( a17498a  and  a17493a );
 a17503a <=( (not A268)  and  (not A266) );
 a17504a <=( (not A265)  and  a17503a );
 a17508a <=( A302  and  A299 );
 a17509a <=( (not A298)  and  a17508a );
 a17510a <=( a17509a  and  a17504a );
 a17514a <=( (not A166)  and  (not A167) );
 a17515a <=( (not A169)  and  a17514a );
 a17519a <=( A203  and  (not A200) );
 a17520a <=( A199  and  a17519a );
 a17521a <=( a17520a  and  a17515a );
 a17525a <=( (not A269)  and  (not A268) );
 a17526a <=( (not A267)  and  a17525a );
 a17530a <=( A302  and  (not A299) );
 a17531a <=( A298  and  a17530a );
 a17532a <=( a17531a  and  a17526a );
 a17536a <=( (not A166)  and  (not A167) );
 a17537a <=( (not A169)  and  a17536a );
 a17541a <=( A203  and  (not A200) );
 a17542a <=( A199  and  a17541a );
 a17543a <=( a17542a  and  a17537a );
 a17547a <=( (not A269)  and  (not A268) );
 a17548a <=( (not A267)  and  a17547a );
 a17552a <=( A302  and  A299 );
 a17553a <=( (not A298)  and  a17552a );
 a17554a <=( a17553a  and  a17548a );
 a17558a <=( (not A166)  and  (not A167) );
 a17559a <=( (not A169)  and  a17558a );
 a17563a <=( A203  and  (not A200) );
 a17564a <=( A199  and  a17563a );
 a17565a <=( a17564a  and  a17559a );
 a17569a <=( (not A267)  and  A266 );
 a17570a <=( A265  and  a17569a );
 a17574a <=( A300  and  A299 );
 a17575a <=( (not A268)  and  a17574a );
 a17576a <=( a17575a  and  a17570a );
 a17580a <=( (not A166)  and  (not A167) );
 a17581a <=( (not A169)  and  a17580a );
 a17585a <=( A203  and  (not A200) );
 a17586a <=( A199  and  a17585a );
 a17587a <=( a17586a  and  a17581a );
 a17591a <=( (not A267)  and  A266 );
 a17592a <=( A265  and  a17591a );
 a17596a <=( A300  and  A298 );
 a17597a <=( (not A268)  and  a17596a );
 a17598a <=( a17597a  and  a17592a );
 a17602a <=( (not A166)  and  (not A167) );
 a17603a <=( (not A169)  and  a17602a );
 a17607a <=( A203  and  (not A200) );
 a17608a <=( A199  and  a17607a );
 a17609a <=( a17608a  and  a17603a );
 a17613a <=( (not A268)  and  (not A266) );
 a17614a <=( (not A265)  and  a17613a );
 a17618a <=( A302  and  (not A299) );
 a17619a <=( A298  and  a17618a );
 a17620a <=( a17619a  and  a17614a );
 a17624a <=( (not A166)  and  (not A167) );
 a17625a <=( (not A169)  and  a17624a );
 a17629a <=( A203  and  (not A200) );
 a17630a <=( A199  and  a17629a );
 a17631a <=( a17630a  and  a17625a );
 a17635a <=( (not A268)  and  (not A266) );
 a17636a <=( (not A265)  and  a17635a );
 a17640a <=( A302  and  A299 );
 a17641a <=( (not A298)  and  a17640a );
 a17642a <=( a17641a  and  a17636a );
 a17646a <=( (not A166)  and  (not A167) );
 a17647a <=( (not A169)  and  a17646a );
 a17651a <=( (not A202)  and  (not A200) );
 a17652a <=( (not A199)  and  a17651a );
 a17653a <=( a17652a  and  a17647a );
 a17657a <=( A298  and  A267 );
 a17658a <=( A265  and  a17657a );
 a17662a <=( (not A301)  and  (not A300) );
 a17663a <=( A299  and  a17662a );
 a17664a <=( a17663a  and  a17658a );
 a17668a <=( (not A166)  and  (not A167) );
 a17669a <=( (not A169)  and  a17668a );
 a17673a <=( (not A202)  and  (not A200) );
 a17674a <=( (not A199)  and  a17673a );
 a17675a <=( a17674a  and  a17669a );
 a17679a <=( A298  and  A267 );
 a17680a <=( A266  and  a17679a );
 a17684a <=( (not A301)  and  (not A300) );
 a17685a <=( A299  and  a17684a );
 a17686a <=( a17685a  and  a17680a );
 a17690a <=( (not A166)  and  (not A167) );
 a17691a <=( (not A169)  and  a17690a );
 a17695a <=( (not A202)  and  (not A200) );
 a17696a <=( (not A199)  and  a17695a );
 a17697a <=( a17696a  and  a17691a );
 a17701a <=( A269  and  A266 );
 a17702a <=( (not A265)  and  a17701a );
 a17706a <=( (not A302)  and  (not A301) );
 a17707a <=( (not A300)  and  a17706a );
 a17708a <=( a17707a  and  a17702a );
 a17712a <=( (not A166)  and  (not A167) );
 a17713a <=( (not A169)  and  a17712a );
 a17717a <=( (not A202)  and  (not A200) );
 a17718a <=( (not A199)  and  a17717a );
 a17719a <=( a17718a  and  a17713a );
 a17723a <=( A269  and  A266 );
 a17724a <=( (not A265)  and  a17723a );
 a17728a <=( (not A301)  and  (not A299) );
 a17729a <=( (not A298)  and  a17728a );
 a17730a <=( a17729a  and  a17724a );
 a17734a <=( (not A166)  and  (not A167) );
 a17735a <=( (not A169)  and  a17734a );
 a17739a <=( (not A202)  and  (not A200) );
 a17740a <=( (not A199)  and  a17739a );
 a17741a <=( a17740a  and  a17735a );
 a17745a <=( A269  and  (not A266) );
 a17746a <=( A265  and  a17745a );
 a17750a <=( (not A302)  and  (not A301) );
 a17751a <=( (not A300)  and  a17750a );
 a17752a <=( a17751a  and  a17746a );
 a17756a <=( (not A166)  and  (not A167) );
 a17757a <=( (not A169)  and  a17756a );
 a17761a <=( (not A202)  and  (not A200) );
 a17762a <=( (not A199)  and  a17761a );
 a17763a <=( a17762a  and  a17757a );
 a17767a <=( A269  and  (not A266) );
 a17768a <=( A265  and  a17767a );
 a17772a <=( (not A301)  and  (not A299) );
 a17773a <=( (not A298)  and  a17772a );
 a17774a <=( a17773a  and  a17768a );
 a17778a <=( A167  and  (not A168) );
 a17779a <=( (not A169)  and  a17778a );
 a17783a <=( A265  and  A202 );
 a17784a <=( A166  and  a17783a );
 a17785a <=( a17784a  and  a17779a );
 a17789a <=( (not A268)  and  (not A267) );
 a17790a <=( A266  and  a17789a );
 a17794a <=( A302  and  (not A299) );
 a17795a <=( A298  and  a17794a );
 a17796a <=( a17795a  and  a17790a );
 a17800a <=( A167  and  (not A168) );
 a17801a <=( (not A169)  and  a17800a );
 a17805a <=( A265  and  A202 );
 a17806a <=( A166  and  a17805a );
 a17807a <=( a17806a  and  a17801a );
 a17811a <=( (not A268)  and  (not A267) );
 a17812a <=( A266  and  a17811a );
 a17816a <=( A302  and  A299 );
 a17817a <=( (not A298)  and  a17816a );
 a17818a <=( a17817a  and  a17812a );
 a17822a <=( A167  and  (not A168) );
 a17823a <=( (not A169)  and  a17822a );
 a17827a <=( (not A202)  and  (not A201) );
 a17828a <=( A166  and  a17827a );
 a17829a <=( a17828a  and  a17823a );
 a17833a <=( A298  and  A268 );
 a17834a <=( (not A203)  and  a17833a );
 a17838a <=( (not A301)  and  (not A300) );
 a17839a <=( A299  and  a17838a );
 a17840a <=( a17839a  and  a17834a );
 a17844a <=( A167  and  (not A168) );
 a17845a <=( (not A169)  and  a17844a );
 a17849a <=( (not A202)  and  (not A201) );
 a17850a <=( A166  and  a17849a );
 a17851a <=( a17850a  and  a17845a );
 a17855a <=( A267  and  A265 );
 a17856a <=( (not A203)  and  a17855a );
 a17860a <=( (not A302)  and  (not A301) );
 a17861a <=( (not A300)  and  a17860a );
 a17862a <=( a17861a  and  a17856a );
 a17866a <=( A167  and  (not A168) );
 a17867a <=( (not A169)  and  a17866a );
 a17871a <=( (not A202)  and  (not A201) );
 a17872a <=( A166  and  a17871a );
 a17873a <=( a17872a  and  a17867a );
 a17877a <=( A267  and  A265 );
 a17878a <=( (not A203)  and  a17877a );
 a17882a <=( (not A301)  and  (not A299) );
 a17883a <=( (not A298)  and  a17882a );
 a17884a <=( a17883a  and  a17878a );
 a17888a <=( A167  and  (not A168) );
 a17889a <=( (not A169)  and  a17888a );
 a17893a <=( (not A202)  and  (not A201) );
 a17894a <=( A166  and  a17893a );
 a17895a <=( a17894a  and  a17889a );
 a17899a <=( A267  and  A266 );
 a17900a <=( (not A203)  and  a17899a );
 a17904a <=( (not A302)  and  (not A301) );
 a17905a <=( (not A300)  and  a17904a );
 a17906a <=( a17905a  and  a17900a );
 a17910a <=( A167  and  (not A168) );
 a17911a <=( (not A169)  and  a17910a );
 a17915a <=( (not A202)  and  (not A201) );
 a17916a <=( A166  and  a17915a );
 a17917a <=( a17916a  and  a17911a );
 a17921a <=( A267  and  A266 );
 a17922a <=( (not A203)  and  a17921a );
 a17926a <=( (not A301)  and  (not A299) );
 a17927a <=( (not A298)  and  a17926a );
 a17928a <=( a17927a  and  a17922a );
 a17932a <=( A167  and  (not A168) );
 a17933a <=( (not A169)  and  a17932a );
 a17937a <=( A201  and  A199 );
 a17938a <=( A166  and  a17937a );
 a17939a <=( a17938a  and  a17933a );
 a17943a <=( (not A269)  and  (not A268) );
 a17944a <=( (not A267)  and  a17943a );
 a17948a <=( A302  and  (not A299) );
 a17949a <=( A298  and  a17948a );
 a17950a <=( a17949a  and  a17944a );
 a17954a <=( A167  and  (not A168) );
 a17955a <=( (not A169)  and  a17954a );
 a17959a <=( A201  and  A199 );
 a17960a <=( A166  and  a17959a );
 a17961a <=( a17960a  and  a17955a );
 a17965a <=( (not A269)  and  (not A268) );
 a17966a <=( (not A267)  and  a17965a );
 a17970a <=( A302  and  A299 );
 a17971a <=( (not A298)  and  a17970a );
 a17972a <=( a17971a  and  a17966a );
 a17976a <=( A167  and  (not A168) );
 a17977a <=( (not A169)  and  a17976a );
 a17981a <=( A201  and  A199 );
 a17982a <=( A166  and  a17981a );
 a17983a <=( a17982a  and  a17977a );
 a17987a <=( (not A267)  and  A266 );
 a17988a <=( A265  and  a17987a );
 a17992a <=( A300  and  A299 );
 a17993a <=( (not A268)  and  a17992a );
 a17994a <=( a17993a  and  a17988a );
 a17998a <=( A167  and  (not A168) );
 a17999a <=( (not A169)  and  a17998a );
 a18003a <=( A201  and  A199 );
 a18004a <=( A166  and  a18003a );
 a18005a <=( a18004a  and  a17999a );
 a18009a <=( (not A267)  and  A266 );
 a18010a <=( A265  and  a18009a );
 a18014a <=( A300  and  A298 );
 a18015a <=( (not A268)  and  a18014a );
 a18016a <=( a18015a  and  a18010a );
 a18020a <=( A167  and  (not A168) );
 a18021a <=( (not A169)  and  a18020a );
 a18025a <=( A201  and  A199 );
 a18026a <=( A166  and  a18025a );
 a18027a <=( a18026a  and  a18021a );
 a18031a <=( (not A268)  and  (not A266) );
 a18032a <=( (not A265)  and  a18031a );
 a18036a <=( A302  and  (not A299) );
 a18037a <=( A298  and  a18036a );
 a18038a <=( a18037a  and  a18032a );
 a18042a <=( A167  and  (not A168) );
 a18043a <=( (not A169)  and  a18042a );
 a18047a <=( A201  and  A199 );
 a18048a <=( A166  and  a18047a );
 a18049a <=( a18048a  and  a18043a );
 a18053a <=( (not A268)  and  (not A266) );
 a18054a <=( (not A265)  and  a18053a );
 a18058a <=( A302  and  A299 );
 a18059a <=( (not A298)  and  a18058a );
 a18060a <=( a18059a  and  a18054a );
 a18064a <=( A167  and  (not A168) );
 a18065a <=( (not A169)  and  a18064a );
 a18069a <=( A201  and  A200 );
 a18070a <=( A166  and  a18069a );
 a18071a <=( a18070a  and  a18065a );
 a18075a <=( (not A269)  and  (not A268) );
 a18076a <=( (not A267)  and  a18075a );
 a18080a <=( A302  and  (not A299) );
 a18081a <=( A298  and  a18080a );
 a18082a <=( a18081a  and  a18076a );
 a18086a <=( A167  and  (not A168) );
 a18087a <=( (not A169)  and  a18086a );
 a18091a <=( A201  and  A200 );
 a18092a <=( A166  and  a18091a );
 a18093a <=( a18092a  and  a18087a );
 a18097a <=( (not A269)  and  (not A268) );
 a18098a <=( (not A267)  and  a18097a );
 a18102a <=( A302  and  A299 );
 a18103a <=( (not A298)  and  a18102a );
 a18104a <=( a18103a  and  a18098a );
 a18108a <=( A167  and  (not A168) );
 a18109a <=( (not A169)  and  a18108a );
 a18113a <=( A201  and  A200 );
 a18114a <=( A166  and  a18113a );
 a18115a <=( a18114a  and  a18109a );
 a18119a <=( (not A267)  and  A266 );
 a18120a <=( A265  and  a18119a );
 a18124a <=( A300  and  A299 );
 a18125a <=( (not A268)  and  a18124a );
 a18126a <=( a18125a  and  a18120a );
 a18130a <=( A167  and  (not A168) );
 a18131a <=( (not A169)  and  a18130a );
 a18135a <=( A201  and  A200 );
 a18136a <=( A166  and  a18135a );
 a18137a <=( a18136a  and  a18131a );
 a18141a <=( (not A267)  and  A266 );
 a18142a <=( A265  and  a18141a );
 a18146a <=( A300  and  A298 );
 a18147a <=( (not A268)  and  a18146a );
 a18148a <=( a18147a  and  a18142a );
 a18152a <=( A167  and  (not A168) );
 a18153a <=( (not A169)  and  a18152a );
 a18157a <=( A201  and  A200 );
 a18158a <=( A166  and  a18157a );
 a18159a <=( a18158a  and  a18153a );
 a18163a <=( (not A268)  and  (not A266) );
 a18164a <=( (not A265)  and  a18163a );
 a18168a <=( A302  and  (not A299) );
 a18169a <=( A298  and  a18168a );
 a18170a <=( a18169a  and  a18164a );
 a18174a <=( A167  and  (not A168) );
 a18175a <=( (not A169)  and  a18174a );
 a18179a <=( A201  and  A200 );
 a18180a <=( A166  and  a18179a );
 a18181a <=( a18180a  and  a18175a );
 a18185a <=( (not A268)  and  (not A266) );
 a18186a <=( (not A265)  and  a18185a );
 a18190a <=( A302  and  A299 );
 a18191a <=( (not A298)  and  a18190a );
 a18192a <=( a18191a  and  a18186a );
 a18196a <=( A167  and  (not A168) );
 a18197a <=( (not A169)  and  a18196a );
 a18201a <=( A200  and  A199 );
 a18202a <=( A166  and  a18201a );
 a18203a <=( a18202a  and  a18197a );
 a18207a <=( A268  and  (not A202) );
 a18208a <=( (not A201)  and  a18207a );
 a18212a <=( (not A302)  and  (not A301) );
 a18213a <=( (not A300)  and  a18212a );
 a18214a <=( a18213a  and  a18208a );
 a18218a <=( A167  and  (not A168) );
 a18219a <=( (not A169)  and  a18218a );
 a18223a <=( A200  and  A199 );
 a18224a <=( A166  and  a18223a );
 a18225a <=( a18224a  and  a18219a );
 a18229a <=( A268  and  (not A202) );
 a18230a <=( (not A201)  and  a18229a );
 a18234a <=( (not A301)  and  (not A299) );
 a18235a <=( (not A298)  and  a18234a );
 a18236a <=( a18235a  and  a18230a );
 a18240a <=( A167  and  (not A168) );
 a18241a <=( (not A169)  and  a18240a );
 a18245a <=( A200  and  (not A199) );
 a18246a <=( A166  and  a18245a );
 a18247a <=( a18246a  and  a18241a );
 a18251a <=( (not A268)  and  (not A267) );
 a18252a <=( A203  and  a18251a );
 a18256a <=( A300  and  A299 );
 a18257a <=( (not A269)  and  a18256a );
 a18258a <=( a18257a  and  a18252a );
 a18262a <=( A167  and  (not A168) );
 a18263a <=( (not A169)  and  a18262a );
 a18267a <=( A200  and  (not A199) );
 a18268a <=( A166  and  a18267a );
 a18269a <=( a18268a  and  a18263a );
 a18273a <=( (not A268)  and  (not A267) );
 a18274a <=( A203  and  a18273a );
 a18278a <=( A300  and  A298 );
 a18279a <=( (not A269)  and  a18278a );
 a18280a <=( a18279a  and  a18274a );
 a18284a <=( A167  and  (not A168) );
 a18285a <=( (not A169)  and  a18284a );
 a18289a <=( A200  and  (not A199) );
 a18290a <=( A166  and  a18289a );
 a18291a <=( a18290a  and  a18285a );
 a18295a <=( A266  and  A265 );
 a18296a <=( A203  and  a18295a );
 a18300a <=( A301  and  (not A268) );
 a18301a <=( (not A267)  and  a18300a );
 a18302a <=( a18301a  and  a18296a );
 a18306a <=( A167  and  (not A168) );
 a18307a <=( (not A169)  and  a18306a );
 a18311a <=( A200  and  (not A199) );
 a18312a <=( A166  and  a18311a );
 a18313a <=( a18312a  and  a18307a );
 a18317a <=( (not A266)  and  (not A265) );
 a18318a <=( A203  and  a18317a );
 a18322a <=( A300  and  A299 );
 a18323a <=( (not A268)  and  a18322a );
 a18324a <=( a18323a  and  a18318a );
 a18328a <=( A167  and  (not A168) );
 a18329a <=( (not A169)  and  a18328a );
 a18333a <=( A200  and  (not A199) );
 a18334a <=( A166  and  a18333a );
 a18335a <=( a18334a  and  a18329a );
 a18339a <=( (not A266)  and  (not A265) );
 a18340a <=( A203  and  a18339a );
 a18344a <=( A300  and  A298 );
 a18345a <=( (not A268)  and  a18344a );
 a18346a <=( a18345a  and  a18340a );
 a18350a <=( A167  and  (not A168) );
 a18351a <=( (not A169)  and  a18350a );
 a18355a <=( (not A200)  and  A199 );
 a18356a <=( A166  and  a18355a );
 a18357a <=( a18356a  and  a18351a );
 a18361a <=( (not A268)  and  (not A267) );
 a18362a <=( A203  and  a18361a );
 a18366a <=( A300  and  A299 );
 a18367a <=( (not A269)  and  a18366a );
 a18368a <=( a18367a  and  a18362a );
 a18372a <=( A167  and  (not A168) );
 a18373a <=( (not A169)  and  a18372a );
 a18377a <=( (not A200)  and  A199 );
 a18378a <=( A166  and  a18377a );
 a18379a <=( a18378a  and  a18373a );
 a18383a <=( (not A268)  and  (not A267) );
 a18384a <=( A203  and  a18383a );
 a18388a <=( A300  and  A298 );
 a18389a <=( (not A269)  and  a18388a );
 a18390a <=( a18389a  and  a18384a );
 a18394a <=( A167  and  (not A168) );
 a18395a <=( (not A169)  and  a18394a );
 a18399a <=( (not A200)  and  A199 );
 a18400a <=( A166  and  a18399a );
 a18401a <=( a18400a  and  a18395a );
 a18405a <=( A266  and  A265 );
 a18406a <=( A203  and  a18405a );
 a18410a <=( A301  and  (not A268) );
 a18411a <=( (not A267)  and  a18410a );
 a18412a <=( a18411a  and  a18406a );
 a18416a <=( A167  and  (not A168) );
 a18417a <=( (not A169)  and  a18416a );
 a18421a <=( (not A200)  and  A199 );
 a18422a <=( A166  and  a18421a );
 a18423a <=( a18422a  and  a18417a );
 a18427a <=( (not A266)  and  (not A265) );
 a18428a <=( A203  and  a18427a );
 a18432a <=( A300  and  A299 );
 a18433a <=( (not A268)  and  a18432a );
 a18434a <=( a18433a  and  a18428a );
 a18438a <=( A167  and  (not A168) );
 a18439a <=( (not A169)  and  a18438a );
 a18443a <=( (not A200)  and  A199 );
 a18444a <=( A166  and  a18443a );
 a18445a <=( a18444a  and  a18439a );
 a18449a <=( (not A266)  and  (not A265) );
 a18450a <=( A203  and  a18449a );
 a18454a <=( A300  and  A298 );
 a18455a <=( (not A268)  and  a18454a );
 a18456a <=( a18455a  and  a18450a );
 a18460a <=( A167  and  (not A168) );
 a18461a <=( (not A169)  and  a18460a );
 a18465a <=( (not A200)  and  (not A199) );
 a18466a <=( A166  and  a18465a );
 a18467a <=( a18466a  and  a18461a );
 a18471a <=( A298  and  A268 );
 a18472a <=( (not A202)  and  a18471a );
 a18476a <=( (not A301)  and  (not A300) );
 a18477a <=( A299  and  a18476a );
 a18478a <=( a18477a  and  a18472a );
 a18482a <=( A167  and  (not A168) );
 a18483a <=( (not A169)  and  a18482a );
 a18487a <=( (not A200)  and  (not A199) );
 a18488a <=( A166  and  a18487a );
 a18489a <=( a18488a  and  a18483a );
 a18493a <=( A267  and  A265 );
 a18494a <=( (not A202)  and  a18493a );
 a18498a <=( (not A302)  and  (not A301) );
 a18499a <=( (not A300)  and  a18498a );
 a18500a <=( a18499a  and  a18494a );
 a18504a <=( A167  and  (not A168) );
 a18505a <=( (not A169)  and  a18504a );
 a18509a <=( (not A200)  and  (not A199) );
 a18510a <=( A166  and  a18509a );
 a18511a <=( a18510a  and  a18505a );
 a18515a <=( A267  and  A265 );
 a18516a <=( (not A202)  and  a18515a );
 a18520a <=( (not A301)  and  (not A299) );
 a18521a <=( (not A298)  and  a18520a );
 a18522a <=( a18521a  and  a18516a );
 a18526a <=( A167  and  (not A168) );
 a18527a <=( (not A169)  and  a18526a );
 a18531a <=( (not A200)  and  (not A199) );
 a18532a <=( A166  and  a18531a );
 a18533a <=( a18532a  and  a18527a );
 a18537a <=( A267  and  A266 );
 a18538a <=( (not A202)  and  a18537a );
 a18542a <=( (not A302)  and  (not A301) );
 a18543a <=( (not A300)  and  a18542a );
 a18544a <=( a18543a  and  a18538a );
 a18548a <=( A167  and  (not A168) );
 a18549a <=( (not A169)  and  a18548a );
 a18553a <=( (not A200)  and  (not A199) );
 a18554a <=( A166  and  a18553a );
 a18555a <=( a18554a  and  a18549a );
 a18559a <=( A267  and  A266 );
 a18560a <=( (not A202)  and  a18559a );
 a18564a <=( (not A301)  and  (not A299) );
 a18565a <=( (not A298)  and  a18564a );
 a18566a <=( a18565a  and  a18560a );
 a18570a <=( (not A168)  and  (not A169) );
 a18571a <=( (not A170)  and  a18570a );
 a18575a <=( (not A203)  and  (not A202) );
 a18576a <=( (not A201)  and  a18575a );
 a18577a <=( a18576a  and  a18571a );
 a18581a <=( A298  and  A267 );
 a18582a <=( A265  and  a18581a );
 a18586a <=( (not A301)  and  (not A300) );
 a18587a <=( A299  and  a18586a );
 a18588a <=( a18587a  and  a18582a );
 a18592a <=( (not A168)  and  (not A169) );
 a18593a <=( (not A170)  and  a18592a );
 a18597a <=( (not A203)  and  (not A202) );
 a18598a <=( (not A201)  and  a18597a );
 a18599a <=( a18598a  and  a18593a );
 a18603a <=( A298  and  A267 );
 a18604a <=( A266  and  a18603a );
 a18608a <=( (not A301)  and  (not A300) );
 a18609a <=( A299  and  a18608a );
 a18610a <=( a18609a  and  a18604a );
 a18614a <=( (not A168)  and  (not A169) );
 a18615a <=( (not A170)  and  a18614a );
 a18619a <=( (not A203)  and  (not A202) );
 a18620a <=( (not A201)  and  a18619a );
 a18621a <=( a18620a  and  a18615a );
 a18625a <=( A269  and  A266 );
 a18626a <=( (not A265)  and  a18625a );
 a18630a <=( (not A302)  and  (not A301) );
 a18631a <=( (not A300)  and  a18630a );
 a18632a <=( a18631a  and  a18626a );
 a18636a <=( (not A168)  and  (not A169) );
 a18637a <=( (not A170)  and  a18636a );
 a18641a <=( (not A203)  and  (not A202) );
 a18642a <=( (not A201)  and  a18641a );
 a18643a <=( a18642a  and  a18637a );
 a18647a <=( A269  and  A266 );
 a18648a <=( (not A265)  and  a18647a );
 a18652a <=( (not A301)  and  (not A299) );
 a18653a <=( (not A298)  and  a18652a );
 a18654a <=( a18653a  and  a18648a );
 a18658a <=( (not A168)  and  (not A169) );
 a18659a <=( (not A170)  and  a18658a );
 a18663a <=( (not A203)  and  (not A202) );
 a18664a <=( (not A201)  and  a18663a );
 a18665a <=( a18664a  and  a18659a );
 a18669a <=( A269  and  (not A266) );
 a18670a <=( A265  and  a18669a );
 a18674a <=( (not A302)  and  (not A301) );
 a18675a <=( (not A300)  and  a18674a );
 a18676a <=( a18675a  and  a18670a );
 a18680a <=( (not A168)  and  (not A169) );
 a18681a <=( (not A170)  and  a18680a );
 a18685a <=( (not A203)  and  (not A202) );
 a18686a <=( (not A201)  and  a18685a );
 a18687a <=( a18686a  and  a18681a );
 a18691a <=( A269  and  (not A266) );
 a18692a <=( A265  and  a18691a );
 a18696a <=( (not A301)  and  (not A299) );
 a18697a <=( (not A298)  and  a18696a );
 a18698a <=( a18697a  and  a18692a );
 a18702a <=( (not A168)  and  (not A169) );
 a18703a <=( (not A170)  and  a18702a );
 a18707a <=( A265  and  A201 );
 a18708a <=( A199  and  a18707a );
 a18709a <=( a18708a  and  a18703a );
 a18713a <=( (not A268)  and  (not A267) );
 a18714a <=( A266  and  a18713a );
 a18718a <=( A302  and  (not A299) );
 a18719a <=( A298  and  a18718a );
 a18720a <=( a18719a  and  a18714a );
 a18724a <=( (not A168)  and  (not A169) );
 a18725a <=( (not A170)  and  a18724a );
 a18729a <=( A265  and  A201 );
 a18730a <=( A199  and  a18729a );
 a18731a <=( a18730a  and  a18725a );
 a18735a <=( (not A268)  and  (not A267) );
 a18736a <=( A266  and  a18735a );
 a18740a <=( A302  and  A299 );
 a18741a <=( (not A298)  and  a18740a );
 a18742a <=( a18741a  and  a18736a );
 a18746a <=( (not A168)  and  (not A169) );
 a18747a <=( (not A170)  and  a18746a );
 a18751a <=( A265  and  A201 );
 a18752a <=( A200  and  a18751a );
 a18753a <=( a18752a  and  a18747a );
 a18757a <=( (not A268)  and  (not A267) );
 a18758a <=( A266  and  a18757a );
 a18762a <=( A302  and  (not A299) );
 a18763a <=( A298  and  a18762a );
 a18764a <=( a18763a  and  a18758a );
 a18768a <=( (not A168)  and  (not A169) );
 a18769a <=( (not A170)  and  a18768a );
 a18773a <=( A265  and  A201 );
 a18774a <=( A200  and  a18773a );
 a18775a <=( a18774a  and  a18769a );
 a18779a <=( (not A268)  and  (not A267) );
 a18780a <=( A266  and  a18779a );
 a18784a <=( A302  and  A299 );
 a18785a <=( (not A298)  and  a18784a );
 a18786a <=( a18785a  and  a18780a );
 a18790a <=( (not A168)  and  (not A169) );
 a18791a <=( (not A170)  and  a18790a );
 a18795a <=( (not A201)  and  A200 );
 a18796a <=( A199  and  a18795a );
 a18797a <=( a18796a  and  a18791a );
 a18801a <=( A298  and  A268 );
 a18802a <=( (not A202)  and  a18801a );
 a18806a <=( (not A301)  and  (not A300) );
 a18807a <=( A299  and  a18806a );
 a18808a <=( a18807a  and  a18802a );
 a18812a <=( (not A168)  and  (not A169) );
 a18813a <=( (not A170)  and  a18812a );
 a18817a <=( (not A201)  and  A200 );
 a18818a <=( A199  and  a18817a );
 a18819a <=( a18818a  and  a18813a );
 a18823a <=( A267  and  A265 );
 a18824a <=( (not A202)  and  a18823a );
 a18828a <=( (not A302)  and  (not A301) );
 a18829a <=( (not A300)  and  a18828a );
 a18830a <=( a18829a  and  a18824a );
 a18834a <=( (not A168)  and  (not A169) );
 a18835a <=( (not A170)  and  a18834a );
 a18839a <=( (not A201)  and  A200 );
 a18840a <=( A199  and  a18839a );
 a18841a <=( a18840a  and  a18835a );
 a18845a <=( A267  and  A265 );
 a18846a <=( (not A202)  and  a18845a );
 a18850a <=( (not A301)  and  (not A299) );
 a18851a <=( (not A298)  and  a18850a );
 a18852a <=( a18851a  and  a18846a );
 a18856a <=( (not A168)  and  (not A169) );
 a18857a <=( (not A170)  and  a18856a );
 a18861a <=( (not A201)  and  A200 );
 a18862a <=( A199  and  a18861a );
 a18863a <=( a18862a  and  a18857a );
 a18867a <=( A267  and  A266 );
 a18868a <=( (not A202)  and  a18867a );
 a18872a <=( (not A302)  and  (not A301) );
 a18873a <=( (not A300)  and  a18872a );
 a18874a <=( a18873a  and  a18868a );
 a18878a <=( (not A168)  and  (not A169) );
 a18879a <=( (not A170)  and  a18878a );
 a18883a <=( (not A201)  and  A200 );
 a18884a <=( A199  and  a18883a );
 a18885a <=( a18884a  and  a18879a );
 a18889a <=( A267  and  A266 );
 a18890a <=( (not A202)  and  a18889a );
 a18894a <=( (not A301)  and  (not A299) );
 a18895a <=( (not A298)  and  a18894a );
 a18896a <=( a18895a  and  a18890a );
 a18900a <=( (not A168)  and  (not A169) );
 a18901a <=( (not A170)  and  a18900a );
 a18905a <=( A203  and  A200 );
 a18906a <=( (not A199)  and  a18905a );
 a18907a <=( a18906a  and  a18901a );
 a18911a <=( (not A269)  and  (not A268) );
 a18912a <=( (not A267)  and  a18911a );
 a18916a <=( A302  and  (not A299) );
 a18917a <=( A298  and  a18916a );
 a18918a <=( a18917a  and  a18912a );
 a18922a <=( (not A168)  and  (not A169) );
 a18923a <=( (not A170)  and  a18922a );
 a18927a <=( A203  and  A200 );
 a18928a <=( (not A199)  and  a18927a );
 a18929a <=( a18928a  and  a18923a );
 a18933a <=( (not A269)  and  (not A268) );
 a18934a <=( (not A267)  and  a18933a );
 a18938a <=( A302  and  A299 );
 a18939a <=( (not A298)  and  a18938a );
 a18940a <=( a18939a  and  a18934a );
 a18944a <=( (not A168)  and  (not A169) );
 a18945a <=( (not A170)  and  a18944a );
 a18949a <=( A203  and  A200 );
 a18950a <=( (not A199)  and  a18949a );
 a18951a <=( a18950a  and  a18945a );
 a18955a <=( (not A267)  and  A266 );
 a18956a <=( A265  and  a18955a );
 a18960a <=( A300  and  A299 );
 a18961a <=( (not A268)  and  a18960a );
 a18962a <=( a18961a  and  a18956a );
 a18966a <=( (not A168)  and  (not A169) );
 a18967a <=( (not A170)  and  a18966a );
 a18971a <=( A203  and  A200 );
 a18972a <=( (not A199)  and  a18971a );
 a18973a <=( a18972a  and  a18967a );
 a18977a <=( (not A267)  and  A266 );
 a18978a <=( A265  and  a18977a );
 a18982a <=( A300  and  A298 );
 a18983a <=( (not A268)  and  a18982a );
 a18984a <=( a18983a  and  a18978a );
 a18988a <=( (not A168)  and  (not A169) );
 a18989a <=( (not A170)  and  a18988a );
 a18993a <=( A203  and  A200 );
 a18994a <=( (not A199)  and  a18993a );
 a18995a <=( a18994a  and  a18989a );
 a18999a <=( (not A268)  and  (not A266) );
 a19000a <=( (not A265)  and  a18999a );
 a19004a <=( A302  and  (not A299) );
 a19005a <=( A298  and  a19004a );
 a19006a <=( a19005a  and  a19000a );
 a19010a <=( (not A168)  and  (not A169) );
 a19011a <=( (not A170)  and  a19010a );
 a19015a <=( A203  and  A200 );
 a19016a <=( (not A199)  and  a19015a );
 a19017a <=( a19016a  and  a19011a );
 a19021a <=( (not A268)  and  (not A266) );
 a19022a <=( (not A265)  and  a19021a );
 a19026a <=( A302  and  A299 );
 a19027a <=( (not A298)  and  a19026a );
 a19028a <=( a19027a  and  a19022a );
 a19032a <=( (not A168)  and  (not A169) );
 a19033a <=( (not A170)  and  a19032a );
 a19037a <=( A203  and  (not A200) );
 a19038a <=( A199  and  a19037a );
 a19039a <=( a19038a  and  a19033a );
 a19043a <=( (not A269)  and  (not A268) );
 a19044a <=( (not A267)  and  a19043a );
 a19048a <=( A302  and  (not A299) );
 a19049a <=( A298  and  a19048a );
 a19050a <=( a19049a  and  a19044a );
 a19054a <=( (not A168)  and  (not A169) );
 a19055a <=( (not A170)  and  a19054a );
 a19059a <=( A203  and  (not A200) );
 a19060a <=( A199  and  a19059a );
 a19061a <=( a19060a  and  a19055a );
 a19065a <=( (not A269)  and  (not A268) );
 a19066a <=( (not A267)  and  a19065a );
 a19070a <=( A302  and  A299 );
 a19071a <=( (not A298)  and  a19070a );
 a19072a <=( a19071a  and  a19066a );
 a19076a <=( (not A168)  and  (not A169) );
 a19077a <=( (not A170)  and  a19076a );
 a19081a <=( A203  and  (not A200) );
 a19082a <=( A199  and  a19081a );
 a19083a <=( a19082a  and  a19077a );
 a19087a <=( (not A267)  and  A266 );
 a19088a <=( A265  and  a19087a );
 a19092a <=( A300  and  A299 );
 a19093a <=( (not A268)  and  a19092a );
 a19094a <=( a19093a  and  a19088a );
 a19098a <=( (not A168)  and  (not A169) );
 a19099a <=( (not A170)  and  a19098a );
 a19103a <=( A203  and  (not A200) );
 a19104a <=( A199  and  a19103a );
 a19105a <=( a19104a  and  a19099a );
 a19109a <=( (not A267)  and  A266 );
 a19110a <=( A265  and  a19109a );
 a19114a <=( A300  and  A298 );
 a19115a <=( (not A268)  and  a19114a );
 a19116a <=( a19115a  and  a19110a );
 a19120a <=( (not A168)  and  (not A169) );
 a19121a <=( (not A170)  and  a19120a );
 a19125a <=( A203  and  (not A200) );
 a19126a <=( A199  and  a19125a );
 a19127a <=( a19126a  and  a19121a );
 a19131a <=( (not A268)  and  (not A266) );
 a19132a <=( (not A265)  and  a19131a );
 a19136a <=( A302  and  (not A299) );
 a19137a <=( A298  and  a19136a );
 a19138a <=( a19137a  and  a19132a );
 a19142a <=( (not A168)  and  (not A169) );
 a19143a <=( (not A170)  and  a19142a );
 a19147a <=( A203  and  (not A200) );
 a19148a <=( A199  and  a19147a );
 a19149a <=( a19148a  and  a19143a );
 a19153a <=( (not A268)  and  (not A266) );
 a19154a <=( (not A265)  and  a19153a );
 a19158a <=( A302  and  A299 );
 a19159a <=( (not A298)  and  a19158a );
 a19160a <=( a19159a  and  a19154a );
 a19164a <=( (not A168)  and  (not A169) );
 a19165a <=( (not A170)  and  a19164a );
 a19169a <=( (not A202)  and  (not A200) );
 a19170a <=( (not A199)  and  a19169a );
 a19171a <=( a19170a  and  a19165a );
 a19175a <=( A298  and  A267 );
 a19176a <=( A265  and  a19175a );
 a19180a <=( (not A301)  and  (not A300) );
 a19181a <=( A299  and  a19180a );
 a19182a <=( a19181a  and  a19176a );
 a19186a <=( (not A168)  and  (not A169) );
 a19187a <=( (not A170)  and  a19186a );
 a19191a <=( (not A202)  and  (not A200) );
 a19192a <=( (not A199)  and  a19191a );
 a19193a <=( a19192a  and  a19187a );
 a19197a <=( A298  and  A267 );
 a19198a <=( A266  and  a19197a );
 a19202a <=( (not A301)  and  (not A300) );
 a19203a <=( A299  and  a19202a );
 a19204a <=( a19203a  and  a19198a );
 a19208a <=( (not A168)  and  (not A169) );
 a19209a <=( (not A170)  and  a19208a );
 a19213a <=( (not A202)  and  (not A200) );
 a19214a <=( (not A199)  and  a19213a );
 a19215a <=( a19214a  and  a19209a );
 a19219a <=( A269  and  A266 );
 a19220a <=( (not A265)  and  a19219a );
 a19224a <=( (not A302)  and  (not A301) );
 a19225a <=( (not A300)  and  a19224a );
 a19226a <=( a19225a  and  a19220a );
 a19230a <=( (not A168)  and  (not A169) );
 a19231a <=( (not A170)  and  a19230a );
 a19235a <=( (not A202)  and  (not A200) );
 a19236a <=( (not A199)  and  a19235a );
 a19237a <=( a19236a  and  a19231a );
 a19241a <=( A269  and  A266 );
 a19242a <=( (not A265)  and  a19241a );
 a19246a <=( (not A301)  and  (not A299) );
 a19247a <=( (not A298)  and  a19246a );
 a19248a <=( a19247a  and  a19242a );
 a19252a <=( (not A168)  and  (not A169) );
 a19253a <=( (not A170)  and  a19252a );
 a19257a <=( (not A202)  and  (not A200) );
 a19258a <=( (not A199)  and  a19257a );
 a19259a <=( a19258a  and  a19253a );
 a19263a <=( A269  and  (not A266) );
 a19264a <=( A265  and  a19263a );
 a19268a <=( (not A302)  and  (not A301) );
 a19269a <=( (not A300)  and  a19268a );
 a19270a <=( a19269a  and  a19264a );
 a19274a <=( (not A168)  and  (not A169) );
 a19275a <=( (not A170)  and  a19274a );
 a19279a <=( (not A202)  and  (not A200) );
 a19280a <=( (not A199)  and  a19279a );
 a19281a <=( a19280a  and  a19275a );
 a19285a <=( A269  and  (not A266) );
 a19286a <=( A265  and  a19285a );
 a19290a <=( (not A301)  and  (not A299) );
 a19291a <=( (not A298)  and  a19290a );
 a19292a <=( a19291a  and  a19286a );
 a19296a <=( A199  and  A166 );
 a19297a <=( A168  and  a19296a );
 a19301a <=( (not A202)  and  (not A201) );
 a19302a <=( A200  and  a19301a );
 a19303a <=( a19302a  and  a19297a );
 a19307a <=( (not A267)  and  A266 );
 a19308a <=( A265  and  a19307a );
 a19311a <=( A298  and  (not A268) );
 a19314a <=( A302  and  (not A299) );
 a19315a <=( a19314a  and  a19311a );
 a19316a <=( a19315a  and  a19308a );
 a19320a <=( A199  and  A166 );
 a19321a <=( A168  and  a19320a );
 a19325a <=( (not A202)  and  (not A201) );
 a19326a <=( A200  and  a19325a );
 a19327a <=( a19326a  and  a19321a );
 a19331a <=( (not A267)  and  A266 );
 a19332a <=( A265  and  a19331a );
 a19335a <=( (not A298)  and  (not A268) );
 a19338a <=( A302  and  A299 );
 a19339a <=( a19338a  and  a19335a );
 a19340a <=( a19339a  and  a19332a );
 a19344a <=( A199  and  A167 );
 a19345a <=( A168  and  a19344a );
 a19349a <=( (not A202)  and  (not A201) );
 a19350a <=( A200  and  a19349a );
 a19351a <=( a19350a  and  a19345a );
 a19355a <=( (not A267)  and  A266 );
 a19356a <=( A265  and  a19355a );
 a19359a <=( A298  and  (not A268) );
 a19362a <=( A302  and  (not A299) );
 a19363a <=( a19362a  and  a19359a );
 a19364a <=( a19363a  and  a19356a );
 a19368a <=( A199  and  A167 );
 a19369a <=( A168  and  a19368a );
 a19373a <=( (not A202)  and  (not A201) );
 a19374a <=( A200  and  a19373a );
 a19375a <=( a19374a  and  a19369a );
 a19379a <=( (not A267)  and  A266 );
 a19380a <=( A265  and  a19379a );
 a19383a <=( (not A298)  and  (not A268) );
 a19386a <=( A302  and  A299 );
 a19387a <=( a19386a  and  a19383a );
 a19388a <=( a19387a  and  a19380a );
 a19392a <=( (not A166)  and  A167 );
 a19393a <=( A170  and  a19392a );
 a19397a <=( (not A203)  and  (not A202) );
 a19398a <=( (not A201)  and  a19397a );
 a19399a <=( a19398a  and  a19393a );
 a19403a <=( (not A267)  and  A266 );
 a19404a <=( A265  and  a19403a );
 a19407a <=( A298  and  (not A268) );
 a19410a <=( A302  and  (not A299) );
 a19411a <=( a19410a  and  a19407a );
 a19412a <=( a19411a  and  a19404a );
 a19416a <=( (not A166)  and  A167 );
 a19417a <=( A170  and  a19416a );
 a19421a <=( (not A203)  and  (not A202) );
 a19422a <=( (not A201)  and  a19421a );
 a19423a <=( a19422a  and  a19417a );
 a19427a <=( (not A267)  and  A266 );
 a19428a <=( A265  and  a19427a );
 a19431a <=( (not A298)  and  (not A268) );
 a19434a <=( A302  and  A299 );
 a19435a <=( a19434a  and  a19431a );
 a19436a <=( a19435a  and  a19428a );
 a19440a <=( (not A166)  and  A167 );
 a19441a <=( A170  and  a19440a );
 a19445a <=( (not A201)  and  A200 );
 a19446a <=( A199  and  a19445a );
 a19447a <=( a19446a  and  a19441a );
 a19451a <=( (not A268)  and  (not A267) );
 a19452a <=( (not A202)  and  a19451a );
 a19455a <=( A298  and  (not A269) );
 a19458a <=( A302  and  (not A299) );
 a19459a <=( a19458a  and  a19455a );
 a19460a <=( a19459a  and  a19452a );
 a19464a <=( (not A166)  and  A167 );
 a19465a <=( A170  and  a19464a );
 a19469a <=( (not A201)  and  A200 );
 a19470a <=( A199  and  a19469a );
 a19471a <=( a19470a  and  a19465a );
 a19475a <=( (not A268)  and  (not A267) );
 a19476a <=( (not A202)  and  a19475a );
 a19479a <=( (not A298)  and  (not A269) );
 a19482a <=( A302  and  A299 );
 a19483a <=( a19482a  and  a19479a );
 a19484a <=( a19483a  and  a19476a );
 a19488a <=( (not A166)  and  A167 );
 a19489a <=( A170  and  a19488a );
 a19493a <=( (not A201)  and  A200 );
 a19494a <=( A199  and  a19493a );
 a19495a <=( a19494a  and  a19489a );
 a19499a <=( A266  and  A265 );
 a19500a <=( (not A202)  and  a19499a );
 a19503a <=( (not A268)  and  (not A267) );
 a19506a <=( A300  and  A299 );
 a19507a <=( a19506a  and  a19503a );
 a19508a <=( a19507a  and  a19500a );
 a19512a <=( (not A166)  and  A167 );
 a19513a <=( A170  and  a19512a );
 a19517a <=( (not A201)  and  A200 );
 a19518a <=( A199  and  a19517a );
 a19519a <=( a19518a  and  a19513a );
 a19523a <=( A266  and  A265 );
 a19524a <=( (not A202)  and  a19523a );
 a19527a <=( (not A268)  and  (not A267) );
 a19530a <=( A300  and  A298 );
 a19531a <=( a19530a  and  a19527a );
 a19532a <=( a19531a  and  a19524a );
 a19536a <=( (not A166)  and  A167 );
 a19537a <=( A170  and  a19536a );
 a19541a <=( (not A201)  and  A200 );
 a19542a <=( A199  and  a19541a );
 a19543a <=( a19542a  and  a19537a );
 a19547a <=( (not A266)  and  (not A265) );
 a19548a <=( (not A202)  and  a19547a );
 a19551a <=( A298  and  (not A268) );
 a19554a <=( A302  and  (not A299) );
 a19555a <=( a19554a  and  a19551a );
 a19556a <=( a19555a  and  a19548a );
 a19560a <=( (not A166)  and  A167 );
 a19561a <=( A170  and  a19560a );
 a19565a <=( (not A201)  and  A200 );
 a19566a <=( A199  and  a19565a );
 a19567a <=( a19566a  and  a19561a );
 a19571a <=( (not A266)  and  (not A265) );
 a19572a <=( (not A202)  and  a19571a );
 a19575a <=( (not A298)  and  (not A268) );
 a19578a <=( A302  and  A299 );
 a19579a <=( a19578a  and  a19575a );
 a19580a <=( a19579a  and  a19572a );
 a19584a <=( (not A166)  and  A167 );
 a19585a <=( A170  and  a19584a );
 a19589a <=( A203  and  A200 );
 a19590a <=( (not A199)  and  a19589a );
 a19591a <=( a19590a  and  a19585a );
 a19595a <=( A269  and  A266 );
 a19596a <=( (not A265)  and  a19595a );
 a19599a <=( A299  and  A298 );
 a19602a <=( (not A301)  and  (not A300) );
 a19603a <=( a19602a  and  a19599a );
 a19604a <=( a19603a  and  a19596a );
 a19608a <=( (not A166)  and  A167 );
 a19609a <=( A170  and  a19608a );
 a19613a <=( A203  and  A200 );
 a19614a <=( (not A199)  and  a19613a );
 a19615a <=( a19614a  and  a19609a );
 a19619a <=( A269  and  (not A266) );
 a19620a <=( A265  and  a19619a );
 a19623a <=( A299  and  A298 );
 a19626a <=( (not A301)  and  (not A300) );
 a19627a <=( a19626a  and  a19623a );
 a19628a <=( a19627a  and  a19620a );
 a19632a <=( (not A166)  and  A167 );
 a19633a <=( A170  and  a19632a );
 a19637a <=( A203  and  (not A200) );
 a19638a <=( A199  and  a19637a );
 a19639a <=( a19638a  and  a19633a );
 a19643a <=( A269  and  A266 );
 a19644a <=( (not A265)  and  a19643a );
 a19647a <=( A299  and  A298 );
 a19650a <=( (not A301)  and  (not A300) );
 a19651a <=( a19650a  and  a19647a );
 a19652a <=( a19651a  and  a19644a );
 a19656a <=( (not A166)  and  A167 );
 a19657a <=( A170  and  a19656a );
 a19661a <=( A203  and  (not A200) );
 a19662a <=( A199  and  a19661a );
 a19663a <=( a19662a  and  a19657a );
 a19667a <=( A269  and  (not A266) );
 a19668a <=( A265  and  a19667a );
 a19671a <=( A299  and  A298 );
 a19674a <=( (not A301)  and  (not A300) );
 a19675a <=( a19674a  and  a19671a );
 a19676a <=( a19675a  and  a19668a );
 a19680a <=( (not A166)  and  A167 );
 a19681a <=( A170  and  a19680a );
 a19685a <=( (not A202)  and  (not A200) );
 a19686a <=( (not A199)  and  a19685a );
 a19687a <=( a19686a  and  a19681a );
 a19691a <=( (not A267)  and  A266 );
 a19692a <=( A265  and  a19691a );
 a19695a <=( A298  and  (not A268) );
 a19698a <=( A302  and  (not A299) );
 a19699a <=( a19698a  and  a19695a );
 a19700a <=( a19699a  and  a19692a );
 a19704a <=( (not A166)  and  A167 );
 a19705a <=( A170  and  a19704a );
 a19709a <=( (not A202)  and  (not A200) );
 a19710a <=( (not A199)  and  a19709a );
 a19711a <=( a19710a  and  a19705a );
 a19715a <=( (not A267)  and  A266 );
 a19716a <=( A265  and  a19715a );
 a19719a <=( (not A298)  and  (not A268) );
 a19722a <=( A302  and  A299 );
 a19723a <=( a19722a  and  a19719a );
 a19724a <=( a19723a  and  a19716a );
 a19728a <=( A166  and  (not A167) );
 a19729a <=( A170  and  a19728a );
 a19733a <=( (not A203)  and  (not A202) );
 a19734a <=( (not A201)  and  a19733a );
 a19735a <=( a19734a  and  a19729a );
 a19739a <=( (not A267)  and  A266 );
 a19740a <=( A265  and  a19739a );
 a19743a <=( A298  and  (not A268) );
 a19746a <=( A302  and  (not A299) );
 a19747a <=( a19746a  and  a19743a );
 a19748a <=( a19747a  and  a19740a );
 a19752a <=( A166  and  (not A167) );
 a19753a <=( A170  and  a19752a );
 a19757a <=( (not A203)  and  (not A202) );
 a19758a <=( (not A201)  and  a19757a );
 a19759a <=( a19758a  and  a19753a );
 a19763a <=( (not A267)  and  A266 );
 a19764a <=( A265  and  a19763a );
 a19767a <=( (not A298)  and  (not A268) );
 a19770a <=( A302  and  A299 );
 a19771a <=( a19770a  and  a19767a );
 a19772a <=( a19771a  and  a19764a );
 a19776a <=( A166  and  (not A167) );
 a19777a <=( A170  and  a19776a );
 a19781a <=( (not A201)  and  A200 );
 a19782a <=( A199  and  a19781a );
 a19783a <=( a19782a  and  a19777a );
 a19787a <=( (not A268)  and  (not A267) );
 a19788a <=( (not A202)  and  a19787a );
 a19791a <=( A298  and  (not A269) );
 a19794a <=( A302  and  (not A299) );
 a19795a <=( a19794a  and  a19791a );
 a19796a <=( a19795a  and  a19788a );
 a19800a <=( A166  and  (not A167) );
 a19801a <=( A170  and  a19800a );
 a19805a <=( (not A201)  and  A200 );
 a19806a <=( A199  and  a19805a );
 a19807a <=( a19806a  and  a19801a );
 a19811a <=( (not A268)  and  (not A267) );
 a19812a <=( (not A202)  and  a19811a );
 a19815a <=( (not A298)  and  (not A269) );
 a19818a <=( A302  and  A299 );
 a19819a <=( a19818a  and  a19815a );
 a19820a <=( a19819a  and  a19812a );
 a19824a <=( A166  and  (not A167) );
 a19825a <=( A170  and  a19824a );
 a19829a <=( (not A201)  and  A200 );
 a19830a <=( A199  and  a19829a );
 a19831a <=( a19830a  and  a19825a );
 a19835a <=( A266  and  A265 );
 a19836a <=( (not A202)  and  a19835a );
 a19839a <=( (not A268)  and  (not A267) );
 a19842a <=( A300  and  A299 );
 a19843a <=( a19842a  and  a19839a );
 a19844a <=( a19843a  and  a19836a );
 a19848a <=( A166  and  (not A167) );
 a19849a <=( A170  and  a19848a );
 a19853a <=( (not A201)  and  A200 );
 a19854a <=( A199  and  a19853a );
 a19855a <=( a19854a  and  a19849a );
 a19859a <=( A266  and  A265 );
 a19860a <=( (not A202)  and  a19859a );
 a19863a <=( (not A268)  and  (not A267) );
 a19866a <=( A300  and  A298 );
 a19867a <=( a19866a  and  a19863a );
 a19868a <=( a19867a  and  a19860a );
 a19872a <=( A166  and  (not A167) );
 a19873a <=( A170  and  a19872a );
 a19877a <=( (not A201)  and  A200 );
 a19878a <=( A199  and  a19877a );
 a19879a <=( a19878a  and  a19873a );
 a19883a <=( (not A266)  and  (not A265) );
 a19884a <=( (not A202)  and  a19883a );
 a19887a <=( A298  and  (not A268) );
 a19890a <=( A302  and  (not A299) );
 a19891a <=( a19890a  and  a19887a );
 a19892a <=( a19891a  and  a19884a );
 a19896a <=( A166  and  (not A167) );
 a19897a <=( A170  and  a19896a );
 a19901a <=( (not A201)  and  A200 );
 a19902a <=( A199  and  a19901a );
 a19903a <=( a19902a  and  a19897a );
 a19907a <=( (not A266)  and  (not A265) );
 a19908a <=( (not A202)  and  a19907a );
 a19911a <=( (not A298)  and  (not A268) );
 a19914a <=( A302  and  A299 );
 a19915a <=( a19914a  and  a19911a );
 a19916a <=( a19915a  and  a19908a );
 a19920a <=( A166  and  (not A167) );
 a19921a <=( A170  and  a19920a );
 a19925a <=( A203  and  A200 );
 a19926a <=( (not A199)  and  a19925a );
 a19927a <=( a19926a  and  a19921a );
 a19931a <=( A269  and  A266 );
 a19932a <=( (not A265)  and  a19931a );
 a19935a <=( A299  and  A298 );
 a19938a <=( (not A301)  and  (not A300) );
 a19939a <=( a19938a  and  a19935a );
 a19940a <=( a19939a  and  a19932a );
 a19944a <=( A166  and  (not A167) );
 a19945a <=( A170  and  a19944a );
 a19949a <=( A203  and  A200 );
 a19950a <=( (not A199)  and  a19949a );
 a19951a <=( a19950a  and  a19945a );
 a19955a <=( A269  and  (not A266) );
 a19956a <=( A265  and  a19955a );
 a19959a <=( A299  and  A298 );
 a19962a <=( (not A301)  and  (not A300) );
 a19963a <=( a19962a  and  a19959a );
 a19964a <=( a19963a  and  a19956a );
 a19968a <=( A166  and  (not A167) );
 a19969a <=( A170  and  a19968a );
 a19973a <=( A203  and  (not A200) );
 a19974a <=( A199  and  a19973a );
 a19975a <=( a19974a  and  a19969a );
 a19979a <=( A269  and  A266 );
 a19980a <=( (not A265)  and  a19979a );
 a19983a <=( A299  and  A298 );
 a19986a <=( (not A301)  and  (not A300) );
 a19987a <=( a19986a  and  a19983a );
 a19988a <=( a19987a  and  a19980a );
 a19992a <=( A166  and  (not A167) );
 a19993a <=( A170  and  a19992a );
 a19997a <=( A203  and  (not A200) );
 a19998a <=( A199  and  a19997a );
 a19999a <=( a19998a  and  a19993a );
 a20003a <=( A269  and  (not A266) );
 a20004a <=( A265  and  a20003a );
 a20007a <=( A299  and  A298 );
 a20010a <=( (not A301)  and  (not A300) );
 a20011a <=( a20010a  and  a20007a );
 a20012a <=( a20011a  and  a20004a );
 a20016a <=( A166  and  (not A167) );
 a20017a <=( A170  and  a20016a );
 a20021a <=( (not A202)  and  (not A200) );
 a20022a <=( (not A199)  and  a20021a );
 a20023a <=( a20022a  and  a20017a );
 a20027a <=( (not A267)  and  A266 );
 a20028a <=( A265  and  a20027a );
 a20031a <=( A298  and  (not A268) );
 a20034a <=( A302  and  (not A299) );
 a20035a <=( a20034a  and  a20031a );
 a20036a <=( a20035a  and  a20028a );
 a20040a <=( A166  and  (not A167) );
 a20041a <=( A170  and  a20040a );
 a20045a <=( (not A202)  and  (not A200) );
 a20046a <=( (not A199)  and  a20045a );
 a20047a <=( a20046a  and  a20041a );
 a20051a <=( (not A267)  and  A266 );
 a20052a <=( A265  and  a20051a );
 a20055a <=( (not A298)  and  (not A268) );
 a20058a <=( A302  and  A299 );
 a20059a <=( a20058a  and  a20055a );
 a20060a <=( a20059a  and  a20052a );
 a20064a <=( (not A166)  and  (not A167) );
 a20065a <=( (not A169)  and  a20064a );
 a20069a <=( (not A203)  and  (not A202) );
 a20070a <=( (not A201)  and  a20069a );
 a20071a <=( a20070a  and  a20065a );
 a20075a <=( A269  and  A266 );
 a20076a <=( (not A265)  and  a20075a );
 a20079a <=( A299  and  A298 );
 a20082a <=( (not A301)  and  (not A300) );
 a20083a <=( a20082a  and  a20079a );
 a20084a <=( a20083a  and  a20076a );
 a20088a <=( (not A166)  and  (not A167) );
 a20089a <=( (not A169)  and  a20088a );
 a20093a <=( (not A203)  and  (not A202) );
 a20094a <=( (not A201)  and  a20093a );
 a20095a <=( a20094a  and  a20089a );
 a20099a <=( A269  and  (not A266) );
 a20100a <=( A265  and  a20099a );
 a20103a <=( A299  and  A298 );
 a20106a <=( (not A301)  and  (not A300) );
 a20107a <=( a20106a  and  a20103a );
 a20108a <=( a20107a  and  a20100a );
 a20112a <=( (not A166)  and  (not A167) );
 a20113a <=( (not A169)  and  a20112a );
 a20117a <=( (not A201)  and  A200 );
 a20118a <=( A199  and  a20117a );
 a20119a <=( a20118a  and  a20113a );
 a20123a <=( A267  and  A265 );
 a20124a <=( (not A202)  and  a20123a );
 a20127a <=( A299  and  A298 );
 a20130a <=( (not A301)  and  (not A300) );
 a20131a <=( a20130a  and  a20127a );
 a20132a <=( a20131a  and  a20124a );
 a20136a <=( (not A166)  and  (not A167) );
 a20137a <=( (not A169)  and  a20136a );
 a20141a <=( (not A201)  and  A200 );
 a20142a <=( A199  and  a20141a );
 a20143a <=( a20142a  and  a20137a );
 a20147a <=( A267  and  A266 );
 a20148a <=( (not A202)  and  a20147a );
 a20151a <=( A299  and  A298 );
 a20154a <=( (not A301)  and  (not A300) );
 a20155a <=( a20154a  and  a20151a );
 a20156a <=( a20155a  and  a20148a );
 a20160a <=( (not A166)  and  (not A167) );
 a20161a <=( (not A169)  and  a20160a );
 a20165a <=( (not A201)  and  A200 );
 a20166a <=( A199  and  a20165a );
 a20167a <=( a20166a  and  a20161a );
 a20171a <=( A266  and  (not A265) );
 a20172a <=( (not A202)  and  a20171a );
 a20175a <=( (not A300)  and  A269 );
 a20178a <=( (not A302)  and  (not A301) );
 a20179a <=( a20178a  and  a20175a );
 a20180a <=( a20179a  and  a20172a );
 a20184a <=( (not A166)  and  (not A167) );
 a20185a <=( (not A169)  and  a20184a );
 a20189a <=( (not A201)  and  A200 );
 a20190a <=( A199  and  a20189a );
 a20191a <=( a20190a  and  a20185a );
 a20195a <=( A266  and  (not A265) );
 a20196a <=( (not A202)  and  a20195a );
 a20199a <=( (not A298)  and  A269 );
 a20202a <=( (not A301)  and  (not A299) );
 a20203a <=( a20202a  and  a20199a );
 a20204a <=( a20203a  and  a20196a );
 a20208a <=( (not A166)  and  (not A167) );
 a20209a <=( (not A169)  and  a20208a );
 a20213a <=( (not A201)  and  A200 );
 a20214a <=( A199  and  a20213a );
 a20215a <=( a20214a  and  a20209a );
 a20219a <=( (not A266)  and  A265 );
 a20220a <=( (not A202)  and  a20219a );
 a20223a <=( (not A300)  and  A269 );
 a20226a <=( (not A302)  and  (not A301) );
 a20227a <=( a20226a  and  a20223a );
 a20228a <=( a20227a  and  a20220a );
 a20232a <=( (not A166)  and  (not A167) );
 a20233a <=( (not A169)  and  a20232a );
 a20237a <=( (not A201)  and  A200 );
 a20238a <=( A199  and  a20237a );
 a20239a <=( a20238a  and  a20233a );
 a20243a <=( (not A266)  and  A265 );
 a20244a <=( (not A202)  and  a20243a );
 a20247a <=( (not A298)  and  A269 );
 a20250a <=( (not A301)  and  (not A299) );
 a20251a <=( a20250a  and  a20247a );
 a20252a <=( a20251a  and  a20244a );
 a20256a <=( (not A166)  and  (not A167) );
 a20257a <=( (not A169)  and  a20256a );
 a20261a <=( A203  and  A200 );
 a20262a <=( (not A199)  and  a20261a );
 a20263a <=( a20262a  and  a20257a );
 a20267a <=( (not A267)  and  A266 );
 a20268a <=( A265  and  a20267a );
 a20271a <=( A298  and  (not A268) );
 a20274a <=( A302  and  (not A299) );
 a20275a <=( a20274a  and  a20271a );
 a20276a <=( a20275a  and  a20268a );
 a20280a <=( (not A166)  and  (not A167) );
 a20281a <=( (not A169)  and  a20280a );
 a20285a <=( A203  and  A200 );
 a20286a <=( (not A199)  and  a20285a );
 a20287a <=( a20286a  and  a20281a );
 a20291a <=( (not A267)  and  A266 );
 a20292a <=( A265  and  a20291a );
 a20295a <=( (not A298)  and  (not A268) );
 a20298a <=( A302  and  A299 );
 a20299a <=( a20298a  and  a20295a );
 a20300a <=( a20299a  and  a20292a );
 a20304a <=( (not A166)  and  (not A167) );
 a20305a <=( (not A169)  and  a20304a );
 a20309a <=( A203  and  (not A200) );
 a20310a <=( A199  and  a20309a );
 a20311a <=( a20310a  and  a20305a );
 a20315a <=( (not A267)  and  A266 );
 a20316a <=( A265  and  a20315a );
 a20319a <=( A298  and  (not A268) );
 a20322a <=( A302  and  (not A299) );
 a20323a <=( a20322a  and  a20319a );
 a20324a <=( a20323a  and  a20316a );
 a20328a <=( (not A166)  and  (not A167) );
 a20329a <=( (not A169)  and  a20328a );
 a20333a <=( A203  and  (not A200) );
 a20334a <=( A199  and  a20333a );
 a20335a <=( a20334a  and  a20329a );
 a20339a <=( (not A267)  and  A266 );
 a20340a <=( A265  and  a20339a );
 a20343a <=( (not A298)  and  (not A268) );
 a20346a <=( A302  and  A299 );
 a20347a <=( a20346a  and  a20343a );
 a20348a <=( a20347a  and  a20340a );
 a20352a <=( (not A166)  and  (not A167) );
 a20353a <=( (not A169)  and  a20352a );
 a20357a <=( (not A202)  and  (not A200) );
 a20358a <=( (not A199)  and  a20357a );
 a20359a <=( a20358a  and  a20353a );
 a20363a <=( A269  and  A266 );
 a20364a <=( (not A265)  and  a20363a );
 a20367a <=( A299  and  A298 );
 a20370a <=( (not A301)  and  (not A300) );
 a20371a <=( a20370a  and  a20367a );
 a20372a <=( a20371a  and  a20364a );
 a20376a <=( (not A166)  and  (not A167) );
 a20377a <=( (not A169)  and  a20376a );
 a20381a <=( (not A202)  and  (not A200) );
 a20382a <=( (not A199)  and  a20381a );
 a20383a <=( a20382a  and  a20377a );
 a20387a <=( A269  and  (not A266) );
 a20388a <=( A265  and  a20387a );
 a20391a <=( A299  and  A298 );
 a20394a <=( (not A301)  and  (not A300) );
 a20395a <=( a20394a  and  a20391a );
 a20396a <=( a20395a  and  a20388a );
 a20400a <=( A167  and  (not A168) );
 a20401a <=( (not A169)  and  a20400a );
 a20405a <=( (not A202)  and  (not A201) );
 a20406a <=( A166  and  a20405a );
 a20407a <=( a20406a  and  a20401a );
 a20411a <=( A267  and  A265 );
 a20412a <=( (not A203)  and  a20411a );
 a20415a <=( A299  and  A298 );
 a20418a <=( (not A301)  and  (not A300) );
 a20419a <=( a20418a  and  a20415a );
 a20420a <=( a20419a  and  a20412a );
 a20424a <=( A167  and  (not A168) );
 a20425a <=( (not A169)  and  a20424a );
 a20429a <=( (not A202)  and  (not A201) );
 a20430a <=( A166  and  a20429a );
 a20431a <=( a20430a  and  a20425a );
 a20435a <=( A267  and  A266 );
 a20436a <=( (not A203)  and  a20435a );
 a20439a <=( A299  and  A298 );
 a20442a <=( (not A301)  and  (not A300) );
 a20443a <=( a20442a  and  a20439a );
 a20444a <=( a20443a  and  a20436a );
 a20448a <=( A167  and  (not A168) );
 a20449a <=( (not A169)  and  a20448a );
 a20453a <=( (not A202)  and  (not A201) );
 a20454a <=( A166  and  a20453a );
 a20455a <=( a20454a  and  a20449a );
 a20459a <=( A266  and  (not A265) );
 a20460a <=( (not A203)  and  a20459a );
 a20463a <=( (not A300)  and  A269 );
 a20466a <=( (not A302)  and  (not A301) );
 a20467a <=( a20466a  and  a20463a );
 a20468a <=( a20467a  and  a20460a );
 a20472a <=( A167  and  (not A168) );
 a20473a <=( (not A169)  and  a20472a );
 a20477a <=( (not A202)  and  (not A201) );
 a20478a <=( A166  and  a20477a );
 a20479a <=( a20478a  and  a20473a );
 a20483a <=( A266  and  (not A265) );
 a20484a <=( (not A203)  and  a20483a );
 a20487a <=( (not A298)  and  A269 );
 a20490a <=( (not A301)  and  (not A299) );
 a20491a <=( a20490a  and  a20487a );
 a20492a <=( a20491a  and  a20484a );
 a20496a <=( A167  and  (not A168) );
 a20497a <=( (not A169)  and  a20496a );
 a20501a <=( (not A202)  and  (not A201) );
 a20502a <=( A166  and  a20501a );
 a20503a <=( a20502a  and  a20497a );
 a20507a <=( (not A266)  and  A265 );
 a20508a <=( (not A203)  and  a20507a );
 a20511a <=( (not A300)  and  A269 );
 a20514a <=( (not A302)  and  (not A301) );
 a20515a <=( a20514a  and  a20511a );
 a20516a <=( a20515a  and  a20508a );
 a20520a <=( A167  and  (not A168) );
 a20521a <=( (not A169)  and  a20520a );
 a20525a <=( (not A202)  and  (not A201) );
 a20526a <=( A166  and  a20525a );
 a20527a <=( a20526a  and  a20521a );
 a20531a <=( (not A266)  and  A265 );
 a20532a <=( (not A203)  and  a20531a );
 a20535a <=( (not A298)  and  A269 );
 a20538a <=( (not A301)  and  (not A299) );
 a20539a <=( a20538a  and  a20535a );
 a20540a <=( a20539a  and  a20532a );
 a20544a <=( A167  and  (not A168) );
 a20545a <=( (not A169)  and  a20544a );
 a20549a <=( A201  and  A199 );
 a20550a <=( A166  and  a20549a );
 a20551a <=( a20550a  and  a20545a );
 a20555a <=( (not A267)  and  A266 );
 a20556a <=( A265  and  a20555a );
 a20559a <=( A298  and  (not A268) );
 a20562a <=( A302  and  (not A299) );
 a20563a <=( a20562a  and  a20559a );
 a20564a <=( a20563a  and  a20556a );
 a20568a <=( A167  and  (not A168) );
 a20569a <=( (not A169)  and  a20568a );
 a20573a <=( A201  and  A199 );
 a20574a <=( A166  and  a20573a );
 a20575a <=( a20574a  and  a20569a );
 a20579a <=( (not A267)  and  A266 );
 a20580a <=( A265  and  a20579a );
 a20583a <=( (not A298)  and  (not A268) );
 a20586a <=( A302  and  A299 );
 a20587a <=( a20586a  and  a20583a );
 a20588a <=( a20587a  and  a20580a );
 a20592a <=( A167  and  (not A168) );
 a20593a <=( (not A169)  and  a20592a );
 a20597a <=( A201  and  A200 );
 a20598a <=( A166  and  a20597a );
 a20599a <=( a20598a  and  a20593a );
 a20603a <=( (not A267)  and  A266 );
 a20604a <=( A265  and  a20603a );
 a20607a <=( A298  and  (not A268) );
 a20610a <=( A302  and  (not A299) );
 a20611a <=( a20610a  and  a20607a );
 a20612a <=( a20611a  and  a20604a );
 a20616a <=( A167  and  (not A168) );
 a20617a <=( (not A169)  and  a20616a );
 a20621a <=( A201  and  A200 );
 a20622a <=( A166  and  a20621a );
 a20623a <=( a20622a  and  a20617a );
 a20627a <=( (not A267)  and  A266 );
 a20628a <=( A265  and  a20627a );
 a20631a <=( (not A298)  and  (not A268) );
 a20634a <=( A302  and  A299 );
 a20635a <=( a20634a  and  a20631a );
 a20636a <=( a20635a  and  a20628a );
 a20640a <=( A167  and  (not A168) );
 a20641a <=( (not A169)  and  a20640a );
 a20645a <=( A200  and  A199 );
 a20646a <=( A166  and  a20645a );
 a20647a <=( a20646a  and  a20641a );
 a20651a <=( A268  and  (not A202) );
 a20652a <=( (not A201)  and  a20651a );
 a20655a <=( A299  and  A298 );
 a20658a <=( (not A301)  and  (not A300) );
 a20659a <=( a20658a  and  a20655a );
 a20660a <=( a20659a  and  a20652a );
 a20664a <=( A167  and  (not A168) );
 a20665a <=( (not A169)  and  a20664a );
 a20669a <=( A200  and  A199 );
 a20670a <=( A166  and  a20669a );
 a20671a <=( a20670a  and  a20665a );
 a20675a <=( A265  and  (not A202) );
 a20676a <=( (not A201)  and  a20675a );
 a20679a <=( (not A300)  and  A267 );
 a20682a <=( (not A302)  and  (not A301) );
 a20683a <=( a20682a  and  a20679a );
 a20684a <=( a20683a  and  a20676a );
 a20688a <=( A167  and  (not A168) );
 a20689a <=( (not A169)  and  a20688a );
 a20693a <=( A200  and  A199 );
 a20694a <=( A166  and  a20693a );
 a20695a <=( a20694a  and  a20689a );
 a20699a <=( A265  and  (not A202) );
 a20700a <=( (not A201)  and  a20699a );
 a20703a <=( (not A298)  and  A267 );
 a20706a <=( (not A301)  and  (not A299) );
 a20707a <=( a20706a  and  a20703a );
 a20708a <=( a20707a  and  a20700a );
 a20712a <=( A167  and  (not A168) );
 a20713a <=( (not A169)  and  a20712a );
 a20717a <=( A200  and  A199 );
 a20718a <=( A166  and  a20717a );
 a20719a <=( a20718a  and  a20713a );
 a20723a <=( A266  and  (not A202) );
 a20724a <=( (not A201)  and  a20723a );
 a20727a <=( (not A300)  and  A267 );
 a20730a <=( (not A302)  and  (not A301) );
 a20731a <=( a20730a  and  a20727a );
 a20732a <=( a20731a  and  a20724a );
 a20736a <=( A167  and  (not A168) );
 a20737a <=( (not A169)  and  a20736a );
 a20741a <=( A200  and  A199 );
 a20742a <=( A166  and  a20741a );
 a20743a <=( a20742a  and  a20737a );
 a20747a <=( A266  and  (not A202) );
 a20748a <=( (not A201)  and  a20747a );
 a20751a <=( (not A298)  and  A267 );
 a20754a <=( (not A301)  and  (not A299) );
 a20755a <=( a20754a  and  a20751a );
 a20756a <=( a20755a  and  a20748a );
 a20760a <=( A167  and  (not A168) );
 a20761a <=( (not A169)  and  a20760a );
 a20765a <=( A200  and  (not A199) );
 a20766a <=( A166  and  a20765a );
 a20767a <=( a20766a  and  a20761a );
 a20771a <=( (not A268)  and  (not A267) );
 a20772a <=( A203  and  a20771a );
 a20775a <=( A298  and  (not A269) );
 a20778a <=( A302  and  (not A299) );
 a20779a <=( a20778a  and  a20775a );
 a20780a <=( a20779a  and  a20772a );
 a20784a <=( A167  and  (not A168) );
 a20785a <=( (not A169)  and  a20784a );
 a20789a <=( A200  and  (not A199) );
 a20790a <=( A166  and  a20789a );
 a20791a <=( a20790a  and  a20785a );
 a20795a <=( (not A268)  and  (not A267) );
 a20796a <=( A203  and  a20795a );
 a20799a <=( (not A298)  and  (not A269) );
 a20802a <=( A302  and  A299 );
 a20803a <=( a20802a  and  a20799a );
 a20804a <=( a20803a  and  a20796a );
 a20808a <=( A167  and  (not A168) );
 a20809a <=( (not A169)  and  a20808a );
 a20813a <=( A200  and  (not A199) );
 a20814a <=( A166  and  a20813a );
 a20815a <=( a20814a  and  a20809a );
 a20819a <=( A266  and  A265 );
 a20820a <=( A203  and  a20819a );
 a20823a <=( (not A268)  and  (not A267) );
 a20826a <=( A300  and  A299 );
 a20827a <=( a20826a  and  a20823a );
 a20828a <=( a20827a  and  a20820a );
 a20832a <=( A167  and  (not A168) );
 a20833a <=( (not A169)  and  a20832a );
 a20837a <=( A200  and  (not A199) );
 a20838a <=( A166  and  a20837a );
 a20839a <=( a20838a  and  a20833a );
 a20843a <=( A266  and  A265 );
 a20844a <=( A203  and  a20843a );
 a20847a <=( (not A268)  and  (not A267) );
 a20850a <=( A300  and  A298 );
 a20851a <=( a20850a  and  a20847a );
 a20852a <=( a20851a  and  a20844a );
 a20856a <=( A167  and  (not A168) );
 a20857a <=( (not A169)  and  a20856a );
 a20861a <=( A200  and  (not A199) );
 a20862a <=( A166  and  a20861a );
 a20863a <=( a20862a  and  a20857a );
 a20867a <=( (not A266)  and  (not A265) );
 a20868a <=( A203  and  a20867a );
 a20871a <=( A298  and  (not A268) );
 a20874a <=( A302  and  (not A299) );
 a20875a <=( a20874a  and  a20871a );
 a20876a <=( a20875a  and  a20868a );
 a20880a <=( A167  and  (not A168) );
 a20881a <=( (not A169)  and  a20880a );
 a20885a <=( A200  and  (not A199) );
 a20886a <=( A166  and  a20885a );
 a20887a <=( a20886a  and  a20881a );
 a20891a <=( (not A266)  and  (not A265) );
 a20892a <=( A203  and  a20891a );
 a20895a <=( (not A298)  and  (not A268) );
 a20898a <=( A302  and  A299 );
 a20899a <=( a20898a  and  a20895a );
 a20900a <=( a20899a  and  a20892a );
 a20904a <=( A167  and  (not A168) );
 a20905a <=( (not A169)  and  a20904a );
 a20909a <=( (not A200)  and  A199 );
 a20910a <=( A166  and  a20909a );
 a20911a <=( a20910a  and  a20905a );
 a20915a <=( (not A268)  and  (not A267) );
 a20916a <=( A203  and  a20915a );
 a20919a <=( A298  and  (not A269) );
 a20922a <=( A302  and  (not A299) );
 a20923a <=( a20922a  and  a20919a );
 a20924a <=( a20923a  and  a20916a );
 a20928a <=( A167  and  (not A168) );
 a20929a <=( (not A169)  and  a20928a );
 a20933a <=( (not A200)  and  A199 );
 a20934a <=( A166  and  a20933a );
 a20935a <=( a20934a  and  a20929a );
 a20939a <=( (not A268)  and  (not A267) );
 a20940a <=( A203  and  a20939a );
 a20943a <=( (not A298)  and  (not A269) );
 a20946a <=( A302  and  A299 );
 a20947a <=( a20946a  and  a20943a );
 a20948a <=( a20947a  and  a20940a );
 a20952a <=( A167  and  (not A168) );
 a20953a <=( (not A169)  and  a20952a );
 a20957a <=( (not A200)  and  A199 );
 a20958a <=( A166  and  a20957a );
 a20959a <=( a20958a  and  a20953a );
 a20963a <=( A266  and  A265 );
 a20964a <=( A203  and  a20963a );
 a20967a <=( (not A268)  and  (not A267) );
 a20970a <=( A300  and  A299 );
 a20971a <=( a20970a  and  a20967a );
 a20972a <=( a20971a  and  a20964a );
 a20976a <=( A167  and  (not A168) );
 a20977a <=( (not A169)  and  a20976a );
 a20981a <=( (not A200)  and  A199 );
 a20982a <=( A166  and  a20981a );
 a20983a <=( a20982a  and  a20977a );
 a20987a <=( A266  and  A265 );
 a20988a <=( A203  and  a20987a );
 a20991a <=( (not A268)  and  (not A267) );
 a20994a <=( A300  and  A298 );
 a20995a <=( a20994a  and  a20991a );
 a20996a <=( a20995a  and  a20988a );
 a21000a <=( A167  and  (not A168) );
 a21001a <=( (not A169)  and  a21000a );
 a21005a <=( (not A200)  and  A199 );
 a21006a <=( A166  and  a21005a );
 a21007a <=( a21006a  and  a21001a );
 a21011a <=( (not A266)  and  (not A265) );
 a21012a <=( A203  and  a21011a );
 a21015a <=( A298  and  (not A268) );
 a21018a <=( A302  and  (not A299) );
 a21019a <=( a21018a  and  a21015a );
 a21020a <=( a21019a  and  a21012a );
 a21024a <=( A167  and  (not A168) );
 a21025a <=( (not A169)  and  a21024a );
 a21029a <=( (not A200)  and  A199 );
 a21030a <=( A166  and  a21029a );
 a21031a <=( a21030a  and  a21025a );
 a21035a <=( (not A266)  and  (not A265) );
 a21036a <=( A203  and  a21035a );
 a21039a <=( (not A298)  and  (not A268) );
 a21042a <=( A302  and  A299 );
 a21043a <=( a21042a  and  a21039a );
 a21044a <=( a21043a  and  a21036a );
 a21048a <=( A167  and  (not A168) );
 a21049a <=( (not A169)  and  a21048a );
 a21053a <=( (not A200)  and  (not A199) );
 a21054a <=( A166  and  a21053a );
 a21055a <=( a21054a  and  a21049a );
 a21059a <=( A267  and  A265 );
 a21060a <=( (not A202)  and  a21059a );
 a21063a <=( A299  and  A298 );
 a21066a <=( (not A301)  and  (not A300) );
 a21067a <=( a21066a  and  a21063a );
 a21068a <=( a21067a  and  a21060a );
 a21072a <=( A167  and  (not A168) );
 a21073a <=( (not A169)  and  a21072a );
 a21077a <=( (not A200)  and  (not A199) );
 a21078a <=( A166  and  a21077a );
 a21079a <=( a21078a  and  a21073a );
 a21083a <=( A267  and  A266 );
 a21084a <=( (not A202)  and  a21083a );
 a21087a <=( A299  and  A298 );
 a21090a <=( (not A301)  and  (not A300) );
 a21091a <=( a21090a  and  a21087a );
 a21092a <=( a21091a  and  a21084a );
 a21096a <=( A167  and  (not A168) );
 a21097a <=( (not A169)  and  a21096a );
 a21101a <=( (not A200)  and  (not A199) );
 a21102a <=( A166  and  a21101a );
 a21103a <=( a21102a  and  a21097a );
 a21107a <=( A266  and  (not A265) );
 a21108a <=( (not A202)  and  a21107a );
 a21111a <=( (not A300)  and  A269 );
 a21114a <=( (not A302)  and  (not A301) );
 a21115a <=( a21114a  and  a21111a );
 a21116a <=( a21115a  and  a21108a );
 a21120a <=( A167  and  (not A168) );
 a21121a <=( (not A169)  and  a21120a );
 a21125a <=( (not A200)  and  (not A199) );
 a21126a <=( A166  and  a21125a );
 a21127a <=( a21126a  and  a21121a );
 a21131a <=( A266  and  (not A265) );
 a21132a <=( (not A202)  and  a21131a );
 a21135a <=( (not A298)  and  A269 );
 a21138a <=( (not A301)  and  (not A299) );
 a21139a <=( a21138a  and  a21135a );
 a21140a <=( a21139a  and  a21132a );
 a21144a <=( A167  and  (not A168) );
 a21145a <=( (not A169)  and  a21144a );
 a21149a <=( (not A200)  and  (not A199) );
 a21150a <=( A166  and  a21149a );
 a21151a <=( a21150a  and  a21145a );
 a21155a <=( (not A266)  and  A265 );
 a21156a <=( (not A202)  and  a21155a );
 a21159a <=( (not A300)  and  A269 );
 a21162a <=( (not A302)  and  (not A301) );
 a21163a <=( a21162a  and  a21159a );
 a21164a <=( a21163a  and  a21156a );
 a21168a <=( A167  and  (not A168) );
 a21169a <=( (not A169)  and  a21168a );
 a21173a <=( (not A200)  and  (not A199) );
 a21174a <=( A166  and  a21173a );
 a21175a <=( a21174a  and  a21169a );
 a21179a <=( (not A266)  and  A265 );
 a21180a <=( (not A202)  and  a21179a );
 a21183a <=( (not A298)  and  A269 );
 a21186a <=( (not A301)  and  (not A299) );
 a21187a <=( a21186a  and  a21183a );
 a21188a <=( a21187a  and  a21180a );
 a21192a <=( (not A168)  and  (not A169) );
 a21193a <=( (not A170)  and  a21192a );
 a21197a <=( (not A203)  and  (not A202) );
 a21198a <=( (not A201)  and  a21197a );
 a21199a <=( a21198a  and  a21193a );
 a21203a <=( A269  and  A266 );
 a21204a <=( (not A265)  and  a21203a );
 a21207a <=( A299  and  A298 );
 a21210a <=( (not A301)  and  (not A300) );
 a21211a <=( a21210a  and  a21207a );
 a21212a <=( a21211a  and  a21204a );
 a21216a <=( (not A168)  and  (not A169) );
 a21217a <=( (not A170)  and  a21216a );
 a21221a <=( (not A203)  and  (not A202) );
 a21222a <=( (not A201)  and  a21221a );
 a21223a <=( a21222a  and  a21217a );
 a21227a <=( A269  and  (not A266) );
 a21228a <=( A265  and  a21227a );
 a21231a <=( A299  and  A298 );
 a21234a <=( (not A301)  and  (not A300) );
 a21235a <=( a21234a  and  a21231a );
 a21236a <=( a21235a  and  a21228a );
 a21240a <=( (not A168)  and  (not A169) );
 a21241a <=( (not A170)  and  a21240a );
 a21245a <=( (not A201)  and  A200 );
 a21246a <=( A199  and  a21245a );
 a21247a <=( a21246a  and  a21241a );
 a21251a <=( A267  and  A265 );
 a21252a <=( (not A202)  and  a21251a );
 a21255a <=( A299  and  A298 );
 a21258a <=( (not A301)  and  (not A300) );
 a21259a <=( a21258a  and  a21255a );
 a21260a <=( a21259a  and  a21252a );
 a21264a <=( (not A168)  and  (not A169) );
 a21265a <=( (not A170)  and  a21264a );
 a21269a <=( (not A201)  and  A200 );
 a21270a <=( A199  and  a21269a );
 a21271a <=( a21270a  and  a21265a );
 a21275a <=( A267  and  A266 );
 a21276a <=( (not A202)  and  a21275a );
 a21279a <=( A299  and  A298 );
 a21282a <=( (not A301)  and  (not A300) );
 a21283a <=( a21282a  and  a21279a );
 a21284a <=( a21283a  and  a21276a );
 a21288a <=( (not A168)  and  (not A169) );
 a21289a <=( (not A170)  and  a21288a );
 a21293a <=( (not A201)  and  A200 );
 a21294a <=( A199  and  a21293a );
 a21295a <=( a21294a  and  a21289a );
 a21299a <=( A266  and  (not A265) );
 a21300a <=( (not A202)  and  a21299a );
 a21303a <=( (not A300)  and  A269 );
 a21306a <=( (not A302)  and  (not A301) );
 a21307a <=( a21306a  and  a21303a );
 a21308a <=( a21307a  and  a21300a );
 a21312a <=( (not A168)  and  (not A169) );
 a21313a <=( (not A170)  and  a21312a );
 a21317a <=( (not A201)  and  A200 );
 a21318a <=( A199  and  a21317a );
 a21319a <=( a21318a  and  a21313a );
 a21323a <=( A266  and  (not A265) );
 a21324a <=( (not A202)  and  a21323a );
 a21327a <=( (not A298)  and  A269 );
 a21330a <=( (not A301)  and  (not A299) );
 a21331a <=( a21330a  and  a21327a );
 a21332a <=( a21331a  and  a21324a );
 a21336a <=( (not A168)  and  (not A169) );
 a21337a <=( (not A170)  and  a21336a );
 a21341a <=( (not A201)  and  A200 );
 a21342a <=( A199  and  a21341a );
 a21343a <=( a21342a  and  a21337a );
 a21347a <=( (not A266)  and  A265 );
 a21348a <=( (not A202)  and  a21347a );
 a21351a <=( (not A300)  and  A269 );
 a21354a <=( (not A302)  and  (not A301) );
 a21355a <=( a21354a  and  a21351a );
 a21356a <=( a21355a  and  a21348a );
 a21360a <=( (not A168)  and  (not A169) );
 a21361a <=( (not A170)  and  a21360a );
 a21365a <=( (not A201)  and  A200 );
 a21366a <=( A199  and  a21365a );
 a21367a <=( a21366a  and  a21361a );
 a21371a <=( (not A266)  and  A265 );
 a21372a <=( (not A202)  and  a21371a );
 a21375a <=( (not A298)  and  A269 );
 a21378a <=( (not A301)  and  (not A299) );
 a21379a <=( a21378a  and  a21375a );
 a21380a <=( a21379a  and  a21372a );
 a21384a <=( (not A168)  and  (not A169) );
 a21385a <=( (not A170)  and  a21384a );
 a21389a <=( A203  and  A200 );
 a21390a <=( (not A199)  and  a21389a );
 a21391a <=( a21390a  and  a21385a );
 a21395a <=( (not A267)  and  A266 );
 a21396a <=( A265  and  a21395a );
 a21399a <=( A298  and  (not A268) );
 a21402a <=( A302  and  (not A299) );
 a21403a <=( a21402a  and  a21399a );
 a21404a <=( a21403a  and  a21396a );
 a21408a <=( (not A168)  and  (not A169) );
 a21409a <=( (not A170)  and  a21408a );
 a21413a <=( A203  and  A200 );
 a21414a <=( (not A199)  and  a21413a );
 a21415a <=( a21414a  and  a21409a );
 a21419a <=( (not A267)  and  A266 );
 a21420a <=( A265  and  a21419a );
 a21423a <=( (not A298)  and  (not A268) );
 a21426a <=( A302  and  A299 );
 a21427a <=( a21426a  and  a21423a );
 a21428a <=( a21427a  and  a21420a );
 a21432a <=( (not A168)  and  (not A169) );
 a21433a <=( (not A170)  and  a21432a );
 a21437a <=( A203  and  (not A200) );
 a21438a <=( A199  and  a21437a );
 a21439a <=( a21438a  and  a21433a );
 a21443a <=( (not A267)  and  A266 );
 a21444a <=( A265  and  a21443a );
 a21447a <=( A298  and  (not A268) );
 a21450a <=( A302  and  (not A299) );
 a21451a <=( a21450a  and  a21447a );
 a21452a <=( a21451a  and  a21444a );
 a21456a <=( (not A168)  and  (not A169) );
 a21457a <=( (not A170)  and  a21456a );
 a21461a <=( A203  and  (not A200) );
 a21462a <=( A199  and  a21461a );
 a21463a <=( a21462a  and  a21457a );
 a21467a <=( (not A267)  and  A266 );
 a21468a <=( A265  and  a21467a );
 a21471a <=( (not A298)  and  (not A268) );
 a21474a <=( A302  and  A299 );
 a21475a <=( a21474a  and  a21471a );
 a21476a <=( a21475a  and  a21468a );
 a21480a <=( (not A168)  and  (not A169) );
 a21481a <=( (not A170)  and  a21480a );
 a21485a <=( (not A202)  and  (not A200) );
 a21486a <=( (not A199)  and  a21485a );
 a21487a <=( a21486a  and  a21481a );
 a21491a <=( A269  and  A266 );
 a21492a <=( (not A265)  and  a21491a );
 a21495a <=( A299  and  A298 );
 a21498a <=( (not A301)  and  (not A300) );
 a21499a <=( a21498a  and  a21495a );
 a21500a <=( a21499a  and  a21492a );
 a21504a <=( (not A168)  and  (not A169) );
 a21505a <=( (not A170)  and  a21504a );
 a21509a <=( (not A202)  and  (not A200) );
 a21510a <=( (not A199)  and  a21509a );
 a21511a <=( a21510a  and  a21505a );
 a21515a <=( A269  and  (not A266) );
 a21516a <=( A265  and  a21515a );
 a21519a <=( A299  and  A298 );
 a21522a <=( (not A301)  and  (not A300) );
 a21523a <=( a21522a  and  a21519a );
 a21524a <=( a21523a  and  a21516a );
 a21528a <=( (not A166)  and  A167 );
 a21529a <=( A170  and  a21528a );
 a21532a <=( A200  and  A199 );
 a21535a <=( (not A202)  and  (not A201) );
 a21536a <=( a21535a  and  a21532a );
 a21537a <=( a21536a  and  a21529a );
 a21541a <=( (not A267)  and  A266 );
 a21542a <=( A265  and  a21541a );
 a21545a <=( A298  and  (not A268) );
 a21548a <=( A302  and  (not A299) );
 a21549a <=( a21548a  and  a21545a );
 a21550a <=( a21549a  and  a21542a );
 a21554a <=( (not A166)  and  A167 );
 a21555a <=( A170  and  a21554a );
 a21558a <=( A200  and  A199 );
 a21561a <=( (not A202)  and  (not A201) );
 a21562a <=( a21561a  and  a21558a );
 a21563a <=( a21562a  and  a21555a );
 a21567a <=( (not A267)  and  A266 );
 a21568a <=( A265  and  a21567a );
 a21571a <=( (not A298)  and  (not A268) );
 a21574a <=( A302  and  A299 );
 a21575a <=( a21574a  and  a21571a );
 a21576a <=( a21575a  and  a21568a );
 a21580a <=( A166  and  (not A167) );
 a21581a <=( A170  and  a21580a );
 a21584a <=( A200  and  A199 );
 a21587a <=( (not A202)  and  (not A201) );
 a21588a <=( a21587a  and  a21584a );
 a21589a <=( a21588a  and  a21581a );
 a21593a <=( (not A267)  and  A266 );
 a21594a <=( A265  and  a21593a );
 a21597a <=( A298  and  (not A268) );
 a21600a <=( A302  and  (not A299) );
 a21601a <=( a21600a  and  a21597a );
 a21602a <=( a21601a  and  a21594a );
 a21606a <=( A166  and  (not A167) );
 a21607a <=( A170  and  a21606a );
 a21610a <=( A200  and  A199 );
 a21613a <=( (not A202)  and  (not A201) );
 a21614a <=( a21613a  and  a21610a );
 a21615a <=( a21614a  and  a21607a );
 a21619a <=( (not A267)  and  A266 );
 a21620a <=( A265  and  a21619a );
 a21623a <=( (not A298)  and  (not A268) );
 a21626a <=( A302  and  A299 );
 a21627a <=( a21626a  and  a21623a );
 a21628a <=( a21627a  and  a21620a );
 a21632a <=( (not A166)  and  (not A167) );
 a21633a <=( (not A169)  and  a21632a );
 a21636a <=( A200  and  A199 );
 a21639a <=( (not A202)  and  (not A201) );
 a21640a <=( a21639a  and  a21636a );
 a21641a <=( a21640a  and  a21633a );
 a21645a <=( A269  and  A266 );
 a21646a <=( (not A265)  and  a21645a );
 a21649a <=( A299  and  A298 );
 a21652a <=( (not A301)  and  (not A300) );
 a21653a <=( a21652a  and  a21649a );
 a21654a <=( a21653a  and  a21646a );
 a21658a <=( (not A166)  and  (not A167) );
 a21659a <=( (not A169)  and  a21658a );
 a21662a <=( A200  and  A199 );
 a21665a <=( (not A202)  and  (not A201) );
 a21666a <=( a21665a  and  a21662a );
 a21667a <=( a21666a  and  a21659a );
 a21671a <=( A269  and  (not A266) );
 a21672a <=( A265  and  a21671a );
 a21675a <=( A299  and  A298 );
 a21678a <=( (not A301)  and  (not A300) );
 a21679a <=( a21678a  and  a21675a );
 a21680a <=( a21679a  and  a21672a );
 a21684a <=( A167  and  (not A168) );
 a21685a <=( (not A169)  and  a21684a );
 a21688a <=( (not A201)  and  A166 );
 a21691a <=( (not A203)  and  (not A202) );
 a21692a <=( a21691a  and  a21688a );
 a21693a <=( a21692a  and  a21685a );
 a21697a <=( A269  and  A266 );
 a21698a <=( (not A265)  and  a21697a );
 a21701a <=( A299  and  A298 );
 a21704a <=( (not A301)  and  (not A300) );
 a21705a <=( a21704a  and  a21701a );
 a21706a <=( a21705a  and  a21698a );
 a21710a <=( A167  and  (not A168) );
 a21711a <=( (not A169)  and  a21710a );
 a21714a <=( (not A201)  and  A166 );
 a21717a <=( (not A203)  and  (not A202) );
 a21718a <=( a21717a  and  a21714a );
 a21719a <=( a21718a  and  a21711a );
 a21723a <=( A269  and  (not A266) );
 a21724a <=( A265  and  a21723a );
 a21727a <=( A299  and  A298 );
 a21730a <=( (not A301)  and  (not A300) );
 a21731a <=( a21730a  and  a21727a );
 a21732a <=( a21731a  and  a21724a );
 a21736a <=( A167  and  (not A168) );
 a21737a <=( (not A169)  and  a21736a );
 a21740a <=( A199  and  A166 );
 a21743a <=( (not A201)  and  A200 );
 a21744a <=( a21743a  and  a21740a );
 a21745a <=( a21744a  and  a21737a );
 a21749a <=( A267  and  A265 );
 a21750a <=( (not A202)  and  a21749a );
 a21753a <=( A299  and  A298 );
 a21756a <=( (not A301)  and  (not A300) );
 a21757a <=( a21756a  and  a21753a );
 a21758a <=( a21757a  and  a21750a );
 a21762a <=( A167  and  (not A168) );
 a21763a <=( (not A169)  and  a21762a );
 a21766a <=( A199  and  A166 );
 a21769a <=( (not A201)  and  A200 );
 a21770a <=( a21769a  and  a21766a );
 a21771a <=( a21770a  and  a21763a );
 a21775a <=( A267  and  A266 );
 a21776a <=( (not A202)  and  a21775a );
 a21779a <=( A299  and  A298 );
 a21782a <=( (not A301)  and  (not A300) );
 a21783a <=( a21782a  and  a21779a );
 a21784a <=( a21783a  and  a21776a );
 a21788a <=( A167  and  (not A168) );
 a21789a <=( (not A169)  and  a21788a );
 a21792a <=( A199  and  A166 );
 a21795a <=( (not A201)  and  A200 );
 a21796a <=( a21795a  and  a21792a );
 a21797a <=( a21796a  and  a21789a );
 a21801a <=( A266  and  (not A265) );
 a21802a <=( (not A202)  and  a21801a );
 a21805a <=( (not A300)  and  A269 );
 a21808a <=( (not A302)  and  (not A301) );
 a21809a <=( a21808a  and  a21805a );
 a21810a <=( a21809a  and  a21802a );
 a21814a <=( A167  and  (not A168) );
 a21815a <=( (not A169)  and  a21814a );
 a21818a <=( A199  and  A166 );
 a21821a <=( (not A201)  and  A200 );
 a21822a <=( a21821a  and  a21818a );
 a21823a <=( a21822a  and  a21815a );
 a21827a <=( A266  and  (not A265) );
 a21828a <=( (not A202)  and  a21827a );
 a21831a <=( (not A298)  and  A269 );
 a21834a <=( (not A301)  and  (not A299) );
 a21835a <=( a21834a  and  a21831a );
 a21836a <=( a21835a  and  a21828a );
 a21840a <=( A167  and  (not A168) );
 a21841a <=( (not A169)  and  a21840a );
 a21844a <=( A199  and  A166 );
 a21847a <=( (not A201)  and  A200 );
 a21848a <=( a21847a  and  a21844a );
 a21849a <=( a21848a  and  a21841a );
 a21853a <=( (not A266)  and  A265 );
 a21854a <=( (not A202)  and  a21853a );
 a21857a <=( (not A300)  and  A269 );
 a21860a <=( (not A302)  and  (not A301) );
 a21861a <=( a21860a  and  a21857a );
 a21862a <=( a21861a  and  a21854a );
 a21866a <=( A167  and  (not A168) );
 a21867a <=( (not A169)  and  a21866a );
 a21870a <=( A199  and  A166 );
 a21873a <=( (not A201)  and  A200 );
 a21874a <=( a21873a  and  a21870a );
 a21875a <=( a21874a  and  a21867a );
 a21879a <=( (not A266)  and  A265 );
 a21880a <=( (not A202)  and  a21879a );
 a21883a <=( (not A298)  and  A269 );
 a21886a <=( (not A301)  and  (not A299) );
 a21887a <=( a21886a  and  a21883a );
 a21888a <=( a21887a  and  a21880a );
 a21892a <=( A167  and  (not A168) );
 a21893a <=( (not A169)  and  a21892a );
 a21896a <=( (not A199)  and  A166 );
 a21899a <=( A203  and  A200 );
 a21900a <=( a21899a  and  a21896a );
 a21901a <=( a21900a  and  a21893a );
 a21905a <=( (not A267)  and  A266 );
 a21906a <=( A265  and  a21905a );
 a21909a <=( A298  and  (not A268) );
 a21912a <=( A302  and  (not A299) );
 a21913a <=( a21912a  and  a21909a );
 a21914a <=( a21913a  and  a21906a );
 a21918a <=( A167  and  (not A168) );
 a21919a <=( (not A169)  and  a21918a );
 a21922a <=( (not A199)  and  A166 );
 a21925a <=( A203  and  A200 );
 a21926a <=( a21925a  and  a21922a );
 a21927a <=( a21926a  and  a21919a );
 a21931a <=( (not A267)  and  A266 );
 a21932a <=( A265  and  a21931a );
 a21935a <=( (not A298)  and  (not A268) );
 a21938a <=( A302  and  A299 );
 a21939a <=( a21938a  and  a21935a );
 a21940a <=( a21939a  and  a21932a );
 a21944a <=( A167  and  (not A168) );
 a21945a <=( (not A169)  and  a21944a );
 a21948a <=( A199  and  A166 );
 a21951a <=( A203  and  (not A200) );
 a21952a <=( a21951a  and  a21948a );
 a21953a <=( a21952a  and  a21945a );
 a21957a <=( (not A267)  and  A266 );
 a21958a <=( A265  and  a21957a );
 a21961a <=( A298  and  (not A268) );
 a21964a <=( A302  and  (not A299) );
 a21965a <=( a21964a  and  a21961a );
 a21966a <=( a21965a  and  a21958a );
 a21970a <=( A167  and  (not A168) );
 a21971a <=( (not A169)  and  a21970a );
 a21974a <=( A199  and  A166 );
 a21977a <=( A203  and  (not A200) );
 a21978a <=( a21977a  and  a21974a );
 a21979a <=( a21978a  and  a21971a );
 a21983a <=( (not A267)  and  A266 );
 a21984a <=( A265  and  a21983a );
 a21987a <=( (not A298)  and  (not A268) );
 a21990a <=( A302  and  A299 );
 a21991a <=( a21990a  and  a21987a );
 a21992a <=( a21991a  and  a21984a );
 a21996a <=( A167  and  (not A168) );
 a21997a <=( (not A169)  and  a21996a );
 a22000a <=( (not A199)  and  A166 );
 a22003a <=( (not A202)  and  (not A200) );
 a22004a <=( a22003a  and  a22000a );
 a22005a <=( a22004a  and  a21997a );
 a22009a <=( A269  and  A266 );
 a22010a <=( (not A265)  and  a22009a );
 a22013a <=( A299  and  A298 );
 a22016a <=( (not A301)  and  (not A300) );
 a22017a <=( a22016a  and  a22013a );
 a22018a <=( a22017a  and  a22010a );
 a22022a <=( A167  and  (not A168) );
 a22023a <=( (not A169)  and  a22022a );
 a22026a <=( (not A199)  and  A166 );
 a22029a <=( (not A202)  and  (not A200) );
 a22030a <=( a22029a  and  a22026a );
 a22031a <=( a22030a  and  a22023a );
 a22035a <=( A269  and  (not A266) );
 a22036a <=( A265  and  a22035a );
 a22039a <=( A299  and  A298 );
 a22042a <=( (not A301)  and  (not A300) );
 a22043a <=( a22042a  and  a22039a );
 a22044a <=( a22043a  and  a22036a );
 a22048a <=( (not A168)  and  (not A169) );
 a22049a <=( (not A170)  and  a22048a );
 a22052a <=( A200  and  A199 );
 a22055a <=( (not A202)  and  (not A201) );
 a22056a <=( a22055a  and  a22052a );
 a22057a <=( a22056a  and  a22049a );
 a22061a <=( A269  and  A266 );
 a22062a <=( (not A265)  and  a22061a );
 a22065a <=( A299  and  A298 );
 a22068a <=( (not A301)  and  (not A300) );
 a22069a <=( a22068a  and  a22065a );
 a22070a <=( a22069a  and  a22062a );
 a22074a <=( (not A168)  and  (not A169) );
 a22075a <=( (not A170)  and  a22074a );
 a22078a <=( A200  and  A199 );
 a22081a <=( (not A202)  and  (not A201) );
 a22082a <=( a22081a  and  a22078a );
 a22083a <=( a22082a  and  a22075a );
 a22087a <=( A269  and  (not A266) );
 a22088a <=( A265  and  a22087a );
 a22091a <=( A299  and  A298 );
 a22094a <=( (not A301)  and  (not A300) );
 a22095a <=( a22094a  and  a22091a );
 a22096a <=( a22095a  and  a22088a );
 a22100a <=( A167  and  (not A168) );
 a22101a <=( (not A169)  and  a22100a );
 a22104a <=( A199  and  A166 );
 a22107a <=( (not A201)  and  A200 );
 a22108a <=( a22107a  and  a22104a );
 a22109a <=( a22108a  and  a22101a );
 a22112a <=( (not A265)  and  (not A202) );
 a22115a <=( A269  and  A266 );
 a22116a <=( a22115a  and  a22112a );
 a22119a <=( A299  and  A298 );
 a22122a <=( (not A301)  and  (not A300) );
 a22123a <=( a22122a  and  a22119a );
 a22124a <=( a22123a  and  a22116a );
 a22128a <=( A167  and  (not A168) );
 a22129a <=( (not A169)  and  a22128a );
 a22132a <=( A199  and  A166 );
 a22135a <=( (not A201)  and  A200 );
 a22136a <=( a22135a  and  a22132a );
 a22137a <=( a22136a  and  a22129a );
 a22140a <=( A265  and  (not A202) );
 a22143a <=( A269  and  (not A266) );
 a22144a <=( a22143a  and  a22140a );
 a22147a <=( A299  and  A298 );
 a22150a <=( (not A301)  and  (not A300) );
 a22151a <=( a22150a  and  a22147a );
 a22152a <=( a22151a  and  a22144a );


end x25_14x_behav;
