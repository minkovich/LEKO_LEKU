Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_3x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A140: buffer std_logic
);
end x25_3x;

architecture x25_3x_behav of x25_3x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a442a,a443a,a447a,a448a,a449a,a453a,a454a,a457a,a460a,a461a,a462a,a463a,a467a,a468a,a471a,a474a,a475a,a476a,a480a,a481a,a484a,a487a,a488a,a489a,a490a,a491a,a495a,a496a,a500a,a501a,a502a,a506a,a507a,a510a,a513a,a514a,a515a,a516a,a520a,a521a,a524a,a527a,a528a,a529a,a533a,a534a,a537a,a540a,a541a,a542a,a543a,a544a,a545a,a549a,a550a,a554a,a555a,a556a,a560a,a561a,a564a,a567a,a568a,a569a,a570a,a574a,a575a,a578a,a581a,a582a,a583a,a587a,a588a,a591a,a594a,a595a,a596a,a597a,a598a,a602a,a603a,a606a,a609a,a610a,a611a,a615a,a616a,a619a,a622a,a623a,a624a,a625a,a629a,a630a,a633a,a636a,a637a,a638a,a642a,a643a,a646a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a659a,a660a,a664a,a665a,a666a,a670a,a671a,a674a,a677a,a678a,a679a,a680a,a684a,a685a,a688a,a691a,a692a,a693a,a697a,a698a,a701a,a704a,a705a,a706a,a707a,a708a,a712a,a713a,a716a,a719a,a720a,a721a,a725a,a726a,a729a,a732a,a733a,a734a,a735a,a739a,a740a,a743a,a746a,a747a,a748a,a752a,a753a,a756a,a759a,a760a,a761a,a762a,a763a,a764a,a768a,a769a,a773a,a774a,a775a,a779a,a780a,a783a,a786a,a787a,a788a,a789a,a793a,a794a,a797a,a800a,a801a,a802a,a806a,a807a,a810a,a813a,a814a,a815a,a816a,a817a,a821a,a822a,a825a,a828a,a829a,a830a,a834a,a835a,a838a,a841a,a842a,a843a,a844a,a848a,a849a,a852a,a855a,a856a,a857a,a861a,a862a,a865a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a879a,a880a,a884a,a885a,a886a,a890a,a891a,a894a,a897a,a898a,a899a,a900a,a904a,a905a,a908a,a911a,a912a,a913a,a917a,a918a,a921a,a924a,a925a,a926a,a927a,a928a,a932a,a933a,a937a,a938a,a939a,a943a,a944a,a947a,a950a,a951a,a952a,a953a,a957a,a958a,a961a,a964a,a965a,a966a,a970a,a971a,a974a,a977a,a978a,a979a,a980a,a981a,a982a,a986a,a987a,a991a,a992a,a993a,a997a,a998a,a1001a,a1004a,a1005a,a1006a,a1007a,a1011a,a1012a,a1015a,a1018a,a1019a,a1020a,a1024a,a1025a,a1028a,a1031a,a1032a,a1033a,a1034a,a1035a,a1039a,a1040a,a1043a,a1046a,a1047a,a1048a,a1052a,a1053a,a1056a,a1059a,a1060a,a1061a,a1062a,a1066a,a1067a,a1070a,a1073a,a1074a,a1075a,a1079a,a1080a,a1083a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1096a,a1097a,a1101a,a1102a,a1103a,a1107a,a1108a,a1111a,a1114a,a1115a,a1116a,a1117a,a1121a,a1122a,a1125a,a1128a,a1129a,a1130a,a1134a,a1135a,a1138a,a1141a,a1142a,a1143a,a1144a,a1145a,a1149a,a1150a,a1153a,a1156a,a1157a,a1158a,a1162a,a1163a,a1166a,a1169a,a1170a,a1171a,a1172a,a1176a,a1177a,a1180a,a1183a,a1184a,a1185a,a1189a,a1190a,a1193a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1205a,a1206a,a1210a,a1211a,a1212a,a1216a,a1217a,a1220a,a1223a,a1224a,a1225a,a1226a,a1230a,a1231a,a1234a,a1237a,a1238a,a1239a,a1243a,a1244a,a1247a,a1250a,a1251a,a1252a,a1253a,a1254a,a1258a,a1259a,a1262a,a1265a,a1266a,a1267a,a1271a,a1272a,a1275a,a1278a,a1279a,a1280a,a1281a,a1285a,a1286a,a1289a,a1292a,a1293a,a1294a,a1298a,a1299a,a1302a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1315a,a1318a,a1321a,a1324a,a1327a,a1330a,a1333a,a1336a,a1339a,a1343a,a1344a,a1347a,a1351a,a1352a,a1355a,a1358a,a1359a,a1362a,a1365a,a1366a,a1369a,a1372a,a1373a,a1376a,a1379a,a1380a,a1383a,a1386a,a1387a,a1390a,a1393a,a1394a,a1397a,a1400a,a1401a,a1404a,a1407a,a1408a,a1411a,a1414a,a1415a,a1418a,a1421a,a1422a,a1425a,a1428a,a1429a,a1432a,a1435a,a1436a,a1439a,a1442a,a1443a,a1446a,a1449a,a1450a,a1453a,a1456a,a1457a,a1460a,a1463a,a1464a,a1467a,a1470a,a1471a,a1474a,a1477a,a1478a,a1481a,a1484a,a1485a,a1488a,a1491a,a1492a,a1495a,a1498a,a1499a,a1502a,a1505a,a1506a,a1509a,a1512a,a1513a,a1516a,a1519a,a1520a,a1523a,a1526a,a1527a,a1530a,a1533a,a1534a,a1537a,a1540a,a1541a,a1544a,a1547a,a1548a,a1551a,a1554a,a1555a,a1558a,a1561a,a1562a,a1565a,a1568a,a1569a,a1572a,a1575a,a1576a,a1579a,a1582a,a1583a,a1586a,a1589a,a1590a,a1593a,a1596a,a1597a,a1600a,a1603a,a1604a,a1607a,a1610a,a1611a,a1614a,a1617a,a1618a,a1621a,a1624a,a1625a,a1628a,a1631a,a1632a,a1635a,a1638a,a1639a,a1642a,a1645a,a1646a,a1649a,a1652a,a1653a,a1656a,a1659a,a1660a,a1663a,a1666a,a1667a,a1670a,a1673a,a1674a,a1677a,a1680a,a1681a,a1684a,a1687a,a1688a,a1691a,a1694a,a1695a,a1698a,a1701a,a1702a,a1705a,a1708a,a1709a,a1712a,a1715a,a1716a,a1719a,a1722a,a1723a,a1726a,a1729a,a1730a,a1733a,a1736a,a1737a,a1740a,a1743a,a1744a,a1747a,a1750a,a1751a,a1754a,a1757a,a1758a,a1761a,a1764a,a1765a,a1768a,a1771a,a1772a,a1775a,a1778a,a1779a,a1782a,a1785a,a1786a,a1789a,a1792a,a1793a,a1796a,a1799a,a1800a,a1803a,a1806a,a1807a,a1810a,a1814a,a1815a,a1816a,a1819a,a1822a,a1823a,a1826a,a1830a,a1831a,a1832a,a1835a,a1838a,a1839a,a1842a,a1846a,a1847a,a1848a,a1851a,a1854a,a1855a,a1858a,a1862a,a1863a,a1864a,a1867a,a1870a,a1871a,a1874a,a1878a,a1879a,a1880a,a1883a,a1886a,a1887a,a1890a,a1894a,a1895a,a1896a,a1899a,a1902a,a1903a,a1906a,a1910a,a1911a,a1912a,a1915a,a1918a,a1919a,a1922a,a1926a,a1927a,a1928a,a1931a,a1934a,a1935a,a1938a,a1942a,a1943a,a1944a,a1947a,a1950a,a1951a,a1954a,a1958a,a1959a,a1960a,a1963a,a1966a,a1967a,a1970a,a1974a,a1975a,a1976a,a1979a,a1982a,a1983a,a1986a,a1990a,a1991a,a1992a,a1995a,a1998a,a1999a,a2002a,a2006a,a2007a,a2008a,a2011a,a2014a,a2015a,a2018a,a2022a,a2023a,a2024a,a2027a,a2030a,a2031a,a2034a,a2038a,a2039a,a2040a,a2043a,a2046a,a2047a,a2050a,a2054a,a2055a,a2056a,a2059a,a2062a,a2063a,a2066a,a2070a,a2071a,a2072a,a2075a,a2078a,a2079a,a2082a,a2086a,a2087a,a2088a,a2091a,a2094a,a2095a,a2098a,a2102a,a2103a,a2104a,a2107a,a2110a,a2111a,a2114a,a2118a,a2119a,a2120a,a2123a,a2126a,a2127a,a2130a,a2134a,a2135a,a2136a,a2139a,a2142a,a2143a,a2146a,a2150a,a2151a,a2152a,a2155a,a2158a,a2159a,a2162a,a2166a,a2167a,a2168a,a2171a,a2174a,a2175a,a2178a,a2182a,a2183a,a2184a,a2187a,a2190a,a2191a,a2194a,a2198a,a2199a,a2200a,a2203a,a2206a,a2207a,a2210a,a2214a,a2215a,a2216a,a2219a,a2222a,a2223a,a2226a,a2230a,a2231a,a2232a,a2235a,a2238a,a2239a,a2242a,a2246a,a2247a,a2248a,a2251a,a2254a,a2255a,a2258a,a2262a,a2263a,a2264a,a2267a,a2270a,a2271a,a2274a,a2278a,a2279a,a2280a,a2283a,a2286a,a2287a,a2290a,a2294a,a2295a,a2296a,a2299a,a2302a,a2303a,a2306a,a2310a,a2311a,a2312a,a2315a,a2319a,a2320a,a2321a,a2324a,a2328a,a2329a,a2330a,a2333a,a2337a,a2338a,a2339a,a2342a,a2346a,a2347a,a2348a,a2351a,a2355a,a2356a,a2357a,a2360a,a2364a,a2365a,a2366a,a2369a,a2373a,a2374a,a2375a,a2378a,a2382a,a2383a,a2384a,a2387a,a2391a,a2392a,a2393a,a2396a,a2400a,a2401a,a2402a,a2405a,a2409a,a2410a,a2411a,a2414a,a2418a,a2419a,a2420a,a2423a,a2427a,a2428a,a2429a,a2432a,a2436a,a2437a,a2438a,a2441a,a2445a,a2446a,a2447a,a2450a,a2454a,a2455a,a2456a,a2459a,a2463a,a2464a,a2465a,a2468a,a2472a,a2473a,a2474a,a2477a,a2481a,a2482a,a2483a,a2486a,a2490a,a2491a,a2492a,a2495a,a2499a,a2500a,a2501a,a2504a,a2508a,a2509a,a2510a,a2513a,a2517a,a2518a,a2519a,a2522a,a2526a,a2527a,a2528a,a2531a,a2535a,a2536a,a2537a,a2540a,a2544a,a2545a,a2546a,a2549a,a2553a,a2554a,a2555a,a2558a,a2562a,a2563a,a2564a,a2567a,a2571a,a2572a,a2573a,a2576a,a2580a,a2581a,a2582a,a2585a,a2589a,a2590a,a2591a,a2594a,a2598a,a2599a,a2600a,a2603a,a2607a,a2608a,a2609a,a2612a,a2616a,a2617a,a2618a,a2621a,a2625a,a2626a,a2627a,a2630a,a2634a,a2635a,a2636a,a2639a,a2643a,a2644a,a2645a,a2648a,a2652a,a2653a,a2654a,a2657a,a2661a,a2662a,a2663a,a2666a,a2670a,a2671a,a2672a,a2675a,a2679a,a2680a,a2681a,a2684a,a2688a,a2689a,a2690a,a2693a,a2697a,a2698a,a2699a,a2702a,a2706a,a2707a,a2708a,a2711a,a2715a,a2716a,a2717a,a2720a,a2724a,a2725a,a2726a,a2729a,a2733a,a2734a,a2735a,a2738a,a2742a,a2743a,a2744a,a2747a,a2751a,a2752a,a2753a,a2756a,a2760a,a2761a,a2762a,a2765a,a2769a,a2770a,a2771a,a2774a,a2778a,a2779a,a2780a,a2783a,a2787a,a2788a,a2789a,a2792a,a2796a,a2797a,a2798a,a2801a,a2805a,a2806a,a2807a,a2810a,a2814a,a2815a,a2816a,a2819a,a2823a,a2824a,a2825a,a2828a,a2832a,a2833a,a2834a,a2837a,a2841a,a2842a,a2843a,a2846a,a2850a,a2851a,a2852a,a2855a,a2859a,a2860a,a2861a,a2864a,a2868a,a2869a,a2870a,a2873a,a2877a,a2878a,a2879a,a2882a,a2886a,a2887a,a2888a,a2891a,a2895a,a2896a,a2897a,a2900a,a2904a,a2905a,a2906a,a2909a,a2913a,a2914a,a2915a,a2918a,a2922a,a2923a,a2924a,a2927a,a2931a,a2932a,a2933a,a2936a,a2940a,a2941a,a2942a,a2945a,a2949a,a2950a,a2951a,a2954a,a2958a,a2959a,a2960a,a2963a,a2967a,a2968a,a2969a,a2972a,a2976a,a2977a,a2978a,a2981a,a2985a,a2986a,a2987a,a2990a,a2994a,a2995a,a2996a,a2999a,a3003a,a3004a,a3005a,a3008a,a3012a,a3013a,a3014a,a3017a,a3021a,a3022a,a3023a,a3026a,a3030a,a3031a,a3032a,a3035a,a3039a,a3040a,a3041a,a3044a,a3048a,a3049a,a3050a,a3053a,a3057a,a3058a,a3059a,a3062a,a3066a,a3067a,a3068a,a3071a,a3075a,a3076a,a3077a,a3080a,a3084a,a3085a,a3086a,a3089a,a3093a,a3094a,a3095a,a3098a,a3102a,a3103a,a3104a,a3107a,a3111a,a3112a,a3113a,a3116a,a3120a,a3121a,a3122a,a3125a,a3129a,a3130a,a3131a,a3134a,a3138a,a3139a,a3140a,a3143a,a3147a,a3148a,a3149a,a3152a,a3156a,a3157a,a3158a,a3161a,a3165a,a3166a,a3167a,a3170a,a3174a,a3175a,a3176a,a3179a,a3183a,a3184a,a3185a,a3188a,a3192a,a3193a,a3194a,a3197a,a3201a,a3202a,a3203a,a3206a,a3210a,a3211a,a3212a,a3215a,a3219a,a3220a,a3221a,a3224a,a3228a,a3229a,a3230a,a3233a,a3237a,a3238a,a3239a,a3242a,a3246a,a3247a,a3248a,a3251a,a3255a,a3256a,a3257a,a3260a,a3264a,a3265a,a3266a,a3269a,a3273a,a3274a,a3275a,a3278a,a3282a,a3283a,a3284a,a3287a,a3291a,a3292a,a3293a,a3296a,a3300a,a3301a,a3302a,a3305a,a3309a,a3310a,a3311a,a3314a,a3318a,a3319a,a3320a,a3323a,a3327a,a3328a,a3329a,a3332a,a3336a,a3337a,a3338a,a3341a,a3345a,a3346a,a3347a,a3350a,a3354a,a3355a,a3356a,a3359a,a3363a,a3364a,a3365a,a3368a,a3372a,a3373a,a3374a,a3377a,a3381a,a3382a,a3383a,a3386a,a3390a,a3391a,a3392a,a3395a,a3399a,a3400a,a3401a,a3404a,a3408a,a3409a,a3410a,a3413a,a3417a,a3418a,a3419a,a3422a,a3426a,a3427a,a3428a,a3431a,a3435a,a3436a,a3437a,a3440a,a3444a,a3445a,a3446a,a3449a,a3453a,a3454a,a3455a,a3458a,a3462a,a3463a,a3464a,a3467a,a3471a,a3472a,a3473a,a3476a,a3480a,a3481a,a3482a,a3485a,a3489a,a3490a,a3491a,a3494a,a3498a,a3499a,a3500a,a3503a,a3507a,a3508a,a3509a,a3512a,a3516a,a3517a,a3518a,a3521a,a3525a,a3526a,a3527a,a3530a,a3534a,a3535a,a3536a,a3539a,a3543a,a3544a,a3545a,a3548a,a3552a,a3553a,a3554a,a3557a,a3561a,a3562a,a3563a,a3566a,a3570a,a3571a,a3572a,a3575a,a3579a,a3580a,a3581a,a3584a,a3588a,a3589a,a3590a,a3593a,a3597a,a3598a,a3599a,a3602a,a3606a,a3607a,a3608a,a3611a,a3615a,a3616a,a3617a,a3620a,a3624a,a3625a,a3626a,a3629a,a3633a,a3634a,a3635a,a3638a,a3642a,a3643a,a3644a,a3647a,a3651a,a3652a,a3653a,a3656a,a3660a,a3661a,a3662a,a3665a,a3669a,a3670a,a3671a,a3674a,a3678a,a3679a,a3680a,a3683a,a3687a,a3688a,a3689a,a3692a,a3696a,a3697a,a3698a,a3701a,a3705a,a3706a,a3707a,a3710a,a3714a,a3715a,a3716a,a3719a,a3723a,a3724a,a3725a,a3728a,a3732a,a3733a,a3734a,a3737a,a3741a,a3742a,a3743a,a3746a,a3750a,a3751a,a3752a,a3755a,a3759a,a3760a,a3761a,a3764a,a3768a,a3769a,a3770a,a3773a,a3777a,a3778a,a3779a,a3782a,a3786a,a3787a,a3788a,a3791a,a3795a,a3796a,a3797a,a3800a,a3804a,a3805a,a3806a,a3809a,a3813a,a3814a,a3815a,a3818a,a3822a,a3823a,a3824a,a3827a,a3831a,a3832a,a3833a,a3836a,a3840a,a3841a,a3842a,a3845a,a3849a,a3850a,a3851a,a3854a,a3858a,a3859a,a3860a,a3863a,a3867a,a3868a,a3869a,a3872a,a3876a,a3877a,a3878a,a3881a,a3885a,a3886a,a3887a,a3890a,a3894a,a3895a,a3896a,a3899a,a3903a,a3904a,a3905a,a3908a,a3912a,a3913a,a3914a,a3917a,a3921a,a3922a,a3923a,a3926a,a3930a,a3931a,a3932a,a3935a,a3939a,a3940a,a3941a,a3944a,a3948a,a3949a,a3950a,a3953a,a3957a,a3958a,a3959a,a3962a,a3966a,a3967a,a3968a,a3971a,a3975a,a3976a,a3977a,a3980a,a3984a,a3985a,a3986a,a3989a,a3993a,a3994a,a3995a,a3998a,a4002a,a4003a,a4004a,a4007a,a4011a,a4012a,a4013a,a4016a,a4020a,a4021a,a4022a,a4025a,a4029a,a4030a,a4031a,a4034a,a4038a,a4039a,a4040a,a4043a,a4047a,a4048a,a4049a,a4052a,a4056a,a4057a,a4058a,a4061a,a4065a,a4066a,a4067a,a4070a,a4074a,a4075a,a4076a,a4079a,a4083a,a4084a,a4085a,a4088a,a4092a,a4093a,a4094a,a4097a,a4101a,a4102a,a4103a,a4106a,a4110a,a4111a,a4112a,a4115a,a4119a,a4120a,a4121a,a4124a,a4128a,a4129a,a4130a,a4133a,a4137a,a4138a,a4139a,a4142a,a4146a,a4147a,a4148a,a4151a,a4155a,a4156a,a4157a,a4160a,a4164a,a4165a,a4166a,a4169a,a4173a,a4174a,a4175a,a4178a,a4182a,a4183a,a4184a,a4187a,a4191a,a4192a,a4193a,a4196a,a4200a,a4201a,a4202a,a4205a,a4209a,a4210a,a4211a,a4214a,a4218a,a4219a,a4220a,a4223a,a4227a,a4228a,a4229a,a4232a,a4236a,a4237a,a4238a,a4241a,a4245a,a4246a,a4247a,a4250a,a4254a,a4255a,a4256a,a4259a,a4263a,a4264a,a4265a,a4268a,a4272a,a4273a,a4274a,a4277a,a4281a,a4282a,a4283a,a4286a,a4290a,a4291a,a4292a,a4295a,a4299a,a4300a,a4301a,a4304a,a4308a,a4309a,a4310a,a4313a,a4317a,a4318a,a4319a,a4322a,a4326a,a4327a,a4328a,a4331a,a4335a,a4336a,a4337a,a4340a,a4344a,a4345a,a4346a,a4349a,a4353a,a4354a,a4355a,a4358a,a4362a,a4363a,a4364a,a4367a,a4371a,a4372a,a4373a,a4376a,a4380a,a4381a,a4382a,a4385a,a4389a,a4390a,a4391a,a4394a,a4398a,a4399a,a4400a,a4403a,a4407a,a4408a,a4409a,a4412a,a4416a,a4417a,a4418a,a4421a,a4425a,a4426a,a4427a,a4430a,a4434a,a4435a,a4436a,a4439a,a4443a,a4444a,a4445a,a4448a,a4452a,a4453a,a4454a,a4457a,a4461a,a4462a,a4463a,a4466a,a4470a,a4471a,a4472a,a4475a,a4479a,a4480a,a4481a,a4484a,a4488a,a4489a,a4490a,a4493a,a4497a,a4498a,a4499a,a4502a,a4506a,a4507a,a4508a,a4511a,a4515a,a4516a,a4517a,a4520a,a4524a,a4525a,a4526a,a4529a,a4533a,a4534a,a4535a,a4538a,a4542a,a4543a,a4544a,a4547a,a4551a,a4552a,a4553a,a4556a,a4560a,a4561a,a4562a,a4565a,a4569a,a4570a,a4571a,a4574a,a4578a,a4579a,a4580a,a4583a,a4587a,a4588a,a4589a,a4592a,a4596a,a4597a,a4598a,a4601a,a4605a,a4606a,a4607a,a4610a,a4614a,a4615a,a4616a,a4619a,a4623a,a4624a,a4625a,a4628a,a4632a,a4633a,a4634a,a4637a,a4641a,a4642a,a4643a,a4646a,a4650a,a4651a,a4652a,a4655a,a4659a,a4660a,a4661a,a4664a,a4668a,a4669a,a4670a,a4673a,a4677a,a4678a,a4679a,a4682a,a4686a,a4687a,a4688a,a4691a,a4695a,a4696a,a4697a,a4700a,a4704a,a4705a,a4706a,a4709a,a4713a,a4714a,a4715a,a4718a,a4722a,a4723a,a4724a,a4727a,a4731a,a4732a,a4733a,a4736a,a4740a,a4741a,a4742a,a4745a,a4749a,a4750a,a4751a,a4754a,a4758a,a4759a,a4760a,a4763a,a4767a,a4768a,a4769a,a4773a,a4774a,a4778a,a4779a,a4780a,a4783a,a4787a,a4788a,a4789a,a4793a,a4794a,a4798a,a4799a,a4800a,a4803a,a4807a,a4808a,a4809a,a4813a,a4814a,a4818a,a4819a,a4820a,a4823a,a4827a,a4828a,a4829a,a4833a,a4834a,a4838a,a4839a,a4840a,a4843a,a4847a,a4848a,a4849a,a4853a,a4854a,a4858a,a4859a,a4860a,a4863a,a4867a,a4868a,a4869a,a4873a,a4874a,a4878a,a4879a,a4880a,a4883a,a4887a,a4888a,a4889a,a4893a,a4894a,a4898a,a4899a,a4900a,a4903a,a4907a,a4908a,a4909a,a4913a,a4914a,a4918a,a4919a,a4920a,a4923a,a4927a,a4928a,a4929a,a4933a,a4934a,a4938a,a4939a,a4940a,a4943a,a4947a,a4948a,a4949a,a4953a,a4954a,a4958a,a4959a,a4960a,a4963a,a4967a,a4968a,a4969a,a4973a,a4974a,a4978a,a4979a,a4980a,a4983a,a4987a,a4988a,a4989a,a4993a,a4994a,a4998a,a4999a,a5000a,a5003a,a5007a,a5008a,a5009a,a5013a,a5014a,a5018a,a5019a,a5020a,a5023a,a5027a,a5028a,a5029a,a5033a,a5034a,a5038a,a5039a,a5040a,a5043a,a5047a,a5048a,a5049a,a5053a,a5054a,a5058a,a5059a,a5060a,a5063a,a5067a,a5068a,a5069a,a5073a,a5074a,a5078a,a5079a,a5080a,a5083a,a5087a,a5088a,a5089a,a5093a,a5094a,a5098a,a5099a,a5100a,a5103a,a5107a,a5108a,a5109a,a5113a,a5114a,a5118a,a5119a,a5120a,a5123a,a5127a,a5128a,a5129a,a5133a,a5134a,a5138a,a5139a,a5140a,a5143a,a5147a,a5148a,a5149a,a5153a,a5154a,a5158a,a5159a,a5160a,a5163a,a5167a,a5168a,a5169a,a5173a,a5174a,a5178a,a5179a,a5180a,a5183a,a5187a,a5188a,a5189a,a5193a,a5194a,a5198a,a5199a,a5200a,a5203a,a5207a,a5208a,a5209a,a5213a,a5214a,a5218a,a5219a,a5220a,a5223a,a5227a,a5228a,a5229a,a5233a,a5234a,a5238a,a5239a,a5240a,a5243a,a5247a,a5248a,a5249a,a5253a,a5254a,a5258a,a5259a,a5260a,a5263a,a5267a,a5268a,a5269a,a5273a,a5274a,a5278a,a5279a,a5280a,a5283a,a5287a,a5288a,a5289a,a5293a,a5294a,a5298a,a5299a,a5300a,a5303a,a5307a,a5308a,a5309a,a5313a,a5314a,a5318a,a5319a,a5320a,a5323a,a5327a,a5328a,a5329a,a5333a,a5334a,a5338a,a5339a,a5340a,a5343a,a5347a,a5348a,a5349a,a5353a,a5354a,a5358a,a5359a,a5360a,a5363a,a5367a,a5368a,a5369a,a5373a,a5374a,a5378a,a5379a,a5380a,a5383a,a5387a,a5388a,a5389a,a5393a,a5394a,a5398a,a5399a,a5400a,a5403a,a5407a,a5408a,a5409a,a5413a,a5414a,a5418a,a5419a,a5420a,a5423a,a5427a,a5428a,a5429a,a5433a,a5434a,a5438a,a5439a,a5440a,a5443a,a5447a,a5448a,a5449a,a5453a,a5454a,a5458a,a5459a,a5460a,a5463a,a5467a,a5468a,a5469a,a5473a,a5474a,a5478a,a5479a,a5480a,a5483a,a5487a,a5488a,a5489a,a5493a,a5494a,a5498a,a5499a,a5500a,a5503a,a5507a,a5508a,a5509a,a5513a,a5514a,a5518a,a5519a,a5520a,a5523a,a5527a,a5528a,a5529a,a5533a,a5534a,a5538a,a5539a,a5540a,a5543a,a5547a,a5548a,a5549a,a5553a,a5554a,a5558a,a5559a,a5560a,a5563a,a5567a,a5568a,a5569a,a5573a,a5574a,a5578a,a5579a,a5580a,a5583a,a5587a,a5588a,a5589a,a5593a,a5594a,a5598a,a5599a,a5600a,a5603a,a5607a,a5608a,a5609a,a5613a,a5614a,a5618a,a5619a,a5620a,a5623a,a5627a,a5628a,a5629a,a5633a,a5634a,a5638a,a5639a,a5640a,a5643a,a5647a,a5648a,a5649a,a5653a,a5654a,a5658a,a5659a,a5660a,a5663a,a5667a,a5668a,a5669a,a5673a,a5674a,a5678a,a5679a,a5680a,a5683a,a5687a,a5688a,a5689a,a5693a,a5694a,a5698a,a5699a,a5700a,a5703a,a5707a,a5708a,a5709a,a5713a,a5714a,a5718a,a5719a,a5720a,a5723a,a5727a,a5728a,a5729a,a5733a,a5734a,a5738a,a5739a,a5740a,a5743a,a5747a,a5748a,a5749a,a5753a,a5754a,a5758a,a5759a,a5760a,a5763a,a5767a,a5768a,a5769a,a5773a,a5774a,a5778a,a5779a,a5780a,a5783a,a5787a,a5788a,a5789a,a5793a,a5794a,a5798a,a5799a,a5800a,a5803a,a5807a,a5808a,a5809a,a5813a,a5814a,a5818a,a5819a,a5820a,a5823a,a5827a,a5828a,a5829a,a5833a,a5834a,a5838a,a5839a,a5840a,a5843a,a5847a,a5848a,a5849a,a5853a,a5854a,a5858a,a5859a,a5860a,a5863a,a5867a,a5868a,a5869a,a5873a,a5874a,a5878a,a5879a,a5880a,a5883a,a5887a,a5888a,a5889a,a5893a,a5894a,a5898a,a5899a,a5900a,a5903a,a5907a,a5908a,a5909a,a5913a,a5914a,a5918a,a5919a,a5920a,a5923a,a5927a,a5928a,a5929a,a5933a,a5934a,a5938a,a5939a,a5940a,a5943a,a5947a,a5948a,a5949a,a5953a,a5954a,a5958a,a5959a,a5960a,a5963a,a5967a,a5968a,a5969a,a5973a,a5974a,a5978a,a5979a,a5980a,a5983a,a5987a,a5988a,a5989a,a5993a,a5994a,a5998a,a5999a,a6000a,a6003a,a6007a,a6008a,a6009a,a6013a,a6014a,a6018a,a6019a,a6020a,a6023a,a6027a,a6028a,a6029a,a6033a,a6034a,a6038a,a6039a,a6040a,a6043a,a6047a,a6048a,a6049a,a6053a,a6054a,a6058a,a6059a,a6060a,a6063a,a6067a,a6068a,a6069a,a6073a,a6074a,a6078a,a6079a,a6080a,a6083a,a6087a,a6088a,a6089a,a6093a,a6094a,a6098a,a6099a,a6100a,a6103a,a6107a,a6108a,a6109a,a6113a,a6114a,a6118a,a6119a,a6120a,a6123a,a6127a,a6128a,a6129a,a6133a,a6134a,a6138a,a6139a,a6140a,a6143a,a6147a,a6148a,a6149a,a6153a,a6154a,a6158a,a6159a,a6160a,a6163a,a6167a,a6168a,a6169a,a6173a,a6174a,a6178a,a6179a,a6180a,a6183a,a6187a,a6188a,a6189a,a6193a,a6194a,a6198a,a6199a,a6200a,a6203a,a6207a,a6208a,a6209a,a6213a,a6214a,a6218a,a6219a,a6220a,a6223a,a6227a,a6228a,a6229a,a6233a,a6234a,a6238a,a6239a,a6240a,a6243a,a6247a,a6248a,a6249a,a6253a,a6254a,a6258a,a6259a,a6260a,a6263a,a6267a,a6268a,a6269a,a6273a,a6274a,a6278a,a6279a,a6280a,a6283a,a6287a,a6288a,a6289a,a6293a,a6294a,a6298a,a6299a,a6300a,a6303a,a6307a,a6308a,a6309a,a6313a,a6314a,a6318a,a6319a,a6320a,a6323a,a6327a,a6328a,a6329a,a6333a,a6334a,a6338a,a6339a,a6340a,a6343a,a6347a,a6348a,a6349a,a6353a,a6354a,a6358a,a6359a,a6360a,a6363a,a6367a,a6368a,a6369a,a6373a,a6374a,a6378a,a6379a,a6380a,a6383a,a6387a,a6388a,a6389a,a6393a,a6394a,a6398a,a6399a,a6400a,a6403a,a6407a,a6408a,a6409a,a6413a,a6414a,a6418a,a6419a,a6420a,a6423a,a6427a,a6428a,a6429a,a6433a,a6434a,a6438a,a6439a,a6440a,a6443a,a6447a,a6448a,a6449a,a6453a,a6454a,a6458a,a6459a,a6460a,a6463a,a6467a,a6468a,a6469a,a6473a,a6474a,a6478a,a6479a,a6480a,a6483a,a6487a,a6488a,a6489a,a6493a,a6494a,a6498a,a6499a,a6500a,a6503a,a6507a,a6508a,a6509a,a6513a,a6514a,a6518a,a6519a,a6520a,a6523a,a6527a,a6528a,a6529a,a6533a,a6534a,a6538a,a6539a,a6540a,a6543a,a6547a,a6548a,a6549a,a6553a,a6554a,a6558a,a6559a,a6560a,a6563a,a6567a,a6568a,a6569a,a6573a,a6574a,a6578a,a6579a,a6580a,a6583a,a6587a,a6588a,a6589a,a6593a,a6594a,a6598a,a6599a,a6600a,a6603a,a6607a,a6608a,a6609a,a6613a,a6614a,a6618a,a6619a,a6620a,a6623a,a6627a,a6628a,a6629a,a6633a,a6634a,a6638a,a6639a,a6640a,a6643a,a6647a,a6648a,a6649a,a6653a,a6654a,a6658a,a6659a,a6660a,a6663a,a6667a,a6668a,a6669a,a6673a,a6674a,a6678a,a6679a,a6680a,a6683a,a6687a,a6688a,a6689a,a6693a,a6694a,a6698a,a6699a,a6700a,a6703a,a6707a,a6708a,a6709a,a6713a,a6714a,a6718a,a6719a,a6720a,a6723a,a6727a,a6728a,a6729a,a6733a,a6734a,a6738a,a6739a,a6740a,a6743a,a6747a,a6748a,a6749a,a6753a,a6754a,a6758a,a6759a,a6760a,a6763a,a6767a,a6768a,a6769a,a6773a,a6774a,a6778a,a6779a,a6780a,a6783a,a6787a,a6788a,a6789a,a6793a,a6794a,a6798a,a6799a,a6800a,a6803a,a6807a,a6808a,a6809a,a6813a,a6814a,a6818a,a6819a,a6820a,a6823a,a6827a,a6828a,a6829a,a6833a,a6834a,a6838a,a6839a,a6840a,a6843a,a6847a,a6848a,a6849a,a6853a,a6854a,a6858a,a6859a,a6860a,a6863a,a6867a,a6868a,a6869a,a6873a,a6874a,a6878a,a6879a,a6880a,a6883a,a6887a,a6888a,a6889a,a6893a,a6894a,a6898a,a6899a,a6900a,a6903a,a6907a,a6908a,a6909a,a6913a,a6914a,a6918a,a6919a,a6920a,a6923a,a6927a,a6928a,a6929a,a6933a,a6934a,a6938a,a6939a,a6940a,a6943a,a6947a,a6948a,a6949a,a6953a,a6954a,a6958a,a6959a,a6960a,a6963a,a6967a,a6968a,a6969a,a6973a,a6974a,a6978a,a6979a,a6980a,a6983a,a6987a,a6988a,a6989a,a6993a,a6994a,a6998a,a6999a,a7000a,a7003a,a7007a,a7008a,a7009a,a7013a,a7014a,a7018a,a7019a,a7020a,a7023a,a7027a,a7028a,a7029a,a7033a,a7034a,a7038a,a7039a,a7040a,a7043a,a7047a,a7048a,a7049a,a7053a,a7054a,a7058a,a7059a,a7060a,a7063a,a7067a,a7068a,a7069a,a7073a,a7074a,a7078a,a7079a,a7080a,a7083a,a7087a,a7088a,a7089a,a7093a,a7094a,a7098a,a7099a,a7100a,a7103a,a7107a,a7108a,a7109a,a7113a,a7114a,a7118a,a7119a,a7120a,a7123a,a7127a,a7128a,a7129a,a7133a,a7134a,a7138a,a7139a,a7140a,a7143a,a7147a,a7148a,a7149a,a7153a,a7154a,a7158a,a7159a,a7160a,a7163a,a7167a,a7168a,a7169a,a7173a,a7174a,a7178a,a7179a,a7180a,a7183a,a7187a,a7188a,a7189a,a7193a,a7194a,a7198a,a7199a,a7200a,a7203a,a7207a,a7208a,a7209a,a7213a,a7214a,a7218a,a7219a,a7220a,a7223a,a7227a,a7228a,a7229a,a7233a,a7234a,a7238a,a7239a,a7240a,a7243a,a7247a,a7248a,a7249a,a7253a,a7254a,a7258a,a7259a,a7260a,a7263a,a7267a,a7268a,a7269a,a7273a,a7274a,a7278a,a7279a,a7280a,a7283a,a7287a,a7288a,a7289a,a7293a,a7294a,a7298a,a7299a,a7300a,a7303a,a7307a,a7308a,a7309a,a7313a,a7314a,a7318a,a7319a,a7320a,a7323a,a7327a,a7328a,a7329a,a7333a,a7334a,a7338a,a7339a,a7340a,a7343a,a7347a,a7348a,a7349a,a7353a,a7354a,a7358a,a7359a,a7360a,a7363a,a7367a,a7368a,a7369a,a7373a,a7374a,a7378a,a7379a,a7380a,a7383a,a7387a,a7388a,a7389a,a7393a,a7394a,a7398a,a7399a,a7400a,a7403a,a7407a,a7408a,a7409a,a7413a,a7414a,a7418a,a7419a,a7420a,a7423a,a7427a,a7428a,a7429a,a7433a,a7434a,a7438a,a7439a,a7440a,a7443a,a7447a,a7448a,a7449a,a7453a,a7454a,a7458a,a7459a,a7460a,a7463a,a7467a,a7468a,a7469a,a7473a,a7474a,a7478a,a7479a,a7480a,a7483a,a7487a,a7488a,a7489a,a7493a,a7494a,a7498a,a7499a,a7500a,a7503a,a7507a,a7508a,a7509a,a7513a,a7514a,a7518a,a7519a,a7520a,a7523a,a7527a,a7528a,a7529a,a7533a,a7534a,a7538a,a7539a,a7540a,a7543a,a7547a,a7548a,a7549a,a7553a,a7554a,a7558a,a7559a,a7560a,a7563a,a7567a,a7568a,a7569a,a7573a,a7574a,a7578a,a7579a,a7580a,a7583a,a7587a,a7588a,a7589a,a7593a,a7594a,a7598a,a7599a,a7600a,a7603a,a7607a,a7608a,a7609a,a7613a,a7614a,a7618a,a7619a,a7620a,a7623a,a7627a,a7628a,a7629a,a7633a,a7634a,a7638a,a7639a,a7640a,a7643a,a7647a,a7648a,a7649a,a7653a,a7654a,a7658a,a7659a,a7660a,a7663a,a7667a,a7668a,a7669a,a7673a,a7674a,a7678a,a7679a,a7680a,a7683a,a7687a,a7688a,a7689a,a7693a,a7694a,a7698a,a7699a,a7700a,a7703a,a7707a,a7708a,a7709a,a7713a,a7714a,a7718a,a7719a,a7720a,a7723a,a7727a,a7728a,a7729a,a7733a,a7734a,a7738a,a7739a,a7740a,a7743a,a7747a,a7748a,a7749a,a7753a,a7754a,a7758a,a7759a,a7760a,a7763a,a7767a,a7768a,a7769a,a7773a,a7774a,a7778a,a7779a,a7780a,a7783a,a7787a,a7788a,a7789a,a7793a,a7794a,a7798a,a7799a,a7800a,a7803a,a7807a,a7808a,a7809a,a7813a,a7814a,a7818a,a7819a,a7820a,a7823a,a7827a,a7828a,a7829a,a7833a,a7834a,a7838a,a7839a,a7840a,a7843a,a7847a,a7848a,a7849a,a7853a,a7854a,a7858a,a7859a,a7860a,a7863a,a7867a,a7868a,a7869a,a7873a,a7874a,a7878a,a7879a,a7880a,a7883a,a7887a,a7888a,a7889a,a7893a,a7894a,a7898a,a7899a,a7900a,a7903a,a7907a,a7908a,a7909a,a7913a,a7914a,a7918a,a7919a,a7920a,a7923a,a7927a,a7928a,a7929a,a7933a,a7934a,a7938a,a7939a,a7940a,a7943a,a7947a,a7948a,a7949a,a7953a,a7954a,a7958a,a7959a,a7960a,a7964a,a7965a,a7969a,a7970a,a7971a,a7975a,a7976a,a7980a,a7981a,a7982a,a7986a,a7987a,a7991a,a7992a,a7993a,a7997a,a7998a,a8002a,a8003a,a8004a,a8008a,a8009a,a8013a,a8014a,a8015a,a8019a,a8020a,a8024a,a8025a,a8026a,a8030a,a8031a,a8035a,a8036a,a8037a,a8041a,a8042a,a8046a,a8047a,a8048a,a8052a,a8053a,a8057a,a8058a,a8059a,a8063a,a8064a,a8068a,a8069a,a8070a,a8074a,a8075a,a8079a,a8080a,a8081a,a8085a,a8086a,a8090a,a8091a,a8092a,a8096a,a8097a,a8101a,a8102a,a8103a,a8107a,a8108a,a8112a,a8113a,a8114a,a8118a,a8119a,a8123a,a8124a,a8125a,a8129a,a8130a,a8134a,a8135a,a8136a,a8140a,a8141a,a8145a,a8146a,a8147a,a8151a,a8152a,a8156a,a8157a,a8158a,a8162a,a8163a,a8167a,a8168a,a8169a,a8173a,a8174a,a8178a,a8179a,a8180a,a8184a,a8185a,a8189a,a8190a,a8191a,a8195a,a8196a,a8200a,a8201a,a8202a,a8206a,a8207a,a8211a,a8212a,a8213a,a8217a,a8218a,a8222a,a8223a,a8224a,a8228a,a8229a,a8233a,a8234a,a8235a,a8239a,a8240a,a8244a,a8245a,a8246a,a8250a,a8251a,a8255a,a8256a,a8257a,a8261a,a8262a,a8266a,a8267a,a8268a,a8272a,a8273a,a8277a,a8278a,a8279a,a8283a,a8284a,a8288a,a8289a,a8290a,a8294a,a8295a,a8299a,a8300a,a8301a,a8305a,a8306a,a8310a,a8311a,a8312a,a8316a,a8317a,a8321a,a8322a,a8323a,a8327a,a8328a,a8332a,a8333a,a8334a,a8338a,a8339a,a8343a,a8344a,a8345a,a8349a,a8350a,a8354a,a8355a,a8356a,a8360a,a8361a,a8365a,a8366a,a8367a,a8371a,a8372a,a8376a,a8377a,a8378a,a8382a,a8383a,a8387a,a8388a,a8389a,a8393a,a8394a,a8398a,a8399a,a8400a,a8404a,a8405a,a8409a,a8410a,a8411a,a8415a,a8416a,a8420a,a8421a,a8422a,a8426a,a8427a,a8431a,a8432a,a8433a,a8437a,a8438a,a8442a,a8443a,a8444a,a8448a,a8449a,a8453a,a8454a,a8455a,a8459a,a8460a,a8464a,a8465a,a8466a,a8470a,a8471a,a8475a,a8476a,a8477a,a8481a,a8482a,a8486a,a8487a,a8488a,a8492a,a8493a,a8497a,a8498a,a8499a,a8503a,a8504a,a8508a,a8509a,a8510a,a8514a,a8515a,a8519a,a8520a,a8521a,a8525a,a8526a,a8530a,a8531a,a8532a,a8536a,a8537a,a8541a,a8542a,a8543a,a8547a,a8548a,a8552a,a8553a,a8554a,a8558a,a8559a,a8563a,a8564a,a8565a,a8569a,a8570a,a8574a,a8575a,a8576a,a8580a,a8581a,a8585a,a8586a,a8587a,a8591a,a8592a,a8596a,a8597a,a8598a,a8602a,a8603a,a8607a,a8608a,a8609a,a8613a,a8614a,a8618a,a8619a,a8620a,a8624a,a8625a,a8629a,a8630a,a8631a,a8635a,a8636a,a8640a,a8641a,a8642a,a8646a,a8647a,a8651a,a8652a,a8653a,a8657a,a8658a,a8662a,a8663a,a8664a,a8668a,a8669a,a8673a,a8674a,a8675a,a8679a,a8680a,a8684a,a8685a,a8686a,a8690a,a8691a,a8695a,a8696a,a8697a,a8701a,a8702a,a8706a,a8707a,a8708a,a8712a,a8713a,a8717a,a8718a,a8719a,a8723a,a8724a,a8728a,a8729a,a8730a,a8734a,a8735a,a8739a,a8740a,a8741a,a8745a,a8746a,a8750a,a8751a,a8752a,a8756a,a8757a,a8761a,a8762a,a8763a,a8767a,a8768a,a8772a,a8773a,a8774a,a8778a,a8779a,a8783a,a8784a,a8785a,a8789a,a8790a,a8794a,a8795a,a8796a,a8800a,a8801a,a8805a,a8806a,a8807a,a8811a,a8812a,a8816a,a8817a,a8818a,a8822a,a8823a,a8827a,a8828a,a8829a,a8833a,a8834a,a8838a,a8839a,a8840a,a8844a,a8845a,a8849a,a8850a,a8851a,a8855a,a8856a,a8860a,a8861a,a8862a,a8866a,a8867a,a8871a,a8872a,a8873a,a8877a,a8878a,a8882a,a8883a,a8884a,a8888a,a8889a,a8893a,a8894a,a8895a,a8899a,a8900a,a8904a,a8905a,a8906a,a8910a,a8911a,a8915a,a8916a,a8917a,a8921a,a8922a,a8926a,a8927a,a8928a,a8932a,a8933a,a8937a,a8938a,a8939a,a8943a,a8944a,a8948a,a8949a,a8950a,a8954a,a8955a,a8959a,a8960a,a8961a,a8965a,a8966a,a8970a,a8971a,a8972a,a8976a,a8977a,a8981a,a8982a,a8983a,a8987a,a8988a,a8992a,a8993a,a8994a,a8998a,a8999a,a9003a,a9004a,a9005a,a9009a,a9010a,a9014a,a9015a,a9016a,a9020a,a9021a,a9025a,a9026a,a9027a,a9031a,a9032a,a9036a,a9037a,a9038a,a9042a,a9043a,a9047a,a9048a,a9049a,a9053a,a9054a,a9058a,a9059a,a9060a,a9064a,a9065a,a9069a,a9070a,a9071a,a9075a,a9076a,a9080a,a9081a,a9082a,a9086a,a9087a,a9091a,a9092a,a9093a,a9097a,a9098a,a9102a,a9103a,a9104a,a9108a,a9109a,a9113a,a9114a,a9115a,a9119a,a9120a,a9124a,a9125a,a9126a,a9130a,a9131a,a9135a,a9136a,a9137a,a9141a,a9142a,a9146a,a9147a,a9148a,a9152a,a9153a,a9157a,a9158a,a9159a,a9163a,a9164a,a9168a,a9169a,a9170a,a9174a,a9175a,a9179a,a9180a,a9181a,a9185a,a9186a,a9190a,a9191a,a9192a,a9196a,a9197a,a9201a,a9202a,a9203a,a9207a,a9208a,a9212a,a9213a,a9214a,a9218a,a9219a,a9223a,a9224a,a9225a,a9229a,a9230a,a9234a,a9235a,a9236a,a9240a,a9241a,a9245a,a9246a,a9247a,a9251a,a9252a,a9256a,a9257a,a9258a,a9262a,a9263a,a9267a,a9268a,a9269a,a9273a,a9274a,a9278a,a9279a,a9280a,a9284a,a9285a,a9289a,a9290a,a9291a,a9295a,a9296a,a9300a,a9301a,a9302a,a9306a,a9307a,a9311a,a9312a,a9313a,a9317a,a9318a,a9322a,a9323a,a9324a,a9328a,a9329a,a9333a,a9334a,a9335a,a9339a,a9340a,a9344a,a9345a,a9346a,a9350a,a9351a,a9355a,a9356a,a9357a,a9361a,a9362a,a9366a,a9367a,a9368a,a9372a,a9373a,a9377a,a9378a,a9379a,a9383a,a9384a,a9387a,a9390a,a9391a,a9392a,a9396a,a9397a,a9401a,a9402a,a9403a,a9407a,a9408a,a9411a,a9414a,a9415a,a9416a,a9420a,a9421a,a9425a,a9426a,a9427a,a9431a,a9432a,a9435a,a9438a,a9439a,a9440a,a9444a,a9445a,a9449a,a9450a,a9451a,a9455a,a9456a,a9459a,a9462a,a9463a,a9464a,a9468a,a9469a,a9473a,a9474a,a9475a,a9479a,a9480a,a9483a,a9486a,a9487a,a9488a,a9492a,a9493a,a9497a,a9498a,a9499a,a9503a,a9504a,a9507a,a9510a,a9511a,a9512a,a9516a,a9517a,a9521a,a9522a,a9523a,a9527a,a9528a,a9531a,a9534a,a9535a,a9536a,a9540a,a9541a,a9545a,a9546a,a9547a,a9551a,a9552a,a9555a,a9558a,a9559a,a9560a: std_logic;
begin

A140 <=( a1312a ) or ( a875a );
 a1a <=( a9560a  and  a9547a );
 a2a <=( a9536a  and  a9523a );
 a3a <=( a9512a  and  a9499a );
 a4a <=( a9488a  and  a9475a );
 a5a <=( a9464a  and  a9451a );
 a6a <=( a9440a  and  a9427a );
 a7a <=( a9416a  and  a9403a );
 a8a <=( a9392a  and  a9379a );
 a9a <=( a9368a  and  a9357a );
 a10a <=( a9346a  and  a9335a );
 a11a <=( a9324a  and  a9313a );
 a12a <=( a9302a  and  a9291a );
 a13a <=( a9280a  and  a9269a );
 a14a <=( a9258a  and  a9247a );
 a15a <=( a9236a  and  a9225a );
 a16a <=( a9214a  and  a9203a );
 a17a <=( a9192a  and  a9181a );
 a18a <=( a9170a  and  a9159a );
 a19a <=( a9148a  and  a9137a );
 a20a <=( a9126a  and  a9115a );
 a21a <=( a9104a  and  a9093a );
 a22a <=( a9082a  and  a9071a );
 a23a <=( a9060a  and  a9049a );
 a24a <=( a9038a  and  a9027a );
 a25a <=( a9016a  and  a9005a );
 a26a <=( a8994a  and  a8983a );
 a27a <=( a8972a  and  a8961a );
 a28a <=( a8950a  and  a8939a );
 a29a <=( a8928a  and  a8917a );
 a30a <=( a8906a  and  a8895a );
 a31a <=( a8884a  and  a8873a );
 a32a <=( a8862a  and  a8851a );
 a33a <=( a8840a  and  a8829a );
 a34a <=( a8818a  and  a8807a );
 a35a <=( a8796a  and  a8785a );
 a36a <=( a8774a  and  a8763a );
 a37a <=( a8752a  and  a8741a );
 a38a <=( a8730a  and  a8719a );
 a39a <=( a8708a  and  a8697a );
 a40a <=( a8686a  and  a8675a );
 a41a <=( a8664a  and  a8653a );
 a42a <=( a8642a  and  a8631a );
 a43a <=( a8620a  and  a8609a );
 a44a <=( a8598a  and  a8587a );
 a45a <=( a8576a  and  a8565a );
 a46a <=( a8554a  and  a8543a );
 a47a <=( a8532a  and  a8521a );
 a48a <=( a8510a  and  a8499a );
 a49a <=( a8488a  and  a8477a );
 a50a <=( a8466a  and  a8455a );
 a51a <=( a8444a  and  a8433a );
 a52a <=( a8422a  and  a8411a );
 a53a <=( a8400a  and  a8389a );
 a54a <=( a8378a  and  a8367a );
 a55a <=( a8356a  and  a8345a );
 a56a <=( a8334a  and  a8323a );
 a57a <=( a8312a  and  a8301a );
 a58a <=( a8290a  and  a8279a );
 a59a <=( a8268a  and  a8257a );
 a60a <=( a8246a  and  a8235a );
 a61a <=( a8224a  and  a8213a );
 a62a <=( a8202a  and  a8191a );
 a63a <=( a8180a  and  a8169a );
 a64a <=( a8158a  and  a8147a );
 a65a <=( a8136a  and  a8125a );
 a66a <=( a8114a  and  a8103a );
 a67a <=( a8092a  and  a8081a );
 a68a <=( a8070a  and  a8059a );
 a69a <=( a8048a  and  a8037a );
 a70a <=( a8026a  and  a8015a );
 a71a <=( a8004a  and  a7993a );
 a72a <=( a7982a  and  a7971a );
 a73a <=( a7960a  and  a7949a );
 a74a <=( a7940a  and  a7929a );
 a75a <=( a7920a  and  a7909a );
 a76a <=( a7900a  and  a7889a );
 a77a <=( a7880a  and  a7869a );
 a78a <=( a7860a  and  a7849a );
 a79a <=( a7840a  and  a7829a );
 a80a <=( a7820a  and  a7809a );
 a81a <=( a7800a  and  a7789a );
 a82a <=( a7780a  and  a7769a );
 a83a <=( a7760a  and  a7749a );
 a84a <=( a7740a  and  a7729a );
 a85a <=( a7720a  and  a7709a );
 a86a <=( a7700a  and  a7689a );
 a87a <=( a7680a  and  a7669a );
 a88a <=( a7660a  and  a7649a );
 a89a <=( a7640a  and  a7629a );
 a90a <=( a7620a  and  a7609a );
 a91a <=( a7600a  and  a7589a );
 a92a <=( a7580a  and  a7569a );
 a93a <=( a7560a  and  a7549a );
 a94a <=( a7540a  and  a7529a );
 a95a <=( a7520a  and  a7509a );
 a96a <=( a7500a  and  a7489a );
 a97a <=( a7480a  and  a7469a );
 a98a <=( a7460a  and  a7449a );
 a99a <=( a7440a  and  a7429a );
 a100a <=( a7420a  and  a7409a );
 a101a <=( a7400a  and  a7389a );
 a102a <=( a7380a  and  a7369a );
 a103a <=( a7360a  and  a7349a );
 a104a <=( a7340a  and  a7329a );
 a105a <=( a7320a  and  a7309a );
 a106a <=( a7300a  and  a7289a );
 a107a <=( a7280a  and  a7269a );
 a108a <=( a7260a  and  a7249a );
 a109a <=( a7240a  and  a7229a );
 a110a <=( a7220a  and  a7209a );
 a111a <=( a7200a  and  a7189a );
 a112a <=( a7180a  and  a7169a );
 a113a <=( a7160a  and  a7149a );
 a114a <=( a7140a  and  a7129a );
 a115a <=( a7120a  and  a7109a );
 a116a <=( a7100a  and  a7089a );
 a117a <=( a7080a  and  a7069a );
 a118a <=( a7060a  and  a7049a );
 a119a <=( a7040a  and  a7029a );
 a120a <=( a7020a  and  a7009a );
 a121a <=( a7000a  and  a6989a );
 a122a <=( a6980a  and  a6969a );
 a123a <=( a6960a  and  a6949a );
 a124a <=( a6940a  and  a6929a );
 a125a <=( a6920a  and  a6909a );
 a126a <=( a6900a  and  a6889a );
 a127a <=( a6880a  and  a6869a );
 a128a <=( a6860a  and  a6849a );
 a129a <=( a6840a  and  a6829a );
 a130a <=( a6820a  and  a6809a );
 a131a <=( a6800a  and  a6789a );
 a132a <=( a6780a  and  a6769a );
 a133a <=( a6760a  and  a6749a );
 a134a <=( a6740a  and  a6729a );
 a135a <=( a6720a  and  a6709a );
 a136a <=( a6700a  and  a6689a );
 a137a <=( a6680a  and  a6669a );
 a138a <=( a6660a  and  a6649a );
 a139a <=( a6640a  and  a6629a );
 a140a <=( a6620a  and  a6609a );
 a141a <=( a6600a  and  a6589a );
 a142a <=( a6580a  and  a6569a );
 a143a <=( a6560a  and  a6549a );
 a144a <=( a6540a  and  a6529a );
 a145a <=( a6520a  and  a6509a );
 a146a <=( a6500a  and  a6489a );
 a147a <=( a6480a  and  a6469a );
 a148a <=( a6460a  and  a6449a );
 a149a <=( a6440a  and  a6429a );
 a150a <=( a6420a  and  a6409a );
 a151a <=( a6400a  and  a6389a );
 a152a <=( a6380a  and  a6369a );
 a153a <=( a6360a  and  a6349a );
 a154a <=( a6340a  and  a6329a );
 a155a <=( a6320a  and  a6309a );
 a156a <=( a6300a  and  a6289a );
 a157a <=( a6280a  and  a6269a );
 a158a <=( a6260a  and  a6249a );
 a159a <=( a6240a  and  a6229a );
 a160a <=( a6220a  and  a6209a );
 a161a <=( a6200a  and  a6189a );
 a162a <=( a6180a  and  a6169a );
 a163a <=( a6160a  and  a6149a );
 a164a <=( a6140a  and  a6129a );
 a165a <=( a6120a  and  a6109a );
 a166a <=( a6100a  and  a6089a );
 a167a <=( a6080a  and  a6069a );
 a168a <=( a6060a  and  a6049a );
 a169a <=( a6040a  and  a6029a );
 a170a <=( a6020a  and  a6009a );
 a171a <=( a6000a  and  a5989a );
 a172a <=( a5980a  and  a5969a );
 a173a <=( a5960a  and  a5949a );
 a174a <=( a5940a  and  a5929a );
 a175a <=( a5920a  and  a5909a );
 a176a <=( a5900a  and  a5889a );
 a177a <=( a5880a  and  a5869a );
 a178a <=( a5860a  and  a5849a );
 a179a <=( a5840a  and  a5829a );
 a180a <=( a5820a  and  a5809a );
 a181a <=( a5800a  and  a5789a );
 a182a <=( a5780a  and  a5769a );
 a183a <=( a5760a  and  a5749a );
 a184a <=( a5740a  and  a5729a );
 a185a <=( a5720a  and  a5709a );
 a186a <=( a5700a  and  a5689a );
 a187a <=( a5680a  and  a5669a );
 a188a <=( a5660a  and  a5649a );
 a189a <=( a5640a  and  a5629a );
 a190a <=( a5620a  and  a5609a );
 a191a <=( a5600a  and  a5589a );
 a192a <=( a5580a  and  a5569a );
 a193a <=( a5560a  and  a5549a );
 a194a <=( a5540a  and  a5529a );
 a195a <=( a5520a  and  a5509a );
 a196a <=( a5500a  and  a5489a );
 a197a <=( a5480a  and  a5469a );
 a198a <=( a5460a  and  a5449a );
 a199a <=( a5440a  and  a5429a );
 a200a <=( a5420a  and  a5409a );
 a201a <=( a5400a  and  a5389a );
 a202a <=( a5380a  and  a5369a );
 a203a <=( a5360a  and  a5349a );
 a204a <=( a5340a  and  a5329a );
 a205a <=( a5320a  and  a5309a );
 a206a <=( a5300a  and  a5289a );
 a207a <=( a5280a  and  a5269a );
 a208a <=( a5260a  and  a5249a );
 a209a <=( a5240a  and  a5229a );
 a210a <=( a5220a  and  a5209a );
 a211a <=( a5200a  and  a5189a );
 a212a <=( a5180a  and  a5169a );
 a213a <=( a5160a  and  a5149a );
 a214a <=( a5140a  and  a5129a );
 a215a <=( a5120a  and  a5109a );
 a216a <=( a5100a  and  a5089a );
 a217a <=( a5080a  and  a5069a );
 a218a <=( a5060a  and  a5049a );
 a219a <=( a5040a  and  a5029a );
 a220a <=( a5020a  and  a5009a );
 a221a <=( a5000a  and  a4989a );
 a222a <=( a4980a  and  a4969a );
 a223a <=( a4960a  and  a4949a );
 a224a <=( a4940a  and  a4929a );
 a225a <=( a4920a  and  a4909a );
 a226a <=( a4900a  and  a4889a );
 a227a <=( a4880a  and  a4869a );
 a228a <=( a4860a  and  a4849a );
 a229a <=( a4840a  and  a4829a );
 a230a <=( a4820a  and  a4809a );
 a231a <=( a4800a  and  a4789a );
 a232a <=( a4780a  and  a4769a );
 a233a <=( a4760a  and  a4751a );
 a234a <=( a4742a  and  a4733a );
 a235a <=( a4724a  and  a4715a );
 a236a <=( a4706a  and  a4697a );
 a237a <=( a4688a  and  a4679a );
 a238a <=( a4670a  and  a4661a );
 a239a <=( a4652a  and  a4643a );
 a240a <=( a4634a  and  a4625a );
 a241a <=( a4616a  and  a4607a );
 a242a <=( a4598a  and  a4589a );
 a243a <=( a4580a  and  a4571a );
 a244a <=( a4562a  and  a4553a );
 a245a <=( a4544a  and  a4535a );
 a246a <=( a4526a  and  a4517a );
 a247a <=( a4508a  and  a4499a );
 a248a <=( a4490a  and  a4481a );
 a249a <=( a4472a  and  a4463a );
 a250a <=( a4454a  and  a4445a );
 a251a <=( a4436a  and  a4427a );
 a252a <=( a4418a  and  a4409a );
 a253a <=( a4400a  and  a4391a );
 a254a <=( a4382a  and  a4373a );
 a255a <=( a4364a  and  a4355a );
 a256a <=( a4346a  and  a4337a );
 a257a <=( a4328a  and  a4319a );
 a258a <=( a4310a  and  a4301a );
 a259a <=( a4292a  and  a4283a );
 a260a <=( a4274a  and  a4265a );
 a261a <=( a4256a  and  a4247a );
 a262a <=( a4238a  and  a4229a );
 a263a <=( a4220a  and  a4211a );
 a264a <=( a4202a  and  a4193a );
 a265a <=( a4184a  and  a4175a );
 a266a <=( a4166a  and  a4157a );
 a267a <=( a4148a  and  a4139a );
 a268a <=( a4130a  and  a4121a );
 a269a <=( a4112a  and  a4103a );
 a270a <=( a4094a  and  a4085a );
 a271a <=( a4076a  and  a4067a );
 a272a <=( a4058a  and  a4049a );
 a273a <=( a4040a  and  a4031a );
 a274a <=( a4022a  and  a4013a );
 a275a <=( a4004a  and  a3995a );
 a276a <=( a3986a  and  a3977a );
 a277a <=( a3968a  and  a3959a );
 a278a <=( a3950a  and  a3941a );
 a279a <=( a3932a  and  a3923a );
 a280a <=( a3914a  and  a3905a );
 a281a <=( a3896a  and  a3887a );
 a282a <=( a3878a  and  a3869a );
 a283a <=( a3860a  and  a3851a );
 a284a <=( a3842a  and  a3833a );
 a285a <=( a3824a  and  a3815a );
 a286a <=( a3806a  and  a3797a );
 a287a <=( a3788a  and  a3779a );
 a288a <=( a3770a  and  a3761a );
 a289a <=( a3752a  and  a3743a );
 a290a <=( a3734a  and  a3725a );
 a291a <=( a3716a  and  a3707a );
 a292a <=( a3698a  and  a3689a );
 a293a <=( a3680a  and  a3671a );
 a294a <=( a3662a  and  a3653a );
 a295a <=( a3644a  and  a3635a );
 a296a <=( a3626a  and  a3617a );
 a297a <=( a3608a  and  a3599a );
 a298a <=( a3590a  and  a3581a );
 a299a <=( a3572a  and  a3563a );
 a300a <=( a3554a  and  a3545a );
 a301a <=( a3536a  and  a3527a );
 a302a <=( a3518a  and  a3509a );
 a303a <=( a3500a  and  a3491a );
 a304a <=( a3482a  and  a3473a );
 a305a <=( a3464a  and  a3455a );
 a306a <=( a3446a  and  a3437a );
 a307a <=( a3428a  and  a3419a );
 a308a <=( a3410a  and  a3401a );
 a309a <=( a3392a  and  a3383a );
 a310a <=( a3374a  and  a3365a );
 a311a <=( a3356a  and  a3347a );
 a312a <=( a3338a  and  a3329a );
 a313a <=( a3320a  and  a3311a );
 a314a <=( a3302a  and  a3293a );
 a315a <=( a3284a  and  a3275a );
 a316a <=( a3266a  and  a3257a );
 a317a <=( a3248a  and  a3239a );
 a318a <=( a3230a  and  a3221a );
 a319a <=( a3212a  and  a3203a );
 a320a <=( a3194a  and  a3185a );
 a321a <=( a3176a  and  a3167a );
 a322a <=( a3158a  and  a3149a );
 a323a <=( a3140a  and  a3131a );
 a324a <=( a3122a  and  a3113a );
 a325a <=( a3104a  and  a3095a );
 a326a <=( a3086a  and  a3077a );
 a327a <=( a3068a  and  a3059a );
 a328a <=( a3050a  and  a3041a );
 a329a <=( a3032a  and  a3023a );
 a330a <=( a3014a  and  a3005a );
 a331a <=( a2996a  and  a2987a );
 a332a <=( a2978a  and  a2969a );
 a333a <=( a2960a  and  a2951a );
 a334a <=( a2942a  and  a2933a );
 a335a <=( a2924a  and  a2915a );
 a336a <=( a2906a  and  a2897a );
 a337a <=( a2888a  and  a2879a );
 a338a <=( a2870a  and  a2861a );
 a339a <=( a2852a  and  a2843a );
 a340a <=( a2834a  and  a2825a );
 a341a <=( a2816a  and  a2807a );
 a342a <=( a2798a  and  a2789a );
 a343a <=( a2780a  and  a2771a );
 a344a <=( a2762a  and  a2753a );
 a345a <=( a2744a  and  a2735a );
 a346a <=( a2726a  and  a2717a );
 a347a <=( a2708a  and  a2699a );
 a348a <=( a2690a  and  a2681a );
 a349a <=( a2672a  and  a2663a );
 a350a <=( a2654a  and  a2645a );
 a351a <=( a2636a  and  a2627a );
 a352a <=( a2618a  and  a2609a );
 a353a <=( a2600a  and  a2591a );
 a354a <=( a2582a  and  a2573a );
 a355a <=( a2564a  and  a2555a );
 a356a <=( a2546a  and  a2537a );
 a357a <=( a2528a  and  a2519a );
 a358a <=( a2510a  and  a2501a );
 a359a <=( a2492a  and  a2483a );
 a360a <=( a2474a  and  a2465a );
 a361a <=( a2456a  and  a2447a );
 a362a <=( a2438a  and  a2429a );
 a363a <=( a2420a  and  a2411a );
 a364a <=( a2402a  and  a2393a );
 a365a <=( a2384a  and  a2375a );
 a366a <=( a2366a  and  a2357a );
 a367a <=( a2348a  and  a2339a );
 a368a <=( a2330a  and  a2321a );
 a369a <=( a2312a  and  a2303a );
 a370a <=( a2296a  and  a2287a );
 a371a <=( a2280a  and  a2271a );
 a372a <=( a2264a  and  a2255a );
 a373a <=( a2248a  and  a2239a );
 a374a <=( a2232a  and  a2223a );
 a375a <=( a2216a  and  a2207a );
 a376a <=( a2200a  and  a2191a );
 a377a <=( a2184a  and  a2175a );
 a378a <=( a2168a  and  a2159a );
 a379a <=( a2152a  and  a2143a );
 a380a <=( a2136a  and  a2127a );
 a381a <=( a2120a  and  a2111a );
 a382a <=( a2104a  and  a2095a );
 a383a <=( a2088a  and  a2079a );
 a384a <=( a2072a  and  a2063a );
 a385a <=( a2056a  and  a2047a );
 a386a <=( a2040a  and  a2031a );
 a387a <=( a2024a  and  a2015a );
 a388a <=( a2008a  and  a1999a );
 a389a <=( a1992a  and  a1983a );
 a390a <=( a1976a  and  a1967a );
 a391a <=( a1960a  and  a1951a );
 a392a <=( a1944a  and  a1935a );
 a393a <=( a1928a  and  a1919a );
 a394a <=( a1912a  and  a1903a );
 a395a <=( a1896a  and  a1887a );
 a396a <=( a1880a  and  a1871a );
 a397a <=( a1864a  and  a1855a );
 a398a <=( a1848a  and  a1839a );
 a399a <=( a1832a  and  a1823a );
 a400a <=( a1816a  and  a1807a );
 a401a <=( a1800a  and  a1793a );
 a402a <=( a1786a  and  a1779a );
 a403a <=( a1772a  and  a1765a );
 a404a <=( a1758a  and  a1751a );
 a405a <=( a1744a  and  a1737a );
 a406a <=( a1730a  and  a1723a );
 a407a <=( a1716a  and  a1709a );
 a408a <=( a1702a  and  a1695a );
 a409a <=( a1688a  and  a1681a );
 a410a <=( a1674a  and  a1667a );
 a411a <=( a1660a  and  a1653a );
 a412a <=( a1646a  and  a1639a );
 a413a <=( a1632a  and  a1625a );
 a414a <=( a1618a  and  a1611a );
 a415a <=( a1604a  and  a1597a );
 a416a <=( a1590a  and  a1583a );
 a417a <=( a1576a  and  a1569a );
 a418a <=( a1562a  and  a1555a );
 a419a <=( a1548a  and  a1541a );
 a420a <=( a1534a  and  a1527a );
 a421a <=( a1520a  and  a1513a );
 a422a <=( a1506a  and  a1499a );
 a423a <=( a1492a  and  a1485a );
 a424a <=( a1478a  and  a1471a );
 a425a <=( a1464a  and  a1457a );
 a426a <=( a1450a  and  a1443a );
 a427a <=( a1436a  and  a1429a );
 a428a <=( a1422a  and  a1415a );
 a429a <=( a1408a  and  a1401a );
 a430a <=( a1394a  and  a1387a );
 a431a <=( a1380a  and  a1373a );
 a432a <=( a1366a  and  a1359a );
 a433a <=( a1352a  and  a1347a );
 a434a <=( a1344a  and  a1339a );
 a435a <=( a1336a  and  a1333a );
 a436a <=( a1330a  and  a1327a );
 a437a <=( a1324a  and  a1321a );
 a438a <=( a1318a  and  a1315a );
 a442a <=( a436a ) or ( a437a );
 a443a <=( a438a ) or ( a442a );
 a447a <=( a433a ) or ( a434a );
 a448a <=( a435a ) or ( a447a );
 a449a <=( a448a ) or ( a443a );
 a453a <=( a430a ) or ( a431a );
 a454a <=( a432a ) or ( a453a );
 a457a <=( a428a ) or ( a429a );
 a460a <=( a426a ) or ( a427a );
 a461a <=( a460a ) or ( a457a );
 a462a <=( a461a ) or ( a454a );
 a463a <=( a462a ) or ( a449a );
 a467a <=( a423a ) or ( a424a );
 a468a <=( a425a ) or ( a467a );
 a471a <=( a421a ) or ( a422a );
 a474a <=( a419a ) or ( a420a );
 a475a <=( a474a ) or ( a471a );
 a476a <=( a475a ) or ( a468a );
 a480a <=( a416a ) or ( a417a );
 a481a <=( a418a ) or ( a480a );
 a484a <=( a414a ) or ( a415a );
 a487a <=( a412a ) or ( a413a );
 a488a <=( a487a ) or ( a484a );
 a489a <=( a488a ) or ( a481a );
 a490a <=( a489a ) or ( a476a );
 a491a <=( a490a ) or ( a463a );
 a495a <=( a409a ) or ( a410a );
 a496a <=( a411a ) or ( a495a );
 a500a <=( a406a ) or ( a407a );
 a501a <=( a408a ) or ( a500a );
 a502a <=( a501a ) or ( a496a );
 a506a <=( a403a ) or ( a404a );
 a507a <=( a405a ) or ( a506a );
 a510a <=( a401a ) or ( a402a );
 a513a <=( a399a ) or ( a400a );
 a514a <=( a513a ) or ( a510a );
 a515a <=( a514a ) or ( a507a );
 a516a <=( a515a ) or ( a502a );
 a520a <=( a396a ) or ( a397a );
 a521a <=( a398a ) or ( a520a );
 a524a <=( a394a ) or ( a395a );
 a527a <=( a392a ) or ( a393a );
 a528a <=( a527a ) or ( a524a );
 a529a <=( a528a ) or ( a521a );
 a533a <=( a389a ) or ( a390a );
 a534a <=( a391a ) or ( a533a );
 a537a <=( a387a ) or ( a388a );
 a540a <=( a385a ) or ( a386a );
 a541a <=( a540a ) or ( a537a );
 a542a <=( a541a ) or ( a534a );
 a543a <=( a542a ) or ( a529a );
 a544a <=( a543a ) or ( a516a );
 a545a <=( a544a ) or ( a491a );
 a549a <=( a382a ) or ( a383a );
 a550a <=( a384a ) or ( a549a );
 a554a <=( a379a ) or ( a380a );
 a555a <=( a381a ) or ( a554a );
 a556a <=( a555a ) or ( a550a );
 a560a <=( a376a ) or ( a377a );
 a561a <=( a378a ) or ( a560a );
 a564a <=( a374a ) or ( a375a );
 a567a <=( a372a ) or ( a373a );
 a568a <=( a567a ) or ( a564a );
 a569a <=( a568a ) or ( a561a );
 a570a <=( a569a ) or ( a556a );
 a574a <=( a369a ) or ( a370a );
 a575a <=( a371a ) or ( a574a );
 a578a <=( a367a ) or ( a368a );
 a581a <=( a365a ) or ( a366a );
 a582a <=( a581a ) or ( a578a );
 a583a <=( a582a ) or ( a575a );
 a587a <=( a362a ) or ( a363a );
 a588a <=( a364a ) or ( a587a );
 a591a <=( a360a ) or ( a361a );
 a594a <=( a358a ) or ( a359a );
 a595a <=( a594a ) or ( a591a );
 a596a <=( a595a ) or ( a588a );
 a597a <=( a596a ) or ( a583a );
 a598a <=( a597a ) or ( a570a );
 a602a <=( a355a ) or ( a356a );
 a603a <=( a357a ) or ( a602a );
 a606a <=( a353a ) or ( a354a );
 a609a <=( a351a ) or ( a352a );
 a610a <=( a609a ) or ( a606a );
 a611a <=( a610a ) or ( a603a );
 a615a <=( a348a ) or ( a349a );
 a616a <=( a350a ) or ( a615a );
 a619a <=( a346a ) or ( a347a );
 a622a <=( a344a ) or ( a345a );
 a623a <=( a622a ) or ( a619a );
 a624a <=( a623a ) or ( a616a );
 a625a <=( a624a ) or ( a611a );
 a629a <=( a341a ) or ( a342a );
 a630a <=( a343a ) or ( a629a );
 a633a <=( a339a ) or ( a340a );
 a636a <=( a337a ) or ( a338a );
 a637a <=( a636a ) or ( a633a );
 a638a <=( a637a ) or ( a630a );
 a642a <=( a334a ) or ( a335a );
 a643a <=( a336a ) or ( a642a );
 a646a <=( a332a ) or ( a333a );
 a649a <=( a330a ) or ( a331a );
 a650a <=( a649a ) or ( a646a );
 a651a <=( a650a ) or ( a643a );
 a652a <=( a651a ) or ( a638a );
 a653a <=( a652a ) or ( a625a );
 a654a <=( a653a ) or ( a598a );
 a655a <=( a654a ) or ( a545a );
 a659a <=( a327a ) or ( a328a );
 a660a <=( a329a ) or ( a659a );
 a664a <=( a324a ) or ( a325a );
 a665a <=( a326a ) or ( a664a );
 a666a <=( a665a ) or ( a660a );
 a670a <=( a321a ) or ( a322a );
 a671a <=( a323a ) or ( a670a );
 a674a <=( a319a ) or ( a320a );
 a677a <=( a317a ) or ( a318a );
 a678a <=( a677a ) or ( a674a );
 a679a <=( a678a ) or ( a671a );
 a680a <=( a679a ) or ( a666a );
 a684a <=( a314a ) or ( a315a );
 a685a <=( a316a ) or ( a684a );
 a688a <=( a312a ) or ( a313a );
 a691a <=( a310a ) or ( a311a );
 a692a <=( a691a ) or ( a688a );
 a693a <=( a692a ) or ( a685a );
 a697a <=( a307a ) or ( a308a );
 a698a <=( a309a ) or ( a697a );
 a701a <=( a305a ) or ( a306a );
 a704a <=( a303a ) or ( a304a );
 a705a <=( a704a ) or ( a701a );
 a706a <=( a705a ) or ( a698a );
 a707a <=( a706a ) or ( a693a );
 a708a <=( a707a ) or ( a680a );
 a712a <=( a300a ) or ( a301a );
 a713a <=( a302a ) or ( a712a );
 a716a <=( a298a ) or ( a299a );
 a719a <=( a296a ) or ( a297a );
 a720a <=( a719a ) or ( a716a );
 a721a <=( a720a ) or ( a713a );
 a725a <=( a293a ) or ( a294a );
 a726a <=( a295a ) or ( a725a );
 a729a <=( a291a ) or ( a292a );
 a732a <=( a289a ) or ( a290a );
 a733a <=( a732a ) or ( a729a );
 a734a <=( a733a ) or ( a726a );
 a735a <=( a734a ) or ( a721a );
 a739a <=( a286a ) or ( a287a );
 a740a <=( a288a ) or ( a739a );
 a743a <=( a284a ) or ( a285a );
 a746a <=( a282a ) or ( a283a );
 a747a <=( a746a ) or ( a743a );
 a748a <=( a747a ) or ( a740a );
 a752a <=( a279a ) or ( a280a );
 a753a <=( a281a ) or ( a752a );
 a756a <=( a277a ) or ( a278a );
 a759a <=( a275a ) or ( a276a );
 a760a <=( a759a ) or ( a756a );
 a761a <=( a760a ) or ( a753a );
 a762a <=( a761a ) or ( a748a );
 a763a <=( a762a ) or ( a735a );
 a764a <=( a763a ) or ( a708a );
 a768a <=( a272a ) or ( a273a );
 a769a <=( a274a ) or ( a768a );
 a773a <=( a269a ) or ( a270a );
 a774a <=( a271a ) or ( a773a );
 a775a <=( a774a ) or ( a769a );
 a779a <=( a266a ) or ( a267a );
 a780a <=( a268a ) or ( a779a );
 a783a <=( a264a ) or ( a265a );
 a786a <=( a262a ) or ( a263a );
 a787a <=( a786a ) or ( a783a );
 a788a <=( a787a ) or ( a780a );
 a789a <=( a788a ) or ( a775a );
 a793a <=( a259a ) or ( a260a );
 a794a <=( a261a ) or ( a793a );
 a797a <=( a257a ) or ( a258a );
 a800a <=( a255a ) or ( a256a );
 a801a <=( a800a ) or ( a797a );
 a802a <=( a801a ) or ( a794a );
 a806a <=( a252a ) or ( a253a );
 a807a <=( a254a ) or ( a806a );
 a810a <=( a250a ) or ( a251a );
 a813a <=( a248a ) or ( a249a );
 a814a <=( a813a ) or ( a810a );
 a815a <=( a814a ) or ( a807a );
 a816a <=( a815a ) or ( a802a );
 a817a <=( a816a ) or ( a789a );
 a821a <=( a245a ) or ( a246a );
 a822a <=( a247a ) or ( a821a );
 a825a <=( a243a ) or ( a244a );
 a828a <=( a241a ) or ( a242a );
 a829a <=( a828a ) or ( a825a );
 a830a <=( a829a ) or ( a822a );
 a834a <=( a238a ) or ( a239a );
 a835a <=( a240a ) or ( a834a );
 a838a <=( a236a ) or ( a237a );
 a841a <=( a234a ) or ( a235a );
 a842a <=( a841a ) or ( a838a );
 a843a <=( a842a ) or ( a835a );
 a844a <=( a843a ) or ( a830a );
 a848a <=( a231a ) or ( a232a );
 a849a <=( a233a ) or ( a848a );
 a852a <=( a229a ) or ( a230a );
 a855a <=( a227a ) or ( a228a );
 a856a <=( a855a ) or ( a852a );
 a857a <=( a856a ) or ( a849a );
 a861a <=( a224a ) or ( a225a );
 a862a <=( a226a ) or ( a861a );
 a865a <=( a222a ) or ( a223a );
 a868a <=( a220a ) or ( a221a );
 a869a <=( a868a ) or ( a865a );
 a870a <=( a869a ) or ( a862a );
 a871a <=( a870a ) or ( a857a );
 a872a <=( a871a ) or ( a844a );
 a873a <=( a872a ) or ( a817a );
 a874a <=( a873a ) or ( a764a );
 a875a <=( a874a ) or ( a655a );
 a879a <=( a217a ) or ( a218a );
 a880a <=( a219a ) or ( a879a );
 a884a <=( a214a ) or ( a215a );
 a885a <=( a216a ) or ( a884a );
 a886a <=( a885a ) or ( a880a );
 a890a <=( a211a ) or ( a212a );
 a891a <=( a213a ) or ( a890a );
 a894a <=( a209a ) or ( a210a );
 a897a <=( a207a ) or ( a208a );
 a898a <=( a897a ) or ( a894a );
 a899a <=( a898a ) or ( a891a );
 a900a <=( a899a ) or ( a886a );
 a904a <=( a204a ) or ( a205a );
 a905a <=( a206a ) or ( a904a );
 a908a <=( a202a ) or ( a203a );
 a911a <=( a200a ) or ( a201a );
 a912a <=( a911a ) or ( a908a );
 a913a <=( a912a ) or ( a905a );
 a917a <=( a197a ) or ( a198a );
 a918a <=( a199a ) or ( a917a );
 a921a <=( a195a ) or ( a196a );
 a924a <=( a193a ) or ( a194a );
 a925a <=( a924a ) or ( a921a );
 a926a <=( a925a ) or ( a918a );
 a927a <=( a926a ) or ( a913a );
 a928a <=( a927a ) or ( a900a );
 a932a <=( a190a ) or ( a191a );
 a933a <=( a192a ) or ( a932a );
 a937a <=( a187a ) or ( a188a );
 a938a <=( a189a ) or ( a937a );
 a939a <=( a938a ) or ( a933a );
 a943a <=( a184a ) or ( a185a );
 a944a <=( a186a ) or ( a943a );
 a947a <=( a182a ) or ( a183a );
 a950a <=( a180a ) or ( a181a );
 a951a <=( a950a ) or ( a947a );
 a952a <=( a951a ) or ( a944a );
 a953a <=( a952a ) or ( a939a );
 a957a <=( a177a ) or ( a178a );
 a958a <=( a179a ) or ( a957a );
 a961a <=( a175a ) or ( a176a );
 a964a <=( a173a ) or ( a174a );
 a965a <=( a964a ) or ( a961a );
 a966a <=( a965a ) or ( a958a );
 a970a <=( a170a ) or ( a171a );
 a971a <=( a172a ) or ( a970a );
 a974a <=( a168a ) or ( a169a );
 a977a <=( a166a ) or ( a167a );
 a978a <=( a977a ) or ( a974a );
 a979a <=( a978a ) or ( a971a );
 a980a <=( a979a ) or ( a966a );
 a981a <=( a980a ) or ( a953a );
 a982a <=( a981a ) or ( a928a );
 a986a <=( a163a ) or ( a164a );
 a987a <=( a165a ) or ( a986a );
 a991a <=( a160a ) or ( a161a );
 a992a <=( a162a ) or ( a991a );
 a993a <=( a992a ) or ( a987a );
 a997a <=( a157a ) or ( a158a );
 a998a <=( a159a ) or ( a997a );
 a1001a <=( a155a ) or ( a156a );
 a1004a <=( a153a ) or ( a154a );
 a1005a <=( a1004a ) or ( a1001a );
 a1006a <=( a1005a ) or ( a998a );
 a1007a <=( a1006a ) or ( a993a );
 a1011a <=( a150a ) or ( a151a );
 a1012a <=( a152a ) or ( a1011a );
 a1015a <=( a148a ) or ( a149a );
 a1018a <=( a146a ) or ( a147a );
 a1019a <=( a1018a ) or ( a1015a );
 a1020a <=( a1019a ) or ( a1012a );
 a1024a <=( a143a ) or ( a144a );
 a1025a <=( a145a ) or ( a1024a );
 a1028a <=( a141a ) or ( a142a );
 a1031a <=( a139a ) or ( a140a );
 a1032a <=( a1031a ) or ( a1028a );
 a1033a <=( a1032a ) or ( a1025a );
 a1034a <=( a1033a ) or ( a1020a );
 a1035a <=( a1034a ) or ( a1007a );
 a1039a <=( a136a ) or ( a137a );
 a1040a <=( a138a ) or ( a1039a );
 a1043a <=( a134a ) or ( a135a );
 a1046a <=( a132a ) or ( a133a );
 a1047a <=( a1046a ) or ( a1043a );
 a1048a <=( a1047a ) or ( a1040a );
 a1052a <=( a129a ) or ( a130a );
 a1053a <=( a131a ) or ( a1052a );
 a1056a <=( a127a ) or ( a128a );
 a1059a <=( a125a ) or ( a126a );
 a1060a <=( a1059a ) or ( a1056a );
 a1061a <=( a1060a ) or ( a1053a );
 a1062a <=( a1061a ) or ( a1048a );
 a1066a <=( a122a ) or ( a123a );
 a1067a <=( a124a ) or ( a1066a );
 a1070a <=( a120a ) or ( a121a );
 a1073a <=( a118a ) or ( a119a );
 a1074a <=( a1073a ) or ( a1070a );
 a1075a <=( a1074a ) or ( a1067a );
 a1079a <=( a115a ) or ( a116a );
 a1080a <=( a117a ) or ( a1079a );
 a1083a <=( a113a ) or ( a114a );
 a1086a <=( a111a ) or ( a112a );
 a1087a <=( a1086a ) or ( a1083a );
 a1088a <=( a1087a ) or ( a1080a );
 a1089a <=( a1088a ) or ( a1075a );
 a1090a <=( a1089a ) or ( a1062a );
 a1091a <=( a1090a ) or ( a1035a );
 a1092a <=( a1091a ) or ( a982a );
 a1096a <=( a108a ) or ( a109a );
 a1097a <=( a110a ) or ( a1096a );
 a1101a <=( a105a ) or ( a106a );
 a1102a <=( a107a ) or ( a1101a );
 a1103a <=( a1102a ) or ( a1097a );
 a1107a <=( a102a ) or ( a103a );
 a1108a <=( a104a ) or ( a1107a );
 a1111a <=( a100a ) or ( a101a );
 a1114a <=( a98a ) or ( a99a );
 a1115a <=( a1114a ) or ( a1111a );
 a1116a <=( a1115a ) or ( a1108a );
 a1117a <=( a1116a ) or ( a1103a );
 a1121a <=( a95a ) or ( a96a );
 a1122a <=( a97a ) or ( a1121a );
 a1125a <=( a93a ) or ( a94a );
 a1128a <=( a91a ) or ( a92a );
 a1129a <=( a1128a ) or ( a1125a );
 a1130a <=( a1129a ) or ( a1122a );
 a1134a <=( a88a ) or ( a89a );
 a1135a <=( a90a ) or ( a1134a );
 a1138a <=( a86a ) or ( a87a );
 a1141a <=( a84a ) or ( a85a );
 a1142a <=( a1141a ) or ( a1138a );
 a1143a <=( a1142a ) or ( a1135a );
 a1144a <=( a1143a ) or ( a1130a );
 a1145a <=( a1144a ) or ( a1117a );
 a1149a <=( a81a ) or ( a82a );
 a1150a <=( a83a ) or ( a1149a );
 a1153a <=( a79a ) or ( a80a );
 a1156a <=( a77a ) or ( a78a );
 a1157a <=( a1156a ) or ( a1153a );
 a1158a <=( a1157a ) or ( a1150a );
 a1162a <=( a74a ) or ( a75a );
 a1163a <=( a76a ) or ( a1162a );
 a1166a <=( a72a ) or ( a73a );
 a1169a <=( a70a ) or ( a71a );
 a1170a <=( a1169a ) or ( a1166a );
 a1171a <=( a1170a ) or ( a1163a );
 a1172a <=( a1171a ) or ( a1158a );
 a1176a <=( a67a ) or ( a68a );
 a1177a <=( a69a ) or ( a1176a );
 a1180a <=( a65a ) or ( a66a );
 a1183a <=( a63a ) or ( a64a );
 a1184a <=( a1183a ) or ( a1180a );
 a1185a <=( a1184a ) or ( a1177a );
 a1189a <=( a60a ) or ( a61a );
 a1190a <=( a62a ) or ( a1189a );
 a1193a <=( a58a ) or ( a59a );
 a1196a <=( a56a ) or ( a57a );
 a1197a <=( a1196a ) or ( a1193a );
 a1198a <=( a1197a ) or ( a1190a );
 a1199a <=( a1198a ) or ( a1185a );
 a1200a <=( a1199a ) or ( a1172a );
 a1201a <=( a1200a ) or ( a1145a );
 a1205a <=( a53a ) or ( a54a );
 a1206a <=( a55a ) or ( a1205a );
 a1210a <=( a50a ) or ( a51a );
 a1211a <=( a52a ) or ( a1210a );
 a1212a <=( a1211a ) or ( a1206a );
 a1216a <=( a47a ) or ( a48a );
 a1217a <=( a49a ) or ( a1216a );
 a1220a <=( a45a ) or ( a46a );
 a1223a <=( a43a ) or ( a44a );
 a1224a <=( a1223a ) or ( a1220a );
 a1225a <=( a1224a ) or ( a1217a );
 a1226a <=( a1225a ) or ( a1212a );
 a1230a <=( a40a ) or ( a41a );
 a1231a <=( a42a ) or ( a1230a );
 a1234a <=( a38a ) or ( a39a );
 a1237a <=( a36a ) or ( a37a );
 a1238a <=( a1237a ) or ( a1234a );
 a1239a <=( a1238a ) or ( a1231a );
 a1243a <=( a33a ) or ( a34a );
 a1244a <=( a35a ) or ( a1243a );
 a1247a <=( a31a ) or ( a32a );
 a1250a <=( a29a ) or ( a30a );
 a1251a <=( a1250a ) or ( a1247a );
 a1252a <=( a1251a ) or ( a1244a );
 a1253a <=( a1252a ) or ( a1239a );
 a1254a <=( a1253a ) or ( a1226a );
 a1258a <=( a26a ) or ( a27a );
 a1259a <=( a28a ) or ( a1258a );
 a1262a <=( a24a ) or ( a25a );
 a1265a <=( a22a ) or ( a23a );
 a1266a <=( a1265a ) or ( a1262a );
 a1267a <=( a1266a ) or ( a1259a );
 a1271a <=( a19a ) or ( a20a );
 a1272a <=( a21a ) or ( a1271a );
 a1275a <=( a17a ) or ( a18a );
 a1278a <=( a15a ) or ( a16a );
 a1279a <=( a1278a ) or ( a1275a );
 a1280a <=( a1279a ) or ( a1272a );
 a1281a <=( a1280a ) or ( a1267a );
 a1285a <=( a12a ) or ( a13a );
 a1286a <=( a14a ) or ( a1285a );
 a1289a <=( a10a ) or ( a11a );
 a1292a <=( a8a ) or ( a9a );
 a1293a <=( a1292a ) or ( a1289a );
 a1294a <=( a1293a ) or ( a1286a );
 a1298a <=( a5a ) or ( a6a );
 a1299a <=( a7a ) or ( a1298a );
 a1302a <=( a3a ) or ( a4a );
 a1305a <=( a1a ) or ( a2a );
 a1306a <=( a1305a ) or ( a1302a );
 a1307a <=( a1306a ) or ( a1299a );
 a1308a <=( a1307a ) or ( a1294a );
 a1309a <=( a1308a ) or ( a1281a );
 a1310a <=( a1309a ) or ( a1254a );
 a1311a <=( a1310a ) or ( a1201a );
 a1312a <=( a1311a ) or ( a1092a );
 a1315a <=( A266  and  (not A265) );
 a1318a <=( A268  and  A267 );
 a1321a <=( A266  and  (not A265) );
 a1324a <=( A269  and  A267 );
 a1327a <=( (not A266)  and  A265 );
 a1330a <=( A268  and  A267 );
 a1333a <=( (not A266)  and  A265 );
 a1336a <=( A269  and  A267 );
 a1339a <=( A266  and  (not A265) );
 a1343a <=( (not A269)  and  (not A268) );
 a1344a <=( (not A267)  and  a1343a );
 a1347a <=( (not A266)  and  A265 );
 a1351a <=( (not A269)  and  (not A268) );
 a1352a <=( (not A267)  and  a1351a );
 a1355a <=( A200  and  (not A199) );
 a1358a <=( A202  and  A201 );
 a1359a <=( a1358a  and  a1355a );
 a1362a <=( A233  and  (not A232) );
 a1365a <=( A235  and  A234 );
 a1366a <=( a1365a  and  a1362a );
 a1369a <=( A200  and  (not A199) );
 a1372a <=( A202  and  A201 );
 a1373a <=( a1372a  and  a1369a );
 a1376a <=( A233  and  (not A232) );
 a1379a <=( A236  and  A234 );
 a1380a <=( a1379a  and  a1376a );
 a1383a <=( A200  and  (not A199) );
 a1386a <=( A202  and  A201 );
 a1387a <=( a1386a  and  a1383a );
 a1390a <=( (not A233)  and  A232 );
 a1393a <=( A235  and  A234 );
 a1394a <=( a1393a  and  a1390a );
 a1397a <=( A200  and  (not A199) );
 a1400a <=( A202  and  A201 );
 a1401a <=( a1400a  and  a1397a );
 a1404a <=( (not A233)  and  A232 );
 a1407a <=( A236  and  A234 );
 a1408a <=( a1407a  and  a1404a );
 a1411a <=( A200  and  (not A199) );
 a1414a <=( A203  and  A201 );
 a1415a <=( a1414a  and  a1411a );
 a1418a <=( A233  and  (not A232) );
 a1421a <=( A235  and  A234 );
 a1422a <=( a1421a  and  a1418a );
 a1425a <=( A200  and  (not A199) );
 a1428a <=( A203  and  A201 );
 a1429a <=( a1428a  and  a1425a );
 a1432a <=( A233  and  (not A232) );
 a1435a <=( A236  and  A234 );
 a1436a <=( a1435a  and  a1432a );
 a1439a <=( A200  and  (not A199) );
 a1442a <=( A203  and  A201 );
 a1443a <=( a1442a  and  a1439a );
 a1446a <=( (not A233)  and  A232 );
 a1449a <=( A235  and  A234 );
 a1450a <=( a1449a  and  a1446a );
 a1453a <=( A200  and  (not A199) );
 a1456a <=( A203  and  A201 );
 a1457a <=( a1456a  and  a1453a );
 a1460a <=( (not A233)  and  A232 );
 a1463a <=( A236  and  A234 );
 a1464a <=( a1463a  and  a1460a );
 a1467a <=( (not A200)  and  A199 );
 a1470a <=( A202  and  A201 );
 a1471a <=( a1470a  and  a1467a );
 a1474a <=( A233  and  (not A232) );
 a1477a <=( A235  and  A234 );
 a1478a <=( a1477a  and  a1474a );
 a1481a <=( (not A200)  and  A199 );
 a1484a <=( A202  and  A201 );
 a1485a <=( a1484a  and  a1481a );
 a1488a <=( A233  and  (not A232) );
 a1491a <=( A236  and  A234 );
 a1492a <=( a1491a  and  a1488a );
 a1495a <=( (not A200)  and  A199 );
 a1498a <=( A202  and  A201 );
 a1499a <=( a1498a  and  a1495a );
 a1502a <=( (not A233)  and  A232 );
 a1505a <=( A235  and  A234 );
 a1506a <=( a1505a  and  a1502a );
 a1509a <=( (not A200)  and  A199 );
 a1512a <=( A202  and  A201 );
 a1513a <=( a1512a  and  a1509a );
 a1516a <=( (not A233)  and  A232 );
 a1519a <=( A236  and  A234 );
 a1520a <=( a1519a  and  a1516a );
 a1523a <=( (not A200)  and  A199 );
 a1526a <=( A203  and  A201 );
 a1527a <=( a1526a  and  a1523a );
 a1530a <=( A233  and  (not A232) );
 a1533a <=( A235  and  A234 );
 a1534a <=( a1533a  and  a1530a );
 a1537a <=( (not A200)  and  A199 );
 a1540a <=( A203  and  A201 );
 a1541a <=( a1540a  and  a1537a );
 a1544a <=( A233  and  (not A232) );
 a1547a <=( A236  and  A234 );
 a1548a <=( a1547a  and  a1544a );
 a1551a <=( (not A200)  and  A199 );
 a1554a <=( A203  and  A201 );
 a1555a <=( a1554a  and  a1551a );
 a1558a <=( (not A233)  and  A232 );
 a1561a <=( A235  and  A234 );
 a1562a <=( a1561a  and  a1558a );
 a1565a <=( (not A200)  and  A199 );
 a1568a <=( A203  and  A201 );
 a1569a <=( a1568a  and  a1565a );
 a1572a <=( (not A233)  and  A232 );
 a1575a <=( A236  and  A234 );
 a1576a <=( a1575a  and  a1572a );
 a1579a <=( A168  and  (not A170) );
 a1582a <=( (not A166)  and  A167 );
 a1583a <=( a1582a  and  a1579a );
 a1586a <=( A233  and  (not A232) );
 a1589a <=( A235  and  A234 );
 a1590a <=( a1589a  and  a1586a );
 a1593a <=( A168  and  (not A170) );
 a1596a <=( (not A166)  and  A167 );
 a1597a <=( a1596a  and  a1593a );
 a1600a <=( A233  and  (not A232) );
 a1603a <=( A236  and  A234 );
 a1604a <=( a1603a  and  a1600a );
 a1607a <=( A168  and  (not A170) );
 a1610a <=( (not A166)  and  A167 );
 a1611a <=( a1610a  and  a1607a );
 a1614a <=( (not A233)  and  A232 );
 a1617a <=( A235  and  A234 );
 a1618a <=( a1617a  and  a1614a );
 a1621a <=( A168  and  (not A170) );
 a1624a <=( (not A166)  and  A167 );
 a1625a <=( a1624a  and  a1621a );
 a1628a <=( (not A233)  and  A232 );
 a1631a <=( A236  and  A234 );
 a1632a <=( a1631a  and  a1628a );
 a1635a <=( A168  and  (not A170) );
 a1638a <=( A166  and  (not A167) );
 a1639a <=( a1638a  and  a1635a );
 a1642a <=( A233  and  (not A232) );
 a1645a <=( A235  and  A234 );
 a1646a <=( a1645a  and  a1642a );
 a1649a <=( A168  and  (not A170) );
 a1652a <=( A166  and  (not A167) );
 a1653a <=( a1652a  and  a1649a );
 a1656a <=( A233  and  (not A232) );
 a1659a <=( A236  and  A234 );
 a1660a <=( a1659a  and  a1656a );
 a1663a <=( A168  and  (not A170) );
 a1666a <=( A166  and  (not A167) );
 a1667a <=( a1666a  and  a1663a );
 a1670a <=( (not A233)  and  A232 );
 a1673a <=( A235  and  A234 );
 a1674a <=( a1673a  and  a1670a );
 a1677a <=( A168  and  (not A170) );
 a1680a <=( A166  and  (not A167) );
 a1681a <=( a1680a  and  a1677a );
 a1684a <=( (not A233)  and  A232 );
 a1687a <=( A236  and  A234 );
 a1688a <=( a1687a  and  a1684a );
 a1691a <=( A168  and  A169 );
 a1694a <=( (not A166)  and  A167 );
 a1695a <=( a1694a  and  a1691a );
 a1698a <=( A233  and  (not A232) );
 a1701a <=( A235  and  A234 );
 a1702a <=( a1701a  and  a1698a );
 a1705a <=( A168  and  A169 );
 a1708a <=( (not A166)  and  A167 );
 a1709a <=( a1708a  and  a1705a );
 a1712a <=( A233  and  (not A232) );
 a1715a <=( A236  and  A234 );
 a1716a <=( a1715a  and  a1712a );
 a1719a <=( A168  and  A169 );
 a1722a <=( (not A166)  and  A167 );
 a1723a <=( a1722a  and  a1719a );
 a1726a <=( (not A233)  and  A232 );
 a1729a <=( A235  and  A234 );
 a1730a <=( a1729a  and  a1726a );
 a1733a <=( A168  and  A169 );
 a1736a <=( (not A166)  and  A167 );
 a1737a <=( a1736a  and  a1733a );
 a1740a <=( (not A233)  and  A232 );
 a1743a <=( A236  and  A234 );
 a1744a <=( a1743a  and  a1740a );
 a1747a <=( A168  and  A169 );
 a1750a <=( A166  and  (not A167) );
 a1751a <=( a1750a  and  a1747a );
 a1754a <=( A233  and  (not A232) );
 a1757a <=( A235  and  A234 );
 a1758a <=( a1757a  and  a1754a );
 a1761a <=( A168  and  A169 );
 a1764a <=( A166  and  (not A167) );
 a1765a <=( a1764a  and  a1761a );
 a1768a <=( A233  and  (not A232) );
 a1771a <=( A236  and  A234 );
 a1772a <=( a1771a  and  a1768a );
 a1775a <=( A168  and  A169 );
 a1778a <=( A166  and  (not A167) );
 a1779a <=( a1778a  and  a1775a );
 a1782a <=( (not A233)  and  A232 );
 a1785a <=( A235  and  A234 );
 a1786a <=( a1785a  and  a1782a );
 a1789a <=( A168  and  A169 );
 a1792a <=( A166  and  (not A167) );
 a1793a <=( a1792a  and  a1789a );
 a1796a <=( (not A233)  and  A232 );
 a1799a <=( A236  and  A234 );
 a1800a <=( a1799a  and  a1796a );
 a1803a <=( A200  and  (not A199) );
 a1806a <=( A202  and  A201 );
 a1807a <=( a1806a  and  a1803a );
 a1810a <=( A233  and  (not A232) );
 a1814a <=( (not A236)  and  (not A235) );
 a1815a <=( (not A234)  and  a1814a );
 a1816a <=( a1815a  and  a1810a );
 a1819a <=( A200  and  (not A199) );
 a1822a <=( A202  and  A201 );
 a1823a <=( a1822a  and  a1819a );
 a1826a <=( (not A233)  and  A232 );
 a1830a <=( (not A236)  and  (not A235) );
 a1831a <=( (not A234)  and  a1830a );
 a1832a <=( a1831a  and  a1826a );
 a1835a <=( A200  and  (not A199) );
 a1838a <=( A203  and  A201 );
 a1839a <=( a1838a  and  a1835a );
 a1842a <=( A233  and  (not A232) );
 a1846a <=( (not A236)  and  (not A235) );
 a1847a <=( (not A234)  and  a1846a );
 a1848a <=( a1847a  and  a1842a );
 a1851a <=( A200  and  (not A199) );
 a1854a <=( A203  and  A201 );
 a1855a <=( a1854a  and  a1851a );
 a1858a <=( (not A233)  and  A232 );
 a1862a <=( (not A236)  and  (not A235) );
 a1863a <=( (not A234)  and  a1862a );
 a1864a <=( a1863a  and  a1858a );
 a1867a <=( A200  and  (not A199) );
 a1870a <=( (not A202)  and  (not A201) );
 a1871a <=( a1870a  and  a1867a );
 a1874a <=( (not A232)  and  (not A203) );
 a1878a <=( A235  and  A234 );
 a1879a <=( A233  and  a1878a );
 a1880a <=( a1879a  and  a1874a );
 a1883a <=( A200  and  (not A199) );
 a1886a <=( (not A202)  and  (not A201) );
 a1887a <=( a1886a  and  a1883a );
 a1890a <=( (not A232)  and  (not A203) );
 a1894a <=( A236  and  A234 );
 a1895a <=( A233  and  a1894a );
 a1896a <=( a1895a  and  a1890a );
 a1899a <=( A200  and  (not A199) );
 a1902a <=( (not A202)  and  (not A201) );
 a1903a <=( a1902a  and  a1899a );
 a1906a <=( A232  and  (not A203) );
 a1910a <=( A235  and  A234 );
 a1911a <=( (not A233)  and  a1910a );
 a1912a <=( a1911a  and  a1906a );
 a1915a <=( A200  and  (not A199) );
 a1918a <=( (not A202)  and  (not A201) );
 a1919a <=( a1918a  and  a1915a );
 a1922a <=( A232  and  (not A203) );
 a1926a <=( A236  and  A234 );
 a1927a <=( (not A233)  and  a1926a );
 a1928a <=( a1927a  and  a1922a );
 a1931a <=( (not A200)  and  A199 );
 a1934a <=( A202  and  A201 );
 a1935a <=( a1934a  and  a1931a );
 a1938a <=( A233  and  (not A232) );
 a1942a <=( (not A236)  and  (not A235) );
 a1943a <=( (not A234)  and  a1942a );
 a1944a <=( a1943a  and  a1938a );
 a1947a <=( (not A200)  and  A199 );
 a1950a <=( A202  and  A201 );
 a1951a <=( a1950a  and  a1947a );
 a1954a <=( (not A233)  and  A232 );
 a1958a <=( (not A236)  and  (not A235) );
 a1959a <=( (not A234)  and  a1958a );
 a1960a <=( a1959a  and  a1954a );
 a1963a <=( (not A200)  and  A199 );
 a1966a <=( A203  and  A201 );
 a1967a <=( a1966a  and  a1963a );
 a1970a <=( A233  and  (not A232) );
 a1974a <=( (not A236)  and  (not A235) );
 a1975a <=( (not A234)  and  a1974a );
 a1976a <=( a1975a  and  a1970a );
 a1979a <=( (not A200)  and  A199 );
 a1982a <=( A203  and  A201 );
 a1983a <=( a1982a  and  a1979a );
 a1986a <=( (not A233)  and  A232 );
 a1990a <=( (not A236)  and  (not A235) );
 a1991a <=( (not A234)  and  a1990a );
 a1992a <=( a1991a  and  a1986a );
 a1995a <=( (not A200)  and  A199 );
 a1998a <=( (not A202)  and  (not A201) );
 a1999a <=( a1998a  and  a1995a );
 a2002a <=( (not A232)  and  (not A203) );
 a2006a <=( A235  and  A234 );
 a2007a <=( A233  and  a2006a );
 a2008a <=( a2007a  and  a2002a );
 a2011a <=( (not A200)  and  A199 );
 a2014a <=( (not A202)  and  (not A201) );
 a2015a <=( a2014a  and  a2011a );
 a2018a <=( (not A232)  and  (not A203) );
 a2022a <=( A236  and  A234 );
 a2023a <=( A233  and  a2022a );
 a2024a <=( a2023a  and  a2018a );
 a2027a <=( (not A200)  and  A199 );
 a2030a <=( (not A202)  and  (not A201) );
 a2031a <=( a2030a  and  a2027a );
 a2034a <=( A232  and  (not A203) );
 a2038a <=( A235  and  A234 );
 a2039a <=( (not A233)  and  a2038a );
 a2040a <=( a2039a  and  a2034a );
 a2043a <=( (not A200)  and  A199 );
 a2046a <=( (not A202)  and  (not A201) );
 a2047a <=( a2046a  and  a2043a );
 a2050a <=( A232  and  (not A203) );
 a2054a <=( A236  and  A234 );
 a2055a <=( (not A233)  and  a2054a );
 a2056a <=( a2055a  and  a2050a );
 a2059a <=( A168  and  (not A170) );
 a2062a <=( (not A166)  and  A167 );
 a2063a <=( a2062a  and  a2059a );
 a2066a <=( A233  and  (not A232) );
 a2070a <=( (not A236)  and  (not A235) );
 a2071a <=( (not A234)  and  a2070a );
 a2072a <=( a2071a  and  a2066a );
 a2075a <=( A168  and  (not A170) );
 a2078a <=( (not A166)  and  A167 );
 a2079a <=( a2078a  and  a2075a );
 a2082a <=( (not A233)  and  A232 );
 a2086a <=( (not A236)  and  (not A235) );
 a2087a <=( (not A234)  and  a2086a );
 a2088a <=( a2087a  and  a2082a );
 a2091a <=( A168  and  (not A170) );
 a2094a <=( A166  and  (not A167) );
 a2095a <=( a2094a  and  a2091a );
 a2098a <=( A233  and  (not A232) );
 a2102a <=( (not A236)  and  (not A235) );
 a2103a <=( (not A234)  and  a2102a );
 a2104a <=( a2103a  and  a2098a );
 a2107a <=( A168  and  (not A170) );
 a2110a <=( A166  and  (not A167) );
 a2111a <=( a2110a  and  a2107a );
 a2114a <=( (not A233)  and  A232 );
 a2118a <=( (not A236)  and  (not A235) );
 a2119a <=( (not A234)  and  a2118a );
 a2120a <=( a2119a  and  a2114a );
 a2123a <=( A168  and  A169 );
 a2126a <=( (not A166)  and  A167 );
 a2127a <=( a2126a  and  a2123a );
 a2130a <=( A233  and  (not A232) );
 a2134a <=( (not A236)  and  (not A235) );
 a2135a <=( (not A234)  and  a2134a );
 a2136a <=( a2135a  and  a2130a );
 a2139a <=( A168  and  A169 );
 a2142a <=( (not A166)  and  A167 );
 a2143a <=( a2142a  and  a2139a );
 a2146a <=( (not A233)  and  A232 );
 a2150a <=( (not A236)  and  (not A235) );
 a2151a <=( (not A234)  and  a2150a );
 a2152a <=( a2151a  and  a2146a );
 a2155a <=( A168  and  A169 );
 a2158a <=( A166  and  (not A167) );
 a2159a <=( a2158a  and  a2155a );
 a2162a <=( A233  and  (not A232) );
 a2166a <=( (not A236)  and  (not A235) );
 a2167a <=( (not A234)  and  a2166a );
 a2168a <=( a2167a  and  a2162a );
 a2171a <=( A168  and  A169 );
 a2174a <=( A166  and  (not A167) );
 a2175a <=( a2174a  and  a2171a );
 a2178a <=( (not A233)  and  A232 );
 a2182a <=( (not A236)  and  (not A235) );
 a2183a <=( (not A234)  and  a2182a );
 a2184a <=( a2183a  and  a2178a );
 a2187a <=( (not A169)  and  A170 );
 a2190a <=( A167  and  (not A168) );
 a2191a <=( a2190a  and  a2187a );
 a2194a <=( (not A232)  and  (not A166) );
 a2198a <=( A235  and  A234 );
 a2199a <=( A233  and  a2198a );
 a2200a <=( a2199a  and  a2194a );
 a2203a <=( (not A169)  and  A170 );
 a2206a <=( A167  and  (not A168) );
 a2207a <=( a2206a  and  a2203a );
 a2210a <=( (not A232)  and  (not A166) );
 a2214a <=( A236  and  A234 );
 a2215a <=( A233  and  a2214a );
 a2216a <=( a2215a  and  a2210a );
 a2219a <=( (not A169)  and  A170 );
 a2222a <=( A167  and  (not A168) );
 a2223a <=( a2222a  and  a2219a );
 a2226a <=( A232  and  (not A166) );
 a2230a <=( A235  and  A234 );
 a2231a <=( (not A233)  and  a2230a );
 a2232a <=( a2231a  and  a2226a );
 a2235a <=( (not A169)  and  A170 );
 a2238a <=( A167  and  (not A168) );
 a2239a <=( a2238a  and  a2235a );
 a2242a <=( A232  and  (not A166) );
 a2246a <=( A236  and  A234 );
 a2247a <=( (not A233)  and  a2246a );
 a2248a <=( a2247a  and  a2242a );
 a2251a <=( (not A169)  and  A170 );
 a2254a <=( (not A167)  and  (not A168) );
 a2255a <=( a2254a  and  a2251a );
 a2258a <=( (not A232)  and  A166 );
 a2262a <=( A235  and  A234 );
 a2263a <=( A233  and  a2262a );
 a2264a <=( a2263a  and  a2258a );
 a2267a <=( (not A169)  and  A170 );
 a2270a <=( (not A167)  and  (not A168) );
 a2271a <=( a2270a  and  a2267a );
 a2274a <=( (not A232)  and  A166 );
 a2278a <=( A236  and  A234 );
 a2279a <=( A233  and  a2278a );
 a2280a <=( a2279a  and  a2274a );
 a2283a <=( (not A169)  and  A170 );
 a2286a <=( (not A167)  and  (not A168) );
 a2287a <=( a2286a  and  a2283a );
 a2290a <=( A232  and  A166 );
 a2294a <=( A235  and  A234 );
 a2295a <=( (not A233)  and  a2294a );
 a2296a <=( a2295a  and  a2290a );
 a2299a <=( (not A169)  and  A170 );
 a2302a <=( (not A167)  and  (not A168) );
 a2303a <=( a2302a  and  a2299a );
 a2306a <=( A232  and  A166 );
 a2310a <=( A236  and  A234 );
 a2311a <=( (not A233)  and  a2310a );
 a2312a <=( a2311a  and  a2306a );
 a2315a <=( A200  and  (not A199) );
 a2319a <=( (not A203)  and  (not A202) );
 a2320a <=( (not A201)  and  a2319a );
 a2321a <=( a2320a  and  a2315a );
 a2324a <=( A233  and  (not A232) );
 a2328a <=( (not A236)  and  (not A235) );
 a2329a <=( (not A234)  and  a2328a );
 a2330a <=( a2329a  and  a2324a );
 a2333a <=( A200  and  (not A199) );
 a2337a <=( (not A203)  and  (not A202) );
 a2338a <=( (not A201)  and  a2337a );
 a2339a <=( a2338a  and  a2333a );
 a2342a <=( (not A233)  and  A232 );
 a2346a <=( (not A236)  and  (not A235) );
 a2347a <=( (not A234)  and  a2346a );
 a2348a <=( a2347a  and  a2342a );
 a2351a <=( (not A200)  and  A199 );
 a2355a <=( (not A203)  and  (not A202) );
 a2356a <=( (not A201)  and  a2355a );
 a2357a <=( a2356a  and  a2351a );
 a2360a <=( A233  and  (not A232) );
 a2364a <=( (not A236)  and  (not A235) );
 a2365a <=( (not A234)  and  a2364a );
 a2366a <=( a2365a  and  a2360a );
 a2369a <=( (not A200)  and  A199 );
 a2373a <=( (not A203)  and  (not A202) );
 a2374a <=( (not A201)  and  a2373a );
 a2375a <=( a2374a  and  a2369a );
 a2378a <=( (not A233)  and  A232 );
 a2382a <=( (not A236)  and  (not A235) );
 a2383a <=( (not A234)  and  a2382a );
 a2384a <=( a2383a  and  a2378a );
 a2387a <=( A166  and  A167 );
 a2391a <=( A201  and  A200 );
 a2392a <=( (not A199)  and  a2391a );
 a2393a <=( a2392a  and  a2387a );
 a2396a <=( A298  and  A202 );
 a2400a <=( A301  and  A300 );
 a2401a <=( (not A299)  and  a2400a );
 a2402a <=( a2401a  and  a2396a );
 a2405a <=( A166  and  A167 );
 a2409a <=( A201  and  A200 );
 a2410a <=( (not A199)  and  a2409a );
 a2411a <=( a2410a  and  a2405a );
 a2414a <=( A298  and  A202 );
 a2418a <=( A302  and  A300 );
 a2419a <=( (not A299)  and  a2418a );
 a2420a <=( a2419a  and  a2414a );
 a2423a <=( A166  and  A167 );
 a2427a <=( A201  and  A200 );
 a2428a <=( (not A199)  and  a2427a );
 a2429a <=( a2428a  and  a2423a );
 a2432a <=( (not A298)  and  A202 );
 a2436a <=( A301  and  A300 );
 a2437a <=( A299  and  a2436a );
 a2438a <=( a2437a  and  a2432a );
 a2441a <=( A166  and  A167 );
 a2445a <=( A201  and  A200 );
 a2446a <=( (not A199)  and  a2445a );
 a2447a <=( a2446a  and  a2441a );
 a2450a <=( (not A298)  and  A202 );
 a2454a <=( A302  and  A300 );
 a2455a <=( A299  and  a2454a );
 a2456a <=( a2455a  and  a2450a );
 a2459a <=( A166  and  A167 );
 a2463a <=( A201  and  A200 );
 a2464a <=( (not A199)  and  a2463a );
 a2465a <=( a2464a  and  a2459a );
 a2468a <=( A298  and  A203 );
 a2472a <=( A301  and  A300 );
 a2473a <=( (not A299)  and  a2472a );
 a2474a <=( a2473a  and  a2468a );
 a2477a <=( A166  and  A167 );
 a2481a <=( A201  and  A200 );
 a2482a <=( (not A199)  and  a2481a );
 a2483a <=( a2482a  and  a2477a );
 a2486a <=( A298  and  A203 );
 a2490a <=( A302  and  A300 );
 a2491a <=( (not A299)  and  a2490a );
 a2492a <=( a2491a  and  a2486a );
 a2495a <=( A166  and  A167 );
 a2499a <=( A201  and  A200 );
 a2500a <=( (not A199)  and  a2499a );
 a2501a <=( a2500a  and  a2495a );
 a2504a <=( (not A298)  and  A203 );
 a2508a <=( A301  and  A300 );
 a2509a <=( A299  and  a2508a );
 a2510a <=( a2509a  and  a2504a );
 a2513a <=( A166  and  A167 );
 a2517a <=( A201  and  A200 );
 a2518a <=( (not A199)  and  a2517a );
 a2519a <=( a2518a  and  a2513a );
 a2522a <=( (not A298)  and  A203 );
 a2526a <=( A302  and  A300 );
 a2527a <=( A299  and  a2526a );
 a2528a <=( a2527a  and  a2522a );
 a2531a <=( A166  and  A167 );
 a2535a <=( A201  and  (not A200) );
 a2536a <=( A199  and  a2535a );
 a2537a <=( a2536a  and  a2531a );
 a2540a <=( A298  and  A202 );
 a2544a <=( A301  and  A300 );
 a2545a <=( (not A299)  and  a2544a );
 a2546a <=( a2545a  and  a2540a );
 a2549a <=( A166  and  A167 );
 a2553a <=( A201  and  (not A200) );
 a2554a <=( A199  and  a2553a );
 a2555a <=( a2554a  and  a2549a );
 a2558a <=( A298  and  A202 );
 a2562a <=( A302  and  A300 );
 a2563a <=( (not A299)  and  a2562a );
 a2564a <=( a2563a  and  a2558a );
 a2567a <=( A166  and  A167 );
 a2571a <=( A201  and  (not A200) );
 a2572a <=( A199  and  a2571a );
 a2573a <=( a2572a  and  a2567a );
 a2576a <=( (not A298)  and  A202 );
 a2580a <=( A301  and  A300 );
 a2581a <=( A299  and  a2580a );
 a2582a <=( a2581a  and  a2576a );
 a2585a <=( A166  and  A167 );
 a2589a <=( A201  and  (not A200) );
 a2590a <=( A199  and  a2589a );
 a2591a <=( a2590a  and  a2585a );
 a2594a <=( (not A298)  and  A202 );
 a2598a <=( A302  and  A300 );
 a2599a <=( A299  and  a2598a );
 a2600a <=( a2599a  and  a2594a );
 a2603a <=( A166  and  A167 );
 a2607a <=( A201  and  (not A200) );
 a2608a <=( A199  and  a2607a );
 a2609a <=( a2608a  and  a2603a );
 a2612a <=( A298  and  A203 );
 a2616a <=( A301  and  A300 );
 a2617a <=( (not A299)  and  a2616a );
 a2618a <=( a2617a  and  a2612a );
 a2621a <=( A166  and  A167 );
 a2625a <=( A201  and  (not A200) );
 a2626a <=( A199  and  a2625a );
 a2627a <=( a2626a  and  a2621a );
 a2630a <=( A298  and  A203 );
 a2634a <=( A302  and  A300 );
 a2635a <=( (not A299)  and  a2634a );
 a2636a <=( a2635a  and  a2630a );
 a2639a <=( A166  and  A167 );
 a2643a <=( A201  and  (not A200) );
 a2644a <=( A199  and  a2643a );
 a2645a <=( a2644a  and  a2639a );
 a2648a <=( (not A298)  and  A203 );
 a2652a <=( A301  and  A300 );
 a2653a <=( A299  and  a2652a );
 a2654a <=( a2653a  and  a2648a );
 a2657a <=( A166  and  A167 );
 a2661a <=( A201  and  (not A200) );
 a2662a <=( A199  and  a2661a );
 a2663a <=( a2662a  and  a2657a );
 a2666a <=( (not A298)  and  A203 );
 a2670a <=( A302  and  A300 );
 a2671a <=( A299  and  a2670a );
 a2672a <=( a2671a  and  a2666a );
 a2675a <=( (not A166)  and  (not A167) );
 a2679a <=( A201  and  A200 );
 a2680a <=( (not A199)  and  a2679a );
 a2681a <=( a2680a  and  a2675a );
 a2684a <=( A298  and  A202 );
 a2688a <=( A301  and  A300 );
 a2689a <=( (not A299)  and  a2688a );
 a2690a <=( a2689a  and  a2684a );
 a2693a <=( (not A166)  and  (not A167) );
 a2697a <=( A201  and  A200 );
 a2698a <=( (not A199)  and  a2697a );
 a2699a <=( a2698a  and  a2693a );
 a2702a <=( A298  and  A202 );
 a2706a <=( A302  and  A300 );
 a2707a <=( (not A299)  and  a2706a );
 a2708a <=( a2707a  and  a2702a );
 a2711a <=( (not A166)  and  (not A167) );
 a2715a <=( A201  and  A200 );
 a2716a <=( (not A199)  and  a2715a );
 a2717a <=( a2716a  and  a2711a );
 a2720a <=( (not A298)  and  A202 );
 a2724a <=( A301  and  A300 );
 a2725a <=( A299  and  a2724a );
 a2726a <=( a2725a  and  a2720a );
 a2729a <=( (not A166)  and  (not A167) );
 a2733a <=( A201  and  A200 );
 a2734a <=( (not A199)  and  a2733a );
 a2735a <=( a2734a  and  a2729a );
 a2738a <=( (not A298)  and  A202 );
 a2742a <=( A302  and  A300 );
 a2743a <=( A299  and  a2742a );
 a2744a <=( a2743a  and  a2738a );
 a2747a <=( (not A166)  and  (not A167) );
 a2751a <=( A201  and  A200 );
 a2752a <=( (not A199)  and  a2751a );
 a2753a <=( a2752a  and  a2747a );
 a2756a <=( A298  and  A203 );
 a2760a <=( A301  and  A300 );
 a2761a <=( (not A299)  and  a2760a );
 a2762a <=( a2761a  and  a2756a );
 a2765a <=( (not A166)  and  (not A167) );
 a2769a <=( A201  and  A200 );
 a2770a <=( (not A199)  and  a2769a );
 a2771a <=( a2770a  and  a2765a );
 a2774a <=( A298  and  A203 );
 a2778a <=( A302  and  A300 );
 a2779a <=( (not A299)  and  a2778a );
 a2780a <=( a2779a  and  a2774a );
 a2783a <=( (not A166)  and  (not A167) );
 a2787a <=( A201  and  A200 );
 a2788a <=( (not A199)  and  a2787a );
 a2789a <=( a2788a  and  a2783a );
 a2792a <=( (not A298)  and  A203 );
 a2796a <=( A301  and  A300 );
 a2797a <=( A299  and  a2796a );
 a2798a <=( a2797a  and  a2792a );
 a2801a <=( (not A166)  and  (not A167) );
 a2805a <=( A201  and  A200 );
 a2806a <=( (not A199)  and  a2805a );
 a2807a <=( a2806a  and  a2801a );
 a2810a <=( (not A298)  and  A203 );
 a2814a <=( A302  and  A300 );
 a2815a <=( A299  and  a2814a );
 a2816a <=( a2815a  and  a2810a );
 a2819a <=( (not A166)  and  (not A167) );
 a2823a <=( A201  and  (not A200) );
 a2824a <=( A199  and  a2823a );
 a2825a <=( a2824a  and  a2819a );
 a2828a <=( A298  and  A202 );
 a2832a <=( A301  and  A300 );
 a2833a <=( (not A299)  and  a2832a );
 a2834a <=( a2833a  and  a2828a );
 a2837a <=( (not A166)  and  (not A167) );
 a2841a <=( A201  and  (not A200) );
 a2842a <=( A199  and  a2841a );
 a2843a <=( a2842a  and  a2837a );
 a2846a <=( A298  and  A202 );
 a2850a <=( A302  and  A300 );
 a2851a <=( (not A299)  and  a2850a );
 a2852a <=( a2851a  and  a2846a );
 a2855a <=( (not A166)  and  (not A167) );
 a2859a <=( A201  and  (not A200) );
 a2860a <=( A199  and  a2859a );
 a2861a <=( a2860a  and  a2855a );
 a2864a <=( (not A298)  and  A202 );
 a2868a <=( A301  and  A300 );
 a2869a <=( A299  and  a2868a );
 a2870a <=( a2869a  and  a2864a );
 a2873a <=( (not A166)  and  (not A167) );
 a2877a <=( A201  and  (not A200) );
 a2878a <=( A199  and  a2877a );
 a2879a <=( a2878a  and  a2873a );
 a2882a <=( (not A298)  and  A202 );
 a2886a <=( A302  and  A300 );
 a2887a <=( A299  and  a2886a );
 a2888a <=( a2887a  and  a2882a );
 a2891a <=( (not A166)  and  (not A167) );
 a2895a <=( A201  and  (not A200) );
 a2896a <=( A199  and  a2895a );
 a2897a <=( a2896a  and  a2891a );
 a2900a <=( A298  and  A203 );
 a2904a <=( A301  and  A300 );
 a2905a <=( (not A299)  and  a2904a );
 a2906a <=( a2905a  and  a2900a );
 a2909a <=( (not A166)  and  (not A167) );
 a2913a <=( A201  and  (not A200) );
 a2914a <=( A199  and  a2913a );
 a2915a <=( a2914a  and  a2909a );
 a2918a <=( A298  and  A203 );
 a2922a <=( A302  and  A300 );
 a2923a <=( (not A299)  and  a2922a );
 a2924a <=( a2923a  and  a2918a );
 a2927a <=( (not A166)  and  (not A167) );
 a2931a <=( A201  and  (not A200) );
 a2932a <=( A199  and  a2931a );
 a2933a <=( a2932a  and  a2927a );
 a2936a <=( (not A298)  and  A203 );
 a2940a <=( A301  and  A300 );
 a2941a <=( A299  and  a2940a );
 a2942a <=( a2941a  and  a2936a );
 a2945a <=( (not A166)  and  (not A167) );
 a2949a <=( A201  and  (not A200) );
 a2950a <=( A199  and  a2949a );
 a2951a <=( a2950a  and  a2945a );
 a2954a <=( (not A298)  and  A203 );
 a2958a <=( A302  and  A300 );
 a2959a <=( A299  and  a2958a );
 a2960a <=( a2959a  and  a2954a );
 a2963a <=( A168  and  (not A170) );
 a2967a <=( (not A201)  and  (not A166) );
 a2968a <=( A167  and  a2967a );
 a2969a <=( a2968a  and  a2963a );
 a2972a <=( A298  and  A202 );
 a2976a <=( A301  and  A300 );
 a2977a <=( (not A299)  and  a2976a );
 a2978a <=( a2977a  and  a2972a );
 a2981a <=( A168  and  (not A170) );
 a2985a <=( (not A201)  and  (not A166) );
 a2986a <=( A167  and  a2985a );
 a2987a <=( a2986a  and  a2981a );
 a2990a <=( A298  and  A202 );
 a2994a <=( A302  and  A300 );
 a2995a <=( (not A299)  and  a2994a );
 a2996a <=( a2995a  and  a2990a );
 a2999a <=( A168  and  (not A170) );
 a3003a <=( (not A201)  and  (not A166) );
 a3004a <=( A167  and  a3003a );
 a3005a <=( a3004a  and  a2999a );
 a3008a <=( (not A298)  and  A202 );
 a3012a <=( A301  and  A300 );
 a3013a <=( A299  and  a3012a );
 a3014a <=( a3013a  and  a3008a );
 a3017a <=( A168  and  (not A170) );
 a3021a <=( (not A201)  and  (not A166) );
 a3022a <=( A167  and  a3021a );
 a3023a <=( a3022a  and  a3017a );
 a3026a <=( (not A298)  and  A202 );
 a3030a <=( A302  and  A300 );
 a3031a <=( A299  and  a3030a );
 a3032a <=( a3031a  and  a3026a );
 a3035a <=( A168  and  (not A170) );
 a3039a <=( (not A201)  and  (not A166) );
 a3040a <=( A167  and  a3039a );
 a3041a <=( a3040a  and  a3035a );
 a3044a <=( A298  and  A203 );
 a3048a <=( A301  and  A300 );
 a3049a <=( (not A299)  and  a3048a );
 a3050a <=( a3049a  and  a3044a );
 a3053a <=( A168  and  (not A170) );
 a3057a <=( (not A201)  and  (not A166) );
 a3058a <=( A167  and  a3057a );
 a3059a <=( a3058a  and  a3053a );
 a3062a <=( A298  and  A203 );
 a3066a <=( A302  and  A300 );
 a3067a <=( (not A299)  and  a3066a );
 a3068a <=( a3067a  and  a3062a );
 a3071a <=( A168  and  (not A170) );
 a3075a <=( (not A201)  and  (not A166) );
 a3076a <=( A167  and  a3075a );
 a3077a <=( a3076a  and  a3071a );
 a3080a <=( (not A298)  and  A203 );
 a3084a <=( A301  and  A300 );
 a3085a <=( A299  and  a3084a );
 a3086a <=( a3085a  and  a3080a );
 a3089a <=( A168  and  (not A170) );
 a3093a <=( (not A201)  and  (not A166) );
 a3094a <=( A167  and  a3093a );
 a3095a <=( a3094a  and  a3089a );
 a3098a <=( (not A298)  and  A203 );
 a3102a <=( A302  and  A300 );
 a3103a <=( A299  and  a3102a );
 a3104a <=( a3103a  and  a3098a );
 a3107a <=( A168  and  (not A170) );
 a3111a <=( A199  and  (not A166) );
 a3112a <=( A167  and  a3111a );
 a3113a <=( a3112a  and  a3107a );
 a3116a <=( A298  and  A200 );
 a3120a <=( A301  and  A300 );
 a3121a <=( (not A299)  and  a3120a );
 a3122a <=( a3121a  and  a3116a );
 a3125a <=( A168  and  (not A170) );
 a3129a <=( A199  and  (not A166) );
 a3130a <=( A167  and  a3129a );
 a3131a <=( a3130a  and  a3125a );
 a3134a <=( A298  and  A200 );
 a3138a <=( A302  and  A300 );
 a3139a <=( (not A299)  and  a3138a );
 a3140a <=( a3139a  and  a3134a );
 a3143a <=( A168  and  (not A170) );
 a3147a <=( A199  and  (not A166) );
 a3148a <=( A167  and  a3147a );
 a3149a <=( a3148a  and  a3143a );
 a3152a <=( (not A298)  and  A200 );
 a3156a <=( A301  and  A300 );
 a3157a <=( A299  and  a3156a );
 a3158a <=( a3157a  and  a3152a );
 a3161a <=( A168  and  (not A170) );
 a3165a <=( A199  and  (not A166) );
 a3166a <=( A167  and  a3165a );
 a3167a <=( a3166a  and  a3161a );
 a3170a <=( (not A298)  and  A200 );
 a3174a <=( A302  and  A300 );
 a3175a <=( A299  and  a3174a );
 a3176a <=( a3175a  and  a3170a );
 a3179a <=( A168  and  (not A170) );
 a3183a <=( (not A199)  and  (not A166) );
 a3184a <=( A167  and  a3183a );
 a3185a <=( a3184a  and  a3179a );
 a3188a <=( A298  and  (not A200) );
 a3192a <=( A301  and  A300 );
 a3193a <=( (not A299)  and  a3192a );
 a3194a <=( a3193a  and  a3188a );
 a3197a <=( A168  and  (not A170) );
 a3201a <=( (not A199)  and  (not A166) );
 a3202a <=( A167  and  a3201a );
 a3203a <=( a3202a  and  a3197a );
 a3206a <=( A298  and  (not A200) );
 a3210a <=( A302  and  A300 );
 a3211a <=( (not A299)  and  a3210a );
 a3212a <=( a3211a  and  a3206a );
 a3215a <=( A168  and  (not A170) );
 a3219a <=( (not A199)  and  (not A166) );
 a3220a <=( A167  and  a3219a );
 a3221a <=( a3220a  and  a3215a );
 a3224a <=( (not A298)  and  (not A200) );
 a3228a <=( A301  and  A300 );
 a3229a <=( A299  and  a3228a );
 a3230a <=( a3229a  and  a3224a );
 a3233a <=( A168  and  (not A170) );
 a3237a <=( (not A199)  and  (not A166) );
 a3238a <=( A167  and  a3237a );
 a3239a <=( a3238a  and  a3233a );
 a3242a <=( (not A298)  and  (not A200) );
 a3246a <=( A302  and  A300 );
 a3247a <=( A299  and  a3246a );
 a3248a <=( a3247a  and  a3242a );
 a3251a <=( A168  and  (not A170) );
 a3255a <=( (not A201)  and  A166 );
 a3256a <=( (not A167)  and  a3255a );
 a3257a <=( a3256a  and  a3251a );
 a3260a <=( A298  and  A202 );
 a3264a <=( A301  and  A300 );
 a3265a <=( (not A299)  and  a3264a );
 a3266a <=( a3265a  and  a3260a );
 a3269a <=( A168  and  (not A170) );
 a3273a <=( (not A201)  and  A166 );
 a3274a <=( (not A167)  and  a3273a );
 a3275a <=( a3274a  and  a3269a );
 a3278a <=( A298  and  A202 );
 a3282a <=( A302  and  A300 );
 a3283a <=( (not A299)  and  a3282a );
 a3284a <=( a3283a  and  a3278a );
 a3287a <=( A168  and  (not A170) );
 a3291a <=( (not A201)  and  A166 );
 a3292a <=( (not A167)  and  a3291a );
 a3293a <=( a3292a  and  a3287a );
 a3296a <=( (not A298)  and  A202 );
 a3300a <=( A301  and  A300 );
 a3301a <=( A299  and  a3300a );
 a3302a <=( a3301a  and  a3296a );
 a3305a <=( A168  and  (not A170) );
 a3309a <=( (not A201)  and  A166 );
 a3310a <=( (not A167)  and  a3309a );
 a3311a <=( a3310a  and  a3305a );
 a3314a <=( (not A298)  and  A202 );
 a3318a <=( A302  and  A300 );
 a3319a <=( A299  and  a3318a );
 a3320a <=( a3319a  and  a3314a );
 a3323a <=( A168  and  (not A170) );
 a3327a <=( (not A201)  and  A166 );
 a3328a <=( (not A167)  and  a3327a );
 a3329a <=( a3328a  and  a3323a );
 a3332a <=( A298  and  A203 );
 a3336a <=( A301  and  A300 );
 a3337a <=( (not A299)  and  a3336a );
 a3338a <=( a3337a  and  a3332a );
 a3341a <=( A168  and  (not A170) );
 a3345a <=( (not A201)  and  A166 );
 a3346a <=( (not A167)  and  a3345a );
 a3347a <=( a3346a  and  a3341a );
 a3350a <=( A298  and  A203 );
 a3354a <=( A302  and  A300 );
 a3355a <=( (not A299)  and  a3354a );
 a3356a <=( a3355a  and  a3350a );
 a3359a <=( A168  and  (not A170) );
 a3363a <=( (not A201)  and  A166 );
 a3364a <=( (not A167)  and  a3363a );
 a3365a <=( a3364a  and  a3359a );
 a3368a <=( (not A298)  and  A203 );
 a3372a <=( A301  and  A300 );
 a3373a <=( A299  and  a3372a );
 a3374a <=( a3373a  and  a3368a );
 a3377a <=( A168  and  (not A170) );
 a3381a <=( (not A201)  and  A166 );
 a3382a <=( (not A167)  and  a3381a );
 a3383a <=( a3382a  and  a3377a );
 a3386a <=( (not A298)  and  A203 );
 a3390a <=( A302  and  A300 );
 a3391a <=( A299  and  a3390a );
 a3392a <=( a3391a  and  a3386a );
 a3395a <=( A168  and  (not A170) );
 a3399a <=( A199  and  A166 );
 a3400a <=( (not A167)  and  a3399a );
 a3401a <=( a3400a  and  a3395a );
 a3404a <=( A298  and  A200 );
 a3408a <=( A301  and  A300 );
 a3409a <=( (not A299)  and  a3408a );
 a3410a <=( a3409a  and  a3404a );
 a3413a <=( A168  and  (not A170) );
 a3417a <=( A199  and  A166 );
 a3418a <=( (not A167)  and  a3417a );
 a3419a <=( a3418a  and  a3413a );
 a3422a <=( A298  and  A200 );
 a3426a <=( A302  and  A300 );
 a3427a <=( (not A299)  and  a3426a );
 a3428a <=( a3427a  and  a3422a );
 a3431a <=( A168  and  (not A170) );
 a3435a <=( A199  and  A166 );
 a3436a <=( (not A167)  and  a3435a );
 a3437a <=( a3436a  and  a3431a );
 a3440a <=( (not A298)  and  A200 );
 a3444a <=( A301  and  A300 );
 a3445a <=( A299  and  a3444a );
 a3446a <=( a3445a  and  a3440a );
 a3449a <=( A168  and  (not A170) );
 a3453a <=( A199  and  A166 );
 a3454a <=( (not A167)  and  a3453a );
 a3455a <=( a3454a  and  a3449a );
 a3458a <=( (not A298)  and  A200 );
 a3462a <=( A302  and  A300 );
 a3463a <=( A299  and  a3462a );
 a3464a <=( a3463a  and  a3458a );
 a3467a <=( A168  and  (not A170) );
 a3471a <=( (not A199)  and  A166 );
 a3472a <=( (not A167)  and  a3471a );
 a3473a <=( a3472a  and  a3467a );
 a3476a <=( A298  and  (not A200) );
 a3480a <=( A301  and  A300 );
 a3481a <=( (not A299)  and  a3480a );
 a3482a <=( a3481a  and  a3476a );
 a3485a <=( A168  and  (not A170) );
 a3489a <=( (not A199)  and  A166 );
 a3490a <=( (not A167)  and  a3489a );
 a3491a <=( a3490a  and  a3485a );
 a3494a <=( A298  and  (not A200) );
 a3498a <=( A302  and  A300 );
 a3499a <=( (not A299)  and  a3498a );
 a3500a <=( a3499a  and  a3494a );
 a3503a <=( A168  and  (not A170) );
 a3507a <=( (not A199)  and  A166 );
 a3508a <=( (not A167)  and  a3507a );
 a3509a <=( a3508a  and  a3503a );
 a3512a <=( (not A298)  and  (not A200) );
 a3516a <=( A301  and  A300 );
 a3517a <=( A299  and  a3516a );
 a3518a <=( a3517a  and  a3512a );
 a3521a <=( A168  and  (not A170) );
 a3525a <=( (not A199)  and  A166 );
 a3526a <=( (not A167)  and  a3525a );
 a3527a <=( a3526a  and  a3521a );
 a3530a <=( (not A298)  and  (not A200) );
 a3534a <=( A302  and  A300 );
 a3535a <=( A299  and  a3534a );
 a3536a <=( a3535a  and  a3530a );
 a3539a <=( (not A168)  and  (not A170) );
 a3543a <=( A201  and  A200 );
 a3544a <=( (not A199)  and  a3543a );
 a3545a <=( a3544a  and  a3539a );
 a3548a <=( A298  and  A202 );
 a3552a <=( A301  and  A300 );
 a3553a <=( (not A299)  and  a3552a );
 a3554a <=( a3553a  and  a3548a );
 a3557a <=( (not A168)  and  (not A170) );
 a3561a <=( A201  and  A200 );
 a3562a <=( (not A199)  and  a3561a );
 a3563a <=( a3562a  and  a3557a );
 a3566a <=( A298  and  A202 );
 a3570a <=( A302  and  A300 );
 a3571a <=( (not A299)  and  a3570a );
 a3572a <=( a3571a  and  a3566a );
 a3575a <=( (not A168)  and  (not A170) );
 a3579a <=( A201  and  A200 );
 a3580a <=( (not A199)  and  a3579a );
 a3581a <=( a3580a  and  a3575a );
 a3584a <=( (not A298)  and  A202 );
 a3588a <=( A301  and  A300 );
 a3589a <=( A299  and  a3588a );
 a3590a <=( a3589a  and  a3584a );
 a3593a <=( (not A168)  and  (not A170) );
 a3597a <=( A201  and  A200 );
 a3598a <=( (not A199)  and  a3597a );
 a3599a <=( a3598a  and  a3593a );
 a3602a <=( (not A298)  and  A202 );
 a3606a <=( A302  and  A300 );
 a3607a <=( A299  and  a3606a );
 a3608a <=( a3607a  and  a3602a );
 a3611a <=( (not A168)  and  (not A170) );
 a3615a <=( A201  and  A200 );
 a3616a <=( (not A199)  and  a3615a );
 a3617a <=( a3616a  and  a3611a );
 a3620a <=( A298  and  A203 );
 a3624a <=( A301  and  A300 );
 a3625a <=( (not A299)  and  a3624a );
 a3626a <=( a3625a  and  a3620a );
 a3629a <=( (not A168)  and  (not A170) );
 a3633a <=( A201  and  A200 );
 a3634a <=( (not A199)  and  a3633a );
 a3635a <=( a3634a  and  a3629a );
 a3638a <=( A298  and  A203 );
 a3642a <=( A302  and  A300 );
 a3643a <=( (not A299)  and  a3642a );
 a3644a <=( a3643a  and  a3638a );
 a3647a <=( (not A168)  and  (not A170) );
 a3651a <=( A201  and  A200 );
 a3652a <=( (not A199)  and  a3651a );
 a3653a <=( a3652a  and  a3647a );
 a3656a <=( (not A298)  and  A203 );
 a3660a <=( A301  and  A300 );
 a3661a <=( A299  and  a3660a );
 a3662a <=( a3661a  and  a3656a );
 a3665a <=( (not A168)  and  (not A170) );
 a3669a <=( A201  and  A200 );
 a3670a <=( (not A199)  and  a3669a );
 a3671a <=( a3670a  and  a3665a );
 a3674a <=( (not A298)  and  A203 );
 a3678a <=( A302  and  A300 );
 a3679a <=( A299  and  a3678a );
 a3680a <=( a3679a  and  a3674a );
 a3683a <=( (not A168)  and  (not A170) );
 a3687a <=( A201  and  (not A200) );
 a3688a <=( A199  and  a3687a );
 a3689a <=( a3688a  and  a3683a );
 a3692a <=( A298  and  A202 );
 a3696a <=( A301  and  A300 );
 a3697a <=( (not A299)  and  a3696a );
 a3698a <=( a3697a  and  a3692a );
 a3701a <=( (not A168)  and  (not A170) );
 a3705a <=( A201  and  (not A200) );
 a3706a <=( A199  and  a3705a );
 a3707a <=( a3706a  and  a3701a );
 a3710a <=( A298  and  A202 );
 a3714a <=( A302  and  A300 );
 a3715a <=( (not A299)  and  a3714a );
 a3716a <=( a3715a  and  a3710a );
 a3719a <=( (not A168)  and  (not A170) );
 a3723a <=( A201  and  (not A200) );
 a3724a <=( A199  and  a3723a );
 a3725a <=( a3724a  and  a3719a );
 a3728a <=( (not A298)  and  A202 );
 a3732a <=( A301  and  A300 );
 a3733a <=( A299  and  a3732a );
 a3734a <=( a3733a  and  a3728a );
 a3737a <=( (not A168)  and  (not A170) );
 a3741a <=( A201  and  (not A200) );
 a3742a <=( A199  and  a3741a );
 a3743a <=( a3742a  and  a3737a );
 a3746a <=( (not A298)  and  A202 );
 a3750a <=( A302  and  A300 );
 a3751a <=( A299  and  a3750a );
 a3752a <=( a3751a  and  a3746a );
 a3755a <=( (not A168)  and  (not A170) );
 a3759a <=( A201  and  (not A200) );
 a3760a <=( A199  and  a3759a );
 a3761a <=( a3760a  and  a3755a );
 a3764a <=( A298  and  A203 );
 a3768a <=( A301  and  A300 );
 a3769a <=( (not A299)  and  a3768a );
 a3770a <=( a3769a  and  a3764a );
 a3773a <=( (not A168)  and  (not A170) );
 a3777a <=( A201  and  (not A200) );
 a3778a <=( A199  and  a3777a );
 a3779a <=( a3778a  and  a3773a );
 a3782a <=( A298  and  A203 );
 a3786a <=( A302  and  A300 );
 a3787a <=( (not A299)  and  a3786a );
 a3788a <=( a3787a  and  a3782a );
 a3791a <=( (not A168)  and  (not A170) );
 a3795a <=( A201  and  (not A200) );
 a3796a <=( A199  and  a3795a );
 a3797a <=( a3796a  and  a3791a );
 a3800a <=( (not A298)  and  A203 );
 a3804a <=( A301  and  A300 );
 a3805a <=( A299  and  a3804a );
 a3806a <=( a3805a  and  a3800a );
 a3809a <=( (not A168)  and  (not A170) );
 a3813a <=( A201  and  (not A200) );
 a3814a <=( A199  and  a3813a );
 a3815a <=( a3814a  and  a3809a );
 a3818a <=( (not A298)  and  A203 );
 a3822a <=( A302  and  A300 );
 a3823a <=( A299  and  a3822a );
 a3824a <=( a3823a  and  a3818a );
 a3827a <=( A168  and  A169 );
 a3831a <=( (not A201)  and  (not A166) );
 a3832a <=( A167  and  a3831a );
 a3833a <=( a3832a  and  a3827a );
 a3836a <=( A298  and  A202 );
 a3840a <=( A301  and  A300 );
 a3841a <=( (not A299)  and  a3840a );
 a3842a <=( a3841a  and  a3836a );
 a3845a <=( A168  and  A169 );
 a3849a <=( (not A201)  and  (not A166) );
 a3850a <=( A167  and  a3849a );
 a3851a <=( a3850a  and  a3845a );
 a3854a <=( A298  and  A202 );
 a3858a <=( A302  and  A300 );
 a3859a <=( (not A299)  and  a3858a );
 a3860a <=( a3859a  and  a3854a );
 a3863a <=( A168  and  A169 );
 a3867a <=( (not A201)  and  (not A166) );
 a3868a <=( A167  and  a3867a );
 a3869a <=( a3868a  and  a3863a );
 a3872a <=( (not A298)  and  A202 );
 a3876a <=( A301  and  A300 );
 a3877a <=( A299  and  a3876a );
 a3878a <=( a3877a  and  a3872a );
 a3881a <=( A168  and  A169 );
 a3885a <=( (not A201)  and  (not A166) );
 a3886a <=( A167  and  a3885a );
 a3887a <=( a3886a  and  a3881a );
 a3890a <=( (not A298)  and  A202 );
 a3894a <=( A302  and  A300 );
 a3895a <=( A299  and  a3894a );
 a3896a <=( a3895a  and  a3890a );
 a3899a <=( A168  and  A169 );
 a3903a <=( (not A201)  and  (not A166) );
 a3904a <=( A167  and  a3903a );
 a3905a <=( a3904a  and  a3899a );
 a3908a <=( A298  and  A203 );
 a3912a <=( A301  and  A300 );
 a3913a <=( (not A299)  and  a3912a );
 a3914a <=( a3913a  and  a3908a );
 a3917a <=( A168  and  A169 );
 a3921a <=( (not A201)  and  (not A166) );
 a3922a <=( A167  and  a3921a );
 a3923a <=( a3922a  and  a3917a );
 a3926a <=( A298  and  A203 );
 a3930a <=( A302  and  A300 );
 a3931a <=( (not A299)  and  a3930a );
 a3932a <=( a3931a  and  a3926a );
 a3935a <=( A168  and  A169 );
 a3939a <=( (not A201)  and  (not A166) );
 a3940a <=( A167  and  a3939a );
 a3941a <=( a3940a  and  a3935a );
 a3944a <=( (not A298)  and  A203 );
 a3948a <=( A301  and  A300 );
 a3949a <=( A299  and  a3948a );
 a3950a <=( a3949a  and  a3944a );
 a3953a <=( A168  and  A169 );
 a3957a <=( (not A201)  and  (not A166) );
 a3958a <=( A167  and  a3957a );
 a3959a <=( a3958a  and  a3953a );
 a3962a <=( (not A298)  and  A203 );
 a3966a <=( A302  and  A300 );
 a3967a <=( A299  and  a3966a );
 a3968a <=( a3967a  and  a3962a );
 a3971a <=( A168  and  A169 );
 a3975a <=( A199  and  (not A166) );
 a3976a <=( A167  and  a3975a );
 a3977a <=( a3976a  and  a3971a );
 a3980a <=( A298  and  A200 );
 a3984a <=( A301  and  A300 );
 a3985a <=( (not A299)  and  a3984a );
 a3986a <=( a3985a  and  a3980a );
 a3989a <=( A168  and  A169 );
 a3993a <=( A199  and  (not A166) );
 a3994a <=( A167  and  a3993a );
 a3995a <=( a3994a  and  a3989a );
 a3998a <=( A298  and  A200 );
 a4002a <=( A302  and  A300 );
 a4003a <=( (not A299)  and  a4002a );
 a4004a <=( a4003a  and  a3998a );
 a4007a <=( A168  and  A169 );
 a4011a <=( A199  and  (not A166) );
 a4012a <=( A167  and  a4011a );
 a4013a <=( a4012a  and  a4007a );
 a4016a <=( (not A298)  and  A200 );
 a4020a <=( A301  and  A300 );
 a4021a <=( A299  and  a4020a );
 a4022a <=( a4021a  and  a4016a );
 a4025a <=( A168  and  A169 );
 a4029a <=( A199  and  (not A166) );
 a4030a <=( A167  and  a4029a );
 a4031a <=( a4030a  and  a4025a );
 a4034a <=( (not A298)  and  A200 );
 a4038a <=( A302  and  A300 );
 a4039a <=( A299  and  a4038a );
 a4040a <=( a4039a  and  a4034a );
 a4043a <=( A168  and  A169 );
 a4047a <=( (not A199)  and  (not A166) );
 a4048a <=( A167  and  a4047a );
 a4049a <=( a4048a  and  a4043a );
 a4052a <=( A298  and  (not A200) );
 a4056a <=( A301  and  A300 );
 a4057a <=( (not A299)  and  a4056a );
 a4058a <=( a4057a  and  a4052a );
 a4061a <=( A168  and  A169 );
 a4065a <=( (not A199)  and  (not A166) );
 a4066a <=( A167  and  a4065a );
 a4067a <=( a4066a  and  a4061a );
 a4070a <=( A298  and  (not A200) );
 a4074a <=( A302  and  A300 );
 a4075a <=( (not A299)  and  a4074a );
 a4076a <=( a4075a  and  a4070a );
 a4079a <=( A168  and  A169 );
 a4083a <=( (not A199)  and  (not A166) );
 a4084a <=( A167  and  a4083a );
 a4085a <=( a4084a  and  a4079a );
 a4088a <=( (not A298)  and  (not A200) );
 a4092a <=( A301  and  A300 );
 a4093a <=( A299  and  a4092a );
 a4094a <=( a4093a  and  a4088a );
 a4097a <=( A168  and  A169 );
 a4101a <=( (not A199)  and  (not A166) );
 a4102a <=( A167  and  a4101a );
 a4103a <=( a4102a  and  a4097a );
 a4106a <=( (not A298)  and  (not A200) );
 a4110a <=( A302  and  A300 );
 a4111a <=( A299  and  a4110a );
 a4112a <=( a4111a  and  a4106a );
 a4115a <=( A168  and  A169 );
 a4119a <=( (not A201)  and  A166 );
 a4120a <=( (not A167)  and  a4119a );
 a4121a <=( a4120a  and  a4115a );
 a4124a <=( A298  and  A202 );
 a4128a <=( A301  and  A300 );
 a4129a <=( (not A299)  and  a4128a );
 a4130a <=( a4129a  and  a4124a );
 a4133a <=( A168  and  A169 );
 a4137a <=( (not A201)  and  A166 );
 a4138a <=( (not A167)  and  a4137a );
 a4139a <=( a4138a  and  a4133a );
 a4142a <=( A298  and  A202 );
 a4146a <=( A302  and  A300 );
 a4147a <=( (not A299)  and  a4146a );
 a4148a <=( a4147a  and  a4142a );
 a4151a <=( A168  and  A169 );
 a4155a <=( (not A201)  and  A166 );
 a4156a <=( (not A167)  and  a4155a );
 a4157a <=( a4156a  and  a4151a );
 a4160a <=( (not A298)  and  A202 );
 a4164a <=( A301  and  A300 );
 a4165a <=( A299  and  a4164a );
 a4166a <=( a4165a  and  a4160a );
 a4169a <=( A168  and  A169 );
 a4173a <=( (not A201)  and  A166 );
 a4174a <=( (not A167)  and  a4173a );
 a4175a <=( a4174a  and  a4169a );
 a4178a <=( (not A298)  and  A202 );
 a4182a <=( A302  and  A300 );
 a4183a <=( A299  and  a4182a );
 a4184a <=( a4183a  and  a4178a );
 a4187a <=( A168  and  A169 );
 a4191a <=( (not A201)  and  A166 );
 a4192a <=( (not A167)  and  a4191a );
 a4193a <=( a4192a  and  a4187a );
 a4196a <=( A298  and  A203 );
 a4200a <=( A301  and  A300 );
 a4201a <=( (not A299)  and  a4200a );
 a4202a <=( a4201a  and  a4196a );
 a4205a <=( A168  and  A169 );
 a4209a <=( (not A201)  and  A166 );
 a4210a <=( (not A167)  and  a4209a );
 a4211a <=( a4210a  and  a4205a );
 a4214a <=( A298  and  A203 );
 a4218a <=( A302  and  A300 );
 a4219a <=( (not A299)  and  a4218a );
 a4220a <=( a4219a  and  a4214a );
 a4223a <=( A168  and  A169 );
 a4227a <=( (not A201)  and  A166 );
 a4228a <=( (not A167)  and  a4227a );
 a4229a <=( a4228a  and  a4223a );
 a4232a <=( (not A298)  and  A203 );
 a4236a <=( A301  and  A300 );
 a4237a <=( A299  and  a4236a );
 a4238a <=( a4237a  and  a4232a );
 a4241a <=( A168  and  A169 );
 a4245a <=( (not A201)  and  A166 );
 a4246a <=( (not A167)  and  a4245a );
 a4247a <=( a4246a  and  a4241a );
 a4250a <=( (not A298)  and  A203 );
 a4254a <=( A302  and  A300 );
 a4255a <=( A299  and  a4254a );
 a4256a <=( a4255a  and  a4250a );
 a4259a <=( A168  and  A169 );
 a4263a <=( A199  and  A166 );
 a4264a <=( (not A167)  and  a4263a );
 a4265a <=( a4264a  and  a4259a );
 a4268a <=( A298  and  A200 );
 a4272a <=( A301  and  A300 );
 a4273a <=( (not A299)  and  a4272a );
 a4274a <=( a4273a  and  a4268a );
 a4277a <=( A168  and  A169 );
 a4281a <=( A199  and  A166 );
 a4282a <=( (not A167)  and  a4281a );
 a4283a <=( a4282a  and  a4277a );
 a4286a <=( A298  and  A200 );
 a4290a <=( A302  and  A300 );
 a4291a <=( (not A299)  and  a4290a );
 a4292a <=( a4291a  and  a4286a );
 a4295a <=( A168  and  A169 );
 a4299a <=( A199  and  A166 );
 a4300a <=( (not A167)  and  a4299a );
 a4301a <=( a4300a  and  a4295a );
 a4304a <=( (not A298)  and  A200 );
 a4308a <=( A301  and  A300 );
 a4309a <=( A299  and  a4308a );
 a4310a <=( a4309a  and  a4304a );
 a4313a <=( A168  and  A169 );
 a4317a <=( A199  and  A166 );
 a4318a <=( (not A167)  and  a4317a );
 a4319a <=( a4318a  and  a4313a );
 a4322a <=( (not A298)  and  A200 );
 a4326a <=( A302  and  A300 );
 a4327a <=( A299  and  a4326a );
 a4328a <=( a4327a  and  a4322a );
 a4331a <=( A168  and  A169 );
 a4335a <=( (not A199)  and  A166 );
 a4336a <=( (not A167)  and  a4335a );
 a4337a <=( a4336a  and  a4331a );
 a4340a <=( A298  and  (not A200) );
 a4344a <=( A301  and  A300 );
 a4345a <=( (not A299)  and  a4344a );
 a4346a <=( a4345a  and  a4340a );
 a4349a <=( A168  and  A169 );
 a4353a <=( (not A199)  and  A166 );
 a4354a <=( (not A167)  and  a4353a );
 a4355a <=( a4354a  and  a4349a );
 a4358a <=( A298  and  (not A200) );
 a4362a <=( A302  and  A300 );
 a4363a <=( (not A299)  and  a4362a );
 a4364a <=( a4363a  and  a4358a );
 a4367a <=( A168  and  A169 );
 a4371a <=( (not A199)  and  A166 );
 a4372a <=( (not A167)  and  a4371a );
 a4373a <=( a4372a  and  a4367a );
 a4376a <=( (not A298)  and  (not A200) );
 a4380a <=( A301  and  A300 );
 a4381a <=( A299  and  a4380a );
 a4382a <=( a4381a  and  a4376a );
 a4385a <=( A168  and  A169 );
 a4389a <=( (not A199)  and  A166 );
 a4390a <=( (not A167)  and  a4389a );
 a4391a <=( a4390a  and  a4385a );
 a4394a <=( (not A298)  and  (not A200) );
 a4398a <=( A302  and  A300 );
 a4399a <=( A299  and  a4398a );
 a4400a <=( a4399a  and  a4394a );
 a4403a <=( (not A168)  and  A169 );
 a4407a <=( A201  and  A200 );
 a4408a <=( (not A199)  and  a4407a );
 a4409a <=( a4408a  and  a4403a );
 a4412a <=( A298  and  A202 );
 a4416a <=( A301  and  A300 );
 a4417a <=( (not A299)  and  a4416a );
 a4418a <=( a4417a  and  a4412a );
 a4421a <=( (not A168)  and  A169 );
 a4425a <=( A201  and  A200 );
 a4426a <=( (not A199)  and  a4425a );
 a4427a <=( a4426a  and  a4421a );
 a4430a <=( A298  and  A202 );
 a4434a <=( A302  and  A300 );
 a4435a <=( (not A299)  and  a4434a );
 a4436a <=( a4435a  and  a4430a );
 a4439a <=( (not A168)  and  A169 );
 a4443a <=( A201  and  A200 );
 a4444a <=( (not A199)  and  a4443a );
 a4445a <=( a4444a  and  a4439a );
 a4448a <=( (not A298)  and  A202 );
 a4452a <=( A301  and  A300 );
 a4453a <=( A299  and  a4452a );
 a4454a <=( a4453a  and  a4448a );
 a4457a <=( (not A168)  and  A169 );
 a4461a <=( A201  and  A200 );
 a4462a <=( (not A199)  and  a4461a );
 a4463a <=( a4462a  and  a4457a );
 a4466a <=( (not A298)  and  A202 );
 a4470a <=( A302  and  A300 );
 a4471a <=( A299  and  a4470a );
 a4472a <=( a4471a  and  a4466a );
 a4475a <=( (not A168)  and  A169 );
 a4479a <=( A201  and  A200 );
 a4480a <=( (not A199)  and  a4479a );
 a4481a <=( a4480a  and  a4475a );
 a4484a <=( A298  and  A203 );
 a4488a <=( A301  and  A300 );
 a4489a <=( (not A299)  and  a4488a );
 a4490a <=( a4489a  and  a4484a );
 a4493a <=( (not A168)  and  A169 );
 a4497a <=( A201  and  A200 );
 a4498a <=( (not A199)  and  a4497a );
 a4499a <=( a4498a  and  a4493a );
 a4502a <=( A298  and  A203 );
 a4506a <=( A302  and  A300 );
 a4507a <=( (not A299)  and  a4506a );
 a4508a <=( a4507a  and  a4502a );
 a4511a <=( (not A168)  and  A169 );
 a4515a <=( A201  and  A200 );
 a4516a <=( (not A199)  and  a4515a );
 a4517a <=( a4516a  and  a4511a );
 a4520a <=( (not A298)  and  A203 );
 a4524a <=( A301  and  A300 );
 a4525a <=( A299  and  a4524a );
 a4526a <=( a4525a  and  a4520a );
 a4529a <=( (not A168)  and  A169 );
 a4533a <=( A201  and  A200 );
 a4534a <=( (not A199)  and  a4533a );
 a4535a <=( a4534a  and  a4529a );
 a4538a <=( (not A298)  and  A203 );
 a4542a <=( A302  and  A300 );
 a4543a <=( A299  and  a4542a );
 a4544a <=( a4543a  and  a4538a );
 a4547a <=( (not A168)  and  A169 );
 a4551a <=( A201  and  (not A200) );
 a4552a <=( A199  and  a4551a );
 a4553a <=( a4552a  and  a4547a );
 a4556a <=( A298  and  A202 );
 a4560a <=( A301  and  A300 );
 a4561a <=( (not A299)  and  a4560a );
 a4562a <=( a4561a  and  a4556a );
 a4565a <=( (not A168)  and  A169 );
 a4569a <=( A201  and  (not A200) );
 a4570a <=( A199  and  a4569a );
 a4571a <=( a4570a  and  a4565a );
 a4574a <=( A298  and  A202 );
 a4578a <=( A302  and  A300 );
 a4579a <=( (not A299)  and  a4578a );
 a4580a <=( a4579a  and  a4574a );
 a4583a <=( (not A168)  and  A169 );
 a4587a <=( A201  and  (not A200) );
 a4588a <=( A199  and  a4587a );
 a4589a <=( a4588a  and  a4583a );
 a4592a <=( (not A298)  and  A202 );
 a4596a <=( A301  and  A300 );
 a4597a <=( A299  and  a4596a );
 a4598a <=( a4597a  and  a4592a );
 a4601a <=( (not A168)  and  A169 );
 a4605a <=( A201  and  (not A200) );
 a4606a <=( A199  and  a4605a );
 a4607a <=( a4606a  and  a4601a );
 a4610a <=( (not A298)  and  A202 );
 a4614a <=( A302  and  A300 );
 a4615a <=( A299  and  a4614a );
 a4616a <=( a4615a  and  a4610a );
 a4619a <=( (not A168)  and  A169 );
 a4623a <=( A201  and  (not A200) );
 a4624a <=( A199  and  a4623a );
 a4625a <=( a4624a  and  a4619a );
 a4628a <=( A298  and  A203 );
 a4632a <=( A301  and  A300 );
 a4633a <=( (not A299)  and  a4632a );
 a4634a <=( a4633a  and  a4628a );
 a4637a <=( (not A168)  and  A169 );
 a4641a <=( A201  and  (not A200) );
 a4642a <=( A199  and  a4641a );
 a4643a <=( a4642a  and  a4637a );
 a4646a <=( A298  and  A203 );
 a4650a <=( A302  and  A300 );
 a4651a <=( (not A299)  and  a4650a );
 a4652a <=( a4651a  and  a4646a );
 a4655a <=( (not A168)  and  A169 );
 a4659a <=( A201  and  (not A200) );
 a4660a <=( A199  and  a4659a );
 a4661a <=( a4660a  and  a4655a );
 a4664a <=( (not A298)  and  A203 );
 a4668a <=( A301  and  A300 );
 a4669a <=( A299  and  a4668a );
 a4670a <=( a4669a  and  a4664a );
 a4673a <=( (not A168)  and  A169 );
 a4677a <=( A201  and  (not A200) );
 a4678a <=( A199  and  a4677a );
 a4679a <=( a4678a  and  a4673a );
 a4682a <=( (not A298)  and  A203 );
 a4686a <=( A302  and  A300 );
 a4687a <=( A299  and  a4686a );
 a4688a <=( a4687a  and  a4682a );
 a4691a <=( (not A169)  and  A170 );
 a4695a <=( (not A166)  and  A167 );
 a4696a <=( (not A168)  and  a4695a );
 a4697a <=( a4696a  and  a4691a );
 a4700a <=( A233  and  (not A232) );
 a4704a <=( (not A236)  and  (not A235) );
 a4705a <=( (not A234)  and  a4704a );
 a4706a <=( a4705a  and  a4700a );
 a4709a <=( (not A169)  and  A170 );
 a4713a <=( (not A166)  and  A167 );
 a4714a <=( (not A168)  and  a4713a );
 a4715a <=( a4714a  and  a4709a );
 a4718a <=( (not A233)  and  A232 );
 a4722a <=( (not A236)  and  (not A235) );
 a4723a <=( (not A234)  and  a4722a );
 a4724a <=( a4723a  and  a4718a );
 a4727a <=( (not A169)  and  A170 );
 a4731a <=( A166  and  (not A167) );
 a4732a <=( (not A168)  and  a4731a );
 a4733a <=( a4732a  and  a4727a );
 a4736a <=( A233  and  (not A232) );
 a4740a <=( (not A236)  and  (not A235) );
 a4741a <=( (not A234)  and  a4740a );
 a4742a <=( a4741a  and  a4736a );
 a4745a <=( (not A169)  and  A170 );
 a4749a <=( A166  and  (not A167) );
 a4750a <=( (not A168)  and  a4749a );
 a4751a <=( a4750a  and  a4745a );
 a4754a <=( (not A233)  and  A232 );
 a4758a <=( (not A236)  and  (not A235) );
 a4759a <=( (not A234)  and  a4758a );
 a4760a <=( a4759a  and  a4754a );
 a4763a <=( A166  and  A167 );
 a4767a <=( A201  and  A200 );
 a4768a <=( (not A199)  and  a4767a );
 a4769a <=( a4768a  and  a4763a );
 a4773a <=( (not A299)  and  A298 );
 a4774a <=( A202  and  a4773a );
 a4778a <=( (not A302)  and  (not A301) );
 a4779a <=( (not A300)  and  a4778a );
 a4780a <=( a4779a  and  a4774a );
 a4783a <=( A166  and  A167 );
 a4787a <=( A201  and  A200 );
 a4788a <=( (not A199)  and  a4787a );
 a4789a <=( a4788a  and  a4783a );
 a4793a <=( A299  and  (not A298) );
 a4794a <=( A202  and  a4793a );
 a4798a <=( (not A302)  and  (not A301) );
 a4799a <=( (not A300)  and  a4798a );
 a4800a <=( a4799a  and  a4794a );
 a4803a <=( A166  and  A167 );
 a4807a <=( A201  and  A200 );
 a4808a <=( (not A199)  and  a4807a );
 a4809a <=( a4808a  and  a4803a );
 a4813a <=( (not A299)  and  A298 );
 a4814a <=( A203  and  a4813a );
 a4818a <=( (not A302)  and  (not A301) );
 a4819a <=( (not A300)  and  a4818a );
 a4820a <=( a4819a  and  a4814a );
 a4823a <=( A166  and  A167 );
 a4827a <=( A201  and  A200 );
 a4828a <=( (not A199)  and  a4827a );
 a4829a <=( a4828a  and  a4823a );
 a4833a <=( A299  and  (not A298) );
 a4834a <=( A203  and  a4833a );
 a4838a <=( (not A302)  and  (not A301) );
 a4839a <=( (not A300)  and  a4838a );
 a4840a <=( a4839a  and  a4834a );
 a4843a <=( A166  and  A167 );
 a4847a <=( (not A201)  and  A200 );
 a4848a <=( (not A199)  and  a4847a );
 a4849a <=( a4848a  and  a4843a );
 a4853a <=( A298  and  (not A203) );
 a4854a <=( (not A202)  and  a4853a );
 a4858a <=( A301  and  A300 );
 a4859a <=( (not A299)  and  a4858a );
 a4860a <=( a4859a  and  a4854a );
 a4863a <=( A166  and  A167 );
 a4867a <=( (not A201)  and  A200 );
 a4868a <=( (not A199)  and  a4867a );
 a4869a <=( a4868a  and  a4863a );
 a4873a <=( A298  and  (not A203) );
 a4874a <=( (not A202)  and  a4873a );
 a4878a <=( A302  and  A300 );
 a4879a <=( (not A299)  and  a4878a );
 a4880a <=( a4879a  and  a4874a );
 a4883a <=( A166  and  A167 );
 a4887a <=( (not A201)  and  A200 );
 a4888a <=( (not A199)  and  a4887a );
 a4889a <=( a4888a  and  a4883a );
 a4893a <=( (not A298)  and  (not A203) );
 a4894a <=( (not A202)  and  a4893a );
 a4898a <=( A301  and  A300 );
 a4899a <=( A299  and  a4898a );
 a4900a <=( a4899a  and  a4894a );
 a4903a <=( A166  and  A167 );
 a4907a <=( (not A201)  and  A200 );
 a4908a <=( (not A199)  and  a4907a );
 a4909a <=( a4908a  and  a4903a );
 a4913a <=( (not A298)  and  (not A203) );
 a4914a <=( (not A202)  and  a4913a );
 a4918a <=( A302  and  A300 );
 a4919a <=( A299  and  a4918a );
 a4920a <=( a4919a  and  a4914a );
 a4923a <=( A166  and  A167 );
 a4927a <=( A201  and  (not A200) );
 a4928a <=( A199  and  a4927a );
 a4929a <=( a4928a  and  a4923a );
 a4933a <=( (not A299)  and  A298 );
 a4934a <=( A202  and  a4933a );
 a4938a <=( (not A302)  and  (not A301) );
 a4939a <=( (not A300)  and  a4938a );
 a4940a <=( a4939a  and  a4934a );
 a4943a <=( A166  and  A167 );
 a4947a <=( A201  and  (not A200) );
 a4948a <=( A199  and  a4947a );
 a4949a <=( a4948a  and  a4943a );
 a4953a <=( A299  and  (not A298) );
 a4954a <=( A202  and  a4953a );
 a4958a <=( (not A302)  and  (not A301) );
 a4959a <=( (not A300)  and  a4958a );
 a4960a <=( a4959a  and  a4954a );
 a4963a <=( A166  and  A167 );
 a4967a <=( A201  and  (not A200) );
 a4968a <=( A199  and  a4967a );
 a4969a <=( a4968a  and  a4963a );
 a4973a <=( (not A299)  and  A298 );
 a4974a <=( A203  and  a4973a );
 a4978a <=( (not A302)  and  (not A301) );
 a4979a <=( (not A300)  and  a4978a );
 a4980a <=( a4979a  and  a4974a );
 a4983a <=( A166  and  A167 );
 a4987a <=( A201  and  (not A200) );
 a4988a <=( A199  and  a4987a );
 a4989a <=( a4988a  and  a4983a );
 a4993a <=( A299  and  (not A298) );
 a4994a <=( A203  and  a4993a );
 a4998a <=( (not A302)  and  (not A301) );
 a4999a <=( (not A300)  and  a4998a );
 a5000a <=( a4999a  and  a4994a );
 a5003a <=( A166  and  A167 );
 a5007a <=( (not A201)  and  (not A200) );
 a5008a <=( A199  and  a5007a );
 a5009a <=( a5008a  and  a5003a );
 a5013a <=( A298  and  (not A203) );
 a5014a <=( (not A202)  and  a5013a );
 a5018a <=( A301  and  A300 );
 a5019a <=( (not A299)  and  a5018a );
 a5020a <=( a5019a  and  a5014a );
 a5023a <=( A166  and  A167 );
 a5027a <=( (not A201)  and  (not A200) );
 a5028a <=( A199  and  a5027a );
 a5029a <=( a5028a  and  a5023a );
 a5033a <=( A298  and  (not A203) );
 a5034a <=( (not A202)  and  a5033a );
 a5038a <=( A302  and  A300 );
 a5039a <=( (not A299)  and  a5038a );
 a5040a <=( a5039a  and  a5034a );
 a5043a <=( A166  and  A167 );
 a5047a <=( (not A201)  and  (not A200) );
 a5048a <=( A199  and  a5047a );
 a5049a <=( a5048a  and  a5043a );
 a5053a <=( (not A298)  and  (not A203) );
 a5054a <=( (not A202)  and  a5053a );
 a5058a <=( A301  and  A300 );
 a5059a <=( A299  and  a5058a );
 a5060a <=( a5059a  and  a5054a );
 a5063a <=( A166  and  A167 );
 a5067a <=( (not A201)  and  (not A200) );
 a5068a <=( A199  and  a5067a );
 a5069a <=( a5068a  and  a5063a );
 a5073a <=( (not A298)  and  (not A203) );
 a5074a <=( (not A202)  and  a5073a );
 a5078a <=( A302  and  A300 );
 a5079a <=( A299  and  a5078a );
 a5080a <=( a5079a  and  a5074a );
 a5083a <=( (not A166)  and  (not A167) );
 a5087a <=( A201  and  A200 );
 a5088a <=( (not A199)  and  a5087a );
 a5089a <=( a5088a  and  a5083a );
 a5093a <=( (not A299)  and  A298 );
 a5094a <=( A202  and  a5093a );
 a5098a <=( (not A302)  and  (not A301) );
 a5099a <=( (not A300)  and  a5098a );
 a5100a <=( a5099a  and  a5094a );
 a5103a <=( (not A166)  and  (not A167) );
 a5107a <=( A201  and  A200 );
 a5108a <=( (not A199)  and  a5107a );
 a5109a <=( a5108a  and  a5103a );
 a5113a <=( A299  and  (not A298) );
 a5114a <=( A202  and  a5113a );
 a5118a <=( (not A302)  and  (not A301) );
 a5119a <=( (not A300)  and  a5118a );
 a5120a <=( a5119a  and  a5114a );
 a5123a <=( (not A166)  and  (not A167) );
 a5127a <=( A201  and  A200 );
 a5128a <=( (not A199)  and  a5127a );
 a5129a <=( a5128a  and  a5123a );
 a5133a <=( (not A299)  and  A298 );
 a5134a <=( A203  and  a5133a );
 a5138a <=( (not A302)  and  (not A301) );
 a5139a <=( (not A300)  and  a5138a );
 a5140a <=( a5139a  and  a5134a );
 a5143a <=( (not A166)  and  (not A167) );
 a5147a <=( A201  and  A200 );
 a5148a <=( (not A199)  and  a5147a );
 a5149a <=( a5148a  and  a5143a );
 a5153a <=( A299  and  (not A298) );
 a5154a <=( A203  and  a5153a );
 a5158a <=( (not A302)  and  (not A301) );
 a5159a <=( (not A300)  and  a5158a );
 a5160a <=( a5159a  and  a5154a );
 a5163a <=( (not A166)  and  (not A167) );
 a5167a <=( (not A201)  and  A200 );
 a5168a <=( (not A199)  and  a5167a );
 a5169a <=( a5168a  and  a5163a );
 a5173a <=( A298  and  (not A203) );
 a5174a <=( (not A202)  and  a5173a );
 a5178a <=( A301  and  A300 );
 a5179a <=( (not A299)  and  a5178a );
 a5180a <=( a5179a  and  a5174a );
 a5183a <=( (not A166)  and  (not A167) );
 a5187a <=( (not A201)  and  A200 );
 a5188a <=( (not A199)  and  a5187a );
 a5189a <=( a5188a  and  a5183a );
 a5193a <=( A298  and  (not A203) );
 a5194a <=( (not A202)  and  a5193a );
 a5198a <=( A302  and  A300 );
 a5199a <=( (not A299)  and  a5198a );
 a5200a <=( a5199a  and  a5194a );
 a5203a <=( (not A166)  and  (not A167) );
 a5207a <=( (not A201)  and  A200 );
 a5208a <=( (not A199)  and  a5207a );
 a5209a <=( a5208a  and  a5203a );
 a5213a <=( (not A298)  and  (not A203) );
 a5214a <=( (not A202)  and  a5213a );
 a5218a <=( A301  and  A300 );
 a5219a <=( A299  and  a5218a );
 a5220a <=( a5219a  and  a5214a );
 a5223a <=( (not A166)  and  (not A167) );
 a5227a <=( (not A201)  and  A200 );
 a5228a <=( (not A199)  and  a5227a );
 a5229a <=( a5228a  and  a5223a );
 a5233a <=( (not A298)  and  (not A203) );
 a5234a <=( (not A202)  and  a5233a );
 a5238a <=( A302  and  A300 );
 a5239a <=( A299  and  a5238a );
 a5240a <=( a5239a  and  a5234a );
 a5243a <=( (not A166)  and  (not A167) );
 a5247a <=( A201  and  (not A200) );
 a5248a <=( A199  and  a5247a );
 a5249a <=( a5248a  and  a5243a );
 a5253a <=( (not A299)  and  A298 );
 a5254a <=( A202  and  a5253a );
 a5258a <=( (not A302)  and  (not A301) );
 a5259a <=( (not A300)  and  a5258a );
 a5260a <=( a5259a  and  a5254a );
 a5263a <=( (not A166)  and  (not A167) );
 a5267a <=( A201  and  (not A200) );
 a5268a <=( A199  and  a5267a );
 a5269a <=( a5268a  and  a5263a );
 a5273a <=( A299  and  (not A298) );
 a5274a <=( A202  and  a5273a );
 a5278a <=( (not A302)  and  (not A301) );
 a5279a <=( (not A300)  and  a5278a );
 a5280a <=( a5279a  and  a5274a );
 a5283a <=( (not A166)  and  (not A167) );
 a5287a <=( A201  and  (not A200) );
 a5288a <=( A199  and  a5287a );
 a5289a <=( a5288a  and  a5283a );
 a5293a <=( (not A299)  and  A298 );
 a5294a <=( A203  and  a5293a );
 a5298a <=( (not A302)  and  (not A301) );
 a5299a <=( (not A300)  and  a5298a );
 a5300a <=( a5299a  and  a5294a );
 a5303a <=( (not A166)  and  (not A167) );
 a5307a <=( A201  and  (not A200) );
 a5308a <=( A199  and  a5307a );
 a5309a <=( a5308a  and  a5303a );
 a5313a <=( A299  and  (not A298) );
 a5314a <=( A203  and  a5313a );
 a5318a <=( (not A302)  and  (not A301) );
 a5319a <=( (not A300)  and  a5318a );
 a5320a <=( a5319a  and  a5314a );
 a5323a <=( (not A166)  and  (not A167) );
 a5327a <=( (not A201)  and  (not A200) );
 a5328a <=( A199  and  a5327a );
 a5329a <=( a5328a  and  a5323a );
 a5333a <=( A298  and  (not A203) );
 a5334a <=( (not A202)  and  a5333a );
 a5338a <=( A301  and  A300 );
 a5339a <=( (not A299)  and  a5338a );
 a5340a <=( a5339a  and  a5334a );
 a5343a <=( (not A166)  and  (not A167) );
 a5347a <=( (not A201)  and  (not A200) );
 a5348a <=( A199  and  a5347a );
 a5349a <=( a5348a  and  a5343a );
 a5353a <=( A298  and  (not A203) );
 a5354a <=( (not A202)  and  a5353a );
 a5358a <=( A302  and  A300 );
 a5359a <=( (not A299)  and  a5358a );
 a5360a <=( a5359a  and  a5354a );
 a5363a <=( (not A166)  and  (not A167) );
 a5367a <=( (not A201)  and  (not A200) );
 a5368a <=( A199  and  a5367a );
 a5369a <=( a5368a  and  a5363a );
 a5373a <=( (not A298)  and  (not A203) );
 a5374a <=( (not A202)  and  a5373a );
 a5378a <=( A301  and  A300 );
 a5379a <=( A299  and  a5378a );
 a5380a <=( a5379a  and  a5374a );
 a5383a <=( (not A166)  and  (not A167) );
 a5387a <=( (not A201)  and  (not A200) );
 a5388a <=( A199  and  a5387a );
 a5389a <=( a5388a  and  a5383a );
 a5393a <=( (not A298)  and  (not A203) );
 a5394a <=( (not A202)  and  a5393a );
 a5398a <=( A302  and  A300 );
 a5399a <=( A299  and  a5398a );
 a5400a <=( a5399a  and  a5394a );
 a5403a <=( A168  and  (not A170) );
 a5407a <=( A201  and  (not A166) );
 a5408a <=( A167  and  a5407a );
 a5409a <=( a5408a  and  a5403a );
 a5413a <=( A298  and  (not A203) );
 a5414a <=( (not A202)  and  a5413a );
 a5418a <=( A301  and  A300 );
 a5419a <=( (not A299)  and  a5418a );
 a5420a <=( a5419a  and  a5414a );
 a5423a <=( A168  and  (not A170) );
 a5427a <=( A201  and  (not A166) );
 a5428a <=( A167  and  a5427a );
 a5429a <=( a5428a  and  a5423a );
 a5433a <=( A298  and  (not A203) );
 a5434a <=( (not A202)  and  a5433a );
 a5438a <=( A302  and  A300 );
 a5439a <=( (not A299)  and  a5438a );
 a5440a <=( a5439a  and  a5434a );
 a5443a <=( A168  and  (not A170) );
 a5447a <=( A201  and  (not A166) );
 a5448a <=( A167  and  a5447a );
 a5449a <=( a5448a  and  a5443a );
 a5453a <=( (not A298)  and  (not A203) );
 a5454a <=( (not A202)  and  a5453a );
 a5458a <=( A301  and  A300 );
 a5459a <=( A299  and  a5458a );
 a5460a <=( a5459a  and  a5454a );
 a5463a <=( A168  and  (not A170) );
 a5467a <=( A201  and  (not A166) );
 a5468a <=( A167  and  a5467a );
 a5469a <=( a5468a  and  a5463a );
 a5473a <=( (not A298)  and  (not A203) );
 a5474a <=( (not A202)  and  a5473a );
 a5478a <=( A302  and  A300 );
 a5479a <=( A299  and  a5478a );
 a5480a <=( a5479a  and  a5474a );
 a5483a <=( A168  and  (not A170) );
 a5487a <=( (not A201)  and  (not A166) );
 a5488a <=( A167  and  a5487a );
 a5489a <=( a5488a  and  a5483a );
 a5493a <=( (not A299)  and  A298 );
 a5494a <=( A202  and  a5493a );
 a5498a <=( (not A302)  and  (not A301) );
 a5499a <=( (not A300)  and  a5498a );
 a5500a <=( a5499a  and  a5494a );
 a5503a <=( A168  and  (not A170) );
 a5507a <=( (not A201)  and  (not A166) );
 a5508a <=( A167  and  a5507a );
 a5509a <=( a5508a  and  a5503a );
 a5513a <=( A299  and  (not A298) );
 a5514a <=( A202  and  a5513a );
 a5518a <=( (not A302)  and  (not A301) );
 a5519a <=( (not A300)  and  a5518a );
 a5520a <=( a5519a  and  a5514a );
 a5523a <=( A168  and  (not A170) );
 a5527a <=( (not A201)  and  (not A166) );
 a5528a <=( A167  and  a5527a );
 a5529a <=( a5528a  and  a5523a );
 a5533a <=( (not A299)  and  A298 );
 a5534a <=( A203  and  a5533a );
 a5538a <=( (not A302)  and  (not A301) );
 a5539a <=( (not A300)  and  a5538a );
 a5540a <=( a5539a  and  a5534a );
 a5543a <=( A168  and  (not A170) );
 a5547a <=( (not A201)  and  (not A166) );
 a5548a <=( A167  and  a5547a );
 a5549a <=( a5548a  and  a5543a );
 a5553a <=( A299  and  (not A298) );
 a5554a <=( A203  and  a5553a );
 a5558a <=( (not A302)  and  (not A301) );
 a5559a <=( (not A300)  and  a5558a );
 a5560a <=( a5559a  and  a5554a );
 a5563a <=( A168  and  (not A170) );
 a5567a <=( A199  and  (not A166) );
 a5568a <=( A167  and  a5567a );
 a5569a <=( a5568a  and  a5563a );
 a5573a <=( (not A299)  and  A298 );
 a5574a <=( A200  and  a5573a );
 a5578a <=( (not A302)  and  (not A301) );
 a5579a <=( (not A300)  and  a5578a );
 a5580a <=( a5579a  and  a5574a );
 a5583a <=( A168  and  (not A170) );
 a5587a <=( A199  and  (not A166) );
 a5588a <=( A167  and  a5587a );
 a5589a <=( a5588a  and  a5583a );
 a5593a <=( A299  and  (not A298) );
 a5594a <=( A200  and  a5593a );
 a5598a <=( (not A302)  and  (not A301) );
 a5599a <=( (not A300)  and  a5598a );
 a5600a <=( a5599a  and  a5594a );
 a5603a <=( A168  and  (not A170) );
 a5607a <=( (not A199)  and  (not A166) );
 a5608a <=( A167  and  a5607a );
 a5609a <=( a5608a  and  a5603a );
 a5613a <=( (not A299)  and  A298 );
 a5614a <=( (not A200)  and  a5613a );
 a5618a <=( (not A302)  and  (not A301) );
 a5619a <=( (not A300)  and  a5618a );
 a5620a <=( a5619a  and  a5614a );
 a5623a <=( A168  and  (not A170) );
 a5627a <=( (not A199)  and  (not A166) );
 a5628a <=( A167  and  a5627a );
 a5629a <=( a5628a  and  a5623a );
 a5633a <=( A299  and  (not A298) );
 a5634a <=( (not A200)  and  a5633a );
 a5638a <=( (not A302)  and  (not A301) );
 a5639a <=( (not A300)  and  a5638a );
 a5640a <=( a5639a  and  a5634a );
 a5643a <=( A168  and  (not A170) );
 a5647a <=( A201  and  A166 );
 a5648a <=( (not A167)  and  a5647a );
 a5649a <=( a5648a  and  a5643a );
 a5653a <=( A298  and  (not A203) );
 a5654a <=( (not A202)  and  a5653a );
 a5658a <=( A301  and  A300 );
 a5659a <=( (not A299)  and  a5658a );
 a5660a <=( a5659a  and  a5654a );
 a5663a <=( A168  and  (not A170) );
 a5667a <=( A201  and  A166 );
 a5668a <=( (not A167)  and  a5667a );
 a5669a <=( a5668a  and  a5663a );
 a5673a <=( A298  and  (not A203) );
 a5674a <=( (not A202)  and  a5673a );
 a5678a <=( A302  and  A300 );
 a5679a <=( (not A299)  and  a5678a );
 a5680a <=( a5679a  and  a5674a );
 a5683a <=( A168  and  (not A170) );
 a5687a <=( A201  and  A166 );
 a5688a <=( (not A167)  and  a5687a );
 a5689a <=( a5688a  and  a5683a );
 a5693a <=( (not A298)  and  (not A203) );
 a5694a <=( (not A202)  and  a5693a );
 a5698a <=( A301  and  A300 );
 a5699a <=( A299  and  a5698a );
 a5700a <=( a5699a  and  a5694a );
 a5703a <=( A168  and  (not A170) );
 a5707a <=( A201  and  A166 );
 a5708a <=( (not A167)  and  a5707a );
 a5709a <=( a5708a  and  a5703a );
 a5713a <=( (not A298)  and  (not A203) );
 a5714a <=( (not A202)  and  a5713a );
 a5718a <=( A302  and  A300 );
 a5719a <=( A299  and  a5718a );
 a5720a <=( a5719a  and  a5714a );
 a5723a <=( A168  and  (not A170) );
 a5727a <=( (not A201)  and  A166 );
 a5728a <=( (not A167)  and  a5727a );
 a5729a <=( a5728a  and  a5723a );
 a5733a <=( (not A299)  and  A298 );
 a5734a <=( A202  and  a5733a );
 a5738a <=( (not A302)  and  (not A301) );
 a5739a <=( (not A300)  and  a5738a );
 a5740a <=( a5739a  and  a5734a );
 a5743a <=( A168  and  (not A170) );
 a5747a <=( (not A201)  and  A166 );
 a5748a <=( (not A167)  and  a5747a );
 a5749a <=( a5748a  and  a5743a );
 a5753a <=( A299  and  (not A298) );
 a5754a <=( A202  and  a5753a );
 a5758a <=( (not A302)  and  (not A301) );
 a5759a <=( (not A300)  and  a5758a );
 a5760a <=( a5759a  and  a5754a );
 a5763a <=( A168  and  (not A170) );
 a5767a <=( (not A201)  and  A166 );
 a5768a <=( (not A167)  and  a5767a );
 a5769a <=( a5768a  and  a5763a );
 a5773a <=( (not A299)  and  A298 );
 a5774a <=( A203  and  a5773a );
 a5778a <=( (not A302)  and  (not A301) );
 a5779a <=( (not A300)  and  a5778a );
 a5780a <=( a5779a  and  a5774a );
 a5783a <=( A168  and  (not A170) );
 a5787a <=( (not A201)  and  A166 );
 a5788a <=( (not A167)  and  a5787a );
 a5789a <=( a5788a  and  a5783a );
 a5793a <=( A299  and  (not A298) );
 a5794a <=( A203  and  a5793a );
 a5798a <=( (not A302)  and  (not A301) );
 a5799a <=( (not A300)  and  a5798a );
 a5800a <=( a5799a  and  a5794a );
 a5803a <=( A168  and  (not A170) );
 a5807a <=( A199  and  A166 );
 a5808a <=( (not A167)  and  a5807a );
 a5809a <=( a5808a  and  a5803a );
 a5813a <=( (not A299)  and  A298 );
 a5814a <=( A200  and  a5813a );
 a5818a <=( (not A302)  and  (not A301) );
 a5819a <=( (not A300)  and  a5818a );
 a5820a <=( a5819a  and  a5814a );
 a5823a <=( A168  and  (not A170) );
 a5827a <=( A199  and  A166 );
 a5828a <=( (not A167)  and  a5827a );
 a5829a <=( a5828a  and  a5823a );
 a5833a <=( A299  and  (not A298) );
 a5834a <=( A200  and  a5833a );
 a5838a <=( (not A302)  and  (not A301) );
 a5839a <=( (not A300)  and  a5838a );
 a5840a <=( a5839a  and  a5834a );
 a5843a <=( A168  and  (not A170) );
 a5847a <=( (not A199)  and  A166 );
 a5848a <=( (not A167)  and  a5847a );
 a5849a <=( a5848a  and  a5843a );
 a5853a <=( (not A299)  and  A298 );
 a5854a <=( (not A200)  and  a5853a );
 a5858a <=( (not A302)  and  (not A301) );
 a5859a <=( (not A300)  and  a5858a );
 a5860a <=( a5859a  and  a5854a );
 a5863a <=( A168  and  (not A170) );
 a5867a <=( (not A199)  and  A166 );
 a5868a <=( (not A167)  and  a5867a );
 a5869a <=( a5868a  and  a5863a );
 a5873a <=( A299  and  (not A298) );
 a5874a <=( (not A200)  and  a5873a );
 a5878a <=( (not A302)  and  (not A301) );
 a5879a <=( (not A300)  and  a5878a );
 a5880a <=( a5879a  and  a5874a );
 a5883a <=( (not A168)  and  (not A170) );
 a5887a <=( A201  and  A200 );
 a5888a <=( (not A199)  and  a5887a );
 a5889a <=( a5888a  and  a5883a );
 a5893a <=( (not A299)  and  A298 );
 a5894a <=( A202  and  a5893a );
 a5898a <=( (not A302)  and  (not A301) );
 a5899a <=( (not A300)  and  a5898a );
 a5900a <=( a5899a  and  a5894a );
 a5903a <=( (not A168)  and  (not A170) );
 a5907a <=( A201  and  A200 );
 a5908a <=( (not A199)  and  a5907a );
 a5909a <=( a5908a  and  a5903a );
 a5913a <=( A299  and  (not A298) );
 a5914a <=( A202  and  a5913a );
 a5918a <=( (not A302)  and  (not A301) );
 a5919a <=( (not A300)  and  a5918a );
 a5920a <=( a5919a  and  a5914a );
 a5923a <=( (not A168)  and  (not A170) );
 a5927a <=( A201  and  A200 );
 a5928a <=( (not A199)  and  a5927a );
 a5929a <=( a5928a  and  a5923a );
 a5933a <=( (not A299)  and  A298 );
 a5934a <=( A203  and  a5933a );
 a5938a <=( (not A302)  and  (not A301) );
 a5939a <=( (not A300)  and  a5938a );
 a5940a <=( a5939a  and  a5934a );
 a5943a <=( (not A168)  and  (not A170) );
 a5947a <=( A201  and  A200 );
 a5948a <=( (not A199)  and  a5947a );
 a5949a <=( a5948a  and  a5943a );
 a5953a <=( A299  and  (not A298) );
 a5954a <=( A203  and  a5953a );
 a5958a <=( (not A302)  and  (not A301) );
 a5959a <=( (not A300)  and  a5958a );
 a5960a <=( a5959a  and  a5954a );
 a5963a <=( (not A168)  and  (not A170) );
 a5967a <=( (not A201)  and  A200 );
 a5968a <=( (not A199)  and  a5967a );
 a5969a <=( a5968a  and  a5963a );
 a5973a <=( A298  and  (not A203) );
 a5974a <=( (not A202)  and  a5973a );
 a5978a <=( A301  and  A300 );
 a5979a <=( (not A299)  and  a5978a );
 a5980a <=( a5979a  and  a5974a );
 a5983a <=( (not A168)  and  (not A170) );
 a5987a <=( (not A201)  and  A200 );
 a5988a <=( (not A199)  and  a5987a );
 a5989a <=( a5988a  and  a5983a );
 a5993a <=( A298  and  (not A203) );
 a5994a <=( (not A202)  and  a5993a );
 a5998a <=( A302  and  A300 );
 a5999a <=( (not A299)  and  a5998a );
 a6000a <=( a5999a  and  a5994a );
 a6003a <=( (not A168)  and  (not A170) );
 a6007a <=( (not A201)  and  A200 );
 a6008a <=( (not A199)  and  a6007a );
 a6009a <=( a6008a  and  a6003a );
 a6013a <=( (not A298)  and  (not A203) );
 a6014a <=( (not A202)  and  a6013a );
 a6018a <=( A301  and  A300 );
 a6019a <=( A299  and  a6018a );
 a6020a <=( a6019a  and  a6014a );
 a6023a <=( (not A168)  and  (not A170) );
 a6027a <=( (not A201)  and  A200 );
 a6028a <=( (not A199)  and  a6027a );
 a6029a <=( a6028a  and  a6023a );
 a6033a <=( (not A298)  and  (not A203) );
 a6034a <=( (not A202)  and  a6033a );
 a6038a <=( A302  and  A300 );
 a6039a <=( A299  and  a6038a );
 a6040a <=( a6039a  and  a6034a );
 a6043a <=( (not A168)  and  (not A170) );
 a6047a <=( A201  and  (not A200) );
 a6048a <=( A199  and  a6047a );
 a6049a <=( a6048a  and  a6043a );
 a6053a <=( (not A299)  and  A298 );
 a6054a <=( A202  and  a6053a );
 a6058a <=( (not A302)  and  (not A301) );
 a6059a <=( (not A300)  and  a6058a );
 a6060a <=( a6059a  and  a6054a );
 a6063a <=( (not A168)  and  (not A170) );
 a6067a <=( A201  and  (not A200) );
 a6068a <=( A199  and  a6067a );
 a6069a <=( a6068a  and  a6063a );
 a6073a <=( A299  and  (not A298) );
 a6074a <=( A202  and  a6073a );
 a6078a <=( (not A302)  and  (not A301) );
 a6079a <=( (not A300)  and  a6078a );
 a6080a <=( a6079a  and  a6074a );
 a6083a <=( (not A168)  and  (not A170) );
 a6087a <=( A201  and  (not A200) );
 a6088a <=( A199  and  a6087a );
 a6089a <=( a6088a  and  a6083a );
 a6093a <=( (not A299)  and  A298 );
 a6094a <=( A203  and  a6093a );
 a6098a <=( (not A302)  and  (not A301) );
 a6099a <=( (not A300)  and  a6098a );
 a6100a <=( a6099a  and  a6094a );
 a6103a <=( (not A168)  and  (not A170) );
 a6107a <=( A201  and  (not A200) );
 a6108a <=( A199  and  a6107a );
 a6109a <=( a6108a  and  a6103a );
 a6113a <=( A299  and  (not A298) );
 a6114a <=( A203  and  a6113a );
 a6118a <=( (not A302)  and  (not A301) );
 a6119a <=( (not A300)  and  a6118a );
 a6120a <=( a6119a  and  a6114a );
 a6123a <=( (not A168)  and  (not A170) );
 a6127a <=( (not A201)  and  (not A200) );
 a6128a <=( A199  and  a6127a );
 a6129a <=( a6128a  and  a6123a );
 a6133a <=( A298  and  (not A203) );
 a6134a <=( (not A202)  and  a6133a );
 a6138a <=( A301  and  A300 );
 a6139a <=( (not A299)  and  a6138a );
 a6140a <=( a6139a  and  a6134a );
 a6143a <=( (not A168)  and  (not A170) );
 a6147a <=( (not A201)  and  (not A200) );
 a6148a <=( A199  and  a6147a );
 a6149a <=( a6148a  and  a6143a );
 a6153a <=( A298  and  (not A203) );
 a6154a <=( (not A202)  and  a6153a );
 a6158a <=( A302  and  A300 );
 a6159a <=( (not A299)  and  a6158a );
 a6160a <=( a6159a  and  a6154a );
 a6163a <=( (not A168)  and  (not A170) );
 a6167a <=( (not A201)  and  (not A200) );
 a6168a <=( A199  and  a6167a );
 a6169a <=( a6168a  and  a6163a );
 a6173a <=( (not A298)  and  (not A203) );
 a6174a <=( (not A202)  and  a6173a );
 a6178a <=( A301  and  A300 );
 a6179a <=( A299  and  a6178a );
 a6180a <=( a6179a  and  a6174a );
 a6183a <=( (not A168)  and  (not A170) );
 a6187a <=( (not A201)  and  (not A200) );
 a6188a <=( A199  and  a6187a );
 a6189a <=( a6188a  and  a6183a );
 a6193a <=( (not A298)  and  (not A203) );
 a6194a <=( (not A202)  and  a6193a );
 a6198a <=( A302  and  A300 );
 a6199a <=( A299  and  a6198a );
 a6200a <=( a6199a  and  a6194a );
 a6203a <=( A168  and  A169 );
 a6207a <=( A201  and  (not A166) );
 a6208a <=( A167  and  a6207a );
 a6209a <=( a6208a  and  a6203a );
 a6213a <=( A298  and  (not A203) );
 a6214a <=( (not A202)  and  a6213a );
 a6218a <=( A301  and  A300 );
 a6219a <=( (not A299)  and  a6218a );
 a6220a <=( a6219a  and  a6214a );
 a6223a <=( A168  and  A169 );
 a6227a <=( A201  and  (not A166) );
 a6228a <=( A167  and  a6227a );
 a6229a <=( a6228a  and  a6223a );
 a6233a <=( A298  and  (not A203) );
 a6234a <=( (not A202)  and  a6233a );
 a6238a <=( A302  and  A300 );
 a6239a <=( (not A299)  and  a6238a );
 a6240a <=( a6239a  and  a6234a );
 a6243a <=( A168  and  A169 );
 a6247a <=( A201  and  (not A166) );
 a6248a <=( A167  and  a6247a );
 a6249a <=( a6248a  and  a6243a );
 a6253a <=( (not A298)  and  (not A203) );
 a6254a <=( (not A202)  and  a6253a );
 a6258a <=( A301  and  A300 );
 a6259a <=( A299  and  a6258a );
 a6260a <=( a6259a  and  a6254a );
 a6263a <=( A168  and  A169 );
 a6267a <=( A201  and  (not A166) );
 a6268a <=( A167  and  a6267a );
 a6269a <=( a6268a  and  a6263a );
 a6273a <=( (not A298)  and  (not A203) );
 a6274a <=( (not A202)  and  a6273a );
 a6278a <=( A302  and  A300 );
 a6279a <=( A299  and  a6278a );
 a6280a <=( a6279a  and  a6274a );
 a6283a <=( A168  and  A169 );
 a6287a <=( (not A201)  and  (not A166) );
 a6288a <=( A167  and  a6287a );
 a6289a <=( a6288a  and  a6283a );
 a6293a <=( (not A299)  and  A298 );
 a6294a <=( A202  and  a6293a );
 a6298a <=( (not A302)  and  (not A301) );
 a6299a <=( (not A300)  and  a6298a );
 a6300a <=( a6299a  and  a6294a );
 a6303a <=( A168  and  A169 );
 a6307a <=( (not A201)  and  (not A166) );
 a6308a <=( A167  and  a6307a );
 a6309a <=( a6308a  and  a6303a );
 a6313a <=( A299  and  (not A298) );
 a6314a <=( A202  and  a6313a );
 a6318a <=( (not A302)  and  (not A301) );
 a6319a <=( (not A300)  and  a6318a );
 a6320a <=( a6319a  and  a6314a );
 a6323a <=( A168  and  A169 );
 a6327a <=( (not A201)  and  (not A166) );
 a6328a <=( A167  and  a6327a );
 a6329a <=( a6328a  and  a6323a );
 a6333a <=( (not A299)  and  A298 );
 a6334a <=( A203  and  a6333a );
 a6338a <=( (not A302)  and  (not A301) );
 a6339a <=( (not A300)  and  a6338a );
 a6340a <=( a6339a  and  a6334a );
 a6343a <=( A168  and  A169 );
 a6347a <=( (not A201)  and  (not A166) );
 a6348a <=( A167  and  a6347a );
 a6349a <=( a6348a  and  a6343a );
 a6353a <=( A299  and  (not A298) );
 a6354a <=( A203  and  a6353a );
 a6358a <=( (not A302)  and  (not A301) );
 a6359a <=( (not A300)  and  a6358a );
 a6360a <=( a6359a  and  a6354a );
 a6363a <=( A168  and  A169 );
 a6367a <=( A199  and  (not A166) );
 a6368a <=( A167  and  a6367a );
 a6369a <=( a6368a  and  a6363a );
 a6373a <=( (not A299)  and  A298 );
 a6374a <=( A200  and  a6373a );
 a6378a <=( (not A302)  and  (not A301) );
 a6379a <=( (not A300)  and  a6378a );
 a6380a <=( a6379a  and  a6374a );
 a6383a <=( A168  and  A169 );
 a6387a <=( A199  and  (not A166) );
 a6388a <=( A167  and  a6387a );
 a6389a <=( a6388a  and  a6383a );
 a6393a <=( A299  and  (not A298) );
 a6394a <=( A200  and  a6393a );
 a6398a <=( (not A302)  and  (not A301) );
 a6399a <=( (not A300)  and  a6398a );
 a6400a <=( a6399a  and  a6394a );
 a6403a <=( A168  and  A169 );
 a6407a <=( (not A199)  and  (not A166) );
 a6408a <=( A167  and  a6407a );
 a6409a <=( a6408a  and  a6403a );
 a6413a <=( (not A299)  and  A298 );
 a6414a <=( (not A200)  and  a6413a );
 a6418a <=( (not A302)  and  (not A301) );
 a6419a <=( (not A300)  and  a6418a );
 a6420a <=( a6419a  and  a6414a );
 a6423a <=( A168  and  A169 );
 a6427a <=( (not A199)  and  (not A166) );
 a6428a <=( A167  and  a6427a );
 a6429a <=( a6428a  and  a6423a );
 a6433a <=( A299  and  (not A298) );
 a6434a <=( (not A200)  and  a6433a );
 a6438a <=( (not A302)  and  (not A301) );
 a6439a <=( (not A300)  and  a6438a );
 a6440a <=( a6439a  and  a6434a );
 a6443a <=( A168  and  A169 );
 a6447a <=( A201  and  A166 );
 a6448a <=( (not A167)  and  a6447a );
 a6449a <=( a6448a  and  a6443a );
 a6453a <=( A298  and  (not A203) );
 a6454a <=( (not A202)  and  a6453a );
 a6458a <=( A301  and  A300 );
 a6459a <=( (not A299)  and  a6458a );
 a6460a <=( a6459a  and  a6454a );
 a6463a <=( A168  and  A169 );
 a6467a <=( A201  and  A166 );
 a6468a <=( (not A167)  and  a6467a );
 a6469a <=( a6468a  and  a6463a );
 a6473a <=( A298  and  (not A203) );
 a6474a <=( (not A202)  and  a6473a );
 a6478a <=( A302  and  A300 );
 a6479a <=( (not A299)  and  a6478a );
 a6480a <=( a6479a  and  a6474a );
 a6483a <=( A168  and  A169 );
 a6487a <=( A201  and  A166 );
 a6488a <=( (not A167)  and  a6487a );
 a6489a <=( a6488a  and  a6483a );
 a6493a <=( (not A298)  and  (not A203) );
 a6494a <=( (not A202)  and  a6493a );
 a6498a <=( A301  and  A300 );
 a6499a <=( A299  and  a6498a );
 a6500a <=( a6499a  and  a6494a );
 a6503a <=( A168  and  A169 );
 a6507a <=( A201  and  A166 );
 a6508a <=( (not A167)  and  a6507a );
 a6509a <=( a6508a  and  a6503a );
 a6513a <=( (not A298)  and  (not A203) );
 a6514a <=( (not A202)  and  a6513a );
 a6518a <=( A302  and  A300 );
 a6519a <=( A299  and  a6518a );
 a6520a <=( a6519a  and  a6514a );
 a6523a <=( A168  and  A169 );
 a6527a <=( (not A201)  and  A166 );
 a6528a <=( (not A167)  and  a6527a );
 a6529a <=( a6528a  and  a6523a );
 a6533a <=( (not A299)  and  A298 );
 a6534a <=( A202  and  a6533a );
 a6538a <=( (not A302)  and  (not A301) );
 a6539a <=( (not A300)  and  a6538a );
 a6540a <=( a6539a  and  a6534a );
 a6543a <=( A168  and  A169 );
 a6547a <=( (not A201)  and  A166 );
 a6548a <=( (not A167)  and  a6547a );
 a6549a <=( a6548a  and  a6543a );
 a6553a <=( A299  and  (not A298) );
 a6554a <=( A202  and  a6553a );
 a6558a <=( (not A302)  and  (not A301) );
 a6559a <=( (not A300)  and  a6558a );
 a6560a <=( a6559a  and  a6554a );
 a6563a <=( A168  and  A169 );
 a6567a <=( (not A201)  and  A166 );
 a6568a <=( (not A167)  and  a6567a );
 a6569a <=( a6568a  and  a6563a );
 a6573a <=( (not A299)  and  A298 );
 a6574a <=( A203  and  a6573a );
 a6578a <=( (not A302)  and  (not A301) );
 a6579a <=( (not A300)  and  a6578a );
 a6580a <=( a6579a  and  a6574a );
 a6583a <=( A168  and  A169 );
 a6587a <=( (not A201)  and  A166 );
 a6588a <=( (not A167)  and  a6587a );
 a6589a <=( a6588a  and  a6583a );
 a6593a <=( A299  and  (not A298) );
 a6594a <=( A203  and  a6593a );
 a6598a <=( (not A302)  and  (not A301) );
 a6599a <=( (not A300)  and  a6598a );
 a6600a <=( a6599a  and  a6594a );
 a6603a <=( A168  and  A169 );
 a6607a <=( A199  and  A166 );
 a6608a <=( (not A167)  and  a6607a );
 a6609a <=( a6608a  and  a6603a );
 a6613a <=( (not A299)  and  A298 );
 a6614a <=( A200  and  a6613a );
 a6618a <=( (not A302)  and  (not A301) );
 a6619a <=( (not A300)  and  a6618a );
 a6620a <=( a6619a  and  a6614a );
 a6623a <=( A168  and  A169 );
 a6627a <=( A199  and  A166 );
 a6628a <=( (not A167)  and  a6627a );
 a6629a <=( a6628a  and  a6623a );
 a6633a <=( A299  and  (not A298) );
 a6634a <=( A200  and  a6633a );
 a6638a <=( (not A302)  and  (not A301) );
 a6639a <=( (not A300)  and  a6638a );
 a6640a <=( a6639a  and  a6634a );
 a6643a <=( A168  and  A169 );
 a6647a <=( (not A199)  and  A166 );
 a6648a <=( (not A167)  and  a6647a );
 a6649a <=( a6648a  and  a6643a );
 a6653a <=( (not A299)  and  A298 );
 a6654a <=( (not A200)  and  a6653a );
 a6658a <=( (not A302)  and  (not A301) );
 a6659a <=( (not A300)  and  a6658a );
 a6660a <=( a6659a  and  a6654a );
 a6663a <=( A168  and  A169 );
 a6667a <=( (not A199)  and  A166 );
 a6668a <=( (not A167)  and  a6667a );
 a6669a <=( a6668a  and  a6663a );
 a6673a <=( A299  and  (not A298) );
 a6674a <=( (not A200)  and  a6673a );
 a6678a <=( (not A302)  and  (not A301) );
 a6679a <=( (not A300)  and  a6678a );
 a6680a <=( a6679a  and  a6674a );
 a6683a <=( (not A168)  and  A169 );
 a6687a <=( A201  and  A200 );
 a6688a <=( (not A199)  and  a6687a );
 a6689a <=( a6688a  and  a6683a );
 a6693a <=( (not A299)  and  A298 );
 a6694a <=( A202  and  a6693a );
 a6698a <=( (not A302)  and  (not A301) );
 a6699a <=( (not A300)  and  a6698a );
 a6700a <=( a6699a  and  a6694a );
 a6703a <=( (not A168)  and  A169 );
 a6707a <=( A201  and  A200 );
 a6708a <=( (not A199)  and  a6707a );
 a6709a <=( a6708a  and  a6703a );
 a6713a <=( A299  and  (not A298) );
 a6714a <=( A202  and  a6713a );
 a6718a <=( (not A302)  and  (not A301) );
 a6719a <=( (not A300)  and  a6718a );
 a6720a <=( a6719a  and  a6714a );
 a6723a <=( (not A168)  and  A169 );
 a6727a <=( A201  and  A200 );
 a6728a <=( (not A199)  and  a6727a );
 a6729a <=( a6728a  and  a6723a );
 a6733a <=( (not A299)  and  A298 );
 a6734a <=( A203  and  a6733a );
 a6738a <=( (not A302)  and  (not A301) );
 a6739a <=( (not A300)  and  a6738a );
 a6740a <=( a6739a  and  a6734a );
 a6743a <=( (not A168)  and  A169 );
 a6747a <=( A201  and  A200 );
 a6748a <=( (not A199)  and  a6747a );
 a6749a <=( a6748a  and  a6743a );
 a6753a <=( A299  and  (not A298) );
 a6754a <=( A203  and  a6753a );
 a6758a <=( (not A302)  and  (not A301) );
 a6759a <=( (not A300)  and  a6758a );
 a6760a <=( a6759a  and  a6754a );
 a6763a <=( (not A168)  and  A169 );
 a6767a <=( (not A201)  and  A200 );
 a6768a <=( (not A199)  and  a6767a );
 a6769a <=( a6768a  and  a6763a );
 a6773a <=( A298  and  (not A203) );
 a6774a <=( (not A202)  and  a6773a );
 a6778a <=( A301  and  A300 );
 a6779a <=( (not A299)  and  a6778a );
 a6780a <=( a6779a  and  a6774a );
 a6783a <=( (not A168)  and  A169 );
 a6787a <=( (not A201)  and  A200 );
 a6788a <=( (not A199)  and  a6787a );
 a6789a <=( a6788a  and  a6783a );
 a6793a <=( A298  and  (not A203) );
 a6794a <=( (not A202)  and  a6793a );
 a6798a <=( A302  and  A300 );
 a6799a <=( (not A299)  and  a6798a );
 a6800a <=( a6799a  and  a6794a );
 a6803a <=( (not A168)  and  A169 );
 a6807a <=( (not A201)  and  A200 );
 a6808a <=( (not A199)  and  a6807a );
 a6809a <=( a6808a  and  a6803a );
 a6813a <=( (not A298)  and  (not A203) );
 a6814a <=( (not A202)  and  a6813a );
 a6818a <=( A301  and  A300 );
 a6819a <=( A299  and  a6818a );
 a6820a <=( a6819a  and  a6814a );
 a6823a <=( (not A168)  and  A169 );
 a6827a <=( (not A201)  and  A200 );
 a6828a <=( (not A199)  and  a6827a );
 a6829a <=( a6828a  and  a6823a );
 a6833a <=( (not A298)  and  (not A203) );
 a6834a <=( (not A202)  and  a6833a );
 a6838a <=( A302  and  A300 );
 a6839a <=( A299  and  a6838a );
 a6840a <=( a6839a  and  a6834a );
 a6843a <=( (not A168)  and  A169 );
 a6847a <=( A201  and  (not A200) );
 a6848a <=( A199  and  a6847a );
 a6849a <=( a6848a  and  a6843a );
 a6853a <=( (not A299)  and  A298 );
 a6854a <=( A202  and  a6853a );
 a6858a <=( (not A302)  and  (not A301) );
 a6859a <=( (not A300)  and  a6858a );
 a6860a <=( a6859a  and  a6854a );
 a6863a <=( (not A168)  and  A169 );
 a6867a <=( A201  and  (not A200) );
 a6868a <=( A199  and  a6867a );
 a6869a <=( a6868a  and  a6863a );
 a6873a <=( A299  and  (not A298) );
 a6874a <=( A202  and  a6873a );
 a6878a <=( (not A302)  and  (not A301) );
 a6879a <=( (not A300)  and  a6878a );
 a6880a <=( a6879a  and  a6874a );
 a6883a <=( (not A168)  and  A169 );
 a6887a <=( A201  and  (not A200) );
 a6888a <=( A199  and  a6887a );
 a6889a <=( a6888a  and  a6883a );
 a6893a <=( (not A299)  and  A298 );
 a6894a <=( A203  and  a6893a );
 a6898a <=( (not A302)  and  (not A301) );
 a6899a <=( (not A300)  and  a6898a );
 a6900a <=( a6899a  and  a6894a );
 a6903a <=( (not A168)  and  A169 );
 a6907a <=( A201  and  (not A200) );
 a6908a <=( A199  and  a6907a );
 a6909a <=( a6908a  and  a6903a );
 a6913a <=( A299  and  (not A298) );
 a6914a <=( A203  and  a6913a );
 a6918a <=( (not A302)  and  (not A301) );
 a6919a <=( (not A300)  and  a6918a );
 a6920a <=( a6919a  and  a6914a );
 a6923a <=( (not A168)  and  A169 );
 a6927a <=( (not A201)  and  (not A200) );
 a6928a <=( A199  and  a6927a );
 a6929a <=( a6928a  and  a6923a );
 a6933a <=( A298  and  (not A203) );
 a6934a <=( (not A202)  and  a6933a );
 a6938a <=( A301  and  A300 );
 a6939a <=( (not A299)  and  a6938a );
 a6940a <=( a6939a  and  a6934a );
 a6943a <=( (not A168)  and  A169 );
 a6947a <=( (not A201)  and  (not A200) );
 a6948a <=( A199  and  a6947a );
 a6949a <=( a6948a  and  a6943a );
 a6953a <=( A298  and  (not A203) );
 a6954a <=( (not A202)  and  a6953a );
 a6958a <=( A302  and  A300 );
 a6959a <=( (not A299)  and  a6958a );
 a6960a <=( a6959a  and  a6954a );
 a6963a <=( (not A168)  and  A169 );
 a6967a <=( (not A201)  and  (not A200) );
 a6968a <=( A199  and  a6967a );
 a6969a <=( a6968a  and  a6963a );
 a6973a <=( (not A298)  and  (not A203) );
 a6974a <=( (not A202)  and  a6973a );
 a6978a <=( A301  and  A300 );
 a6979a <=( A299  and  a6978a );
 a6980a <=( a6979a  and  a6974a );
 a6983a <=( (not A168)  and  A169 );
 a6987a <=( (not A201)  and  (not A200) );
 a6988a <=( A199  and  a6987a );
 a6989a <=( a6988a  and  a6983a );
 a6993a <=( (not A298)  and  (not A203) );
 a6994a <=( (not A202)  and  a6993a );
 a6998a <=( A302  and  A300 );
 a6999a <=( A299  and  a6998a );
 a7000a <=( a6999a  and  a6994a );
 a7003a <=( (not A169)  and  A170 );
 a7007a <=( A200  and  (not A199) );
 a7008a <=( A168  and  a7007a );
 a7009a <=( a7008a  and  a7003a );
 a7013a <=( A298  and  A202 );
 a7014a <=( A201  and  a7013a );
 a7018a <=( A301  and  A300 );
 a7019a <=( (not A299)  and  a7018a );
 a7020a <=( a7019a  and  a7014a );
 a7023a <=( (not A169)  and  A170 );
 a7027a <=( A200  and  (not A199) );
 a7028a <=( A168  and  a7027a );
 a7029a <=( a7028a  and  a7023a );
 a7033a <=( A298  and  A202 );
 a7034a <=( A201  and  a7033a );
 a7038a <=( A302  and  A300 );
 a7039a <=( (not A299)  and  a7038a );
 a7040a <=( a7039a  and  a7034a );
 a7043a <=( (not A169)  and  A170 );
 a7047a <=( A200  and  (not A199) );
 a7048a <=( A168  and  a7047a );
 a7049a <=( a7048a  and  a7043a );
 a7053a <=( (not A298)  and  A202 );
 a7054a <=( A201  and  a7053a );
 a7058a <=( A301  and  A300 );
 a7059a <=( A299  and  a7058a );
 a7060a <=( a7059a  and  a7054a );
 a7063a <=( (not A169)  and  A170 );
 a7067a <=( A200  and  (not A199) );
 a7068a <=( A168  and  a7067a );
 a7069a <=( a7068a  and  a7063a );
 a7073a <=( (not A298)  and  A202 );
 a7074a <=( A201  and  a7073a );
 a7078a <=( A302  and  A300 );
 a7079a <=( A299  and  a7078a );
 a7080a <=( a7079a  and  a7074a );
 a7083a <=( (not A169)  and  A170 );
 a7087a <=( A200  and  (not A199) );
 a7088a <=( A168  and  a7087a );
 a7089a <=( a7088a  and  a7083a );
 a7093a <=( A298  and  A203 );
 a7094a <=( A201  and  a7093a );
 a7098a <=( A301  and  A300 );
 a7099a <=( (not A299)  and  a7098a );
 a7100a <=( a7099a  and  a7094a );
 a7103a <=( (not A169)  and  A170 );
 a7107a <=( A200  and  (not A199) );
 a7108a <=( A168  and  a7107a );
 a7109a <=( a7108a  and  a7103a );
 a7113a <=( A298  and  A203 );
 a7114a <=( A201  and  a7113a );
 a7118a <=( A302  and  A300 );
 a7119a <=( (not A299)  and  a7118a );
 a7120a <=( a7119a  and  a7114a );
 a7123a <=( (not A169)  and  A170 );
 a7127a <=( A200  and  (not A199) );
 a7128a <=( A168  and  a7127a );
 a7129a <=( a7128a  and  a7123a );
 a7133a <=( (not A298)  and  A203 );
 a7134a <=( A201  and  a7133a );
 a7138a <=( A301  and  A300 );
 a7139a <=( A299  and  a7138a );
 a7140a <=( a7139a  and  a7134a );
 a7143a <=( (not A169)  and  A170 );
 a7147a <=( A200  and  (not A199) );
 a7148a <=( A168  and  a7147a );
 a7149a <=( a7148a  and  a7143a );
 a7153a <=( (not A298)  and  A203 );
 a7154a <=( A201  and  a7153a );
 a7158a <=( A302  and  A300 );
 a7159a <=( A299  and  a7158a );
 a7160a <=( a7159a  and  a7154a );
 a7163a <=( (not A169)  and  A170 );
 a7167a <=( (not A200)  and  A199 );
 a7168a <=( A168  and  a7167a );
 a7169a <=( a7168a  and  a7163a );
 a7173a <=( A298  and  A202 );
 a7174a <=( A201  and  a7173a );
 a7178a <=( A301  and  A300 );
 a7179a <=( (not A299)  and  a7178a );
 a7180a <=( a7179a  and  a7174a );
 a7183a <=( (not A169)  and  A170 );
 a7187a <=( (not A200)  and  A199 );
 a7188a <=( A168  and  a7187a );
 a7189a <=( a7188a  and  a7183a );
 a7193a <=( A298  and  A202 );
 a7194a <=( A201  and  a7193a );
 a7198a <=( A302  and  A300 );
 a7199a <=( (not A299)  and  a7198a );
 a7200a <=( a7199a  and  a7194a );
 a7203a <=( (not A169)  and  A170 );
 a7207a <=( (not A200)  and  A199 );
 a7208a <=( A168  and  a7207a );
 a7209a <=( a7208a  and  a7203a );
 a7213a <=( (not A298)  and  A202 );
 a7214a <=( A201  and  a7213a );
 a7218a <=( A301  and  A300 );
 a7219a <=( A299  and  a7218a );
 a7220a <=( a7219a  and  a7214a );
 a7223a <=( (not A169)  and  A170 );
 a7227a <=( (not A200)  and  A199 );
 a7228a <=( A168  and  a7227a );
 a7229a <=( a7228a  and  a7223a );
 a7233a <=( (not A298)  and  A202 );
 a7234a <=( A201  and  a7233a );
 a7238a <=( A302  and  A300 );
 a7239a <=( A299  and  a7238a );
 a7240a <=( a7239a  and  a7234a );
 a7243a <=( (not A169)  and  A170 );
 a7247a <=( (not A200)  and  A199 );
 a7248a <=( A168  and  a7247a );
 a7249a <=( a7248a  and  a7243a );
 a7253a <=( A298  and  A203 );
 a7254a <=( A201  and  a7253a );
 a7258a <=( A301  and  A300 );
 a7259a <=( (not A299)  and  a7258a );
 a7260a <=( a7259a  and  a7254a );
 a7263a <=( (not A169)  and  A170 );
 a7267a <=( (not A200)  and  A199 );
 a7268a <=( A168  and  a7267a );
 a7269a <=( a7268a  and  a7263a );
 a7273a <=( A298  and  A203 );
 a7274a <=( A201  and  a7273a );
 a7278a <=( A302  and  A300 );
 a7279a <=( (not A299)  and  a7278a );
 a7280a <=( a7279a  and  a7274a );
 a7283a <=( (not A169)  and  A170 );
 a7287a <=( (not A200)  and  A199 );
 a7288a <=( A168  and  a7287a );
 a7289a <=( a7288a  and  a7283a );
 a7293a <=( (not A298)  and  A203 );
 a7294a <=( A201  and  a7293a );
 a7298a <=( A301  and  A300 );
 a7299a <=( A299  and  a7298a );
 a7300a <=( a7299a  and  a7294a );
 a7303a <=( (not A169)  and  A170 );
 a7307a <=( (not A200)  and  A199 );
 a7308a <=( A168  and  a7307a );
 a7309a <=( a7308a  and  a7303a );
 a7313a <=( (not A298)  and  A203 );
 a7314a <=( A201  and  a7313a );
 a7318a <=( A302  and  A300 );
 a7319a <=( A299  and  a7318a );
 a7320a <=( a7319a  and  a7314a );
 a7323a <=( (not A169)  and  A170 );
 a7327a <=( (not A166)  and  A167 );
 a7328a <=( (not A168)  and  a7327a );
 a7329a <=( a7328a  and  a7323a );
 a7333a <=( A298  and  A202 );
 a7334a <=( (not A201)  and  a7333a );
 a7338a <=( A301  and  A300 );
 a7339a <=( (not A299)  and  a7338a );
 a7340a <=( a7339a  and  a7334a );
 a7343a <=( (not A169)  and  A170 );
 a7347a <=( (not A166)  and  A167 );
 a7348a <=( (not A168)  and  a7347a );
 a7349a <=( a7348a  and  a7343a );
 a7353a <=( A298  and  A202 );
 a7354a <=( (not A201)  and  a7353a );
 a7358a <=( A302  and  A300 );
 a7359a <=( (not A299)  and  a7358a );
 a7360a <=( a7359a  and  a7354a );
 a7363a <=( (not A169)  and  A170 );
 a7367a <=( (not A166)  and  A167 );
 a7368a <=( (not A168)  and  a7367a );
 a7369a <=( a7368a  and  a7363a );
 a7373a <=( (not A298)  and  A202 );
 a7374a <=( (not A201)  and  a7373a );
 a7378a <=( A301  and  A300 );
 a7379a <=( A299  and  a7378a );
 a7380a <=( a7379a  and  a7374a );
 a7383a <=( (not A169)  and  A170 );
 a7387a <=( (not A166)  and  A167 );
 a7388a <=( (not A168)  and  a7387a );
 a7389a <=( a7388a  and  a7383a );
 a7393a <=( (not A298)  and  A202 );
 a7394a <=( (not A201)  and  a7393a );
 a7398a <=( A302  and  A300 );
 a7399a <=( A299  and  a7398a );
 a7400a <=( a7399a  and  a7394a );
 a7403a <=( (not A169)  and  A170 );
 a7407a <=( (not A166)  and  A167 );
 a7408a <=( (not A168)  and  a7407a );
 a7409a <=( a7408a  and  a7403a );
 a7413a <=( A298  and  A203 );
 a7414a <=( (not A201)  and  a7413a );
 a7418a <=( A301  and  A300 );
 a7419a <=( (not A299)  and  a7418a );
 a7420a <=( a7419a  and  a7414a );
 a7423a <=( (not A169)  and  A170 );
 a7427a <=( (not A166)  and  A167 );
 a7428a <=( (not A168)  and  a7427a );
 a7429a <=( a7428a  and  a7423a );
 a7433a <=( A298  and  A203 );
 a7434a <=( (not A201)  and  a7433a );
 a7438a <=( A302  and  A300 );
 a7439a <=( (not A299)  and  a7438a );
 a7440a <=( a7439a  and  a7434a );
 a7443a <=( (not A169)  and  A170 );
 a7447a <=( (not A166)  and  A167 );
 a7448a <=( (not A168)  and  a7447a );
 a7449a <=( a7448a  and  a7443a );
 a7453a <=( (not A298)  and  A203 );
 a7454a <=( (not A201)  and  a7453a );
 a7458a <=( A301  and  A300 );
 a7459a <=( A299  and  a7458a );
 a7460a <=( a7459a  and  a7454a );
 a7463a <=( (not A169)  and  A170 );
 a7467a <=( (not A166)  and  A167 );
 a7468a <=( (not A168)  and  a7467a );
 a7469a <=( a7468a  and  a7463a );
 a7473a <=( (not A298)  and  A203 );
 a7474a <=( (not A201)  and  a7473a );
 a7478a <=( A302  and  A300 );
 a7479a <=( A299  and  a7478a );
 a7480a <=( a7479a  and  a7474a );
 a7483a <=( (not A169)  and  A170 );
 a7487a <=( (not A166)  and  A167 );
 a7488a <=( (not A168)  and  a7487a );
 a7489a <=( a7488a  and  a7483a );
 a7493a <=( A298  and  A200 );
 a7494a <=( A199  and  a7493a );
 a7498a <=( A301  and  A300 );
 a7499a <=( (not A299)  and  a7498a );
 a7500a <=( a7499a  and  a7494a );
 a7503a <=( (not A169)  and  A170 );
 a7507a <=( (not A166)  and  A167 );
 a7508a <=( (not A168)  and  a7507a );
 a7509a <=( a7508a  and  a7503a );
 a7513a <=( A298  and  A200 );
 a7514a <=( A199  and  a7513a );
 a7518a <=( A302  and  A300 );
 a7519a <=( (not A299)  and  a7518a );
 a7520a <=( a7519a  and  a7514a );
 a7523a <=( (not A169)  and  A170 );
 a7527a <=( (not A166)  and  A167 );
 a7528a <=( (not A168)  and  a7527a );
 a7529a <=( a7528a  and  a7523a );
 a7533a <=( (not A298)  and  A200 );
 a7534a <=( A199  and  a7533a );
 a7538a <=( A301  and  A300 );
 a7539a <=( A299  and  a7538a );
 a7540a <=( a7539a  and  a7534a );
 a7543a <=( (not A169)  and  A170 );
 a7547a <=( (not A166)  and  A167 );
 a7548a <=( (not A168)  and  a7547a );
 a7549a <=( a7548a  and  a7543a );
 a7553a <=( (not A298)  and  A200 );
 a7554a <=( A199  and  a7553a );
 a7558a <=( A302  and  A300 );
 a7559a <=( A299  and  a7558a );
 a7560a <=( a7559a  and  a7554a );
 a7563a <=( (not A169)  and  A170 );
 a7567a <=( (not A166)  and  A167 );
 a7568a <=( (not A168)  and  a7567a );
 a7569a <=( a7568a  and  a7563a );
 a7573a <=( A298  and  (not A200) );
 a7574a <=( (not A199)  and  a7573a );
 a7578a <=( A301  and  A300 );
 a7579a <=( (not A299)  and  a7578a );
 a7580a <=( a7579a  and  a7574a );
 a7583a <=( (not A169)  and  A170 );
 a7587a <=( (not A166)  and  A167 );
 a7588a <=( (not A168)  and  a7587a );
 a7589a <=( a7588a  and  a7583a );
 a7593a <=( A298  and  (not A200) );
 a7594a <=( (not A199)  and  a7593a );
 a7598a <=( A302  and  A300 );
 a7599a <=( (not A299)  and  a7598a );
 a7600a <=( a7599a  and  a7594a );
 a7603a <=( (not A169)  and  A170 );
 a7607a <=( (not A166)  and  A167 );
 a7608a <=( (not A168)  and  a7607a );
 a7609a <=( a7608a  and  a7603a );
 a7613a <=( (not A298)  and  (not A200) );
 a7614a <=( (not A199)  and  a7613a );
 a7618a <=( A301  and  A300 );
 a7619a <=( A299  and  a7618a );
 a7620a <=( a7619a  and  a7614a );
 a7623a <=( (not A169)  and  A170 );
 a7627a <=( (not A166)  and  A167 );
 a7628a <=( (not A168)  and  a7627a );
 a7629a <=( a7628a  and  a7623a );
 a7633a <=( (not A298)  and  (not A200) );
 a7634a <=( (not A199)  and  a7633a );
 a7638a <=( A302  and  A300 );
 a7639a <=( A299  and  a7638a );
 a7640a <=( a7639a  and  a7634a );
 a7643a <=( (not A169)  and  A170 );
 a7647a <=( A166  and  (not A167) );
 a7648a <=( (not A168)  and  a7647a );
 a7649a <=( a7648a  and  a7643a );
 a7653a <=( A298  and  A202 );
 a7654a <=( (not A201)  and  a7653a );
 a7658a <=( A301  and  A300 );
 a7659a <=( (not A299)  and  a7658a );
 a7660a <=( a7659a  and  a7654a );
 a7663a <=( (not A169)  and  A170 );
 a7667a <=( A166  and  (not A167) );
 a7668a <=( (not A168)  and  a7667a );
 a7669a <=( a7668a  and  a7663a );
 a7673a <=( A298  and  A202 );
 a7674a <=( (not A201)  and  a7673a );
 a7678a <=( A302  and  A300 );
 a7679a <=( (not A299)  and  a7678a );
 a7680a <=( a7679a  and  a7674a );
 a7683a <=( (not A169)  and  A170 );
 a7687a <=( A166  and  (not A167) );
 a7688a <=( (not A168)  and  a7687a );
 a7689a <=( a7688a  and  a7683a );
 a7693a <=( (not A298)  and  A202 );
 a7694a <=( (not A201)  and  a7693a );
 a7698a <=( A301  and  A300 );
 a7699a <=( A299  and  a7698a );
 a7700a <=( a7699a  and  a7694a );
 a7703a <=( (not A169)  and  A170 );
 a7707a <=( A166  and  (not A167) );
 a7708a <=( (not A168)  and  a7707a );
 a7709a <=( a7708a  and  a7703a );
 a7713a <=( (not A298)  and  A202 );
 a7714a <=( (not A201)  and  a7713a );
 a7718a <=( A302  and  A300 );
 a7719a <=( A299  and  a7718a );
 a7720a <=( a7719a  and  a7714a );
 a7723a <=( (not A169)  and  A170 );
 a7727a <=( A166  and  (not A167) );
 a7728a <=( (not A168)  and  a7727a );
 a7729a <=( a7728a  and  a7723a );
 a7733a <=( A298  and  A203 );
 a7734a <=( (not A201)  and  a7733a );
 a7738a <=( A301  and  A300 );
 a7739a <=( (not A299)  and  a7738a );
 a7740a <=( a7739a  and  a7734a );
 a7743a <=( (not A169)  and  A170 );
 a7747a <=( A166  and  (not A167) );
 a7748a <=( (not A168)  and  a7747a );
 a7749a <=( a7748a  and  a7743a );
 a7753a <=( A298  and  A203 );
 a7754a <=( (not A201)  and  a7753a );
 a7758a <=( A302  and  A300 );
 a7759a <=( (not A299)  and  a7758a );
 a7760a <=( a7759a  and  a7754a );
 a7763a <=( (not A169)  and  A170 );
 a7767a <=( A166  and  (not A167) );
 a7768a <=( (not A168)  and  a7767a );
 a7769a <=( a7768a  and  a7763a );
 a7773a <=( (not A298)  and  A203 );
 a7774a <=( (not A201)  and  a7773a );
 a7778a <=( A301  and  A300 );
 a7779a <=( A299  and  a7778a );
 a7780a <=( a7779a  and  a7774a );
 a7783a <=( (not A169)  and  A170 );
 a7787a <=( A166  and  (not A167) );
 a7788a <=( (not A168)  and  a7787a );
 a7789a <=( a7788a  and  a7783a );
 a7793a <=( (not A298)  and  A203 );
 a7794a <=( (not A201)  and  a7793a );
 a7798a <=( A302  and  A300 );
 a7799a <=( A299  and  a7798a );
 a7800a <=( a7799a  and  a7794a );
 a7803a <=( (not A169)  and  A170 );
 a7807a <=( A166  and  (not A167) );
 a7808a <=( (not A168)  and  a7807a );
 a7809a <=( a7808a  and  a7803a );
 a7813a <=( A298  and  A200 );
 a7814a <=( A199  and  a7813a );
 a7818a <=( A301  and  A300 );
 a7819a <=( (not A299)  and  a7818a );
 a7820a <=( a7819a  and  a7814a );
 a7823a <=( (not A169)  and  A170 );
 a7827a <=( A166  and  (not A167) );
 a7828a <=( (not A168)  and  a7827a );
 a7829a <=( a7828a  and  a7823a );
 a7833a <=( A298  and  A200 );
 a7834a <=( A199  and  a7833a );
 a7838a <=( A302  and  A300 );
 a7839a <=( (not A299)  and  a7838a );
 a7840a <=( a7839a  and  a7834a );
 a7843a <=( (not A169)  and  A170 );
 a7847a <=( A166  and  (not A167) );
 a7848a <=( (not A168)  and  a7847a );
 a7849a <=( a7848a  and  a7843a );
 a7853a <=( (not A298)  and  A200 );
 a7854a <=( A199  and  a7853a );
 a7858a <=( A301  and  A300 );
 a7859a <=( A299  and  a7858a );
 a7860a <=( a7859a  and  a7854a );
 a7863a <=( (not A169)  and  A170 );
 a7867a <=( A166  and  (not A167) );
 a7868a <=( (not A168)  and  a7867a );
 a7869a <=( a7868a  and  a7863a );
 a7873a <=( (not A298)  and  A200 );
 a7874a <=( A199  and  a7873a );
 a7878a <=( A302  and  A300 );
 a7879a <=( A299  and  a7878a );
 a7880a <=( a7879a  and  a7874a );
 a7883a <=( (not A169)  and  A170 );
 a7887a <=( A166  and  (not A167) );
 a7888a <=( (not A168)  and  a7887a );
 a7889a <=( a7888a  and  a7883a );
 a7893a <=( A298  and  (not A200) );
 a7894a <=( (not A199)  and  a7893a );
 a7898a <=( A301  and  A300 );
 a7899a <=( (not A299)  and  a7898a );
 a7900a <=( a7899a  and  a7894a );
 a7903a <=( (not A169)  and  A170 );
 a7907a <=( A166  and  (not A167) );
 a7908a <=( (not A168)  and  a7907a );
 a7909a <=( a7908a  and  a7903a );
 a7913a <=( A298  and  (not A200) );
 a7914a <=( (not A199)  and  a7913a );
 a7918a <=( A302  and  A300 );
 a7919a <=( (not A299)  and  a7918a );
 a7920a <=( a7919a  and  a7914a );
 a7923a <=( (not A169)  and  A170 );
 a7927a <=( A166  and  (not A167) );
 a7928a <=( (not A168)  and  a7927a );
 a7929a <=( a7928a  and  a7923a );
 a7933a <=( (not A298)  and  (not A200) );
 a7934a <=( (not A199)  and  a7933a );
 a7938a <=( A301  and  A300 );
 a7939a <=( A299  and  a7938a );
 a7940a <=( a7939a  and  a7934a );
 a7943a <=( (not A169)  and  A170 );
 a7947a <=( A166  and  (not A167) );
 a7948a <=( (not A168)  and  a7947a );
 a7949a <=( a7948a  and  a7943a );
 a7953a <=( (not A298)  and  (not A200) );
 a7954a <=( (not A199)  and  a7953a );
 a7958a <=( A302  and  A300 );
 a7959a <=( A299  and  a7958a );
 a7960a <=( a7959a  and  a7954a );
 a7964a <=( (not A199)  and  A166 );
 a7965a <=( A167  and  a7964a );
 a7969a <=( (not A202)  and  (not A201) );
 a7970a <=( A200  and  a7969a );
 a7971a <=( a7970a  and  a7965a );
 a7975a <=( (not A299)  and  A298 );
 a7976a <=( (not A203)  and  a7975a );
 a7980a <=( (not A302)  and  (not A301) );
 a7981a <=( (not A300)  and  a7980a );
 a7982a <=( a7981a  and  a7976a );
 a7986a <=( (not A199)  and  A166 );
 a7987a <=( A167  and  a7986a );
 a7991a <=( (not A202)  and  (not A201) );
 a7992a <=( A200  and  a7991a );
 a7993a <=( a7992a  and  a7987a );
 a7997a <=( A299  and  (not A298) );
 a7998a <=( (not A203)  and  a7997a );
 a8002a <=( (not A302)  and  (not A301) );
 a8003a <=( (not A300)  and  a8002a );
 a8004a <=( a8003a  and  a7998a );
 a8008a <=( A199  and  A166 );
 a8009a <=( A167  and  a8008a );
 a8013a <=( (not A202)  and  (not A201) );
 a8014a <=( (not A200)  and  a8013a );
 a8015a <=( a8014a  and  a8009a );
 a8019a <=( (not A299)  and  A298 );
 a8020a <=( (not A203)  and  a8019a );
 a8024a <=( (not A302)  and  (not A301) );
 a8025a <=( (not A300)  and  a8024a );
 a8026a <=( a8025a  and  a8020a );
 a8030a <=( A199  and  A166 );
 a8031a <=( A167  and  a8030a );
 a8035a <=( (not A202)  and  (not A201) );
 a8036a <=( (not A200)  and  a8035a );
 a8037a <=( a8036a  and  a8031a );
 a8041a <=( A299  and  (not A298) );
 a8042a <=( (not A203)  and  a8041a );
 a8046a <=( (not A302)  and  (not A301) );
 a8047a <=( (not A300)  and  a8046a );
 a8048a <=( a8047a  and  a8042a );
 a8052a <=( (not A199)  and  (not A166) );
 a8053a <=( (not A167)  and  a8052a );
 a8057a <=( (not A202)  and  (not A201) );
 a8058a <=( A200  and  a8057a );
 a8059a <=( a8058a  and  a8053a );
 a8063a <=( (not A299)  and  A298 );
 a8064a <=( (not A203)  and  a8063a );
 a8068a <=( (not A302)  and  (not A301) );
 a8069a <=( (not A300)  and  a8068a );
 a8070a <=( a8069a  and  a8064a );
 a8074a <=( (not A199)  and  (not A166) );
 a8075a <=( (not A167)  and  a8074a );
 a8079a <=( (not A202)  and  (not A201) );
 a8080a <=( A200  and  a8079a );
 a8081a <=( a8080a  and  a8075a );
 a8085a <=( A299  and  (not A298) );
 a8086a <=( (not A203)  and  a8085a );
 a8090a <=( (not A302)  and  (not A301) );
 a8091a <=( (not A300)  and  a8090a );
 a8092a <=( a8091a  and  a8086a );
 a8096a <=( A199  and  (not A166) );
 a8097a <=( (not A167)  and  a8096a );
 a8101a <=( (not A202)  and  (not A201) );
 a8102a <=( (not A200)  and  a8101a );
 a8103a <=( a8102a  and  a8097a );
 a8107a <=( (not A299)  and  A298 );
 a8108a <=( (not A203)  and  a8107a );
 a8112a <=( (not A302)  and  (not A301) );
 a8113a <=( (not A300)  and  a8112a );
 a8114a <=( a8113a  and  a8108a );
 a8118a <=( A199  and  (not A166) );
 a8119a <=( (not A167)  and  a8118a );
 a8123a <=( (not A202)  and  (not A201) );
 a8124a <=( (not A200)  and  a8123a );
 a8125a <=( a8124a  and  a8119a );
 a8129a <=( A299  and  (not A298) );
 a8130a <=( (not A203)  and  a8129a );
 a8134a <=( (not A302)  and  (not A301) );
 a8135a <=( (not A300)  and  a8134a );
 a8136a <=( a8135a  and  a8130a );
 a8140a <=( A167  and  A168 );
 a8141a <=( (not A170)  and  a8140a );
 a8145a <=( (not A202)  and  A201 );
 a8146a <=( (not A166)  and  a8145a );
 a8147a <=( a8146a  and  a8141a );
 a8151a <=( (not A299)  and  A298 );
 a8152a <=( (not A203)  and  a8151a );
 a8156a <=( (not A302)  and  (not A301) );
 a8157a <=( (not A300)  and  a8156a );
 a8158a <=( a8157a  and  a8152a );
 a8162a <=( A167  and  A168 );
 a8163a <=( (not A170)  and  a8162a );
 a8167a <=( (not A202)  and  A201 );
 a8168a <=( (not A166)  and  a8167a );
 a8169a <=( a8168a  and  a8163a );
 a8173a <=( A299  and  (not A298) );
 a8174a <=( (not A203)  and  a8173a );
 a8178a <=( (not A302)  and  (not A301) );
 a8179a <=( (not A300)  and  a8178a );
 a8180a <=( a8179a  and  a8174a );
 a8184a <=( (not A167)  and  A168 );
 a8185a <=( (not A170)  and  a8184a );
 a8189a <=( (not A202)  and  A201 );
 a8190a <=( A166  and  a8189a );
 a8191a <=( a8190a  and  a8185a );
 a8195a <=( (not A299)  and  A298 );
 a8196a <=( (not A203)  and  a8195a );
 a8200a <=( (not A302)  and  (not A301) );
 a8201a <=( (not A300)  and  a8200a );
 a8202a <=( a8201a  and  a8196a );
 a8206a <=( (not A167)  and  A168 );
 a8207a <=( (not A170)  and  a8206a );
 a8211a <=( (not A202)  and  A201 );
 a8212a <=( A166  and  a8211a );
 a8213a <=( a8212a  and  a8207a );
 a8217a <=( A299  and  (not A298) );
 a8218a <=( (not A203)  and  a8217a );
 a8222a <=( (not A302)  and  (not A301) );
 a8223a <=( (not A300)  and  a8222a );
 a8224a <=( a8223a  and  a8218a );
 a8228a <=( (not A199)  and  (not A168) );
 a8229a <=( (not A170)  and  a8228a );
 a8233a <=( (not A202)  and  (not A201) );
 a8234a <=( A200  and  a8233a );
 a8235a <=( a8234a  and  a8229a );
 a8239a <=( (not A299)  and  A298 );
 a8240a <=( (not A203)  and  a8239a );
 a8244a <=( (not A302)  and  (not A301) );
 a8245a <=( (not A300)  and  a8244a );
 a8246a <=( a8245a  and  a8240a );
 a8250a <=( (not A199)  and  (not A168) );
 a8251a <=( (not A170)  and  a8250a );
 a8255a <=( (not A202)  and  (not A201) );
 a8256a <=( A200  and  a8255a );
 a8257a <=( a8256a  and  a8251a );
 a8261a <=( A299  and  (not A298) );
 a8262a <=( (not A203)  and  a8261a );
 a8266a <=( (not A302)  and  (not A301) );
 a8267a <=( (not A300)  and  a8266a );
 a8268a <=( a8267a  and  a8262a );
 a8272a <=( A199  and  (not A168) );
 a8273a <=( (not A170)  and  a8272a );
 a8277a <=( (not A202)  and  (not A201) );
 a8278a <=( (not A200)  and  a8277a );
 a8279a <=( a8278a  and  a8273a );
 a8283a <=( (not A299)  and  A298 );
 a8284a <=( (not A203)  and  a8283a );
 a8288a <=( (not A302)  and  (not A301) );
 a8289a <=( (not A300)  and  a8288a );
 a8290a <=( a8289a  and  a8284a );
 a8294a <=( A199  and  (not A168) );
 a8295a <=( (not A170)  and  a8294a );
 a8299a <=( (not A202)  and  (not A201) );
 a8300a <=( (not A200)  and  a8299a );
 a8301a <=( a8300a  and  a8295a );
 a8305a <=( A299  and  (not A298) );
 a8306a <=( (not A203)  and  a8305a );
 a8310a <=( (not A302)  and  (not A301) );
 a8311a <=( (not A300)  and  a8310a );
 a8312a <=( a8311a  and  a8306a );
 a8316a <=( A167  and  A168 );
 a8317a <=( A169  and  a8316a );
 a8321a <=( (not A202)  and  A201 );
 a8322a <=( (not A166)  and  a8321a );
 a8323a <=( a8322a  and  a8317a );
 a8327a <=( (not A299)  and  A298 );
 a8328a <=( (not A203)  and  a8327a );
 a8332a <=( (not A302)  and  (not A301) );
 a8333a <=( (not A300)  and  a8332a );
 a8334a <=( a8333a  and  a8328a );
 a8338a <=( A167  and  A168 );
 a8339a <=( A169  and  a8338a );
 a8343a <=( (not A202)  and  A201 );
 a8344a <=( (not A166)  and  a8343a );
 a8345a <=( a8344a  and  a8339a );
 a8349a <=( A299  and  (not A298) );
 a8350a <=( (not A203)  and  a8349a );
 a8354a <=( (not A302)  and  (not A301) );
 a8355a <=( (not A300)  and  a8354a );
 a8356a <=( a8355a  and  a8350a );
 a8360a <=( (not A167)  and  A168 );
 a8361a <=( A169  and  a8360a );
 a8365a <=( (not A202)  and  A201 );
 a8366a <=( A166  and  a8365a );
 a8367a <=( a8366a  and  a8361a );
 a8371a <=( (not A299)  and  A298 );
 a8372a <=( (not A203)  and  a8371a );
 a8376a <=( (not A302)  and  (not A301) );
 a8377a <=( (not A300)  and  a8376a );
 a8378a <=( a8377a  and  a8372a );
 a8382a <=( (not A167)  and  A168 );
 a8383a <=( A169  and  a8382a );
 a8387a <=( (not A202)  and  A201 );
 a8388a <=( A166  and  a8387a );
 a8389a <=( a8388a  and  a8383a );
 a8393a <=( A299  and  (not A298) );
 a8394a <=( (not A203)  and  a8393a );
 a8398a <=( (not A302)  and  (not A301) );
 a8399a <=( (not A300)  and  a8398a );
 a8400a <=( a8399a  and  a8394a );
 a8404a <=( (not A199)  and  (not A168) );
 a8405a <=( A169  and  a8404a );
 a8409a <=( (not A202)  and  (not A201) );
 a8410a <=( A200  and  a8409a );
 a8411a <=( a8410a  and  a8405a );
 a8415a <=( (not A299)  and  A298 );
 a8416a <=( (not A203)  and  a8415a );
 a8420a <=( (not A302)  and  (not A301) );
 a8421a <=( (not A300)  and  a8420a );
 a8422a <=( a8421a  and  a8416a );
 a8426a <=( (not A199)  and  (not A168) );
 a8427a <=( A169  and  a8426a );
 a8431a <=( (not A202)  and  (not A201) );
 a8432a <=( A200  and  a8431a );
 a8433a <=( a8432a  and  a8427a );
 a8437a <=( A299  and  (not A298) );
 a8438a <=( (not A203)  and  a8437a );
 a8442a <=( (not A302)  and  (not A301) );
 a8443a <=( (not A300)  and  a8442a );
 a8444a <=( a8443a  and  a8438a );
 a8448a <=( A199  and  (not A168) );
 a8449a <=( A169  and  a8448a );
 a8453a <=( (not A202)  and  (not A201) );
 a8454a <=( (not A200)  and  a8453a );
 a8455a <=( a8454a  and  a8449a );
 a8459a <=( (not A299)  and  A298 );
 a8460a <=( (not A203)  and  a8459a );
 a8464a <=( (not A302)  and  (not A301) );
 a8465a <=( (not A300)  and  a8464a );
 a8466a <=( a8465a  and  a8460a );
 a8470a <=( A199  and  (not A168) );
 a8471a <=( A169  and  a8470a );
 a8475a <=( (not A202)  and  (not A201) );
 a8476a <=( (not A200)  and  a8475a );
 a8477a <=( a8476a  and  a8471a );
 a8481a <=( A299  and  (not A298) );
 a8482a <=( (not A203)  and  a8481a );
 a8486a <=( (not A302)  and  (not A301) );
 a8487a <=( (not A300)  and  a8486a );
 a8488a <=( a8487a  and  a8482a );
 a8492a <=( A168  and  (not A169) );
 a8493a <=( A170  and  a8492a );
 a8497a <=( A201  and  A200 );
 a8498a <=( (not A199)  and  a8497a );
 a8499a <=( a8498a  and  a8493a );
 a8503a <=( (not A299)  and  A298 );
 a8504a <=( A202  and  a8503a );
 a8508a <=( (not A302)  and  (not A301) );
 a8509a <=( (not A300)  and  a8508a );
 a8510a <=( a8509a  and  a8504a );
 a8514a <=( A168  and  (not A169) );
 a8515a <=( A170  and  a8514a );
 a8519a <=( A201  and  A200 );
 a8520a <=( (not A199)  and  a8519a );
 a8521a <=( a8520a  and  a8515a );
 a8525a <=( A299  and  (not A298) );
 a8526a <=( A202  and  a8525a );
 a8530a <=( (not A302)  and  (not A301) );
 a8531a <=( (not A300)  and  a8530a );
 a8532a <=( a8531a  and  a8526a );
 a8536a <=( A168  and  (not A169) );
 a8537a <=( A170  and  a8536a );
 a8541a <=( A201  and  A200 );
 a8542a <=( (not A199)  and  a8541a );
 a8543a <=( a8542a  and  a8537a );
 a8547a <=( (not A299)  and  A298 );
 a8548a <=( A203  and  a8547a );
 a8552a <=( (not A302)  and  (not A301) );
 a8553a <=( (not A300)  and  a8552a );
 a8554a <=( a8553a  and  a8548a );
 a8558a <=( A168  and  (not A169) );
 a8559a <=( A170  and  a8558a );
 a8563a <=( A201  and  A200 );
 a8564a <=( (not A199)  and  a8563a );
 a8565a <=( a8564a  and  a8559a );
 a8569a <=( A299  and  (not A298) );
 a8570a <=( A203  and  a8569a );
 a8574a <=( (not A302)  and  (not A301) );
 a8575a <=( (not A300)  and  a8574a );
 a8576a <=( a8575a  and  a8570a );
 a8580a <=( A168  and  (not A169) );
 a8581a <=( A170  and  a8580a );
 a8585a <=( (not A201)  and  A200 );
 a8586a <=( (not A199)  and  a8585a );
 a8587a <=( a8586a  and  a8581a );
 a8591a <=( A298  and  (not A203) );
 a8592a <=( (not A202)  and  a8591a );
 a8596a <=( A301  and  A300 );
 a8597a <=( (not A299)  and  a8596a );
 a8598a <=( a8597a  and  a8592a );
 a8602a <=( A168  and  (not A169) );
 a8603a <=( A170  and  a8602a );
 a8607a <=( (not A201)  and  A200 );
 a8608a <=( (not A199)  and  a8607a );
 a8609a <=( a8608a  and  a8603a );
 a8613a <=( A298  and  (not A203) );
 a8614a <=( (not A202)  and  a8613a );
 a8618a <=( A302  and  A300 );
 a8619a <=( (not A299)  and  a8618a );
 a8620a <=( a8619a  and  a8614a );
 a8624a <=( A168  and  (not A169) );
 a8625a <=( A170  and  a8624a );
 a8629a <=( (not A201)  and  A200 );
 a8630a <=( (not A199)  and  a8629a );
 a8631a <=( a8630a  and  a8625a );
 a8635a <=( (not A298)  and  (not A203) );
 a8636a <=( (not A202)  and  a8635a );
 a8640a <=( A301  and  A300 );
 a8641a <=( A299  and  a8640a );
 a8642a <=( a8641a  and  a8636a );
 a8646a <=( A168  and  (not A169) );
 a8647a <=( A170  and  a8646a );
 a8651a <=( (not A201)  and  A200 );
 a8652a <=( (not A199)  and  a8651a );
 a8653a <=( a8652a  and  a8647a );
 a8657a <=( (not A298)  and  (not A203) );
 a8658a <=( (not A202)  and  a8657a );
 a8662a <=( A302  and  A300 );
 a8663a <=( A299  and  a8662a );
 a8664a <=( a8663a  and  a8658a );
 a8668a <=( A168  and  (not A169) );
 a8669a <=( A170  and  a8668a );
 a8673a <=( A201  and  (not A200) );
 a8674a <=( A199  and  a8673a );
 a8675a <=( a8674a  and  a8669a );
 a8679a <=( (not A299)  and  A298 );
 a8680a <=( A202  and  a8679a );
 a8684a <=( (not A302)  and  (not A301) );
 a8685a <=( (not A300)  and  a8684a );
 a8686a <=( a8685a  and  a8680a );
 a8690a <=( A168  and  (not A169) );
 a8691a <=( A170  and  a8690a );
 a8695a <=( A201  and  (not A200) );
 a8696a <=( A199  and  a8695a );
 a8697a <=( a8696a  and  a8691a );
 a8701a <=( A299  and  (not A298) );
 a8702a <=( A202  and  a8701a );
 a8706a <=( (not A302)  and  (not A301) );
 a8707a <=( (not A300)  and  a8706a );
 a8708a <=( a8707a  and  a8702a );
 a8712a <=( A168  and  (not A169) );
 a8713a <=( A170  and  a8712a );
 a8717a <=( A201  and  (not A200) );
 a8718a <=( A199  and  a8717a );
 a8719a <=( a8718a  and  a8713a );
 a8723a <=( (not A299)  and  A298 );
 a8724a <=( A203  and  a8723a );
 a8728a <=( (not A302)  and  (not A301) );
 a8729a <=( (not A300)  and  a8728a );
 a8730a <=( a8729a  and  a8724a );
 a8734a <=( A168  and  (not A169) );
 a8735a <=( A170  and  a8734a );
 a8739a <=( A201  and  (not A200) );
 a8740a <=( A199  and  a8739a );
 a8741a <=( a8740a  and  a8735a );
 a8745a <=( A299  and  (not A298) );
 a8746a <=( A203  and  a8745a );
 a8750a <=( (not A302)  and  (not A301) );
 a8751a <=( (not A300)  and  a8750a );
 a8752a <=( a8751a  and  a8746a );
 a8756a <=( A168  and  (not A169) );
 a8757a <=( A170  and  a8756a );
 a8761a <=( (not A201)  and  (not A200) );
 a8762a <=( A199  and  a8761a );
 a8763a <=( a8762a  and  a8757a );
 a8767a <=( A298  and  (not A203) );
 a8768a <=( (not A202)  and  a8767a );
 a8772a <=( A301  and  A300 );
 a8773a <=( (not A299)  and  a8772a );
 a8774a <=( a8773a  and  a8768a );
 a8778a <=( A168  and  (not A169) );
 a8779a <=( A170  and  a8778a );
 a8783a <=( (not A201)  and  (not A200) );
 a8784a <=( A199  and  a8783a );
 a8785a <=( a8784a  and  a8779a );
 a8789a <=( A298  and  (not A203) );
 a8790a <=( (not A202)  and  a8789a );
 a8794a <=( A302  and  A300 );
 a8795a <=( (not A299)  and  a8794a );
 a8796a <=( a8795a  and  a8790a );
 a8800a <=( A168  and  (not A169) );
 a8801a <=( A170  and  a8800a );
 a8805a <=( (not A201)  and  (not A200) );
 a8806a <=( A199  and  a8805a );
 a8807a <=( a8806a  and  a8801a );
 a8811a <=( (not A298)  and  (not A203) );
 a8812a <=( (not A202)  and  a8811a );
 a8816a <=( A301  and  A300 );
 a8817a <=( A299  and  a8816a );
 a8818a <=( a8817a  and  a8812a );
 a8822a <=( A168  and  (not A169) );
 a8823a <=( A170  and  a8822a );
 a8827a <=( (not A201)  and  (not A200) );
 a8828a <=( A199  and  a8827a );
 a8829a <=( a8828a  and  a8823a );
 a8833a <=( (not A298)  and  (not A203) );
 a8834a <=( (not A202)  and  a8833a );
 a8838a <=( A302  and  A300 );
 a8839a <=( A299  and  a8838a );
 a8840a <=( a8839a  and  a8834a );
 a8844a <=( (not A168)  and  (not A169) );
 a8845a <=( A170  and  a8844a );
 a8849a <=( A201  and  (not A166) );
 a8850a <=( A167  and  a8849a );
 a8851a <=( a8850a  and  a8845a );
 a8855a <=( A298  and  (not A203) );
 a8856a <=( (not A202)  and  a8855a );
 a8860a <=( A301  and  A300 );
 a8861a <=( (not A299)  and  a8860a );
 a8862a <=( a8861a  and  a8856a );
 a8866a <=( (not A168)  and  (not A169) );
 a8867a <=( A170  and  a8866a );
 a8871a <=( A201  and  (not A166) );
 a8872a <=( A167  and  a8871a );
 a8873a <=( a8872a  and  a8867a );
 a8877a <=( A298  and  (not A203) );
 a8878a <=( (not A202)  and  a8877a );
 a8882a <=( A302  and  A300 );
 a8883a <=( (not A299)  and  a8882a );
 a8884a <=( a8883a  and  a8878a );
 a8888a <=( (not A168)  and  (not A169) );
 a8889a <=( A170  and  a8888a );
 a8893a <=( A201  and  (not A166) );
 a8894a <=( A167  and  a8893a );
 a8895a <=( a8894a  and  a8889a );
 a8899a <=( (not A298)  and  (not A203) );
 a8900a <=( (not A202)  and  a8899a );
 a8904a <=( A301  and  A300 );
 a8905a <=( A299  and  a8904a );
 a8906a <=( a8905a  and  a8900a );
 a8910a <=( (not A168)  and  (not A169) );
 a8911a <=( A170  and  a8910a );
 a8915a <=( A201  and  (not A166) );
 a8916a <=( A167  and  a8915a );
 a8917a <=( a8916a  and  a8911a );
 a8921a <=( (not A298)  and  (not A203) );
 a8922a <=( (not A202)  and  a8921a );
 a8926a <=( A302  and  A300 );
 a8927a <=( A299  and  a8926a );
 a8928a <=( a8927a  and  a8922a );
 a8932a <=( (not A168)  and  (not A169) );
 a8933a <=( A170  and  a8932a );
 a8937a <=( (not A201)  and  (not A166) );
 a8938a <=( A167  and  a8937a );
 a8939a <=( a8938a  and  a8933a );
 a8943a <=( (not A299)  and  A298 );
 a8944a <=( A202  and  a8943a );
 a8948a <=( (not A302)  and  (not A301) );
 a8949a <=( (not A300)  and  a8948a );
 a8950a <=( a8949a  and  a8944a );
 a8954a <=( (not A168)  and  (not A169) );
 a8955a <=( A170  and  a8954a );
 a8959a <=( (not A201)  and  (not A166) );
 a8960a <=( A167  and  a8959a );
 a8961a <=( a8960a  and  a8955a );
 a8965a <=( A299  and  (not A298) );
 a8966a <=( A202  and  a8965a );
 a8970a <=( (not A302)  and  (not A301) );
 a8971a <=( (not A300)  and  a8970a );
 a8972a <=( a8971a  and  a8966a );
 a8976a <=( (not A168)  and  (not A169) );
 a8977a <=( A170  and  a8976a );
 a8981a <=( (not A201)  and  (not A166) );
 a8982a <=( A167  and  a8981a );
 a8983a <=( a8982a  and  a8977a );
 a8987a <=( (not A299)  and  A298 );
 a8988a <=( A203  and  a8987a );
 a8992a <=( (not A302)  and  (not A301) );
 a8993a <=( (not A300)  and  a8992a );
 a8994a <=( a8993a  and  a8988a );
 a8998a <=( (not A168)  and  (not A169) );
 a8999a <=( A170  and  a8998a );
 a9003a <=( (not A201)  and  (not A166) );
 a9004a <=( A167  and  a9003a );
 a9005a <=( a9004a  and  a8999a );
 a9009a <=( A299  and  (not A298) );
 a9010a <=( A203  and  a9009a );
 a9014a <=( (not A302)  and  (not A301) );
 a9015a <=( (not A300)  and  a9014a );
 a9016a <=( a9015a  and  a9010a );
 a9020a <=( (not A168)  and  (not A169) );
 a9021a <=( A170  and  a9020a );
 a9025a <=( A199  and  (not A166) );
 a9026a <=( A167  and  a9025a );
 a9027a <=( a9026a  and  a9021a );
 a9031a <=( (not A299)  and  A298 );
 a9032a <=( A200  and  a9031a );
 a9036a <=( (not A302)  and  (not A301) );
 a9037a <=( (not A300)  and  a9036a );
 a9038a <=( a9037a  and  a9032a );
 a9042a <=( (not A168)  and  (not A169) );
 a9043a <=( A170  and  a9042a );
 a9047a <=( A199  and  (not A166) );
 a9048a <=( A167  and  a9047a );
 a9049a <=( a9048a  and  a9043a );
 a9053a <=( A299  and  (not A298) );
 a9054a <=( A200  and  a9053a );
 a9058a <=( (not A302)  and  (not A301) );
 a9059a <=( (not A300)  and  a9058a );
 a9060a <=( a9059a  and  a9054a );
 a9064a <=( (not A168)  and  (not A169) );
 a9065a <=( A170  and  a9064a );
 a9069a <=( (not A199)  and  (not A166) );
 a9070a <=( A167  and  a9069a );
 a9071a <=( a9070a  and  a9065a );
 a9075a <=( (not A299)  and  A298 );
 a9076a <=( (not A200)  and  a9075a );
 a9080a <=( (not A302)  and  (not A301) );
 a9081a <=( (not A300)  and  a9080a );
 a9082a <=( a9081a  and  a9076a );
 a9086a <=( (not A168)  and  (not A169) );
 a9087a <=( A170  and  a9086a );
 a9091a <=( (not A199)  and  (not A166) );
 a9092a <=( A167  and  a9091a );
 a9093a <=( a9092a  and  a9087a );
 a9097a <=( A299  and  (not A298) );
 a9098a <=( (not A200)  and  a9097a );
 a9102a <=( (not A302)  and  (not A301) );
 a9103a <=( (not A300)  and  a9102a );
 a9104a <=( a9103a  and  a9098a );
 a9108a <=( (not A168)  and  (not A169) );
 a9109a <=( A170  and  a9108a );
 a9113a <=( A201  and  A166 );
 a9114a <=( (not A167)  and  a9113a );
 a9115a <=( a9114a  and  a9109a );
 a9119a <=( A298  and  (not A203) );
 a9120a <=( (not A202)  and  a9119a );
 a9124a <=( A301  and  A300 );
 a9125a <=( (not A299)  and  a9124a );
 a9126a <=( a9125a  and  a9120a );
 a9130a <=( (not A168)  and  (not A169) );
 a9131a <=( A170  and  a9130a );
 a9135a <=( A201  and  A166 );
 a9136a <=( (not A167)  and  a9135a );
 a9137a <=( a9136a  and  a9131a );
 a9141a <=( A298  and  (not A203) );
 a9142a <=( (not A202)  and  a9141a );
 a9146a <=( A302  and  A300 );
 a9147a <=( (not A299)  and  a9146a );
 a9148a <=( a9147a  and  a9142a );
 a9152a <=( (not A168)  and  (not A169) );
 a9153a <=( A170  and  a9152a );
 a9157a <=( A201  and  A166 );
 a9158a <=( (not A167)  and  a9157a );
 a9159a <=( a9158a  and  a9153a );
 a9163a <=( (not A298)  and  (not A203) );
 a9164a <=( (not A202)  and  a9163a );
 a9168a <=( A301  and  A300 );
 a9169a <=( A299  and  a9168a );
 a9170a <=( a9169a  and  a9164a );
 a9174a <=( (not A168)  and  (not A169) );
 a9175a <=( A170  and  a9174a );
 a9179a <=( A201  and  A166 );
 a9180a <=( (not A167)  and  a9179a );
 a9181a <=( a9180a  and  a9175a );
 a9185a <=( (not A298)  and  (not A203) );
 a9186a <=( (not A202)  and  a9185a );
 a9190a <=( A302  and  A300 );
 a9191a <=( A299  and  a9190a );
 a9192a <=( a9191a  and  a9186a );
 a9196a <=( (not A168)  and  (not A169) );
 a9197a <=( A170  and  a9196a );
 a9201a <=( (not A201)  and  A166 );
 a9202a <=( (not A167)  and  a9201a );
 a9203a <=( a9202a  and  a9197a );
 a9207a <=( (not A299)  and  A298 );
 a9208a <=( A202  and  a9207a );
 a9212a <=( (not A302)  and  (not A301) );
 a9213a <=( (not A300)  and  a9212a );
 a9214a <=( a9213a  and  a9208a );
 a9218a <=( (not A168)  and  (not A169) );
 a9219a <=( A170  and  a9218a );
 a9223a <=( (not A201)  and  A166 );
 a9224a <=( (not A167)  and  a9223a );
 a9225a <=( a9224a  and  a9219a );
 a9229a <=( A299  and  (not A298) );
 a9230a <=( A202  and  a9229a );
 a9234a <=( (not A302)  and  (not A301) );
 a9235a <=( (not A300)  and  a9234a );
 a9236a <=( a9235a  and  a9230a );
 a9240a <=( (not A168)  and  (not A169) );
 a9241a <=( A170  and  a9240a );
 a9245a <=( (not A201)  and  A166 );
 a9246a <=( (not A167)  and  a9245a );
 a9247a <=( a9246a  and  a9241a );
 a9251a <=( (not A299)  and  A298 );
 a9252a <=( A203  and  a9251a );
 a9256a <=( (not A302)  and  (not A301) );
 a9257a <=( (not A300)  and  a9256a );
 a9258a <=( a9257a  and  a9252a );
 a9262a <=( (not A168)  and  (not A169) );
 a9263a <=( A170  and  a9262a );
 a9267a <=( (not A201)  and  A166 );
 a9268a <=( (not A167)  and  a9267a );
 a9269a <=( a9268a  and  a9263a );
 a9273a <=( A299  and  (not A298) );
 a9274a <=( A203  and  a9273a );
 a9278a <=( (not A302)  and  (not A301) );
 a9279a <=( (not A300)  and  a9278a );
 a9280a <=( a9279a  and  a9274a );
 a9284a <=( (not A168)  and  (not A169) );
 a9285a <=( A170  and  a9284a );
 a9289a <=( A199  and  A166 );
 a9290a <=( (not A167)  and  a9289a );
 a9291a <=( a9290a  and  a9285a );
 a9295a <=( (not A299)  and  A298 );
 a9296a <=( A200  and  a9295a );
 a9300a <=( (not A302)  and  (not A301) );
 a9301a <=( (not A300)  and  a9300a );
 a9302a <=( a9301a  and  a9296a );
 a9306a <=( (not A168)  and  (not A169) );
 a9307a <=( A170  and  a9306a );
 a9311a <=( A199  and  A166 );
 a9312a <=( (not A167)  and  a9311a );
 a9313a <=( a9312a  and  a9307a );
 a9317a <=( A299  and  (not A298) );
 a9318a <=( A200  and  a9317a );
 a9322a <=( (not A302)  and  (not A301) );
 a9323a <=( (not A300)  and  a9322a );
 a9324a <=( a9323a  and  a9318a );
 a9328a <=( (not A168)  and  (not A169) );
 a9329a <=( A170  and  a9328a );
 a9333a <=( (not A199)  and  A166 );
 a9334a <=( (not A167)  and  a9333a );
 a9335a <=( a9334a  and  a9329a );
 a9339a <=( (not A299)  and  A298 );
 a9340a <=( (not A200)  and  a9339a );
 a9344a <=( (not A302)  and  (not A301) );
 a9345a <=( (not A300)  and  a9344a );
 a9346a <=( a9345a  and  a9340a );
 a9350a <=( (not A168)  and  (not A169) );
 a9351a <=( A170  and  a9350a );
 a9355a <=( (not A199)  and  A166 );
 a9356a <=( (not A167)  and  a9355a );
 a9357a <=( a9356a  and  a9351a );
 a9361a <=( A299  and  (not A298) );
 a9362a <=( (not A200)  and  a9361a );
 a9366a <=( (not A302)  and  (not A301) );
 a9367a <=( (not A300)  and  a9366a );
 a9368a <=( a9367a  and  a9362a );
 a9372a <=( A168  and  (not A169) );
 a9373a <=( A170  and  a9372a );
 a9377a <=( (not A201)  and  A200 );
 a9378a <=( (not A199)  and  a9377a );
 a9379a <=( a9378a  and  a9373a );
 a9383a <=( A298  and  (not A203) );
 a9384a <=( (not A202)  and  a9383a );
 a9387a <=( (not A300)  and  (not A299) );
 a9390a <=( (not A302)  and  (not A301) );
 a9391a <=( a9390a  and  a9387a );
 a9392a <=( a9391a  and  a9384a );
 a9396a <=( A168  and  (not A169) );
 a9397a <=( A170  and  a9396a );
 a9401a <=( (not A201)  and  A200 );
 a9402a <=( (not A199)  and  a9401a );
 a9403a <=( a9402a  and  a9397a );
 a9407a <=( (not A298)  and  (not A203) );
 a9408a <=( (not A202)  and  a9407a );
 a9411a <=( (not A300)  and  A299 );
 a9414a <=( (not A302)  and  (not A301) );
 a9415a <=( a9414a  and  a9411a );
 a9416a <=( a9415a  and  a9408a );
 a9420a <=( A168  and  (not A169) );
 a9421a <=( A170  and  a9420a );
 a9425a <=( (not A201)  and  (not A200) );
 a9426a <=( A199  and  a9425a );
 a9427a <=( a9426a  and  a9421a );
 a9431a <=( A298  and  (not A203) );
 a9432a <=( (not A202)  and  a9431a );
 a9435a <=( (not A300)  and  (not A299) );
 a9438a <=( (not A302)  and  (not A301) );
 a9439a <=( a9438a  and  a9435a );
 a9440a <=( a9439a  and  a9432a );
 a9444a <=( A168  and  (not A169) );
 a9445a <=( A170  and  a9444a );
 a9449a <=( (not A201)  and  (not A200) );
 a9450a <=( A199  and  a9449a );
 a9451a <=( a9450a  and  a9445a );
 a9455a <=( (not A298)  and  (not A203) );
 a9456a <=( (not A202)  and  a9455a );
 a9459a <=( (not A300)  and  A299 );
 a9462a <=( (not A302)  and  (not A301) );
 a9463a <=( a9462a  and  a9459a );
 a9464a <=( a9463a  and  a9456a );
 a9468a <=( (not A168)  and  (not A169) );
 a9469a <=( A170  and  a9468a );
 a9473a <=( A201  and  (not A166) );
 a9474a <=( A167  and  a9473a );
 a9475a <=( a9474a  and  a9469a );
 a9479a <=( A298  and  (not A203) );
 a9480a <=( (not A202)  and  a9479a );
 a9483a <=( (not A300)  and  (not A299) );
 a9486a <=( (not A302)  and  (not A301) );
 a9487a <=( a9486a  and  a9483a );
 a9488a <=( a9487a  and  a9480a );
 a9492a <=( (not A168)  and  (not A169) );
 a9493a <=( A170  and  a9492a );
 a9497a <=( A201  and  (not A166) );
 a9498a <=( A167  and  a9497a );
 a9499a <=( a9498a  and  a9493a );
 a9503a <=( (not A298)  and  (not A203) );
 a9504a <=( (not A202)  and  a9503a );
 a9507a <=( (not A300)  and  A299 );
 a9510a <=( (not A302)  and  (not A301) );
 a9511a <=( a9510a  and  a9507a );
 a9512a <=( a9511a  and  a9504a );
 a9516a <=( (not A168)  and  (not A169) );
 a9517a <=( A170  and  a9516a );
 a9521a <=( A201  and  A166 );
 a9522a <=( (not A167)  and  a9521a );
 a9523a <=( a9522a  and  a9517a );
 a9527a <=( A298  and  (not A203) );
 a9528a <=( (not A202)  and  a9527a );
 a9531a <=( (not A300)  and  (not A299) );
 a9534a <=( (not A302)  and  (not A301) );
 a9535a <=( a9534a  and  a9531a );
 a9536a <=( a9535a  and  a9528a );
 a9540a <=( (not A168)  and  (not A169) );
 a9541a <=( A170  and  a9540a );
 a9545a <=( A201  and  A166 );
 a9546a <=( (not A167)  and  a9545a );
 a9547a <=( a9546a  and  a9541a );
 a9551a <=( (not A298)  and  (not A203) );
 a9552a <=( (not A202)  and  a9551a );
 a9555a <=( (not A300)  and  A299 );
 a9558a <=( (not A302)  and  (not A301) );
 a9559a <=( a9558a  and  a9555a );
 a9560a <=( a9559a  and  a9552a );


end x25_3x_behav;
