Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_15x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A72: buffer std_logic
);
end x25_15x;

architecture x25_15x_behav of x25_15x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1753a,a1754a,a1755a,a1756a,a1757a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1765a,a1766a,a1767a,a1768a,a1769a,a1770a,a1771a,a1772a,a1773a,a1774a,a1775a,a1776a,a1777a,a1778a,a1779a,a1780a,a1781a,a1782a,a1783a,a1784a,a1785a,a1786a,a1787a,a1788a,a1789a,a1790a,a1791a,a1792a,a1793a,a1794a,a1795a,a1796a,a1797a,a1798a,a1799a,a1800a,a1801a,a1802a,a1803a,a1804a,a1805a,a1806a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1816a,a1817a,a1818a,a1819a,a1820a,a1821a,a1822a,a1823a,a1824a,a1825a,a1826a,a1827a,a1828a,a1829a,a1830a,a1831a,a1832a,a1833a,a1834a,a1835a,a1836a,a1837a,a1838a,a1839a,a1840a,a1841a,a1842a,a1843a,a1844a,a1845a,a1846a,a1847a,a1848a,a1849a,a1850a,a1851a,a1852a,a1853a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1860a,a1861a,a1862a,a1863a,a1864a,a1865a,a1866a,a1867a,a1868a,a1869a,a1870a,a1871a,a1872a,a1873a,a1874a,a1875a,a1876a,a1877a,a1878a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1890a,a1891a,a1892a,a1893a,a1894a,a1895a,a1896a,a1897a,a1898a,a1899a,a1900a,a1901a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1910a,a1911a,a1912a,a1913a,a1914a,a1915a,a1916a,a1917a,a1918a,a1919a,a1920a,a1921a,a1922a,a1923a,a1924a,a1925a,a1926a,a1927a,a1928a,a1929a,a1930a,a1931a,a1932a,a1933a,a1934a,a1935a,a1936a,a1937a,a1938a,a1939a,a1940a,a1941a,a1942a,a1943a,a1944a,a1945a,a1946a,a1947a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1956a,a1957a,a1958a,a1959a,a1960a,a1961a,a1962a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1970a,a1971a,a1972a,a1973a,a1974a,a1975a,a1976a,a1977a,a1978a,a1979a,a1980a,a1981a,a1982a,a1983a,a1984a,a1985a,a1986a,a1987a,a1988a,a1989a,a1990a,a1991a,a1992a,a1993a,a1994a,a1995a,a1996a,a1997a,a1998a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2005a,a2006a,a2007a,a2008a,a2009a,a2010a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2025a,a2026a,a2027a,a2028a,a2029a,a2030a,a2031a,a2032a,a2033a,a2034a,a2035a,a2036a,a2037a,a2038a,a2039a,a2040a,a2041a,a2042a,a2043a,a2044a,a2045a,a2046a,a2047a,a2048a,a2049a,a2050a,a2051a,a2052a,a2053a,a2054a,a2055a,a2056a,a2057a,a2058a,a2059a,a2060a,a2061a,a2062a,a2063a,a2064a,a2065a,a2066a,a2067a,a2068a,a2069a,a2070a,a2071a,a2072a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2079a,a2080a,a2081a,a2082a,a2083a,a2084a,a2085a,a2086a,a2087a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2101a,a2102a,a2103a,a2104a,a2105a,a2106a,a2107a,a2108a,a2109a,a2110a,a2111a,a2112a,a2113a,a2114a,a2115a,a2116a,a2117a,a2118a,a2119a,a2120a,a2121a,a2122a,a2123a,a2124a,a2125a,a2126a,a2127a,a2128a,a2129a,a2130a,a2131a,a2132a,a2133a,a2134a,a2135a,a2136a,a2137a,a2138a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2145a,a2146a,a2147a,a2148a,a2149a,a2150a,a2151a,a2152a,a2153a,a2154a,a2155a,a2156a,a2157a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2164a,a2165a,a2166a,a2167a,a2168a,a2169a,a2170a,a2171a,a2172a,a2173a,a2174a,a2175a,a2176a,a2177a,a2178a,a2179a,a2180a,a2181a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2190a,a2191a,a2192a,a2193a,a2194a,a2195a,a2196a,a2197a,a2198a,a2199a,a2200a,a2201a,a2202a,a2203a,a2204a,a2205a,a2206a,a2207a,a2208a,a2209a,a2210a,a2211a,a2212a,a2213a,a2214a,a2215a,a2216a,a2217a,a2218a,a2219a,a2220a,a2221a,a2222a,a2223a,a2224a,a2225a,a2226a,a2227a,a2228a,a2229a,a2230a,a2231a,a2232a,a2233a,a2234a,a2235a,a2236a,a2237a,a2238a,a2239a,a2240a,a2241a,a2242a,a2243a,a2244a,a2245a,a2246a,a2247a,a2248a,a2249a,a2250a,a2251a,a2252a,a2253a,a2254a,a2255a,a2256a,a2257a,a2258a,a2259a,a2260a,a2261a,a2262a,a2263a,a2264a,a2265a,a2266a,a2267a,a2268a,a2269a,a2270a,a2271a,a2272a,a2273a,a2274a,a2275a,a2276a,a2277a,a2278a,a2279a,a2280a,a2281a,a2282a,a2283a,a2284a,a2285a,a2286a,a2287a,a2288a,a2289a,a2290a,a2291a,a2292a,a2293a,a2294a,a2295a,a2296a,a2297a,a2298a,a2299a,a2300a,a2301a,a2302a,a2303a,a2304a,a2305a,a2306a,a2307a,a2308a,a2309a,a2310a,a2311a,a2312a,a2313a,a2314a,a2315a,a2316a,a2317a,a2318a,a2319a,a2320a,a2321a,a2322a,a2323a,a2324a,a2325a,a2326a,a2327a,a2328a,a2329a,a2330a,a2331a,a2332a,a2333a,a2334a,a2335a,a2336a,a2337a,a2338a,a2339a,a2340a,a2341a,a2342a,a2343a,a2344a,a2345a,a2346a,a2347a,a2348a,a2349a,a2350a,a2351a,a2352a,a2353a,a2354a,a2355a,a2356a,a2357a,a2358a,a2359a,a2360a,a2361a,a2362a,a2363a,a2364a,a2365a,a2366a,a2367a,a2368a,a2369a,a2370a,a2371a,a2372a,a2373a,a2374a,a2375a,a2376a,a2377a,a2378a,a2379a,a2380a,a2381a,a2382a,a2383a,a2384a,a2385a,a2386a,a2387a,a2388a,a2389a,a2390a,a2391a,a2392a,a2393a,a2394a,a2395a,a2396a,a2397a,a2398a,a2399a,a2400a,a2401a,a2402a,a2403a,a2404a,a2405a,a2406a,a2407a,a2408a,a2409a,a2410a,a2411a,a2412a,a2413a,a2414a,a2415a,a2416a,a2417a,a2418a,a2419a,a2420a,a2421a,a2422a,a2423a,a2424a,a2425a,a2426a,a2427a,a2428a,a2429a,a2430a,a2431a,a2432a,a2433a,a2434a,a2435a,a2436a,a2437a,a2438a,a2439a,a2440a,a2441a,a2442a,a2443a,a2444a,a2445a,a2446a,a2447a,a2448a,a2449a,a2450a,a2451a,a2452a,a2453a,a2454a,a2455a,a2456a,a2457a,a2458a,a2459a,a2460a,a2461a,a2462a,a2463a,a2464a,a2465a,a2466a,a2467a,a2468a,a2469a,a2470a,a2471a,a2472a,a2473a,a2474a,a2475a,a2476a,a2477a,a2478a,a2479a,a2480a,a2481a,a2482a,a2483a,a2484a,a2485a,a2486a,a2487a,a2488a,a2489a,a2490a,a2491a,a2492a,a2493a,a2494a,a2495a,a2496a,a2497a,a2498a,a2499a,a2500a,a2501a,a2502a,a2503a,a2504a,a2505a,a2506a,a2507a,a2508a,a2509a,a2510a,a2511a,a2512a,a2513a,a2514a,a2515a,a2516a,a2517a,a2518a,a2519a,a2520a,a2521a,a2522a,a2523a,a2524a,a2525a,a2526a,a2527a,a2528a,a2529a,a2530a,a2531a,a2532a,a2533a,a2534a,a2535a,a2536a,a2537a,a2538a,a2539a,a2540a,a2541a,a2542a,a2543a,a2544a,a2545a,a2546a,a2547a,a2548a,a2549a,a2550a,a2553a,a2556a,a2557a,a2560a,a2564a,a2565a,a2566a,a2567a,a2570a,a2574a,a2575a,a2576a,a2579a,a2583a,a2584a,a2585a,a2586a,a2587a,a2590a,a2594a,a2595a,a2596a,a2599a,a2603a,a2604a,a2605a,a2606a,a2609a,a2613a,a2614a,a2615a,a2618a,a2622a,a2623a,a2624a,a2625a,a2626a,a2627a,a2630a,a2634a,a2635a,a2636a,a2639a,a2643a,a2644a,a2645a,a2646a,a2649a,a2653a,a2654a,a2655a,a2658a,a2662a,a2663a,a2664a,a2665a,a2666a,a2669a,a2673a,a2674a,a2675a,a2678a,a2682a,a2683a,a2684a,a2685a,a2688a,a2692a,a2693a,a2694a,a2697a,a2701a,a2702a,a2703a,a2704a,a2705a,a2706a,a2707a,a2710a,a2714a,a2715a,a2716a,a2719a,a2723a,a2724a,a2725a,a2726a,a2729a,a2733a,a2734a,a2735a,a2738a,a2742a,a2743a,a2744a,a2745a,a2746a,a2749a,a2753a,a2754a,a2755a,a2758a,a2762a,a2763a,a2764a,a2765a,a2768a,a2772a,a2773a,a2774a,a2777a,a2781a,a2782a,a2783a,a2784a,a2785a,a2786a,a2789a,a2793a,a2794a,a2795a,a2798a,a2802a,a2803a,a2804a,a2805a,a2808a,a2812a,a2813a,a2814a,a2817a,a2821a,a2822a,a2823a,a2824a,a2825a,a2828a,a2832a,a2833a,a2834a,a2837a,a2841a,a2842a,a2843a,a2844a,a2847a,a2851a,a2852a,a2853a,a2856a,a2860a,a2861a,a2862a,a2863a,a2864a,a2865a,a2866a,a2867a,a2870a,a2873a,a2874a,a2877a,a2881a,a2882a,a2883a,a2884a,a2887a,a2891a,a2892a,a2893a,a2896a,a2900a,a2901a,a2902a,a2903a,a2904a,a2907a,a2911a,a2912a,a2913a,a2916a,a2920a,a2921a,a2922a,a2923a,a2926a,a2930a,a2931a,a2932a,a2935a,a2939a,a2940a,a2941a,a2942a,a2943a,a2944a,a2947a,a2951a,a2952a,a2953a,a2956a,a2960a,a2961a,a2962a,a2963a,a2966a,a2970a,a2971a,a2972a,a2975a,a2979a,a2980a,a2981a,a2982a,a2983a,a2986a,a2990a,a2991a,a2992a,a2995a,a2999a,a3000a,a3001a,a3002a,a3005a,a3009a,a3010a,a3011a,a3014a,a3018a,a3019a,a3020a,a3021a,a3022a,a3023a,a3024a,a3027a,a3031a,a3032a,a3033a,a3036a,a3040a,a3041a,a3042a,a3043a,a3046a,a3050a,a3051a,a3052a,a3055a,a3059a,a3060a,a3061a,a3062a,a3063a,a3066a,a3070a,a3071a,a3072a,a3075a,a3079a,a3080a,a3081a,a3082a,a3085a,a3089a,a3090a,a3091a,a3094a,a3098a,a3099a,a3100a,a3101a,a3102a,a3103a,a3106a,a3110a,a3111a,a3112a,a3115a,a3119a,a3120a,a3121a,a3122a,a3125a,a3129a,a3130a,a3131a,a3134a,a3138a,a3139a,a3140a,a3141a,a3142a,a3145a,a3149a,a3150a,a3151a,a3154a,a3158a,a3159a,a3160a,a3161a,a3164a,a3168a,a3169a,a3170a,a3173a,a3177a,a3178a,a3179a,a3180a,a3181a,a3182a,a3183a,a3184a,a3185a,a3188a,a3191a,a3192a,a3195a,a3199a,a3200a,a3201a,a3202a,a3205a,a3209a,a3210a,a3211a,a3214a,a3218a,a3219a,a3220a,a3221a,a3222a,a3225a,a3229a,a3230a,a3231a,a3234a,a3238a,a3239a,a3240a,a3241a,a3244a,a3248a,a3249a,a3250a,a3253a,a3257a,a3258a,a3259a,a3260a,a3261a,a3262a,a3265a,a3269a,a3270a,a3271a,a3274a,a3278a,a3279a,a3280a,a3281a,a3284a,a3288a,a3289a,a3290a,a3293a,a3297a,a3298a,a3299a,a3300a,a3301a,a3304a,a3308a,a3309a,a3310a,a3313a,a3317a,a3318a,a3319a,a3320a,a3323a,a3327a,a3328a,a3329a,a3332a,a3336a,a3337a,a3338a,a3339a,a3340a,a3341a,a3342a,a3345a,a3349a,a3350a,a3351a,a3354a,a3358a,a3359a,a3360a,a3361a,a3364a,a3368a,a3369a,a3370a,a3373a,a3377a,a3378a,a3379a,a3380a,a3381a,a3384a,a3388a,a3389a,a3390a,a3393a,a3397a,a3398a,a3399a,a3400a,a3403a,a3407a,a3408a,a3409a,a3412a,a3416a,a3417a,a3418a,a3419a,a3420a,a3421a,a3424a,a3428a,a3429a,a3430a,a3433a,a3437a,a3438a,a3439a,a3440a,a3443a,a3447a,a3448a,a3449a,a3452a,a3456a,a3457a,a3458a,a3459a,a3460a,a3463a,a3467a,a3468a,a3469a,a3472a,a3476a,a3477a,a3478a,a3479a,a3482a,a3486a,a3487a,a3488a,a3491a,a3495a,a3496a,a3497a,a3498a,a3499a,a3500a,a3501a,a3502a,a3505a,a3509a,a3510a,a3511a,a3514a,a3518a,a3519a,a3520a,a3521a,a3524a,a3528a,a3529a,a3530a,a3533a,a3537a,a3538a,a3539a,a3540a,a3541a,a3544a,a3548a,a3549a,a3550a,a3553a,a3557a,a3558a,a3559a,a3560a,a3563a,a3567a,a3568a,a3569a,a3572a,a3576a,a3577a,a3578a,a3579a,a3580a,a3581a,a3584a,a3588a,a3589a,a3590a,a3593a,a3597a,a3598a,a3599a,a3600a,a3603a,a3607a,a3608a,a3609a,a3612a,a3616a,a3617a,a3618a,a3619a,a3620a,a3623a,a3627a,a3628a,a3629a,a3632a,a3636a,a3637a,a3638a,a3639a,a3642a,a3646a,a3647a,a3648a,a3651a,a3655a,a3656a,a3657a,a3658a,a3659a,a3660a,a3661a,a3664a,a3668a,a3669a,a3670a,a3673a,a3677a,a3678a,a3679a,a3680a,a3683a,a3687a,a3688a,a3689a,a3692a,a3696a,a3697a,a3698a,a3699a,a3700a,a3703a,a3707a,a3708a,a3709a,a3712a,a3716a,a3717a,a3718a,a3719a,a3722a,a3726a,a3727a,a3728a,a3731a,a3735a,a3736a,a3737a,a3738a,a3739a,a3740a,a3743a,a3747a,a3748a,a3749a,a3752a,a3756a,a3757a,a3758a,a3759a,a3762a,a3766a,a3767a,a3768a,a3771a,a3775a,a3776a,a3777a,a3778a,a3779a,a3782a,a3786a,a3787a,a3788a,a3791a,a3795a,a3796a,a3797a,a3798a,a3801a,a3805a,a3806a,a3807a,a3810a,a3814a,a3815a,a3816a,a3817a,a3818a,a3819a,a3820a,a3821a,a3822a,a3823a,a3826a,a3829a,a3830a,a3833a,a3837a,a3838a,a3839a,a3840a,a3843a,a3847a,a3848a,a3849a,a3852a,a3856a,a3857a,a3858a,a3859a,a3860a,a3863a,a3867a,a3868a,a3869a,a3872a,a3876a,a3877a,a3878a,a3879a,a3882a,a3886a,a3887a,a3888a,a3891a,a3895a,a3896a,a3897a,a3898a,a3899a,a3900a,a3903a,a3907a,a3908a,a3909a,a3912a,a3916a,a3917a,a3918a,a3919a,a3922a,a3926a,a3927a,a3928a,a3931a,a3935a,a3936a,a3937a,a3938a,a3939a,a3942a,a3946a,a3947a,a3948a,a3951a,a3955a,a3956a,a3957a,a3958a,a3961a,a3965a,a3966a,a3967a,a3970a,a3974a,a3975a,a3976a,a3977a,a3978a,a3979a,a3980a,a3983a,a3987a,a3988a,a3989a,a3992a,a3996a,a3997a,a3998a,a3999a,a4002a,a4006a,a4007a,a4008a,a4011a,a4015a,a4016a,a4017a,a4018a,a4019a,a4022a,a4026a,a4027a,a4028a,a4031a,a4035a,a4036a,a4037a,a4038a,a4041a,a4045a,a4046a,a4047a,a4050a,a4054a,a4055a,a4056a,a4057a,a4058a,a4059a,a4062a,a4066a,a4067a,a4068a,a4071a,a4075a,a4076a,a4077a,a4078a,a4081a,a4085a,a4086a,a4087a,a4090a,a4094a,a4095a,a4096a,a4097a,a4098a,a4101a,a4105a,a4106a,a4107a,a4110a,a4114a,a4115a,a4116a,a4117a,a4120a,a4124a,a4125a,a4126a,a4129a,a4133a,a4134a,a4135a,a4136a,a4137a,a4138a,a4139a,a4140a,a4143a,a4147a,a4148a,a4149a,a4152a,a4156a,a4157a,a4158a,a4159a,a4162a,a4166a,a4167a,a4168a,a4171a,a4175a,a4176a,a4177a,a4178a,a4179a,a4182a,a4186a,a4187a,a4188a,a4191a,a4195a,a4196a,a4197a,a4198a,a4201a,a4205a,a4206a,a4207a,a4210a,a4214a,a4215a,a4216a,a4217a,a4218a,a4219a,a4222a,a4226a,a4227a,a4228a,a4231a,a4235a,a4236a,a4237a,a4238a,a4241a,a4245a,a4246a,a4247a,a4250a,a4254a,a4255a,a4256a,a4257a,a4258a,a4261a,a4265a,a4266a,a4267a,a4270a,a4274a,a4275a,a4276a,a4277a,a4280a,a4284a,a4285a,a4286a,a4289a,a4293a,a4294a,a4295a,a4296a,a4297a,a4298a,a4299a,a4302a,a4306a,a4307a,a4308a,a4311a,a4315a,a4316a,a4317a,a4318a,a4321a,a4325a,a4326a,a4327a,a4330a,a4334a,a4335a,a4336a,a4337a,a4338a,a4341a,a4345a,a4346a,a4347a,a4350a,a4354a,a4355a,a4356a,a4357a,a4360a,a4364a,a4365a,a4366a,a4369a,a4373a,a4374a,a4375a,a4376a,a4377a,a4378a,a4381a,a4385a,a4386a,a4387a,a4390a,a4394a,a4395a,a4396a,a4397a,a4400a,a4404a,a4405a,a4406a,a4409a,a4413a,a4414a,a4415a,a4416a,a4417a,a4420a,a4424a,a4425a,a4426a,a4429a,a4433a,a4434a,a4435a,a4436a,a4439a,a4443a,a4444a,a4445a,a4448a,a4452a,a4453a,a4454a,a4455a,a4456a,a4457a,a4458a,a4459a,a4460a,a4463a,a4466a,a4467a,a4470a,a4474a,a4475a,a4476a,a4477a,a4480a,a4484a,a4485a,a4486a,a4489a,a4493a,a4494a,a4495a,a4496a,a4497a,a4500a,a4504a,a4505a,a4506a,a4509a,a4513a,a4514a,a4515a,a4516a,a4519a,a4523a,a4524a,a4525a,a4528a,a4532a,a4533a,a4534a,a4535a,a4536a,a4537a,a4540a,a4544a,a4545a,a4546a,a4549a,a4553a,a4554a,a4555a,a4556a,a4559a,a4563a,a4564a,a4565a,a4568a,a4572a,a4573a,a4574a,a4575a,a4576a,a4579a,a4583a,a4584a,a4585a,a4588a,a4592a,a4593a,a4594a,a4595a,a4598a,a4602a,a4603a,a4604a,a4607a,a4611a,a4612a,a4613a,a4614a,a4615a,a4616a,a4617a,a4620a,a4624a,a4625a,a4626a,a4629a,a4633a,a4634a,a4635a,a4636a,a4639a,a4643a,a4644a,a4645a,a4648a,a4652a,a4653a,a4654a,a4655a,a4656a,a4659a,a4663a,a4664a,a4665a,a4668a,a4672a,a4673a,a4674a,a4675a,a4678a,a4682a,a4683a,a4684a,a4687a,a4691a,a4692a,a4693a,a4694a,a4695a,a4696a,a4699a,a4703a,a4704a,a4705a,a4708a,a4712a,a4713a,a4714a,a4715a,a4718a,a4722a,a4723a,a4724a,a4727a,a4731a,a4732a,a4733a,a4734a,a4735a,a4738a,a4742a,a4743a,a4744a,a4747a,a4751a,a4752a,a4753a,a4754a,a4757a,a4761a,a4762a,a4763a,a4766a,a4770a,a4771a,a4772a,a4773a,a4774a,a4775a,a4776a,a4777a,a4780a,a4784a,a4785a,a4786a,a4789a,a4793a,a4794a,a4795a,a4796a,a4799a,a4803a,a4804a,a4805a,a4808a,a4812a,a4813a,a4814a,a4815a,a4816a,a4819a,a4823a,a4824a,a4825a,a4828a,a4832a,a4833a,a4834a,a4835a,a4838a,a4842a,a4843a,a4844a,a4847a,a4851a,a4852a,a4853a,a4854a,a4855a,a4856a,a4859a,a4863a,a4864a,a4865a,a4868a,a4872a,a4873a,a4874a,a4875a,a4878a,a4882a,a4883a,a4884a,a4887a,a4891a,a4892a,a4893a,a4894a,a4895a,a4898a,a4902a,a4903a,a4904a,a4907a,a4911a,a4912a,a4913a,a4914a,a4917a,a4921a,a4922a,a4923a,a4926a,a4930a,a4931a,a4932a,a4933a,a4934a,a4935a,a4936a,a4939a,a4943a,a4944a,a4945a,a4948a,a4952a,a4953a,a4954a,a4955a,a4958a,a4962a,a4963a,a4964a,a4967a,a4971a,a4972a,a4973a,a4974a,a4975a,a4978a,a4982a,a4983a,a4984a,a4987a,a4991a,a4992a,a4993a,a4994a,a4997a,a5001a,a5002a,a5003a,a5006a,a5010a,a5011a,a5012a,a5013a,a5014a,a5015a,a5018a,a5022a,a5023a,a5024a,a5027a,a5031a,a5032a,a5033a,a5034a,a5037a,a5041a,a5042a,a5043a,a5046a,a5050a,a5051a,a5052a,a5053a,a5054a,a5057a,a5061a,a5062a,a5063a,a5066a,a5070a,a5071a,a5072a,a5073a,a5076a,a5080a,a5081a,a5082a,a5085a,a5089a,a5090a,a5091a,a5092a,a5093a,a5094a,a5095a,a5096a,a5097a,a5098a,a5099a,a5102a,a5105a,a5106a,a5109a,a5113a,a5114a,a5115a,a5116a,a5119a,a5123a,a5124a,a5125a,a5128a,a5132a,a5133a,a5134a,a5135a,a5136a,a5139a,a5143a,a5144a,a5145a,a5148a,a5152a,a5153a,a5154a,a5155a,a5158a,a5162a,a5163a,a5164a,a5167a,a5171a,a5172a,a5173a,a5174a,a5175a,a5176a,a5179a,a5183a,a5184a,a5185a,a5188a,a5192a,a5193a,a5194a,a5195a,a5198a,a5202a,a5203a,a5204a,a5207a,a5211a,a5212a,a5213a,a5214a,a5215a,a5218a,a5222a,a5223a,a5224a,a5227a,a5231a,a5232a,a5233a,a5234a,a5237a,a5241a,a5242a,a5243a,a5246a,a5250a,a5251a,a5252a,a5253a,a5254a,a5255a,a5256a,a5259a,a5263a,a5264a,a5265a,a5268a,a5272a,a5273a,a5274a,a5275a,a5278a,a5282a,a5283a,a5284a,a5287a,a5291a,a5292a,a5293a,a5294a,a5295a,a5298a,a5302a,a5303a,a5304a,a5307a,a5311a,a5312a,a5313a,a5314a,a5317a,a5321a,a5322a,a5323a,a5326a,a5330a,a5331a,a5332a,a5333a,a5334a,a5335a,a5338a,a5342a,a5343a,a5344a,a5347a,a5351a,a5352a,a5353a,a5354a,a5357a,a5361a,a5362a,a5363a,a5366a,a5370a,a5371a,a5372a,a5373a,a5374a,a5377a,a5381a,a5382a,a5383a,a5386a,a5390a,a5391a,a5392a,a5393a,a5396a,a5400a,a5401a,a5402a,a5405a,a5409a,a5410a,a5411a,a5412a,a5413a,a5414a,a5415a,a5416a,a5419a,a5422a,a5423a,a5426a,a5430a,a5431a,a5432a,a5433a,a5436a,a5440a,a5441a,a5442a,a5445a,a5449a,a5450a,a5451a,a5452a,a5453a,a5456a,a5460a,a5461a,a5462a,a5465a,a5469a,a5470a,a5471a,a5472a,a5475a,a5479a,a5480a,a5481a,a5484a,a5488a,a5489a,a5490a,a5491a,a5492a,a5493a,a5496a,a5500a,a5501a,a5502a,a5505a,a5509a,a5510a,a5511a,a5512a,a5515a,a5519a,a5520a,a5521a,a5524a,a5528a,a5529a,a5530a,a5531a,a5532a,a5535a,a5539a,a5540a,a5541a,a5544a,a5548a,a5549a,a5550a,a5551a,a5554a,a5558a,a5559a,a5560a,a5563a,a5567a,a5568a,a5569a,a5570a,a5571a,a5572a,a5573a,a5576a,a5580a,a5581a,a5582a,a5585a,a5589a,a5590a,a5591a,a5592a,a5595a,a5599a,a5600a,a5601a,a5604a,a5608a,a5609a,a5610a,a5611a,a5612a,a5615a,a5619a,a5620a,a5621a,a5624a,a5628a,a5629a,a5630a,a5631a,a5634a,a5638a,a5639a,a5640a,a5643a,a5647a,a5648a,a5649a,a5650a,a5651a,a5652a,a5655a,a5659a,a5660a,a5661a,a5664a,a5668a,a5669a,a5670a,a5671a,a5674a,a5678a,a5679a,a5680a,a5683a,a5687a,a5688a,a5689a,a5690a,a5691a,a5694a,a5698a,a5699a,a5700a,a5703a,a5707a,a5708a,a5709a,a5710a,a5713a,a5717a,a5718a,a5719a,a5722a,a5726a,a5727a,a5728a,a5729a,a5730a,a5731a,a5732a,a5733a,a5734a,a5737a,a5740a,a5741a,a5744a,a5748a,a5749a,a5750a,a5751a,a5754a,a5758a,a5759a,a5760a,a5763a,a5767a,a5768a,a5769a,a5770a,a5771a,a5774a,a5778a,a5779a,a5780a,a5783a,a5787a,a5788a,a5789a,a5790a,a5793a,a5797a,a5798a,a5799a,a5802a,a5806a,a5807a,a5808a,a5809a,a5810a,a5811a,a5814a,a5818a,a5819a,a5820a,a5823a,a5827a,a5828a,a5829a,a5830a,a5833a,a5837a,a5838a,a5839a,a5842a,a5846a,a5847a,a5848a,a5849a,a5850a,a5853a,a5857a,a5858a,a5859a,a5862a,a5866a,a5867a,a5868a,a5869a,a5872a,a5876a,a5877a,a5878a,a5881a,a5885a,a5886a,a5887a,a5888a,a5889a,a5890a,a5891a,a5894a,a5898a,a5899a,a5900a,a5903a,a5907a,a5908a,a5909a,a5910a,a5913a,a5917a,a5918a,a5919a,a5922a,a5926a,a5927a,a5928a,a5929a,a5930a,a5933a,a5937a,a5938a,a5939a,a5942a,a5946a,a5947a,a5948a,a5949a,a5952a,a5956a,a5957a,a5958a,a5961a,a5965a,a5966a,a5967a,a5968a,a5969a,a5970a,a5973a,a5977a,a5978a,a5979a,a5982a,a5986a,a5987a,a5988a,a5989a,a5992a,a5996a,a5997a,a5998a,a6001a,a6005a,a6006a,a6007a,a6008a,a6009a,a6012a,a6016a,a6017a,a6018a,a6021a,a6025a,a6026a,a6027a,a6028a,a6031a,a6035a,a6036a,a6037a,a6040a,a6044a,a6045a,a6046a,a6047a,a6048a,a6049a,a6050a,a6051a,a6054a,a6058a,a6059a,a6060a,a6063a,a6067a,a6068a,a6069a,a6070a,a6073a,a6077a,a6078a,a6079a,a6082a,a6086a,a6087a,a6088a,a6089a,a6090a,a6093a,a6097a,a6098a,a6099a,a6102a,a6106a,a6107a,a6108a,a6109a,a6112a,a6116a,a6117a,a6118a,a6121a,a6125a,a6126a,a6127a,a6128a,a6129a,a6130a,a6133a,a6137a,a6138a,a6139a,a6142a,a6146a,a6147a,a6148a,a6149a,a6152a,a6156a,a6157a,a6158a,a6161a,a6165a,a6166a,a6167a,a6168a,a6169a,a6172a,a6176a,a6177a,a6178a,a6181a,a6185a,a6186a,a6187a,a6188a,a6191a,a6195a,a6196a,a6197a,a6200a,a6204a,a6205a,a6206a,a6207a,a6208a,a6209a,a6210a,a6213a,a6217a,a6218a,a6219a,a6222a,a6226a,a6227a,a6228a,a6229a,a6232a,a6236a,a6237a,a6238a,a6241a,a6245a,a6246a,a6247a,a6248a,a6249a,a6252a,a6256a,a6257a,a6258a,a6261a,a6265a,a6266a,a6267a,a6268a,a6271a,a6275a,a6276a,a6277a,a6280a,a6284a,a6285a,a6286a,a6287a,a6288a,a6289a,a6292a,a6296a,a6297a,a6298a,a6301a,a6305a,a6306a,a6307a,a6308a,a6311a,a6315a,a6316a,a6317a,a6320a,a6324a,a6325a,a6326a,a6327a,a6328a,a6331a,a6335a,a6336a,a6337a,a6340a,a6344a,a6345a,a6346a,a6347a,a6350a,a6354a,a6355a,a6356a,a6359a,a6363a,a6364a,a6365a,a6366a,a6367a,a6368a,a6369a,a6370a,a6371a,a6372a,a6375a,a6378a,a6379a,a6382a,a6386a,a6387a,a6388a,a6389a,a6392a,a6396a,a6397a,a6398a,a6401a,a6405a,a6406a,a6407a,a6408a,a6409a,a6412a,a6416a,a6417a,a6418a,a6421a,a6425a,a6426a,a6427a,a6428a,a6431a,a6435a,a6436a,a6437a,a6440a,a6444a,a6445a,a6446a,a6447a,a6448a,a6449a,a6452a,a6456a,a6457a,a6458a,a6461a,a6465a,a6466a,a6467a,a6468a,a6471a,a6475a,a6476a,a6477a,a6480a,a6484a,a6485a,a6486a,a6487a,a6488a,a6491a,a6495a,a6496a,a6497a,a6500a,a6504a,a6505a,a6506a,a6507a,a6510a,a6514a,a6515a,a6516a,a6519a,a6523a,a6524a,a6525a,a6526a,a6527a,a6528a,a6529a,a6532a,a6536a,a6537a,a6538a,a6541a,a6545a,a6546a,a6547a,a6548a,a6551a,a6555a,a6556a,a6557a,a6560a,a6564a,a6565a,a6566a,a6567a,a6568a,a6571a,a6575a,a6576a,a6577a,a6580a,a6584a,a6585a,a6586a,a6587a,a6590a,a6594a,a6595a,a6596a,a6599a,a6603a,a6604a,a6605a,a6606a,a6607a,a6608a,a6611a,a6615a,a6616a,a6617a,a6620a,a6624a,a6625a,a6626a,a6627a,a6630a,a6634a,a6635a,a6636a,a6639a,a6643a,a6644a,a6645a,a6646a,a6647a,a6650a,a6654a,a6655a,a6656a,a6659a,a6663a,a6664a,a6665a,a6666a,a6669a,a6673a,a6674a,a6675a,a6678a,a6682a,a6683a,a6684a,a6685a,a6686a,a6687a,a6688a,a6689a,a6692a,a6696a,a6697a,a6698a,a6701a,a6705a,a6706a,a6707a,a6708a,a6711a,a6715a,a6716a,a6717a,a6720a,a6724a,a6725a,a6726a,a6727a,a6728a,a6731a,a6735a,a6736a,a6737a,a6740a,a6744a,a6745a,a6746a,a6747a,a6750a,a6754a,a6755a,a6756a,a6759a,a6763a,a6764a,a6765a,a6766a,a6767a,a6768a,a6771a,a6775a,a6776a,a6777a,a6780a,a6784a,a6785a,a6786a,a6787a,a6790a,a6794a,a6795a,a6796a,a6799a,a6803a,a6804a,a6805a,a6806a,a6807a,a6810a,a6814a,a6815a,a6816a,a6819a,a6823a,a6824a,a6825a,a6826a,a6829a,a6833a,a6834a,a6835a,a6838a,a6842a,a6843a,a6844a,a6845a,a6846a,a6847a,a6848a,a6851a,a6855a,a6856a,a6857a,a6860a,a6864a,a6865a,a6866a,a6867a,a6870a,a6874a,a6875a,a6876a,a6879a,a6883a,a6884a,a6885a,a6886a,a6887a,a6890a,a6894a,a6895a,a6896a,a6899a,a6903a,a6904a,a6905a,a6906a,a6909a,a6913a,a6914a,a6915a,a6918a,a6922a,a6923a,a6924a,a6925a,a6926a,a6927a,a6930a,a6934a,a6935a,a6936a,a6939a,a6943a,a6944a,a6945a,a6946a,a6949a,a6953a,a6954a,a6955a,a6958a,a6962a,a6963a,a6964a,a6965a,a6966a,a6969a,a6973a,a6974a,a6975a,a6978a,a6982a,a6983a,a6984a,a6985a,a6988a,a6992a,a6993a,a6994a,a6997a,a7001a,a7002a,a7003a,a7004a,a7005a,a7006a,a7007a,a7008a,a7009a,a7012a,a7015a,a7016a,a7019a,a7023a,a7024a,a7025a,a7026a,a7029a,a7033a,a7034a,a7035a,a7038a,a7042a,a7043a,a7044a,a7045a,a7046a,a7049a,a7053a,a7054a,a7055a,a7058a,a7062a,a7063a,a7064a,a7065a,a7068a,a7072a,a7073a,a7074a,a7077a,a7081a,a7082a,a7083a,a7084a,a7085a,a7086a,a7089a,a7093a,a7094a,a7095a,a7098a,a7102a,a7103a,a7104a,a7105a,a7108a,a7112a,a7113a,a7114a,a7117a,a7121a,a7122a,a7123a,a7124a,a7125a,a7128a,a7132a,a7133a,a7134a,a7137a,a7141a,a7142a,a7143a,a7144a,a7147a,a7151a,a7152a,a7153a,a7156a,a7160a,a7161a,a7162a,a7163a,a7164a,a7165a,a7166a,a7169a,a7173a,a7174a,a7175a,a7178a,a7182a,a7183a,a7184a,a7185a,a7188a,a7192a,a7193a,a7194a,a7197a,a7201a,a7202a,a7203a,a7204a,a7205a,a7208a,a7212a,a7213a,a7214a,a7217a,a7221a,a7222a,a7223a,a7224a,a7227a,a7231a,a7232a,a7233a,a7236a,a7240a,a7241a,a7242a,a7243a,a7244a,a7245a,a7248a,a7252a,a7253a,a7254a,a7257a,a7261a,a7262a,a7263a,a7264a,a7267a,a7271a,a7272a,a7273a,a7276a,a7280a,a7281a,a7282a,a7283a,a7284a,a7287a,a7291a,a7292a,a7293a,a7296a,a7300a,a7301a,a7302a,a7303a,a7306a,a7310a,a7311a,a7312a,a7315a,a7319a,a7320a,a7321a,a7322a,a7323a,a7324a,a7325a,a7326a,a7329a,a7333a,a7334a,a7335a,a7338a,a7342a,a7343a,a7344a,a7345a,a7348a,a7352a,a7353a,a7354a,a7357a,a7361a,a7362a,a7363a,a7364a,a7365a,a7368a,a7372a,a7373a,a7374a,a7377a,a7381a,a7382a,a7383a,a7384a,a7387a,a7391a,a7392a,a7393a,a7396a,a7400a,a7401a,a7402a,a7403a,a7404a,a7405a,a7408a,a7412a,a7413a,a7414a,a7417a,a7421a,a7422a,a7423a,a7424a,a7427a,a7431a,a7432a,a7433a,a7436a,a7440a,a7441a,a7442a,a7443a,a7444a,a7447a,a7451a,a7452a,a7453a,a7456a,a7460a,a7461a,a7462a,a7463a,a7466a,a7470a,a7471a,a7472a,a7475a,a7479a,a7480a,a7481a,a7482a,a7483a,a7484a,a7485a,a7488a,a7492a,a7493a,a7494a,a7497a,a7501a,a7502a,a7503a,a7504a,a7507a,a7511a,a7512a,a7513a,a7516a,a7520a,a7521a,a7522a,a7523a,a7524a,a7527a,a7531a,a7532a,a7533a,a7536a,a7540a,a7541a,a7542a,a7543a,a7546a,a7550a,a7551a,a7552a,a7555a,a7559a,a7560a,a7561a,a7562a,a7563a,a7564a,a7567a,a7571a,a7572a,a7573a,a7576a,a7580a,a7581a,a7582a,a7583a,a7586a,a7590a,a7591a,a7592a,a7595a,a7599a,a7600a,a7601a,a7602a,a7603a,a7606a,a7610a,a7611a,a7612a,a7615a,a7619a,a7620a,a7621a,a7622a,a7625a,a7629a,a7630a,a7631a,a7634a,a7638a,a7639a,a7640a,a7641a,a7642a,a7643a,a7644a,a7645a,a7646a,a7647a,a7648a,a7652a,a7653a,a7657a,a7658a,a7662a,a7663a,a7667a,a7668a,a7672a,a7673a,a7677a,a7678a,a7682a,a7683a,a7687a,a7688a,a7692a,a7693a,a7696a,a7699a,a7700a,a7704a,a7705a,a7708a,a7711a,a7712a,a7716a,a7717a,a7720a,a7723a,a7724a,a7728a,a7729a,a7732a,a7735a,a7736a,a7740a,a7741a,a7744a,a7747a,a7748a,a7752a,a7753a,a7756a,a7759a,a7760a,a7764a,a7765a,a7768a,a7771a,a7772a,a7776a,a7777a,a7780a,a7783a,a7784a,a7788a,a7789a,a7792a,a7795a,a7796a,a7800a,a7801a,a7804a,a7807a,a7808a,a7812a,a7813a,a7816a,a7819a,a7820a,a7824a,a7825a,a7828a,a7831a,a7832a,a7836a,a7837a,a7840a,a7843a,a7844a,a7848a,a7849a,a7852a,a7855a,a7856a,a7860a,a7861a,a7864a,a7867a,a7868a,a7872a,a7873a,a7876a,a7879a,a7880a,a7884a,a7885a,a7888a,a7891a,a7892a,a7896a,a7897a,a7900a,a7903a,a7904a,a7908a,a7909a,a7912a,a7915a,a7916a,a7920a,a7921a,a7924a,a7927a,a7928a,a7932a,a7933a,a7936a,a7939a,a7940a,a7944a,a7945a,a7948a,a7951a,a7952a,a7956a,a7957a,a7960a,a7963a,a7964a,a7968a,a7969a,a7972a,a7975a,a7976a,a7980a,a7981a,a7984a,a7987a,a7988a,a7992a,a7993a,a7996a,a7999a,a8000a,a8003a,a8006a,a8007a,a8010a,a8013a,a8014a,a8017a,a8020a,a8021a,a8024a,a8027a,a8028a,a8031a,a8034a,a8035a,a8038a,a8041a,a8042a,a8045a,a8048a,a8049a,a8052a,a8055a,a8056a,a8059a,a8062a,a8063a,a8066a,a8069a,a8070a,a8073a,a8076a,a8077a,a8080a,a8083a,a8084a,a8087a,a8090a,a8091a,a8094a,a8097a,a8098a,a8101a,a8104a,a8105a,a8108a,a8111a,a8112a,a8115a,a8118a,a8119a,a8122a,a8125a,a8126a,a8129a,a8132a,a8133a,a8136a,a8139a,a8140a,a8143a,a8146a,a8147a,a8150a,a8153a,a8154a,a8157a,a8160a,a8161a,a8164a,a8167a,a8168a,a8171a,a8174a,a8175a,a8178a,a8181a,a8182a,a8185a,a8188a,a8189a,a8192a,a8195a,a8196a,a8199a,a8202a,a8203a,a8206a,a8209a,a8210a,a8213a,a8216a,a8217a,a8220a,a8223a,a8224a,a8227a,a8230a,a8231a,a8234a,a8237a,a8238a,a8241a,a8244a,a8245a,a8248a,a8251a,a8252a,a8255a,a8258a,a8259a,a8262a,a8265a,a8266a,a8269a,a8272a,a8273a,a8276a,a8279a,a8280a,a8283a,a8286a,a8287a,a8290a,a8293a,a8294a,a8297a,a8300a,a8301a,a8304a,a8307a,a8308a,a8311a,a8314a,a8315a,a8318a,a8321a,a8322a,a8325a,a8328a,a8329a,a8332a,a8335a,a8336a,a8339a,a8342a,a8343a,a8346a,a8349a,a8350a,a8353a,a8356a,a8357a,a8360a,a8363a,a8364a,a8367a,a8370a,a8371a,a8374a,a8377a,a8378a,a8381a,a8384a,a8385a,a8388a,a8391a,a8392a,a8395a,a8398a,a8399a,a8402a,a8405a,a8406a,a8409a,a8412a,a8413a,a8416a,a8419a,a8420a,a8423a,a8426a,a8427a,a8430a,a8433a,a8434a,a8437a,a8440a,a8441a,a8444a,a8447a,a8448a,a8451a,a8454a,a8455a,a8458a,a8461a,a8462a,a8465a,a8468a,a8469a,a8472a,a8475a,a8476a,a8479a,a8482a,a8483a,a8486a,a8489a,a8490a,a8493a,a8496a,a8497a,a8500a,a8503a,a8504a,a8507a,a8510a,a8511a,a8514a,a8517a,a8518a,a8521a,a8524a,a8525a,a8528a,a8531a,a8532a,a8535a,a8538a,a8539a,a8542a,a8545a,a8546a,a8549a,a8552a,a8553a,a8556a,a8559a,a8560a,a8563a,a8566a,a8567a,a8570a,a8573a,a8574a,a8577a,a8580a,a8581a,a8584a,a8587a,a8588a,a8591a,a8594a,a8595a,a8598a,a8601a,a8602a,a8605a,a8608a,a8609a,a8612a,a8615a,a8616a,a8619a,a8622a,a8623a,a8626a,a8629a,a8630a,a8633a,a8636a,a8637a,a8640a,a8643a,a8644a,a8647a,a8650a,a8651a,a8654a,a8657a,a8658a,a8661a,a8664a,a8665a,a8668a,a8671a,a8672a,a8675a,a8678a,a8679a,a8682a,a8685a,a8686a,a8689a,a8692a,a8693a,a8696a,a8699a,a8700a,a8703a,a8706a,a8707a,a8710a,a8713a,a8714a,a8717a,a8720a,a8721a,a8724a,a8727a,a8728a,a8731a,a8734a,a8735a,a8738a,a8741a,a8742a,a8745a,a8748a,a8749a,a8752a,a8755a,a8756a,a8759a,a8762a,a8763a,a8766a,a8769a,a8770a,a8773a,a8776a,a8777a,a8780a,a8783a,a8784a,a8787a,a8790a,a8791a,a8794a,a8797a,a8798a,a8801a,a8804a,a8805a,a8808a,a8811a,a8812a,a8815a,a8818a,a8819a,a8822a,a8825a,a8826a,a8829a,a8832a,a8833a,a8836a,a8839a,a8840a,a8843a,a8846a,a8847a,a8850a,a8853a,a8854a,a8857a,a8860a,a8861a,a8864a,a8867a,a8868a,a8871a,a8874a,a8875a,a8878a,a8881a,a8882a,a8885a,a8888a,a8889a,a8892a,a8895a,a8896a,a8899a,a8902a,a8903a,a8906a,a8909a,a8910a,a8913a,a8916a,a8917a,a8920a,a8923a,a8924a,a8927a,a8930a,a8931a,a8934a,a8937a,a8938a,a8941a,a8944a,a8945a,a8948a,a8951a,a8952a,a8955a,a8958a,a8959a,a8962a,a8965a,a8966a,a8969a,a8972a,a8973a,a8976a,a8979a,a8980a,a8983a,a8986a,a8987a,a8990a,a8993a,a8994a,a8997a,a9000a,a9001a,a9004a,a9007a,a9008a,a9011a,a9014a,a9015a,a9018a,a9021a,a9022a,a9025a,a9028a,a9029a,a9032a,a9035a,a9036a,a9039a,a9042a,a9043a,a9046a,a9049a,a9050a,a9053a,a9056a,a9057a,a9060a,a9063a,a9064a,a9067a,a9070a,a9071a,a9074a,a9077a,a9078a,a9081a,a9084a,a9085a,a9088a,a9091a,a9092a,a9095a,a9098a,a9099a,a9102a,a9105a,a9106a,a9109a,a9112a,a9113a,a9116a,a9119a,a9120a,a9123a,a9126a,a9127a,a9130a,a9133a,a9134a,a9137a,a9140a,a9141a,a9144a,a9147a,a9148a,a9151a,a9154a,a9155a,a9158a,a9161a,a9162a,a9165a,a9168a,a9169a,a9172a,a9175a,a9176a,a9179a,a9182a,a9183a,a9186a,a9189a,a9190a,a9193a,a9196a,a9197a,a9200a,a9203a,a9204a,a9207a,a9210a,a9211a,a9214a,a9217a,a9218a,a9221a,a9224a,a9225a,a9228a,a9231a,a9232a,a9235a,a9238a,a9239a,a9242a,a9245a,a9246a,a9249a,a9252a,a9253a,a9256a,a9259a,a9260a,a9263a,a9266a,a9267a,a9270a,a9273a,a9274a,a9277a,a9280a,a9281a,a9284a,a9287a,a9288a,a9291a,a9294a,a9295a,a9298a,a9302a,a9303a,a9304a,a9307a,a9310a,a9311a,a9314a,a9318a,a9319a,a9320a,a9323a,a9326a,a9327a,a9330a,a9334a,a9335a,a9336a,a9339a,a9342a,a9343a,a9346a,a9350a,a9351a,a9352a,a9355a,a9358a,a9359a,a9362a,a9366a,a9367a,a9368a,a9371a,a9374a,a9375a,a9378a,a9382a,a9383a,a9384a,a9387a,a9390a,a9391a,a9394a,a9398a,a9399a,a9400a,a9403a,a9406a,a9407a,a9410a,a9414a,a9415a,a9416a,a9419a,a9422a,a9423a,a9426a,a9430a,a9431a,a9432a,a9435a,a9438a,a9439a,a9442a,a9446a,a9447a,a9448a,a9451a,a9454a,a9455a,a9458a,a9462a,a9463a,a9464a,a9467a,a9470a,a9471a,a9474a,a9478a,a9479a,a9480a,a9483a,a9486a,a9487a,a9490a,a9494a,a9495a,a9496a,a9499a,a9502a,a9503a,a9506a,a9510a,a9511a,a9512a,a9515a,a9518a,a9519a,a9522a,a9526a,a9527a,a9528a,a9531a,a9534a,a9535a,a9538a,a9542a,a9543a,a9544a,a9547a,a9550a,a9551a,a9554a,a9558a,a9559a,a9560a,a9563a,a9566a,a9567a,a9570a,a9574a,a9575a,a9576a,a9579a,a9582a,a9583a,a9586a,a9590a,a9591a,a9592a,a9595a,a9598a,a9599a,a9602a,a9606a,a9607a,a9608a,a9611a,a9614a,a9615a,a9618a,a9622a,a9623a,a9624a,a9627a,a9630a,a9631a,a9634a,a9638a,a9639a,a9640a,a9643a,a9646a,a9647a,a9650a,a9654a,a9655a,a9656a,a9659a,a9662a,a9663a,a9666a,a9670a,a9671a,a9672a,a9675a,a9678a,a9679a,a9682a,a9686a,a9687a,a9688a,a9691a,a9694a,a9695a,a9698a,a9702a,a9703a,a9704a,a9707a,a9710a,a9711a,a9714a,a9718a,a9719a,a9720a,a9723a,a9726a,a9727a,a9730a,a9734a,a9735a,a9736a,a9739a,a9742a,a9743a,a9746a,a9750a,a9751a,a9752a,a9755a,a9758a,a9759a,a9762a,a9766a,a9767a,a9768a,a9771a,a9774a,a9775a,a9778a,a9782a,a9783a,a9784a,a9787a,a9790a,a9791a,a9794a,a9798a,a9799a,a9800a,a9803a,a9806a,a9807a,a9810a,a9814a,a9815a,a9816a,a9819a,a9822a,a9823a,a9826a,a9830a,a9831a,a9832a,a9835a,a9838a,a9839a,a9842a,a9846a,a9847a,a9848a,a9851a,a9854a,a9855a,a9858a,a9862a,a9863a,a9864a,a9867a,a9870a,a9871a,a9874a,a9878a,a9879a,a9880a,a9883a,a9886a,a9887a,a9890a,a9894a,a9895a,a9896a,a9899a,a9902a,a9903a,a9906a,a9910a,a9911a,a9912a,a9915a,a9918a,a9919a,a9922a,a9926a,a9927a,a9928a,a9931a,a9934a,a9935a,a9938a,a9942a,a9943a,a9944a,a9947a,a9950a,a9951a,a9954a,a9958a,a9959a,a9960a,a9963a,a9966a,a9967a,a9970a,a9974a,a9975a,a9976a,a9979a,a9982a,a9983a,a9986a,a9990a,a9991a,a9992a,a9995a,a9998a,a9999a,a10002a,a10006a,a10007a,a10008a,a10011a,a10014a,a10015a,a10018a,a10022a,a10023a,a10024a,a10027a,a10030a,a10031a,a10034a,a10038a,a10039a,a10040a,a10043a,a10046a,a10047a,a10050a,a10054a,a10055a,a10056a,a10059a,a10062a,a10063a,a10066a,a10070a,a10071a,a10072a,a10075a,a10078a,a10079a,a10082a,a10086a,a10087a,a10088a,a10091a,a10094a,a10095a,a10098a,a10102a,a10103a,a10104a,a10107a,a10110a,a10111a,a10114a,a10118a,a10119a,a10120a,a10123a,a10126a,a10127a,a10130a,a10134a,a10135a,a10136a,a10139a,a10142a,a10143a,a10146a,a10150a,a10151a,a10152a,a10155a,a10158a,a10159a,a10162a,a10166a,a10167a,a10168a,a10171a,a10174a,a10175a,a10178a,a10182a,a10183a,a10184a,a10187a,a10190a,a10191a,a10194a,a10198a,a10199a,a10200a,a10203a,a10206a,a10207a,a10210a,a10214a,a10215a,a10216a,a10219a,a10222a,a10223a,a10226a,a10230a,a10231a,a10232a,a10235a,a10238a,a10239a,a10242a,a10246a,a10247a,a10248a,a10251a,a10254a,a10255a,a10258a,a10262a,a10263a,a10264a,a10267a,a10270a,a10271a,a10274a,a10278a,a10279a,a10280a,a10283a,a10286a,a10287a,a10290a,a10294a,a10295a,a10296a,a10299a,a10302a,a10303a,a10306a,a10310a,a10311a,a10312a,a10315a,a10318a,a10319a,a10322a,a10326a,a10327a,a10328a,a10331a,a10334a,a10335a,a10338a,a10342a,a10343a,a10344a,a10347a,a10350a,a10351a,a10354a,a10358a,a10359a,a10360a,a10363a,a10366a,a10367a,a10370a,a10374a,a10375a,a10376a,a10379a,a10382a,a10383a,a10386a,a10390a,a10391a,a10392a,a10395a,a10398a,a10399a,a10402a,a10406a,a10407a,a10408a,a10411a,a10414a,a10415a,a10418a,a10422a,a10423a,a10424a,a10427a,a10430a,a10431a,a10434a,a10438a,a10439a,a10440a,a10443a,a10446a,a10447a,a10450a,a10454a,a10455a,a10456a,a10459a,a10462a,a10463a,a10466a,a10470a,a10471a,a10472a,a10475a,a10478a,a10479a,a10482a,a10486a,a10487a,a10488a,a10491a,a10494a,a10495a,a10498a,a10502a,a10503a,a10504a,a10507a,a10510a,a10511a,a10514a,a10518a,a10519a,a10520a,a10523a,a10526a,a10527a,a10530a,a10534a,a10535a,a10536a,a10539a,a10542a,a10543a,a10546a,a10550a,a10551a,a10552a,a10555a,a10558a,a10559a,a10562a,a10566a,a10567a,a10568a,a10571a,a10574a,a10575a,a10578a,a10582a,a10583a,a10584a,a10587a,a10590a,a10591a,a10594a,a10598a,a10599a,a10600a,a10603a,a10606a,a10607a,a10610a,a10614a,a10615a,a10616a,a10619a,a10622a,a10623a,a10626a,a10630a,a10631a,a10632a,a10635a,a10638a,a10639a,a10642a,a10646a,a10647a,a10648a,a10651a,a10654a,a10655a,a10658a,a10662a,a10663a,a10664a,a10667a,a10670a,a10671a,a10674a,a10678a,a10679a,a10680a,a10683a,a10686a,a10687a,a10690a,a10694a,a10695a,a10696a,a10699a,a10702a,a10703a,a10706a,a10710a,a10711a,a10712a,a10715a,a10718a,a10719a,a10722a,a10726a,a10727a,a10728a,a10731a,a10734a,a10735a,a10738a,a10742a,a10743a,a10744a,a10747a,a10750a,a10751a,a10754a,a10758a,a10759a,a10760a,a10763a,a10766a,a10767a,a10770a,a10774a,a10775a,a10776a,a10779a,a10782a,a10783a,a10786a,a10790a,a10791a,a10792a,a10795a,a10798a,a10799a,a10802a,a10806a,a10807a,a10808a,a10811a,a10814a,a10815a,a10818a,a10822a,a10823a,a10824a,a10827a,a10830a,a10831a,a10834a,a10838a,a10839a,a10840a,a10843a,a10846a,a10847a,a10850a,a10854a,a10855a,a10856a,a10859a,a10862a,a10863a,a10866a,a10870a,a10871a,a10872a,a10875a,a10878a,a10879a,a10882a,a10886a,a10887a,a10888a,a10891a,a10894a,a10895a,a10898a,a10902a,a10903a,a10904a,a10907a,a10910a,a10911a,a10914a,a10918a,a10919a,a10920a,a10923a,a10926a,a10927a,a10930a,a10934a,a10935a,a10936a,a10939a,a10942a,a10943a,a10946a,a10950a,a10951a,a10952a,a10955a,a10958a,a10959a,a10962a,a10966a,a10967a,a10968a,a10971a,a10974a,a10975a,a10978a,a10982a,a10983a,a10984a,a10987a,a10990a,a10991a,a10994a,a10998a,a10999a,a11000a,a11003a,a11006a,a11007a,a11010a,a11014a,a11015a,a11016a,a11019a,a11022a,a11023a,a11026a,a11030a,a11031a,a11032a,a11035a,a11038a,a11039a,a11042a,a11046a,a11047a,a11048a,a11051a,a11054a,a11055a,a11058a,a11062a,a11063a,a11064a,a11067a,a11070a,a11071a,a11074a,a11078a,a11079a,a11080a,a11083a,a11086a,a11087a,a11090a,a11094a,a11095a,a11096a,a11099a,a11102a,a11103a,a11106a,a11110a,a11111a,a11112a,a11115a,a11118a,a11119a,a11122a,a11126a,a11127a,a11128a,a11131a,a11134a,a11135a,a11138a,a11142a,a11143a,a11144a,a11147a,a11150a,a11151a,a11154a,a11158a,a11159a,a11160a,a11163a,a11166a,a11167a,a11170a,a11174a,a11175a,a11176a,a11179a,a11182a,a11183a,a11186a,a11190a,a11191a,a11192a,a11195a,a11198a,a11199a,a11202a,a11206a,a11207a,a11208a,a11211a,a11214a,a11215a,a11218a,a11222a,a11223a,a11224a,a11227a,a11230a,a11231a,a11234a,a11238a,a11239a,a11240a,a11243a,a11246a,a11247a,a11250a,a11254a,a11255a,a11256a,a11259a,a11262a,a11263a,a11266a,a11270a,a11271a,a11272a,a11275a,a11278a,a11279a,a11282a,a11286a,a11287a,a11288a,a11291a,a11294a,a11295a,a11298a,a11302a,a11303a,a11304a,a11307a,a11310a,a11311a,a11314a,a11318a,a11319a,a11320a,a11323a,a11326a,a11327a,a11330a,a11334a,a11335a,a11336a,a11339a,a11342a,a11343a,a11346a,a11350a,a11351a,a11352a,a11355a,a11358a,a11359a,a11362a,a11366a,a11367a,a11368a,a11371a,a11374a,a11375a,a11378a,a11382a,a11383a,a11384a,a11387a,a11390a,a11391a,a11394a,a11398a,a11399a,a11400a,a11403a,a11406a,a11407a,a11410a,a11414a,a11415a,a11416a,a11419a,a11422a,a11423a,a11426a,a11430a,a11431a,a11432a,a11435a,a11438a,a11439a,a11442a,a11446a,a11447a,a11448a,a11451a,a11454a,a11455a,a11458a,a11462a,a11463a,a11464a,a11467a,a11470a,a11471a,a11474a,a11478a,a11479a,a11480a,a11483a,a11486a,a11487a,a11490a,a11494a,a11495a,a11496a,a11499a,a11502a,a11503a,a11506a,a11510a,a11511a,a11512a,a11515a,a11518a,a11519a,a11522a,a11526a,a11527a,a11528a,a11531a,a11534a,a11535a,a11538a,a11542a,a11543a,a11544a,a11547a,a11550a,a11551a,a11554a,a11558a,a11559a,a11560a,a11563a,a11566a,a11567a,a11570a,a11574a,a11575a,a11576a,a11579a,a11582a,a11583a,a11586a,a11590a,a11591a,a11592a,a11595a,a11598a,a11599a,a11602a,a11606a,a11607a,a11608a,a11611a,a11614a,a11615a,a11618a,a11622a,a11623a,a11624a,a11627a,a11630a,a11631a,a11634a,a11638a,a11639a,a11640a,a11643a,a11646a,a11647a,a11650a,a11654a,a11655a,a11656a,a11659a,a11662a,a11663a,a11666a,a11670a,a11671a,a11672a,a11675a,a11678a,a11679a,a11682a,a11686a,a11687a,a11688a,a11691a,a11694a,a11695a,a11698a,a11702a,a11703a,a11704a,a11707a,a11710a,a11711a,a11714a,a11718a,a11719a,a11720a,a11723a,a11726a,a11727a,a11730a,a11734a,a11735a,a11736a,a11739a,a11742a,a11743a,a11746a,a11750a,a11751a,a11752a,a11755a,a11758a,a11759a,a11762a,a11766a,a11767a,a11768a,a11771a,a11774a,a11775a,a11778a,a11782a,a11783a,a11784a,a11787a,a11790a,a11791a,a11794a,a11798a,a11799a,a11800a,a11803a,a11806a,a11807a,a11810a,a11814a,a11815a,a11816a,a11819a,a11822a,a11823a,a11826a,a11830a,a11831a,a11832a,a11835a,a11838a,a11839a,a11842a,a11846a,a11847a,a11848a,a11851a,a11854a,a11855a,a11858a,a11862a,a11863a,a11864a,a11867a,a11870a,a11871a,a11874a,a11878a,a11879a,a11880a,a11883a,a11886a,a11887a,a11890a,a11894a,a11895a,a11896a,a11899a,a11902a,a11903a,a11906a,a11910a,a11911a,a11912a,a11915a,a11918a,a11919a,a11922a,a11926a,a11927a,a11928a,a11931a,a11934a,a11935a,a11938a,a11942a,a11943a,a11944a,a11947a,a11950a,a11951a,a11954a,a11958a,a11959a,a11960a,a11963a,a11966a,a11967a,a11970a,a11974a,a11975a,a11976a,a11979a,a11982a,a11983a,a11986a,a11990a,a11991a,a11992a,a11995a,a11998a,a11999a,a12002a,a12006a,a12007a,a12008a,a12011a,a12014a,a12015a,a12018a,a12022a,a12023a,a12024a,a12027a,a12030a,a12031a,a12034a,a12038a,a12039a,a12040a,a12043a,a12046a,a12047a,a12050a,a12054a,a12055a,a12056a,a12059a,a12062a,a12063a,a12066a,a12070a,a12071a,a12072a,a12075a,a12078a,a12079a,a12082a,a12086a,a12087a,a12088a,a12091a,a12094a,a12095a,a12098a,a12102a,a12103a,a12104a,a12107a,a12110a,a12111a,a12114a,a12118a,a12119a,a12120a,a12123a,a12126a,a12127a,a12130a,a12134a,a12135a,a12136a,a12139a,a12142a,a12143a,a12146a,a12150a,a12151a,a12152a,a12155a,a12158a,a12159a,a12162a,a12166a,a12167a,a12168a,a12171a,a12174a,a12175a,a12178a,a12182a,a12183a,a12184a,a12187a,a12190a,a12191a,a12194a,a12198a,a12199a,a12200a,a12203a,a12206a,a12207a,a12210a,a12214a,a12215a,a12216a,a12219a,a12222a,a12223a,a12226a,a12230a,a12231a,a12232a,a12235a,a12238a,a12239a,a12242a,a12246a,a12247a,a12248a,a12251a,a12254a,a12255a,a12258a,a12262a,a12263a,a12264a,a12267a,a12270a,a12271a,a12274a,a12278a,a12279a,a12280a,a12283a,a12286a,a12287a,a12290a,a12294a,a12295a,a12296a,a12299a,a12302a,a12303a,a12306a,a12310a,a12311a,a12312a,a12315a,a12318a,a12319a,a12322a,a12326a,a12327a,a12328a,a12331a,a12334a,a12335a,a12338a,a12342a,a12343a,a12344a,a12347a,a12350a,a12351a,a12354a,a12358a,a12359a,a12360a,a12363a,a12366a,a12367a,a12370a,a12374a,a12375a,a12376a,a12379a,a12382a,a12383a,a12386a,a12390a,a12391a,a12392a,a12395a,a12398a,a12399a,a12402a,a12406a,a12407a,a12408a,a12411a,a12414a,a12415a,a12418a,a12422a,a12423a,a12424a,a12427a,a12430a,a12431a,a12434a,a12438a,a12439a,a12440a,a12443a,a12446a,a12447a,a12450a,a12454a,a12455a,a12456a,a12459a,a12462a,a12463a,a12466a,a12470a,a12471a,a12472a,a12475a,a12478a,a12479a,a12482a,a12486a,a12487a,a12488a,a12491a,a12494a,a12495a,a12498a,a12502a,a12503a,a12504a,a12507a,a12510a,a12511a,a12514a,a12518a,a12519a,a12520a,a12523a,a12526a,a12527a,a12530a,a12534a,a12535a,a12536a,a12539a,a12542a,a12543a,a12546a,a12550a,a12551a,a12552a,a12555a,a12559a,a12560a,a12561a,a12564a,a12568a,a12569a,a12570a,a12573a,a12577a,a12578a,a12579a,a12582a,a12586a,a12587a,a12588a,a12591a,a12595a,a12596a,a12597a,a12600a,a12604a,a12605a,a12606a,a12609a,a12613a,a12614a,a12615a,a12618a,a12622a,a12623a,a12624a,a12627a,a12631a,a12632a,a12633a,a12636a,a12640a,a12641a,a12642a,a12645a,a12649a,a12650a,a12651a,a12654a,a12658a,a12659a,a12660a,a12663a,a12667a,a12668a,a12669a,a12672a,a12676a,a12677a,a12678a,a12681a,a12685a,a12686a,a12687a,a12690a,a12694a,a12695a,a12696a,a12699a,a12703a,a12704a,a12705a,a12708a,a12712a,a12713a,a12714a,a12717a,a12721a,a12722a,a12723a,a12726a,a12730a,a12731a,a12732a,a12735a,a12739a,a12740a,a12741a,a12744a,a12748a,a12749a,a12750a,a12753a,a12757a,a12758a,a12759a,a12762a,a12766a,a12767a,a12768a,a12771a,a12775a,a12776a,a12777a,a12780a,a12784a,a12785a,a12786a,a12789a,a12793a,a12794a,a12795a,a12798a,a12802a,a12803a,a12804a,a12807a,a12811a,a12812a,a12813a,a12816a,a12820a,a12821a,a12822a,a12825a,a12829a,a12830a,a12831a,a12834a,a12838a,a12839a,a12840a,a12843a,a12847a,a12848a,a12849a,a12852a,a12856a,a12857a,a12858a,a12861a,a12865a,a12866a,a12867a,a12870a,a12874a,a12875a,a12876a,a12879a,a12883a,a12884a,a12885a,a12888a,a12892a,a12893a,a12894a,a12897a,a12901a,a12902a,a12903a,a12906a,a12910a,a12911a,a12912a,a12915a,a12919a,a12920a,a12921a,a12924a,a12928a,a12929a,a12930a,a12933a,a12937a,a12938a,a12939a,a12942a,a12946a,a12947a,a12948a,a12951a,a12955a,a12956a,a12957a,a12960a,a12964a,a12965a,a12966a,a12969a,a12973a,a12974a,a12975a,a12978a,a12982a,a12983a,a12984a,a12987a,a12991a,a12992a,a12993a,a12996a,a13000a,a13001a,a13002a,a13005a,a13009a,a13010a,a13011a,a13014a,a13018a,a13019a,a13020a,a13023a,a13027a,a13028a,a13029a,a13032a,a13036a,a13037a,a13038a,a13041a,a13045a,a13046a,a13047a,a13050a,a13054a,a13055a,a13056a,a13059a,a13063a,a13064a,a13065a,a13068a,a13072a,a13073a,a13074a,a13077a,a13081a,a13082a,a13083a,a13086a,a13090a,a13091a,a13092a,a13095a,a13099a,a13100a,a13101a,a13104a,a13108a,a13109a,a13110a,a13113a,a13117a,a13118a,a13119a,a13122a,a13126a,a13127a,a13128a,a13131a,a13135a,a13136a,a13137a,a13140a,a13144a,a13145a,a13146a,a13149a,a13153a,a13154a,a13155a,a13158a,a13162a,a13163a,a13164a,a13167a,a13171a,a13172a,a13173a,a13176a,a13180a,a13181a,a13182a,a13185a,a13189a,a13190a,a13191a,a13194a,a13198a,a13199a,a13200a,a13203a,a13207a,a13208a,a13209a,a13212a,a13216a,a13217a,a13218a,a13221a,a13225a,a13226a,a13227a,a13230a,a13234a,a13235a,a13236a,a13239a,a13243a,a13244a,a13245a,a13248a,a13252a,a13253a,a13254a,a13257a,a13261a,a13262a,a13263a,a13266a,a13270a,a13271a,a13272a,a13275a,a13279a,a13280a,a13281a,a13284a,a13288a,a13289a,a13290a,a13293a,a13297a,a13298a,a13299a,a13302a,a13306a,a13307a,a13308a,a13311a,a13315a,a13316a,a13317a,a13320a,a13324a,a13325a,a13326a,a13329a,a13333a,a13334a,a13335a,a13338a,a13342a,a13343a,a13344a,a13347a,a13351a,a13352a,a13353a,a13356a,a13360a,a13361a,a13362a,a13365a,a13369a,a13370a,a13371a,a13374a,a13378a,a13379a,a13380a,a13383a,a13387a,a13388a,a13389a,a13392a,a13396a,a13397a,a13398a,a13401a,a13405a,a13406a,a13407a,a13410a,a13414a,a13415a,a13416a,a13419a,a13423a,a13424a,a13425a,a13428a,a13432a,a13433a,a13434a,a13437a,a13441a,a13442a,a13443a,a13446a,a13450a,a13451a,a13452a,a13455a,a13459a,a13460a,a13461a,a13464a,a13468a,a13469a,a13470a,a13473a,a13477a,a13478a,a13479a,a13482a,a13486a,a13487a,a13488a,a13491a,a13495a,a13496a,a13497a,a13500a,a13504a,a13505a,a13506a,a13509a,a13513a,a13514a,a13515a,a13518a,a13522a,a13523a,a13524a,a13527a,a13531a,a13532a,a13533a,a13536a,a13540a,a13541a,a13542a,a13545a,a13549a,a13550a,a13551a,a13554a,a13558a,a13559a,a13560a,a13563a,a13567a,a13568a,a13569a,a13572a,a13576a,a13577a,a13578a,a13581a,a13585a,a13586a,a13587a,a13590a,a13594a,a13595a,a13596a,a13599a,a13603a,a13604a,a13605a,a13608a,a13612a,a13613a,a13614a,a13617a,a13621a,a13622a,a13623a,a13626a,a13630a,a13631a,a13632a,a13635a,a13639a,a13640a,a13641a,a13644a,a13648a,a13649a,a13650a,a13653a,a13657a,a13658a,a13659a,a13662a,a13666a,a13667a,a13668a,a13671a,a13675a,a13676a,a13677a,a13680a,a13684a,a13685a,a13686a,a13689a,a13693a,a13694a,a13695a,a13698a,a13702a,a13703a,a13704a,a13707a,a13711a,a13712a,a13713a,a13716a,a13720a,a13721a,a13722a,a13725a,a13729a,a13730a,a13731a,a13734a,a13738a,a13739a,a13740a,a13743a,a13747a,a13748a,a13749a,a13752a,a13756a,a13757a,a13758a,a13761a,a13765a,a13766a,a13767a,a13770a,a13774a,a13775a,a13776a,a13779a,a13783a,a13784a,a13785a,a13788a,a13792a,a13793a,a13794a,a13797a,a13801a,a13802a,a13803a,a13806a,a13810a,a13811a,a13812a,a13815a,a13819a,a13820a,a13821a,a13824a,a13828a,a13829a,a13830a,a13833a,a13837a,a13838a,a13839a,a13842a,a13846a,a13847a,a13848a,a13851a,a13855a,a13856a,a13857a,a13860a,a13864a,a13865a,a13866a,a13869a,a13873a,a13874a,a13875a,a13878a,a13882a,a13883a,a13884a,a13887a,a13891a,a13892a,a13893a,a13896a,a13900a,a13901a,a13902a,a13905a,a13909a,a13910a,a13911a,a13914a,a13918a,a13919a,a13920a,a13923a,a13927a,a13928a,a13929a,a13932a,a13936a,a13937a,a13938a,a13941a,a13945a,a13946a,a13947a,a13950a,a13954a,a13955a,a13956a,a13959a,a13963a,a13964a,a13965a,a13968a,a13972a,a13973a,a13974a,a13977a,a13981a,a13982a,a13983a,a13986a,a13990a,a13991a,a13992a,a13995a,a13999a,a14000a,a14001a,a14004a,a14008a,a14009a,a14010a,a14013a,a14017a,a14018a,a14019a,a14022a,a14026a,a14027a,a14028a,a14031a,a14035a,a14036a,a14037a,a14040a,a14044a,a14045a,a14046a,a14049a,a14053a,a14054a,a14055a,a14058a,a14062a,a14063a,a14064a,a14067a,a14071a,a14072a,a14073a,a14076a,a14080a,a14081a,a14082a,a14085a,a14089a,a14090a,a14091a,a14094a,a14098a,a14099a,a14100a,a14103a,a14107a,a14108a,a14109a,a14112a,a14116a,a14117a,a14118a,a14121a,a14125a,a14126a,a14127a,a14130a,a14134a,a14135a,a14136a,a14139a,a14143a,a14144a,a14145a,a14148a,a14152a,a14153a,a14154a,a14157a,a14161a,a14162a,a14163a,a14166a,a14170a,a14171a,a14172a,a14175a,a14179a,a14180a,a14181a,a14184a,a14188a,a14189a,a14190a,a14193a,a14197a,a14198a,a14199a,a14202a,a14206a,a14207a,a14208a,a14211a,a14215a,a14216a,a14217a,a14220a,a14224a,a14225a,a14226a,a14229a,a14233a,a14234a,a14235a,a14238a,a14242a,a14243a,a14244a,a14247a,a14251a,a14252a,a14253a,a14256a,a14260a,a14261a,a14262a,a14265a,a14269a,a14270a,a14271a,a14274a,a14278a,a14279a,a14280a,a14283a,a14287a,a14288a,a14289a,a14292a,a14296a,a14297a,a14298a,a14301a,a14305a,a14306a,a14307a,a14310a,a14314a,a14315a,a14316a,a14319a,a14323a,a14324a,a14325a,a14328a,a14332a,a14333a,a14334a,a14337a,a14341a,a14342a,a14343a,a14346a,a14350a,a14351a,a14352a,a14355a,a14359a,a14360a,a14361a,a14364a,a14368a,a14369a,a14370a,a14373a,a14377a,a14378a,a14379a,a14382a,a14386a,a14387a,a14388a,a14391a,a14395a,a14396a,a14397a,a14400a,a14404a,a14405a,a14406a,a14409a,a14413a,a14414a,a14415a,a14418a,a14422a,a14423a,a14424a,a14427a,a14431a,a14432a,a14433a,a14436a,a14440a,a14441a,a14442a,a14445a,a14449a,a14450a,a14451a,a14454a,a14458a,a14459a,a14460a,a14463a,a14467a,a14468a,a14469a,a14472a,a14476a,a14477a,a14478a,a14481a,a14485a,a14486a,a14487a,a14490a,a14494a,a14495a,a14496a,a14499a,a14503a,a14504a,a14505a,a14508a,a14512a,a14513a,a14514a,a14517a,a14521a,a14522a,a14523a,a14526a,a14530a,a14531a,a14532a,a14535a,a14539a,a14540a,a14541a,a14544a,a14548a,a14549a,a14550a,a14553a,a14557a,a14558a,a14559a,a14562a,a14566a,a14567a,a14568a,a14571a,a14575a,a14576a,a14577a,a14580a,a14584a,a14585a,a14586a,a14589a,a14593a,a14594a,a14595a,a14598a,a14602a,a14603a,a14604a,a14607a,a14611a,a14612a,a14613a,a14616a,a14620a,a14621a,a14622a,a14625a,a14629a,a14630a,a14631a,a14634a,a14638a,a14639a,a14640a,a14643a,a14647a,a14648a,a14649a,a14652a,a14656a,a14657a,a14658a,a14661a,a14665a,a14666a,a14667a,a14670a,a14674a,a14675a,a14676a,a14679a,a14683a,a14684a,a14685a,a14688a,a14692a,a14693a,a14694a,a14697a,a14701a,a14702a,a14703a,a14706a,a14710a,a14711a,a14712a,a14715a,a14719a,a14720a,a14721a,a14724a,a14728a,a14729a,a14730a,a14733a,a14737a,a14738a,a14739a,a14742a,a14746a,a14747a,a14748a,a14751a,a14755a,a14756a,a14757a,a14760a,a14764a,a14765a,a14766a,a14769a,a14773a,a14774a,a14775a,a14778a,a14782a,a14783a,a14784a,a14787a,a14791a,a14792a,a14793a,a14796a,a14800a,a14801a,a14802a,a14805a,a14809a,a14810a,a14811a,a14814a,a14818a,a14819a,a14820a,a14823a,a14827a,a14828a,a14829a,a14832a,a14836a,a14837a,a14838a,a14841a,a14845a,a14846a,a14847a,a14850a,a14854a,a14855a,a14856a,a14859a,a14863a,a14864a,a14865a,a14868a,a14872a,a14873a,a14874a,a14877a,a14881a,a14882a,a14883a,a14886a,a14890a,a14891a,a14892a,a14895a,a14899a,a14900a,a14901a,a14904a,a14908a,a14909a,a14910a,a14913a,a14917a,a14918a,a14919a,a14922a,a14926a,a14927a,a14928a,a14931a,a14935a,a14936a,a14937a,a14940a,a14944a,a14945a,a14946a,a14949a,a14953a,a14954a,a14955a,a14958a,a14962a,a14963a,a14964a,a14967a,a14971a,a14972a,a14973a,a14976a,a14980a,a14981a,a14982a,a14985a,a14989a,a14990a,a14991a,a14994a,a14998a,a14999a,a15000a,a15003a,a15007a,a15008a,a15009a,a15012a,a15016a,a15017a,a15018a,a15021a,a15025a,a15026a,a15027a,a15030a,a15034a,a15035a,a15036a,a15039a,a15043a,a15044a,a15045a,a15048a,a15052a,a15053a,a15054a,a15057a,a15061a,a15062a,a15063a,a15066a,a15070a,a15071a,a15072a,a15075a,a15079a,a15080a,a15081a,a15084a,a15088a,a15089a,a15090a,a15093a,a15097a,a15098a,a15099a,a15102a,a15106a,a15107a,a15108a,a15111a,a15115a,a15116a,a15117a,a15120a,a15124a,a15125a,a15126a,a15129a,a15133a,a15134a,a15135a,a15138a,a15142a,a15143a,a15144a,a15147a,a15151a,a15152a,a15153a,a15156a,a15160a,a15161a,a15162a,a15165a,a15169a,a15170a,a15171a,a15174a,a15178a,a15179a,a15180a,a15183a,a15187a,a15188a,a15189a,a15192a,a15196a,a15197a,a15198a,a15201a,a15205a,a15206a,a15207a,a15210a,a15214a,a15215a,a15216a,a15219a,a15223a,a15224a,a15225a,a15228a,a15232a,a15233a,a15234a,a15237a,a15241a,a15242a,a15243a,a15246a,a15250a,a15251a,a15252a,a15255a,a15259a,a15260a,a15261a,a15264a,a15268a,a15269a,a15270a,a15273a,a15277a,a15278a,a15279a,a15282a,a15286a,a15287a,a15288a,a15291a,a15295a,a15296a,a15297a,a15300a,a15304a,a15305a,a15306a,a15309a,a15313a,a15314a,a15315a,a15318a,a15322a,a15323a,a15324a,a15327a,a15331a,a15332a,a15333a,a15336a,a15340a,a15341a,a15342a,a15345a,a15349a,a15350a,a15351a,a15354a,a15358a,a15359a,a15360a,a15363a,a15367a,a15368a,a15369a,a15372a,a15376a,a15377a,a15378a,a15381a,a15385a,a15386a,a15387a,a15390a,a15394a,a15395a,a15396a,a15399a,a15403a,a15404a,a15405a,a15408a,a15412a,a15413a,a15414a,a15417a,a15421a,a15422a,a15423a,a15426a,a15430a,a15431a,a15432a,a15435a,a15439a,a15440a,a15441a,a15444a,a15448a,a15449a,a15450a,a15453a,a15457a,a15458a,a15459a,a15462a,a15466a,a15467a,a15468a,a15471a,a15475a,a15476a,a15477a,a15480a,a15484a,a15485a,a15486a,a15489a,a15493a,a15494a,a15495a,a15498a,a15502a,a15503a,a15504a,a15507a,a15511a,a15512a,a15513a,a15516a,a15520a,a15521a,a15522a,a15525a,a15529a,a15530a,a15531a,a15534a,a15538a,a15539a,a15540a,a15543a,a15547a,a15548a,a15549a,a15552a,a15556a,a15557a,a15558a,a15561a,a15565a,a15566a,a15567a,a15570a,a15574a,a15575a,a15576a,a15579a,a15583a,a15584a,a15585a,a15588a,a15592a,a15593a,a15594a,a15597a,a15601a,a15602a,a15603a,a15606a,a15610a,a15611a,a15612a,a15615a,a15619a,a15620a,a15621a,a15624a,a15628a,a15629a,a15630a,a15633a,a15637a,a15638a,a15639a,a15642a,a15646a,a15647a,a15648a,a15651a,a15655a,a15656a,a15657a,a15660a,a15664a,a15665a,a15666a,a15669a,a15673a,a15674a,a15675a,a15678a,a15682a,a15683a,a15684a,a15687a,a15691a,a15692a,a15693a,a15696a,a15700a,a15701a,a15702a,a15705a,a15709a,a15710a,a15711a,a15714a,a15718a,a15719a,a15720a,a15723a,a15727a,a15728a,a15729a,a15732a,a15736a,a15737a,a15738a,a15741a,a15745a,a15746a,a15747a,a15750a,a15754a,a15755a,a15756a,a15759a,a15763a,a15764a,a15765a,a15768a,a15772a,a15773a,a15774a,a15777a,a15781a,a15782a,a15783a,a15786a,a15790a,a15791a,a15792a,a15795a,a15799a,a15800a,a15801a,a15804a,a15808a,a15809a,a15810a,a15813a,a15817a,a15818a,a15819a,a15822a,a15826a,a15827a,a15828a,a15831a,a15835a,a15836a,a15837a,a15840a,a15844a,a15845a,a15846a,a15849a,a15853a,a15854a,a15855a,a15858a,a15862a,a15863a,a15864a,a15867a,a15871a,a15872a,a15873a,a15876a,a15880a,a15881a,a15882a,a15885a,a15889a,a15890a,a15891a,a15894a,a15898a,a15899a,a15900a,a15903a,a15907a,a15908a,a15909a,a15912a,a15916a,a15917a,a15918a,a15921a,a15925a,a15926a,a15927a,a15930a,a15934a,a15935a,a15936a,a15939a,a15943a,a15944a,a15945a,a15948a,a15952a,a15953a,a15954a,a15957a,a15961a,a15962a,a15963a,a15966a,a15970a,a15971a,a15972a,a15975a,a15979a,a15980a,a15981a,a15984a,a15988a,a15989a,a15990a,a15993a,a15997a,a15998a,a15999a,a16002a,a16006a,a16007a,a16008a,a16011a,a16015a,a16016a,a16017a,a16020a,a16024a,a16025a,a16026a,a16029a,a16033a,a16034a,a16035a,a16038a,a16042a,a16043a,a16044a,a16047a,a16051a,a16052a,a16053a,a16056a,a16060a,a16061a,a16062a,a16065a,a16069a,a16070a,a16071a,a16074a,a16078a,a16079a,a16080a,a16083a,a16087a,a16088a,a16089a,a16092a,a16096a,a16097a,a16098a,a16101a,a16105a,a16106a,a16107a,a16110a,a16114a,a16115a,a16116a,a16119a,a16123a,a16124a,a16125a,a16128a,a16132a,a16133a,a16134a,a16137a,a16141a,a16142a,a16143a,a16146a,a16150a,a16151a,a16152a,a16155a,a16159a,a16160a,a16161a,a16164a,a16168a,a16169a,a16170a,a16173a,a16177a,a16178a,a16179a,a16182a,a16186a,a16187a,a16188a,a16191a,a16195a,a16196a,a16197a,a16200a,a16204a,a16205a,a16206a,a16209a,a16213a,a16214a,a16215a,a16218a,a16222a,a16223a,a16224a,a16227a,a16231a,a16232a,a16233a,a16236a,a16240a,a16241a,a16242a,a16245a,a16249a,a16250a,a16251a,a16254a,a16258a,a16259a,a16260a,a16263a,a16267a,a16268a,a16269a,a16272a,a16276a,a16277a,a16278a,a16281a,a16285a,a16286a,a16287a,a16290a,a16294a,a16295a,a16296a,a16299a,a16303a,a16304a,a16305a,a16308a,a16312a,a16313a,a16314a,a16317a,a16321a,a16322a,a16323a,a16326a,a16330a,a16331a,a16332a,a16335a,a16339a,a16340a,a16341a,a16344a,a16348a,a16349a,a16350a,a16353a,a16357a,a16358a,a16359a,a16362a,a16366a,a16367a,a16368a,a16371a,a16375a,a16376a,a16377a,a16380a,a16384a,a16385a,a16386a,a16389a,a16393a,a16394a,a16395a,a16398a,a16402a,a16403a,a16404a,a16407a,a16411a,a16412a,a16413a,a16416a,a16420a,a16421a,a16422a,a16425a,a16429a,a16430a,a16431a,a16434a,a16438a,a16439a,a16440a,a16443a,a16447a,a16448a,a16449a,a16452a,a16456a,a16457a,a16458a,a16461a,a16465a,a16466a,a16467a,a16470a,a16474a,a16475a,a16476a,a16479a,a16483a,a16484a,a16485a,a16488a,a16492a,a16493a,a16494a,a16497a,a16501a,a16502a,a16503a,a16506a,a16510a,a16511a,a16512a,a16515a,a16519a,a16520a,a16521a,a16524a,a16528a,a16529a,a16530a,a16533a,a16537a,a16538a,a16539a,a16542a,a16546a,a16547a,a16548a,a16551a,a16555a,a16556a,a16557a,a16560a,a16564a,a16565a,a16566a,a16569a,a16573a,a16574a,a16575a,a16578a,a16582a,a16583a,a16584a,a16587a,a16591a,a16592a,a16593a,a16596a,a16600a,a16601a,a16602a,a16605a,a16609a,a16610a,a16611a,a16614a,a16618a,a16619a,a16620a,a16623a,a16627a,a16628a,a16629a,a16632a,a16636a,a16637a,a16638a,a16641a,a16645a,a16646a,a16647a,a16650a,a16654a,a16655a,a16656a,a16659a,a16663a,a16664a,a16665a,a16668a,a16672a,a16673a,a16674a,a16677a,a16681a,a16682a,a16683a,a16686a,a16690a,a16691a,a16692a,a16695a,a16699a,a16700a,a16701a,a16704a,a16708a,a16709a,a16710a,a16713a,a16717a,a16718a,a16719a,a16722a,a16726a,a16727a,a16728a,a16731a,a16735a,a16736a,a16737a,a16740a,a16744a,a16745a,a16746a,a16749a,a16753a,a16754a,a16755a,a16758a,a16762a,a16763a,a16764a,a16767a,a16771a,a16772a,a16773a,a16776a,a16780a,a16781a,a16782a,a16785a,a16789a,a16790a,a16791a,a16794a,a16798a,a16799a,a16800a,a16803a,a16807a,a16808a,a16809a,a16812a,a16816a,a16817a,a16818a,a16821a,a16825a,a16826a,a16827a,a16830a,a16834a,a16835a,a16836a,a16839a,a16843a,a16844a,a16845a,a16848a,a16852a,a16853a,a16854a,a16857a,a16861a,a16862a,a16863a,a16866a,a16870a,a16871a,a16872a,a16875a,a16879a,a16880a,a16881a,a16884a,a16888a,a16889a,a16890a,a16893a,a16897a,a16898a,a16899a,a16902a,a16906a,a16907a,a16908a,a16911a,a16915a,a16916a,a16917a,a16920a,a16924a,a16925a,a16926a,a16929a,a16933a,a16934a,a16935a,a16938a,a16942a,a16943a,a16944a,a16947a,a16951a,a16952a,a16953a,a16956a,a16960a,a16961a,a16962a,a16965a,a16969a,a16970a,a16971a,a16974a,a16978a,a16979a,a16980a,a16983a,a16987a,a16988a,a16989a,a16992a,a16996a,a16997a,a16998a,a17001a,a17005a,a17006a,a17007a,a17010a,a17014a,a17015a,a17016a,a17019a,a17023a,a17024a,a17025a,a17028a,a17032a,a17033a,a17034a,a17037a,a17041a,a17042a,a17043a,a17046a,a17050a,a17051a,a17052a,a17055a,a17059a,a17060a,a17061a,a17064a,a17068a,a17069a,a17070a,a17073a,a17077a,a17078a,a17079a,a17082a,a17086a,a17087a,a17088a,a17091a,a17095a,a17096a,a17097a,a17100a,a17104a,a17105a,a17106a,a17109a,a17113a,a17114a,a17115a,a17118a,a17122a,a17123a,a17124a,a17127a,a17131a,a17132a,a17133a,a17136a,a17140a,a17141a,a17142a,a17145a,a17149a,a17150a,a17151a,a17154a,a17158a,a17159a,a17160a,a17163a,a17167a,a17168a,a17169a,a17172a,a17176a,a17177a,a17178a,a17181a,a17185a,a17186a,a17187a,a17190a,a17194a,a17195a,a17196a,a17199a,a17203a,a17204a,a17205a,a17208a,a17212a,a17213a,a17214a,a17217a,a17221a,a17222a,a17223a,a17226a,a17230a,a17231a,a17232a,a17235a,a17239a,a17240a,a17241a,a17244a,a17248a,a17249a,a17250a,a17253a,a17257a,a17258a,a17259a,a17262a,a17266a,a17267a,a17268a,a17271a,a17275a,a17276a,a17277a,a17280a,a17284a,a17285a,a17286a,a17289a,a17293a,a17294a,a17295a,a17298a,a17302a,a17303a,a17304a,a17307a,a17311a,a17312a,a17313a,a17316a,a17320a,a17321a,a17322a,a17325a,a17329a,a17330a,a17331a,a17334a,a17338a,a17339a,a17340a,a17343a,a17347a,a17348a,a17349a,a17352a,a17356a,a17357a,a17358a,a17361a,a17365a,a17366a,a17367a,a17370a,a17374a,a17375a,a17376a,a17379a,a17383a,a17384a,a17385a,a17388a,a17392a,a17393a,a17394a,a17397a,a17401a,a17402a,a17403a,a17406a,a17410a,a17411a,a17412a,a17415a,a17419a,a17420a,a17421a,a17424a,a17428a,a17429a,a17430a,a17433a,a17437a,a17438a,a17439a,a17442a,a17446a,a17447a,a17448a,a17451a,a17455a,a17456a,a17457a,a17460a,a17464a,a17465a,a17466a,a17469a,a17473a,a17474a,a17475a,a17478a,a17482a,a17483a,a17484a,a17487a,a17491a,a17492a,a17493a,a17496a,a17500a,a17501a,a17502a,a17505a,a17509a,a17510a,a17511a,a17514a,a17518a,a17519a,a17520a,a17523a,a17527a,a17528a,a17529a,a17532a,a17536a,a17537a,a17538a,a17541a,a17545a,a17546a,a17547a,a17550a,a17554a,a17555a,a17556a,a17559a,a17563a,a17564a,a17565a,a17568a,a17572a,a17573a,a17574a,a17577a,a17581a,a17582a,a17583a,a17586a,a17590a,a17591a,a17592a,a17595a,a17599a,a17600a,a17601a,a17604a,a17608a,a17609a,a17610a,a17613a,a17617a,a17618a,a17619a,a17622a,a17626a,a17627a,a17628a,a17631a,a17635a,a17636a,a17637a,a17640a,a17644a,a17645a,a17646a,a17649a,a17653a,a17654a,a17655a,a17658a,a17662a,a17663a,a17664a,a17667a,a17671a,a17672a,a17673a,a17676a,a17680a,a17681a,a17682a,a17685a,a17689a,a17690a,a17691a,a17694a,a17698a,a17699a,a17700a,a17703a,a17707a,a17708a,a17709a,a17712a,a17716a,a17717a,a17718a,a17721a,a17725a,a17726a,a17727a,a17730a,a17734a,a17735a,a17736a,a17739a,a17743a,a17744a,a17745a,a17748a,a17752a,a17753a,a17754a,a17757a,a17761a,a17762a,a17763a,a17766a,a17770a,a17771a,a17772a,a17775a,a17779a,a17780a,a17781a,a17784a,a17788a,a17789a,a17790a,a17793a,a17797a,a17798a,a17799a,a17802a,a17806a,a17807a,a17808a,a17811a,a17815a,a17816a,a17817a,a17820a,a17824a,a17825a,a17826a,a17829a,a17833a,a17834a,a17835a,a17838a,a17842a,a17843a,a17844a,a17847a,a17851a,a17852a,a17853a,a17856a,a17860a,a17861a,a17862a,a17865a,a17869a,a17870a,a17871a,a17874a,a17878a,a17879a,a17880a,a17883a,a17887a,a17888a,a17889a,a17892a,a17896a,a17897a,a17898a,a17901a,a17905a,a17906a,a17907a,a17910a,a17914a,a17915a,a17916a,a17919a,a17923a,a17924a,a17925a,a17928a,a17932a,a17933a,a17934a,a17937a,a17941a,a17942a,a17943a,a17946a,a17950a,a17951a,a17952a,a17955a,a17959a,a17960a,a17961a,a17964a,a17968a,a17969a,a17970a,a17973a,a17977a,a17978a,a17979a,a17982a,a17986a,a17987a,a17988a,a17991a,a17995a,a17996a,a17997a,a18000a,a18004a,a18005a,a18006a,a18009a,a18013a,a18014a,a18015a,a18018a,a18022a,a18023a,a18024a,a18027a,a18031a,a18032a,a18033a,a18036a,a18040a,a18041a,a18042a,a18045a,a18049a,a18050a,a18051a,a18054a,a18058a,a18059a,a18060a,a18063a,a18067a,a18068a,a18069a,a18073a,a18074a,a18078a,a18079a,a18080a,a18083a,a18087a,a18088a,a18089a,a18093a,a18094a,a18098a,a18099a,a18100a,a18103a,a18107a,a18108a,a18109a,a18113a,a18114a,a18118a,a18119a,a18120a,a18123a,a18127a,a18128a,a18129a,a18133a,a18134a,a18138a,a18139a,a18140a,a18143a,a18147a,a18148a,a18149a,a18153a,a18154a,a18158a,a18159a,a18160a,a18163a,a18167a,a18168a,a18169a,a18173a,a18174a,a18178a,a18179a,a18180a,a18183a,a18187a,a18188a,a18189a,a18193a,a18194a,a18198a,a18199a,a18200a,a18203a,a18207a,a18208a,a18209a,a18213a,a18214a,a18218a,a18219a,a18220a,a18223a,a18227a,a18228a,a18229a,a18233a,a18234a,a18238a,a18239a,a18240a,a18243a,a18247a,a18248a,a18249a,a18253a,a18254a,a18258a,a18259a,a18260a,a18263a,a18267a,a18268a,a18269a,a18273a,a18274a,a18278a,a18279a,a18280a,a18283a,a18287a,a18288a,a18289a,a18293a,a18294a,a18298a,a18299a,a18300a,a18303a,a18307a,a18308a,a18309a,a18313a,a18314a,a18318a,a18319a,a18320a,a18323a,a18327a,a18328a,a18329a,a18333a,a18334a,a18338a,a18339a,a18340a,a18343a,a18347a,a18348a,a18349a,a18353a,a18354a,a18358a,a18359a,a18360a,a18363a,a18367a,a18368a,a18369a,a18373a,a18374a,a18378a,a18379a,a18380a,a18383a,a18387a,a18388a,a18389a,a18393a,a18394a,a18398a,a18399a,a18400a,a18403a,a18407a,a18408a,a18409a,a18413a,a18414a,a18418a,a18419a,a18420a,a18423a,a18427a,a18428a,a18429a,a18433a,a18434a,a18438a,a18439a,a18440a,a18443a,a18447a,a18448a,a18449a,a18453a,a18454a,a18458a,a18459a,a18460a,a18463a,a18467a,a18468a,a18469a,a18473a,a18474a,a18478a,a18479a,a18480a,a18483a,a18487a,a18488a,a18489a,a18493a,a18494a,a18498a,a18499a,a18500a,a18503a,a18507a,a18508a,a18509a,a18513a,a18514a,a18518a,a18519a,a18520a,a18523a,a18527a,a18528a,a18529a,a18533a,a18534a,a18538a,a18539a,a18540a,a18543a,a18547a,a18548a,a18549a,a18553a,a18554a,a18558a,a18559a,a18560a,a18563a,a18567a,a18568a,a18569a,a18573a,a18574a,a18578a,a18579a,a18580a,a18583a,a18587a,a18588a,a18589a,a18593a,a18594a,a18598a,a18599a,a18600a,a18603a,a18607a,a18608a,a18609a,a18613a,a18614a,a18618a,a18619a,a18620a,a18623a,a18627a,a18628a,a18629a,a18633a,a18634a,a18638a,a18639a,a18640a,a18643a,a18647a,a18648a,a18649a,a18653a,a18654a,a18658a,a18659a,a18660a,a18663a,a18667a,a18668a,a18669a,a18673a,a18674a,a18678a,a18679a,a18680a,a18683a,a18687a,a18688a,a18689a,a18693a,a18694a,a18698a,a18699a,a18700a,a18703a,a18707a,a18708a,a18709a,a18713a,a18714a,a18718a,a18719a,a18720a,a18723a,a18727a,a18728a,a18729a,a18733a,a18734a,a18738a,a18739a,a18740a,a18743a,a18747a,a18748a,a18749a,a18753a,a18754a,a18758a,a18759a,a18760a,a18763a,a18767a,a18768a,a18769a,a18773a,a18774a,a18778a,a18779a,a18780a,a18783a,a18787a,a18788a,a18789a,a18793a,a18794a,a18798a,a18799a,a18800a,a18803a,a18807a,a18808a,a18809a,a18813a,a18814a,a18818a,a18819a,a18820a,a18823a,a18827a,a18828a,a18829a,a18833a,a18834a,a18838a,a18839a,a18840a,a18843a,a18847a,a18848a,a18849a,a18853a,a18854a,a18858a,a18859a,a18860a,a18863a,a18867a,a18868a,a18869a,a18873a,a18874a,a18878a,a18879a,a18880a,a18883a,a18887a,a18888a,a18889a,a18893a,a18894a,a18898a,a18899a,a18900a,a18903a,a18907a,a18908a,a18909a,a18913a,a18914a,a18918a,a18919a,a18920a,a18923a,a18927a,a18928a,a18929a,a18933a,a18934a,a18938a,a18939a,a18940a,a18943a,a18947a,a18948a,a18949a,a18953a,a18954a,a18958a,a18959a,a18960a,a18963a,a18967a,a18968a,a18969a,a18973a,a18974a,a18978a,a18979a,a18980a,a18983a,a18987a,a18988a,a18989a,a18993a,a18994a,a18998a,a18999a,a19000a,a19003a,a19007a,a19008a,a19009a,a19013a,a19014a,a19018a,a19019a,a19020a,a19023a,a19027a,a19028a,a19029a,a19033a,a19034a,a19038a,a19039a,a19040a,a19043a,a19047a,a19048a,a19049a,a19053a,a19054a,a19058a,a19059a,a19060a,a19063a,a19067a,a19068a,a19069a,a19073a,a19074a,a19078a,a19079a,a19080a,a19083a,a19087a,a19088a,a19089a,a19093a,a19094a,a19098a,a19099a,a19100a,a19103a,a19107a,a19108a,a19109a,a19113a,a19114a,a19118a,a19119a,a19120a,a19123a,a19127a,a19128a,a19129a,a19133a,a19134a,a19138a,a19139a,a19140a,a19143a,a19147a,a19148a,a19149a,a19153a,a19154a,a19158a,a19159a,a19160a,a19163a,a19167a,a19168a,a19169a,a19173a,a19174a,a19178a,a19179a,a19180a,a19183a,a19187a,a19188a,a19189a,a19193a,a19194a,a19198a,a19199a,a19200a,a19203a,a19207a,a19208a,a19209a,a19213a,a19214a,a19218a,a19219a,a19220a,a19223a,a19227a,a19228a,a19229a,a19233a,a19234a,a19238a,a19239a,a19240a,a19243a,a19247a,a19248a,a19249a,a19253a,a19254a,a19258a,a19259a,a19260a,a19263a,a19267a,a19268a,a19269a,a19273a,a19274a,a19278a,a19279a,a19280a,a19283a,a19287a,a19288a,a19289a,a19293a,a19294a,a19298a,a19299a,a19300a,a19303a,a19307a,a19308a,a19309a,a19313a,a19314a,a19318a,a19319a,a19320a,a19323a,a19327a,a19328a,a19329a,a19333a,a19334a,a19338a,a19339a,a19340a,a19343a,a19347a,a19348a,a19349a,a19353a,a19354a,a19358a,a19359a,a19360a,a19363a,a19367a,a19368a,a19369a,a19373a,a19374a,a19378a,a19379a,a19380a,a19383a,a19387a,a19388a,a19389a,a19393a,a19394a,a19398a,a19399a,a19400a,a19403a,a19407a,a19408a,a19409a,a19413a,a19414a,a19418a,a19419a,a19420a,a19423a,a19427a,a19428a,a19429a,a19433a,a19434a,a19438a,a19439a,a19440a,a19443a,a19447a,a19448a,a19449a,a19453a,a19454a,a19458a,a19459a,a19460a,a19463a,a19467a,a19468a,a19469a,a19473a,a19474a,a19478a,a19479a,a19480a,a19483a,a19487a,a19488a,a19489a,a19493a,a19494a,a19498a,a19499a,a19500a,a19503a,a19507a,a19508a,a19509a,a19513a,a19514a,a19518a,a19519a,a19520a,a19523a,a19527a,a19528a,a19529a,a19533a,a19534a,a19538a,a19539a,a19540a,a19543a,a19547a,a19548a,a19549a,a19553a,a19554a,a19558a,a19559a,a19560a,a19563a,a19567a,a19568a,a19569a,a19573a,a19574a,a19578a,a19579a,a19580a,a19583a,a19587a,a19588a,a19589a,a19593a,a19594a,a19598a,a19599a,a19600a,a19603a,a19607a,a19608a,a19609a,a19613a,a19614a,a19618a,a19619a,a19620a,a19623a,a19627a,a19628a,a19629a,a19633a,a19634a,a19638a,a19639a,a19640a,a19643a,a19647a,a19648a,a19649a,a19653a,a19654a,a19658a,a19659a,a19660a,a19663a,a19667a,a19668a,a19669a,a19673a,a19674a,a19678a,a19679a,a19680a,a19683a,a19687a,a19688a,a19689a,a19693a,a19694a,a19698a,a19699a,a19700a,a19703a,a19707a,a19708a,a19709a,a19713a,a19714a,a19718a,a19719a,a19720a,a19723a,a19727a,a19728a,a19729a,a19733a,a19734a,a19738a,a19739a,a19740a,a19743a,a19747a,a19748a,a19749a,a19753a,a19754a,a19758a,a19759a,a19760a,a19763a,a19767a,a19768a,a19769a,a19773a,a19774a,a19778a,a19779a,a19780a,a19783a,a19787a,a19788a,a19789a,a19793a,a19794a,a19798a,a19799a,a19800a,a19803a,a19807a,a19808a,a19809a,a19813a,a19814a,a19818a,a19819a,a19820a,a19823a,a19827a,a19828a,a19829a,a19833a,a19834a,a19838a,a19839a,a19840a,a19843a,a19847a,a19848a,a19849a,a19853a,a19854a,a19858a,a19859a,a19860a,a19863a,a19867a,a19868a,a19869a,a19873a,a19874a,a19878a,a19879a,a19880a,a19883a,a19887a,a19888a,a19889a,a19893a,a19894a,a19898a,a19899a,a19900a,a19903a,a19907a,a19908a,a19909a,a19913a,a19914a,a19918a,a19919a,a19920a,a19923a,a19927a,a19928a,a19929a,a19933a,a19934a,a19938a,a19939a,a19940a,a19943a,a19947a,a19948a,a19949a,a19953a,a19954a,a19958a,a19959a,a19960a,a19963a,a19967a,a19968a,a19969a,a19973a,a19974a,a19978a,a19979a,a19980a,a19983a,a19987a,a19988a,a19989a,a19993a,a19994a,a19998a,a19999a,a20000a,a20003a,a20007a,a20008a,a20009a,a20013a,a20014a,a20018a,a20019a,a20020a,a20023a,a20027a,a20028a,a20029a,a20033a,a20034a,a20038a,a20039a,a20040a,a20043a,a20047a,a20048a,a20049a,a20053a,a20054a,a20058a,a20059a,a20060a,a20063a,a20067a,a20068a,a20069a,a20073a,a20074a,a20078a,a20079a,a20080a,a20083a,a20087a,a20088a,a20089a,a20093a,a20094a,a20098a,a20099a,a20100a,a20103a,a20107a,a20108a,a20109a,a20113a,a20114a,a20118a,a20119a,a20120a,a20123a,a20127a,a20128a,a20129a,a20133a,a20134a,a20138a,a20139a,a20140a,a20143a,a20147a,a20148a,a20149a,a20153a,a20154a,a20158a,a20159a,a20160a,a20163a,a20167a,a20168a,a20169a,a20173a,a20174a,a20178a,a20179a,a20180a,a20183a,a20187a,a20188a,a20189a,a20193a,a20194a,a20198a,a20199a,a20200a,a20203a,a20207a,a20208a,a20209a,a20213a,a20214a,a20218a,a20219a,a20220a,a20223a,a20227a,a20228a,a20229a,a20233a,a20234a,a20238a,a20239a,a20240a,a20243a,a20247a,a20248a,a20249a,a20253a,a20254a,a20258a,a20259a,a20260a,a20263a,a20267a,a20268a,a20269a,a20273a,a20274a,a20278a,a20279a,a20280a,a20283a,a20287a,a20288a,a20289a,a20293a,a20294a,a20298a,a20299a,a20300a,a20303a,a20307a,a20308a,a20309a,a20313a,a20314a,a20318a,a20319a,a20320a,a20323a,a20327a,a20328a,a20329a,a20333a,a20334a,a20338a,a20339a,a20340a,a20343a,a20347a,a20348a,a20349a,a20353a,a20354a,a20358a,a20359a,a20360a,a20363a,a20367a,a20368a,a20369a,a20373a,a20374a,a20378a,a20379a,a20380a,a20383a,a20387a,a20388a,a20389a,a20393a,a20394a,a20398a,a20399a,a20400a,a20403a,a20407a,a20408a,a20409a,a20413a,a20414a,a20418a,a20419a,a20420a,a20423a,a20427a,a20428a,a20429a,a20433a,a20434a,a20438a,a20439a,a20440a,a20443a,a20447a,a20448a,a20449a,a20453a,a20454a,a20458a,a20459a,a20460a,a20463a,a20467a,a20468a,a20469a,a20473a,a20474a,a20478a,a20479a,a20480a,a20483a,a20487a,a20488a,a20489a,a20493a,a20494a,a20498a,a20499a,a20500a,a20503a,a20507a,a20508a,a20509a,a20513a,a20514a,a20518a,a20519a,a20520a,a20523a,a20527a,a20528a,a20529a,a20533a,a20534a,a20538a,a20539a,a20540a,a20543a,a20547a,a20548a,a20549a,a20553a,a20554a,a20558a,a20559a,a20560a,a20563a,a20567a,a20568a,a20569a,a20573a,a20574a,a20578a,a20579a,a20580a,a20583a,a20587a,a20588a,a20589a,a20593a,a20594a,a20598a,a20599a,a20600a,a20603a,a20607a,a20608a,a20609a,a20613a,a20614a,a20618a,a20619a,a20620a,a20623a,a20627a,a20628a,a20629a,a20633a,a20634a,a20638a,a20639a,a20640a,a20643a,a20647a,a20648a,a20649a,a20653a,a20654a,a20658a,a20659a,a20660a,a20663a,a20667a,a20668a,a20669a,a20673a,a20674a,a20678a,a20679a,a20680a,a20683a,a20687a,a20688a,a20689a,a20693a,a20694a,a20698a,a20699a,a20700a,a20703a,a20707a,a20708a,a20709a,a20713a,a20714a,a20718a,a20719a,a20720a,a20723a,a20727a,a20728a,a20729a,a20733a,a20734a,a20738a,a20739a,a20740a,a20743a,a20747a,a20748a,a20749a,a20753a,a20754a,a20758a,a20759a,a20760a,a20763a,a20767a,a20768a,a20769a,a20773a,a20774a,a20778a,a20779a,a20780a,a20783a,a20787a,a20788a,a20789a,a20793a,a20794a,a20798a,a20799a,a20800a,a20803a,a20807a,a20808a,a20809a,a20813a,a20814a,a20818a,a20819a,a20820a,a20823a,a20827a,a20828a,a20829a,a20833a,a20834a,a20838a,a20839a,a20840a,a20843a,a20847a,a20848a,a20849a,a20853a,a20854a,a20858a,a20859a,a20860a,a20863a,a20867a,a20868a,a20869a,a20873a,a20874a,a20878a,a20879a,a20880a,a20883a,a20887a,a20888a,a20889a,a20893a,a20894a,a20898a,a20899a,a20900a,a20903a,a20907a,a20908a,a20909a,a20913a,a20914a,a20918a,a20919a,a20920a,a20923a,a20927a,a20928a,a20929a,a20933a,a20934a,a20938a,a20939a,a20940a,a20943a,a20947a,a20948a,a20949a,a20953a,a20954a,a20958a,a20959a,a20960a,a20963a,a20967a,a20968a,a20969a,a20973a,a20974a,a20978a,a20979a,a20980a,a20983a,a20987a,a20988a,a20989a,a20993a,a20994a,a20998a,a20999a,a21000a,a21003a,a21007a,a21008a,a21009a,a21013a,a21014a,a21018a,a21019a,a21020a,a21023a,a21027a,a21028a,a21029a,a21033a,a21034a,a21038a,a21039a,a21040a,a21043a,a21047a,a21048a,a21049a,a21053a,a21054a,a21058a,a21059a,a21060a,a21063a,a21067a,a21068a,a21069a,a21073a,a21074a,a21078a,a21079a,a21080a,a21083a,a21087a,a21088a,a21089a,a21093a,a21094a,a21098a,a21099a,a21100a,a21103a,a21107a,a21108a,a21109a,a21113a,a21114a,a21118a,a21119a,a21120a,a21123a,a21127a,a21128a,a21129a,a21133a,a21134a,a21138a,a21139a,a21140a,a21143a,a21147a,a21148a,a21149a,a21153a,a21154a,a21158a,a21159a,a21160a,a21163a,a21167a,a21168a,a21169a,a21173a,a21174a,a21178a,a21179a,a21180a,a21183a,a21187a,a21188a,a21189a,a21193a,a21194a,a21198a,a21199a,a21200a,a21203a,a21207a,a21208a,a21209a,a21213a,a21214a,a21218a,a21219a,a21220a,a21223a,a21227a,a21228a,a21229a,a21233a,a21234a,a21238a,a21239a,a21240a,a21243a,a21247a,a21248a,a21249a,a21253a,a21254a,a21258a,a21259a,a21260a,a21263a,a21267a,a21268a,a21269a,a21273a,a21274a,a21278a,a21279a,a21280a,a21283a,a21287a,a21288a,a21289a,a21293a,a21294a,a21298a,a21299a,a21300a,a21303a,a21307a,a21308a,a21309a,a21313a,a21314a,a21318a,a21319a,a21320a,a21323a,a21327a,a21328a,a21329a,a21333a,a21334a,a21338a,a21339a,a21340a,a21343a,a21347a,a21348a,a21349a,a21353a,a21354a,a21358a,a21359a,a21360a,a21363a,a21367a,a21368a,a21369a,a21373a,a21374a,a21378a,a21379a,a21380a,a21383a,a21387a,a21388a,a21389a,a21393a,a21394a,a21398a,a21399a,a21400a,a21403a,a21407a,a21408a,a21409a,a21413a,a21414a,a21418a,a21419a,a21420a,a21423a,a21427a,a21428a,a21429a,a21433a,a21434a,a21438a,a21439a,a21440a,a21443a,a21447a,a21448a,a21449a,a21453a,a21454a,a21458a,a21459a,a21460a,a21463a,a21467a,a21468a,a21469a,a21473a,a21474a,a21478a,a21479a,a21480a,a21483a,a21487a,a21488a,a21489a,a21493a,a21494a,a21498a,a21499a,a21500a,a21503a,a21507a,a21508a,a21509a,a21513a,a21514a,a21518a,a21519a,a21520a,a21523a,a21527a,a21528a,a21529a,a21533a,a21534a,a21538a,a21539a,a21540a,a21543a,a21547a,a21548a,a21549a,a21553a,a21554a,a21558a,a21559a,a21560a,a21563a,a21567a,a21568a,a21569a,a21573a,a21574a,a21578a,a21579a,a21580a,a21583a,a21587a,a21588a,a21589a,a21593a,a21594a,a21598a,a21599a,a21600a,a21603a,a21607a,a21608a,a21609a,a21613a,a21614a,a21618a,a21619a,a21620a,a21623a,a21627a,a21628a,a21629a,a21633a,a21634a,a21638a,a21639a,a21640a,a21643a,a21647a,a21648a,a21649a,a21653a,a21654a,a21658a,a21659a,a21660a,a21663a,a21667a,a21668a,a21669a,a21673a,a21674a,a21678a,a21679a,a21680a,a21683a,a21687a,a21688a,a21689a,a21693a,a21694a,a21698a,a21699a,a21700a,a21703a,a21707a,a21708a,a21709a,a21713a,a21714a,a21718a,a21719a,a21720a,a21723a,a21727a,a21728a,a21729a,a21733a,a21734a,a21738a,a21739a,a21740a,a21743a,a21747a,a21748a,a21749a,a21753a,a21754a,a21758a,a21759a,a21760a,a21763a,a21767a,a21768a,a21769a,a21773a,a21774a,a21778a,a21779a,a21780a,a21783a,a21787a,a21788a,a21789a,a21793a,a21794a,a21798a,a21799a,a21800a,a21803a,a21807a,a21808a,a21809a,a21813a,a21814a,a21818a,a21819a,a21820a,a21823a,a21827a,a21828a,a21829a,a21833a,a21834a,a21838a,a21839a,a21840a,a21843a,a21847a,a21848a,a21849a,a21853a,a21854a,a21858a,a21859a,a21860a,a21863a,a21867a,a21868a,a21869a,a21873a,a21874a,a21878a,a21879a,a21880a,a21883a,a21887a,a21888a,a21889a,a21893a,a21894a,a21898a,a21899a,a21900a,a21903a,a21907a,a21908a,a21909a,a21913a,a21914a,a21918a,a21919a,a21920a,a21923a,a21927a,a21928a,a21929a,a21933a,a21934a,a21938a,a21939a,a21940a,a21943a,a21947a,a21948a,a21949a,a21953a,a21954a,a21958a,a21959a,a21960a,a21963a,a21967a,a21968a,a21969a,a21973a,a21974a,a21978a,a21979a,a21980a,a21983a,a21987a,a21988a,a21989a,a21993a,a21994a,a21998a,a21999a,a22000a,a22003a,a22007a,a22008a,a22009a,a22013a,a22014a,a22018a,a22019a,a22020a,a22023a,a22027a,a22028a,a22029a,a22033a,a22034a,a22038a,a22039a,a22040a,a22043a,a22047a,a22048a,a22049a,a22053a,a22054a,a22058a,a22059a,a22060a,a22063a,a22067a,a22068a,a22069a,a22073a,a22074a,a22078a,a22079a,a22080a,a22083a,a22087a,a22088a,a22089a,a22093a,a22094a,a22098a,a22099a,a22100a,a22103a,a22107a,a22108a,a22109a,a22113a,a22114a,a22118a,a22119a,a22120a,a22123a,a22127a,a22128a,a22129a,a22133a,a22134a,a22138a,a22139a,a22140a,a22143a,a22147a,a22148a,a22149a,a22153a,a22154a,a22158a,a22159a,a22160a,a22163a,a22167a,a22168a,a22169a,a22173a,a22174a,a22178a,a22179a,a22180a,a22183a,a22187a,a22188a,a22189a,a22193a,a22194a,a22198a,a22199a,a22200a,a22203a,a22207a,a22208a,a22209a,a22213a,a22214a,a22218a,a22219a,a22220a,a22223a,a22227a,a22228a,a22229a,a22233a,a22234a,a22238a,a22239a,a22240a,a22243a,a22247a,a22248a,a22249a,a22253a,a22254a,a22258a,a22259a,a22260a,a22263a,a22267a,a22268a,a22269a,a22273a,a22274a,a22278a,a22279a,a22280a,a22283a,a22287a,a22288a,a22289a,a22293a,a22294a,a22298a,a22299a,a22300a,a22303a,a22307a,a22308a,a22309a,a22313a,a22314a,a22318a,a22319a,a22320a,a22323a,a22327a,a22328a,a22329a,a22333a,a22334a,a22338a,a22339a,a22340a,a22343a,a22347a,a22348a,a22349a,a22353a,a22354a,a22358a,a22359a,a22360a,a22363a,a22367a,a22368a,a22369a,a22373a,a22374a,a22378a,a22379a,a22380a,a22383a,a22387a,a22388a,a22389a,a22393a,a22394a,a22398a,a22399a,a22400a,a22403a,a22407a,a22408a,a22409a,a22413a,a22414a,a22418a,a22419a,a22420a,a22423a,a22427a,a22428a,a22429a,a22433a,a22434a,a22438a,a22439a,a22440a,a22443a,a22447a,a22448a,a22449a,a22453a,a22454a,a22458a,a22459a,a22460a,a22463a,a22467a,a22468a,a22469a,a22473a,a22474a,a22478a,a22479a,a22480a,a22483a,a22487a,a22488a,a22489a,a22493a,a22494a,a22498a,a22499a,a22500a,a22503a,a22507a,a22508a,a22509a,a22513a,a22514a,a22518a,a22519a,a22520a,a22523a,a22527a,a22528a,a22529a,a22533a,a22534a,a22538a,a22539a,a22540a,a22543a,a22547a,a22548a,a22549a,a22553a,a22554a,a22558a,a22559a,a22560a,a22563a,a22567a,a22568a,a22569a,a22573a,a22574a,a22578a,a22579a,a22580a,a22583a,a22587a,a22588a,a22589a,a22593a,a22594a,a22598a,a22599a,a22600a,a22603a,a22607a,a22608a,a22609a,a22613a,a22614a,a22618a,a22619a,a22620a,a22623a,a22627a,a22628a,a22629a,a22633a,a22634a,a22638a,a22639a,a22640a,a22643a,a22647a,a22648a,a22649a,a22653a,a22654a,a22658a,a22659a,a22660a,a22663a,a22667a,a22668a,a22669a,a22673a,a22674a,a22678a,a22679a,a22680a,a22683a,a22687a,a22688a,a22689a,a22693a,a22694a,a22698a,a22699a,a22700a,a22703a,a22707a,a22708a,a22709a,a22713a,a22714a,a22718a,a22719a,a22720a,a22723a,a22727a,a22728a,a22729a,a22733a,a22734a,a22738a,a22739a,a22740a,a22743a,a22747a,a22748a,a22749a,a22753a,a22754a,a22758a,a22759a,a22760a,a22763a,a22767a,a22768a,a22769a,a22773a,a22774a,a22778a,a22779a,a22780a,a22783a,a22787a,a22788a,a22789a,a22793a,a22794a,a22798a,a22799a,a22800a,a22803a,a22807a,a22808a,a22809a,a22813a,a22814a,a22818a,a22819a,a22820a,a22823a,a22827a,a22828a,a22829a,a22833a,a22834a,a22838a,a22839a,a22840a,a22843a,a22847a,a22848a,a22849a,a22853a,a22854a,a22858a,a22859a,a22860a,a22863a,a22867a,a22868a,a22869a,a22873a,a22874a,a22878a,a22879a,a22880a,a22883a,a22887a,a22888a,a22889a,a22893a,a22894a,a22898a,a22899a,a22900a,a22903a,a22907a,a22908a,a22909a,a22913a,a22914a,a22918a,a22919a,a22920a,a22923a,a22927a,a22928a,a22929a,a22933a,a22934a,a22938a,a22939a,a22940a,a22943a,a22947a,a22948a,a22949a,a22953a,a22954a,a22958a,a22959a,a22960a,a22963a,a22967a,a22968a,a22969a,a22973a,a22974a,a22978a,a22979a,a22980a,a22983a,a22987a,a22988a,a22989a,a22993a,a22994a,a22998a,a22999a,a23000a,a23003a,a23007a,a23008a,a23009a,a23013a,a23014a,a23018a,a23019a,a23020a,a23023a,a23027a,a23028a,a23029a,a23033a,a23034a,a23038a,a23039a,a23040a,a23043a,a23047a,a23048a,a23049a,a23053a,a23054a,a23058a,a23059a,a23060a,a23063a,a23067a,a23068a,a23069a,a23073a,a23074a,a23078a,a23079a,a23080a,a23083a,a23087a,a23088a,a23089a,a23093a,a23094a,a23098a,a23099a,a23100a,a23103a,a23107a,a23108a,a23109a,a23113a,a23114a,a23118a,a23119a,a23120a,a23123a,a23127a,a23128a,a23129a,a23133a,a23134a,a23138a,a23139a,a23140a,a23143a,a23147a,a23148a,a23149a,a23153a,a23154a,a23158a,a23159a,a23160a,a23163a,a23167a,a23168a,a23169a,a23173a,a23174a,a23178a,a23179a,a23180a,a23183a,a23187a,a23188a,a23189a,a23193a,a23194a,a23198a,a23199a,a23200a,a23203a,a23207a,a23208a,a23209a,a23213a,a23214a,a23218a,a23219a,a23220a,a23223a,a23227a,a23228a,a23229a,a23233a,a23234a,a23238a,a23239a,a23240a,a23243a,a23247a,a23248a,a23249a,a23253a,a23254a,a23258a,a23259a,a23260a,a23263a,a23267a,a23268a,a23269a,a23273a,a23274a,a23278a,a23279a,a23280a,a23283a,a23287a,a23288a,a23289a,a23293a,a23294a,a23298a,a23299a,a23300a,a23303a,a23307a,a23308a,a23309a,a23313a,a23314a,a23318a,a23319a,a23320a,a23323a,a23327a,a23328a,a23329a,a23333a,a23334a,a23338a,a23339a,a23340a,a23343a,a23347a,a23348a,a23349a,a23353a,a23354a,a23358a,a23359a,a23360a,a23363a,a23367a,a23368a,a23369a,a23373a,a23374a,a23378a,a23379a,a23380a,a23383a,a23387a,a23388a,a23389a,a23393a,a23394a,a23398a,a23399a,a23400a,a23403a,a23407a,a23408a,a23409a,a23413a,a23414a,a23418a,a23419a,a23420a,a23423a,a23427a,a23428a,a23429a,a23433a,a23434a,a23438a,a23439a,a23440a,a23443a,a23447a,a23448a,a23449a,a23453a,a23454a,a23458a,a23459a,a23460a,a23463a,a23467a,a23468a,a23469a,a23473a,a23474a,a23478a,a23479a,a23480a,a23483a,a23487a,a23488a,a23489a,a23493a,a23494a,a23498a,a23499a,a23500a,a23503a,a23507a,a23508a,a23509a,a23513a,a23514a,a23518a,a23519a,a23520a,a23523a,a23527a,a23528a,a23529a,a23533a,a23534a,a23538a,a23539a,a23540a,a23543a,a23547a,a23548a,a23549a,a23553a,a23554a,a23558a,a23559a,a23560a,a23563a,a23567a,a23568a,a23569a,a23573a,a23574a,a23578a,a23579a,a23580a,a23583a,a23587a,a23588a,a23589a,a23593a,a23594a,a23598a,a23599a,a23600a,a23603a,a23607a,a23608a,a23609a,a23613a,a23614a,a23618a,a23619a,a23620a,a23623a,a23627a,a23628a,a23629a,a23633a,a23634a,a23638a,a23639a,a23640a,a23643a,a23647a,a23648a,a23649a,a23653a,a23654a,a23658a,a23659a,a23660a,a23663a,a23667a,a23668a,a23669a,a23673a,a23674a,a23678a,a23679a,a23680a,a23683a,a23687a,a23688a,a23689a,a23693a,a23694a,a23698a,a23699a,a23700a,a23703a,a23707a,a23708a,a23709a,a23713a,a23714a,a23718a,a23719a,a23720a,a23723a,a23727a,a23728a,a23729a,a23733a,a23734a,a23738a,a23739a,a23740a,a23743a,a23747a,a23748a,a23749a,a23753a,a23754a,a23758a,a23759a,a23760a,a23763a,a23767a,a23768a,a23769a,a23773a,a23774a,a23778a,a23779a,a23780a,a23783a,a23787a,a23788a,a23789a,a23793a,a23794a,a23798a,a23799a,a23800a,a23803a,a23807a,a23808a,a23809a,a23813a,a23814a,a23818a,a23819a,a23820a,a23823a,a23827a,a23828a,a23829a,a23833a,a23834a,a23838a,a23839a,a23840a,a23843a,a23847a,a23848a,a23849a,a23853a,a23854a,a23858a,a23859a,a23860a,a23863a,a23867a,a23868a,a23869a,a23873a,a23874a,a23878a,a23879a,a23880a,a23883a,a23887a,a23888a,a23889a,a23893a,a23894a,a23898a,a23899a,a23900a,a23903a,a23907a,a23908a,a23909a,a23913a,a23914a,a23918a,a23919a,a23920a,a23923a,a23927a,a23928a,a23929a,a23933a,a23934a,a23938a,a23939a,a23940a,a23943a,a23947a,a23948a,a23949a,a23953a,a23954a,a23958a,a23959a,a23960a,a23963a,a23967a,a23968a,a23969a,a23973a,a23974a,a23978a,a23979a,a23980a,a23983a,a23987a,a23988a,a23989a,a23993a,a23994a,a23998a,a23999a,a24000a,a24003a,a24007a,a24008a,a24009a,a24013a,a24014a,a24018a,a24019a,a24020a,a24023a,a24027a,a24028a,a24029a,a24033a,a24034a,a24038a,a24039a,a24040a,a24043a,a24047a,a24048a,a24049a,a24053a,a24054a,a24058a,a24059a,a24060a,a24063a,a24067a,a24068a,a24069a,a24073a,a24074a,a24078a,a24079a,a24080a,a24083a,a24087a,a24088a,a24089a,a24093a,a24094a,a24098a,a24099a,a24100a,a24103a,a24107a,a24108a,a24109a,a24113a,a24114a,a24118a,a24119a,a24120a,a24123a,a24127a,a24128a,a24129a,a24133a,a24134a,a24138a,a24139a,a24140a,a24143a,a24147a,a24148a,a24149a,a24153a,a24154a,a24158a,a24159a,a24160a,a24163a,a24167a,a24168a,a24169a,a24173a,a24174a,a24178a,a24179a,a24180a,a24183a,a24187a,a24188a,a24189a,a24193a,a24194a,a24198a,a24199a,a24200a,a24203a,a24207a,a24208a,a24209a,a24213a,a24214a,a24218a,a24219a,a24220a,a24223a,a24227a,a24228a,a24229a,a24233a,a24234a,a24238a,a24239a,a24240a,a24243a,a24247a,a24248a,a24249a,a24253a,a24254a,a24258a,a24259a,a24260a,a24263a,a24267a,a24268a,a24269a,a24273a,a24274a,a24278a,a24279a,a24280a,a24283a,a24287a,a24288a,a24289a,a24293a,a24294a,a24298a,a24299a,a24300a,a24303a,a24307a,a24308a,a24309a,a24313a,a24314a,a24318a,a24319a,a24320a,a24323a,a24327a,a24328a,a24329a,a24333a,a24334a,a24338a,a24339a,a24340a,a24343a,a24347a,a24348a,a24349a,a24353a,a24354a,a24358a,a24359a,a24360a,a24363a,a24367a,a24368a,a24369a,a24373a,a24374a,a24378a,a24379a,a24380a,a24383a,a24387a,a24388a,a24389a,a24393a,a24394a,a24398a,a24399a,a24400a,a24403a,a24407a,a24408a,a24409a,a24413a,a24414a,a24418a,a24419a,a24420a,a24423a,a24427a,a24428a,a24429a,a24433a,a24434a,a24438a,a24439a,a24440a,a24443a,a24447a,a24448a,a24449a,a24453a,a24454a,a24458a,a24459a,a24460a,a24464a,a24465a,a24469a,a24470a,a24471a,a24475a,a24476a,a24480a,a24481a,a24482a,a24486a,a24487a,a24491a,a24492a,a24493a,a24497a,a24498a,a24502a,a24503a,a24504a,a24508a,a24509a,a24513a,a24514a,a24515a,a24519a,a24520a,a24524a,a24525a,a24526a,a24530a,a24531a,a24535a,a24536a,a24537a,a24541a,a24542a,a24546a,a24547a,a24548a,a24552a,a24553a,a24557a,a24558a,a24559a,a24563a,a24564a,a24568a,a24569a,a24570a,a24574a,a24575a,a24579a,a24580a,a24581a,a24585a,a24586a,a24590a,a24591a,a24592a,a24596a,a24597a,a24601a,a24602a,a24603a,a24607a,a24608a,a24612a,a24613a,a24614a,a24618a,a24619a,a24623a,a24624a,a24625a,a24629a,a24630a,a24634a,a24635a,a24636a,a24640a,a24641a,a24645a,a24646a,a24647a,a24651a,a24652a,a24656a,a24657a,a24658a,a24662a,a24663a,a24667a,a24668a,a24669a,a24673a,a24674a,a24678a,a24679a,a24680a,a24684a,a24685a,a24689a,a24690a,a24691a,a24695a,a24696a,a24700a,a24701a,a24702a,a24706a,a24707a,a24711a,a24712a,a24713a,a24717a,a24718a,a24722a,a24723a,a24724a,a24728a,a24729a,a24733a,a24734a,a24735a,a24739a,a24740a,a24744a,a24745a,a24746a,a24750a,a24751a,a24755a,a24756a,a24757a,a24761a,a24762a,a24766a,a24767a,a24768a,a24772a,a24773a,a24777a,a24778a,a24779a,a24783a,a24784a,a24788a,a24789a,a24790a,a24794a,a24795a,a24799a,a24800a,a24801a,a24805a,a24806a,a24810a,a24811a,a24812a,a24816a,a24817a,a24821a,a24822a,a24823a,a24827a,a24828a,a24832a,a24833a,a24834a,a24838a,a24839a,a24843a,a24844a,a24845a,a24849a,a24850a,a24854a,a24855a,a24856a,a24860a,a24861a,a24865a,a24866a,a24867a,a24871a,a24872a,a24876a,a24877a,a24878a,a24882a,a24883a,a24887a,a24888a,a24889a,a24893a,a24894a,a24898a,a24899a,a24900a,a24904a,a24905a,a24909a,a24910a,a24911a,a24915a,a24916a,a24920a,a24921a,a24922a,a24926a,a24927a,a24931a,a24932a,a24933a,a24937a,a24938a,a24942a,a24943a,a24944a,a24948a,a24949a,a24953a,a24954a,a24955a,a24959a,a24960a,a24964a,a24965a,a24966a,a24970a,a24971a,a24975a,a24976a,a24977a,a24981a,a24982a,a24986a,a24987a,a24988a,a24992a,a24993a,a24997a,a24998a,a24999a,a25003a,a25004a,a25008a,a25009a,a25010a,a25014a,a25015a,a25019a,a25020a,a25021a,a25025a,a25026a,a25030a,a25031a,a25032a,a25036a,a25037a,a25041a,a25042a,a25043a,a25047a,a25048a,a25052a,a25053a,a25054a,a25058a,a25059a,a25063a,a25064a,a25065a,a25069a,a25070a,a25074a,a25075a,a25076a,a25080a,a25081a,a25085a,a25086a,a25087a,a25091a,a25092a,a25096a,a25097a,a25098a,a25102a,a25103a,a25107a,a25108a,a25109a,a25113a,a25114a,a25118a,a25119a,a25120a,a25124a,a25125a,a25129a,a25130a,a25131a,a25135a,a25136a,a25140a,a25141a,a25142a,a25146a,a25147a,a25151a,a25152a,a25153a,a25157a,a25158a,a25162a,a25163a,a25164a,a25168a,a25169a,a25173a,a25174a,a25175a,a25179a,a25180a,a25184a,a25185a,a25186a,a25190a,a25191a,a25195a,a25196a,a25197a,a25201a,a25202a,a25206a,a25207a,a25208a,a25212a,a25213a,a25217a,a25218a,a25219a,a25223a,a25224a,a25228a,a25229a,a25230a,a25234a,a25235a,a25239a,a25240a,a25241a,a25245a,a25246a,a25250a,a25251a,a25252a,a25256a,a25257a,a25261a,a25262a,a25263a,a25267a,a25268a,a25272a,a25273a,a25274a,a25278a,a25279a,a25283a,a25284a,a25285a,a25289a,a25290a,a25294a,a25295a,a25296a,a25300a,a25301a,a25305a,a25306a,a25307a,a25311a,a25312a,a25316a,a25317a,a25318a,a25322a,a25323a,a25327a,a25328a,a25329a,a25333a,a25334a,a25338a,a25339a,a25340a,a25344a,a25345a,a25349a,a25350a,a25351a,a25355a,a25356a,a25360a,a25361a,a25362a,a25366a,a25367a,a25371a,a25372a,a25373a,a25377a,a25378a,a25382a,a25383a,a25384a,a25388a,a25389a,a25393a,a25394a,a25395a,a25399a,a25400a,a25404a,a25405a,a25406a,a25410a,a25411a,a25415a,a25416a,a25417a,a25421a,a25422a,a25426a,a25427a,a25428a,a25432a,a25433a,a25437a,a25438a,a25439a,a25443a,a25444a,a25448a,a25449a,a25450a,a25454a,a25455a,a25459a,a25460a,a25461a,a25465a,a25466a,a25470a,a25471a,a25472a,a25476a,a25477a,a25481a,a25482a,a25483a,a25487a,a25488a,a25492a,a25493a,a25494a,a25498a,a25499a,a25503a,a25504a,a25505a,a25509a,a25510a,a25514a,a25515a,a25516a,a25520a,a25521a,a25525a,a25526a,a25527a,a25531a,a25532a,a25536a,a25537a,a25538a,a25542a,a25543a,a25547a,a25548a,a25549a,a25553a,a25554a,a25558a,a25559a,a25560a,a25564a,a25565a,a25569a,a25570a,a25571a,a25575a,a25576a,a25580a,a25581a,a25582a,a25586a,a25587a,a25591a,a25592a,a25593a,a25597a,a25598a,a25602a,a25603a,a25604a,a25608a,a25609a,a25613a,a25614a,a25615a,a25619a,a25620a,a25624a,a25625a,a25626a,a25630a,a25631a,a25635a,a25636a,a25637a,a25641a,a25642a,a25646a,a25647a,a25648a,a25652a,a25653a,a25657a,a25658a,a25659a,a25663a,a25664a,a25668a,a25669a,a25670a,a25674a,a25675a,a25679a,a25680a,a25681a,a25685a,a25686a,a25690a,a25691a,a25692a,a25696a,a25697a,a25701a,a25702a,a25703a,a25707a,a25708a,a25712a,a25713a,a25714a,a25718a,a25719a,a25723a,a25724a,a25725a,a25729a,a25730a,a25734a,a25735a,a25736a,a25740a,a25741a,a25745a,a25746a,a25747a,a25751a,a25752a,a25756a,a25757a,a25758a,a25762a,a25763a,a25767a,a25768a,a25769a,a25773a,a25774a,a25778a,a25779a,a25780a,a25784a,a25785a,a25789a,a25790a,a25791a,a25795a,a25796a,a25800a,a25801a,a25802a,a25806a,a25807a,a25811a,a25812a,a25813a,a25817a,a25818a,a25822a,a25823a,a25824a,a25828a,a25829a,a25833a,a25834a,a25835a,a25839a,a25840a,a25844a,a25845a,a25846a,a25850a,a25851a,a25855a,a25856a,a25857a,a25861a,a25862a,a25866a,a25867a,a25868a,a25872a,a25873a,a25877a,a25878a,a25879a,a25883a,a25884a,a25888a,a25889a,a25890a,a25894a,a25895a,a25899a,a25900a,a25901a,a25905a,a25906a,a25910a,a25911a,a25912a,a25916a,a25917a,a25921a,a25922a,a25923a,a25927a,a25928a,a25932a,a25933a,a25934a,a25938a,a25939a,a25943a,a25944a,a25945a,a25949a,a25950a,a25954a,a25955a,a25956a,a25960a,a25961a,a25965a,a25966a,a25967a,a25971a,a25972a,a25976a,a25977a,a25978a,a25982a,a25983a,a25987a,a25988a,a25989a,a25993a,a25994a,a25998a,a25999a,a26000a,a26004a,a26005a,a26009a,a26010a,a26011a,a26015a,a26016a,a26020a,a26021a,a26022a,a26026a,a26027a,a26031a,a26032a,a26033a,a26037a,a26038a,a26042a,a26043a,a26044a,a26048a,a26049a,a26053a,a26054a,a26055a,a26059a,a26060a,a26064a,a26065a,a26066a,a26070a,a26071a,a26075a,a26076a,a26077a,a26081a,a26082a,a26086a,a26087a,a26088a,a26092a,a26093a,a26097a,a26098a,a26099a,a26103a,a26104a,a26108a,a26109a,a26110a,a26114a,a26115a,a26119a,a26120a,a26121a,a26125a,a26126a,a26130a,a26131a,a26132a,a26136a,a26137a,a26141a,a26142a,a26143a,a26147a,a26148a,a26152a,a26153a,a26154a,a26158a,a26159a,a26163a,a26164a,a26165a,a26169a,a26170a,a26174a,a26175a,a26176a,a26180a,a26181a,a26185a,a26186a,a26187a,a26191a,a26192a,a26196a,a26197a,a26198a,a26202a,a26203a,a26207a,a26208a,a26209a,a26213a,a26214a,a26218a,a26219a,a26220a,a26224a,a26225a,a26229a,a26230a,a26231a,a26235a,a26236a,a26240a,a26241a,a26242a,a26246a,a26247a,a26251a,a26252a,a26253a,a26257a,a26258a,a26262a,a26263a,a26264a,a26268a,a26269a,a26273a,a26274a,a26275a,a26279a,a26280a,a26284a,a26285a,a26286a,a26290a,a26291a,a26295a,a26296a,a26297a,a26301a,a26302a,a26306a,a26307a,a26308a,a26312a,a26313a,a26317a,a26318a,a26319a,a26323a,a26324a,a26328a,a26329a,a26330a,a26334a,a26335a,a26339a,a26340a,a26341a,a26345a,a26346a,a26350a,a26351a,a26352a,a26356a,a26357a,a26361a,a26362a,a26363a,a26367a,a26368a,a26372a,a26373a,a26374a,a26378a,a26379a,a26383a,a26384a,a26385a,a26389a,a26390a,a26394a,a26395a,a26396a,a26400a,a26401a,a26405a,a26406a,a26407a,a26411a,a26412a,a26416a,a26417a,a26418a,a26422a,a26423a,a26427a,a26428a,a26429a,a26433a,a26434a,a26438a,a26439a,a26440a,a26444a,a26445a,a26449a,a26450a,a26451a,a26455a,a26456a,a26460a,a26461a,a26462a,a26466a,a26467a,a26471a,a26472a,a26473a,a26477a,a26478a,a26482a,a26483a,a26484a,a26488a,a26489a,a26493a,a26494a,a26495a,a26499a,a26500a,a26504a,a26505a,a26506a,a26510a,a26511a,a26515a,a26516a,a26517a,a26521a,a26522a,a26526a,a26527a,a26528a,a26532a,a26533a,a26537a,a26538a,a26539a,a26543a,a26544a,a26548a,a26549a,a26550a,a26554a,a26555a,a26559a,a26560a,a26561a,a26565a,a26566a,a26570a,a26571a,a26572a,a26576a,a26577a,a26581a,a26582a,a26583a,a26587a,a26588a,a26592a,a26593a,a26594a,a26598a,a26599a,a26603a,a26604a,a26605a,a26609a,a26610a,a26614a,a26615a,a26616a,a26620a,a26621a,a26625a,a26626a,a26627a,a26631a,a26632a,a26636a,a26637a,a26638a,a26642a,a26643a,a26647a,a26648a,a26649a,a26653a,a26654a,a26658a,a26659a,a26660a,a26664a,a26665a,a26669a,a26670a,a26671a,a26675a,a26676a,a26680a,a26681a,a26682a,a26686a,a26687a,a26691a,a26692a,a26693a,a26697a,a26698a,a26702a,a26703a,a26704a,a26708a,a26709a,a26713a,a26714a,a26715a,a26719a,a26720a,a26724a,a26725a,a26726a,a26730a,a26731a,a26735a,a26736a,a26737a,a26741a,a26742a,a26746a,a26747a,a26748a,a26752a,a26753a,a26757a,a26758a,a26759a,a26763a,a26764a,a26768a,a26769a,a26770a,a26774a,a26775a,a26779a,a26780a,a26781a,a26785a,a26786a,a26790a,a26791a,a26792a,a26796a,a26797a,a26801a,a26802a,a26803a,a26807a,a26808a,a26812a,a26813a,a26814a,a26818a,a26819a,a26823a,a26824a,a26825a,a26829a,a26830a,a26834a,a26835a,a26836a,a26840a,a26841a,a26845a,a26846a,a26847a,a26851a,a26852a,a26856a,a26857a,a26858a,a26862a,a26863a,a26867a,a26868a,a26869a,a26873a,a26874a,a26878a,a26879a,a26880a,a26884a,a26885a,a26889a,a26890a,a26891a,a26895a,a26896a,a26900a,a26901a,a26902a,a26906a,a26907a,a26911a,a26912a,a26913a,a26917a,a26918a,a26922a,a26923a,a26924a,a26928a,a26929a,a26933a,a26934a,a26935a,a26939a,a26940a,a26944a,a26945a,a26946a,a26950a,a26951a,a26955a,a26956a,a26957a,a26961a,a26962a,a26966a,a26967a,a26968a,a26972a,a26973a,a26977a,a26978a,a26979a,a26983a,a26984a,a26988a,a26989a,a26990a,a26994a,a26995a,a26999a,a27000a,a27001a,a27005a,a27006a,a27010a,a27011a,a27012a,a27016a,a27017a,a27021a,a27022a,a27023a,a27027a,a27028a,a27032a,a27033a,a27034a,a27038a,a27039a,a27043a,a27044a,a27045a,a27049a,a27050a,a27054a,a27055a,a27056a,a27060a,a27061a,a27065a,a27066a,a27067a,a27071a,a27072a,a27076a,a27077a,a27078a,a27082a,a27083a,a27087a,a27088a,a27089a,a27093a,a27094a,a27098a,a27099a,a27100a,a27104a,a27105a,a27109a,a27110a,a27111a,a27115a,a27116a,a27120a,a27121a,a27122a,a27126a,a27127a,a27131a,a27132a,a27133a,a27137a,a27138a,a27142a,a27143a,a27144a,a27148a,a27149a,a27153a,a27154a,a27155a,a27159a,a27160a,a27164a,a27165a,a27166a,a27170a,a27171a,a27175a,a27176a,a27177a,a27181a,a27182a,a27186a,a27187a,a27188a,a27192a,a27193a,a27197a,a27198a,a27199a,a27203a,a27204a,a27208a,a27209a,a27210a,a27214a,a27215a,a27219a,a27220a,a27221a,a27225a,a27226a,a27230a,a27231a,a27232a,a27236a,a27237a,a27241a,a27242a,a27243a,a27247a,a27248a,a27252a,a27253a,a27254a,a27258a,a27259a,a27263a,a27264a,a27265a,a27269a,a27270a,a27274a,a27275a,a27276a,a27280a,a27281a,a27285a,a27286a,a27287a,a27291a,a27292a,a27296a,a27297a,a27298a,a27302a,a27303a,a27307a,a27308a,a27309a,a27313a,a27314a,a27318a,a27319a,a27320a,a27324a,a27325a,a27329a,a27330a,a27331a,a27335a,a27336a,a27340a,a27341a,a27342a,a27346a,a27347a,a27351a,a27352a,a27353a,a27357a,a27358a,a27362a,a27363a,a27364a,a27368a,a27369a,a27373a,a27374a,a27375a,a27379a,a27380a,a27384a,a27385a,a27386a,a27390a,a27391a,a27395a,a27396a,a27397a,a27401a,a27402a,a27406a,a27407a,a27408a,a27412a,a27413a,a27417a,a27418a,a27419a,a27423a,a27424a,a27428a,a27429a,a27430a,a27434a,a27435a,a27439a,a27440a,a27441a,a27445a,a27446a,a27450a,a27451a,a27452a,a27456a,a27457a,a27461a,a27462a,a27463a,a27467a,a27468a,a27472a,a27473a,a27474a,a27478a,a27479a,a27483a,a27484a,a27485a,a27489a,a27490a,a27494a,a27495a,a27496a,a27500a,a27501a,a27505a,a27506a,a27507a,a27511a,a27512a,a27516a,a27517a,a27518a,a27522a,a27523a,a27527a,a27528a,a27529a,a27533a,a27534a,a27538a,a27539a,a27540a,a27544a,a27545a,a27549a,a27550a,a27551a,a27555a,a27556a,a27560a,a27561a,a27562a,a27566a,a27567a,a27571a,a27572a,a27573a,a27577a,a27578a,a27582a,a27583a,a27584a,a27588a,a27589a,a27593a,a27594a,a27595a,a27599a,a27600a,a27604a,a27605a,a27606a,a27610a,a27611a,a27615a,a27616a,a27617a,a27621a,a27622a,a27626a,a27627a,a27628a,a27632a,a27633a,a27637a,a27638a,a27639a,a27643a,a27644a,a27648a,a27649a,a27650a,a27654a,a27655a,a27659a,a27660a,a27661a,a27665a,a27666a,a27670a,a27671a,a27672a,a27676a,a27677a,a27681a,a27682a,a27683a,a27687a,a27688a,a27692a,a27693a,a27694a,a27698a,a27699a,a27703a,a27704a,a27705a,a27709a,a27710a,a27714a,a27715a,a27716a,a27720a,a27721a,a27725a,a27726a,a27727a,a27731a,a27732a,a27736a,a27737a,a27738a,a27742a,a27743a,a27747a,a27748a,a27749a,a27753a,a27754a,a27758a,a27759a,a27760a,a27764a,a27765a,a27769a,a27770a,a27771a,a27775a,a27776a,a27780a,a27781a,a27782a,a27786a,a27787a,a27791a,a27792a,a27793a,a27797a,a27798a,a27802a,a27803a,a27804a,a27808a,a27809a,a27813a,a27814a,a27815a,a27819a,a27820a,a27824a,a27825a,a27826a,a27830a,a27831a,a27835a,a27836a,a27837a,a27841a,a27842a,a27846a,a27847a,a27848a,a27852a,a27853a,a27857a,a27858a,a27859a,a27863a,a27864a,a27868a,a27869a,a27870a,a27874a,a27875a,a27879a,a27880a,a27881a,a27885a,a27886a,a27890a,a27891a,a27892a,a27896a,a27897a,a27901a,a27902a,a27903a,a27907a,a27908a,a27912a,a27913a,a27914a,a27918a,a27919a,a27923a,a27924a,a27925a,a27929a,a27930a,a27934a,a27935a,a27936a,a27940a,a27941a,a27945a,a27946a,a27947a,a27951a,a27952a,a27956a,a27957a,a27958a,a27962a,a27963a,a27967a,a27968a,a27969a,a27973a,a27974a,a27978a,a27979a,a27980a,a27984a,a27985a,a27989a,a27990a,a27991a,a27995a,a27996a,a28000a,a28001a,a28002a,a28006a,a28007a,a28011a,a28012a,a28013a,a28017a,a28018a,a28022a,a28023a,a28024a,a28028a,a28029a,a28033a,a28034a,a28035a,a28039a,a28040a,a28044a,a28045a,a28046a,a28050a,a28051a,a28055a,a28056a,a28057a,a28061a,a28062a,a28066a,a28067a,a28068a,a28072a,a28073a,a28077a,a28078a,a28079a,a28083a,a28084a,a28088a,a28089a,a28090a,a28094a,a28095a,a28099a,a28100a,a28101a,a28105a,a28106a,a28110a,a28111a,a28112a,a28116a,a28117a,a28121a,a28122a,a28123a,a28127a,a28128a,a28132a,a28133a,a28134a,a28138a,a28139a,a28143a,a28144a,a28145a,a28149a,a28150a,a28154a,a28155a,a28156a,a28160a,a28161a,a28165a,a28166a,a28167a,a28171a,a28172a,a28176a,a28177a,a28178a,a28182a,a28183a,a28187a,a28188a,a28189a,a28193a,a28194a,a28198a,a28199a,a28200a,a28204a,a28205a,a28209a,a28210a,a28211a,a28215a,a28216a,a28220a,a28221a,a28222a,a28226a,a28227a,a28231a,a28232a,a28233a,a28237a,a28238a,a28242a,a28243a,a28244a,a28248a,a28249a,a28253a,a28254a,a28255a,a28259a,a28260a,a28264a,a28265a,a28266a,a28270a,a28271a,a28275a,a28276a,a28277a,a28281a,a28282a,a28286a,a28287a,a28288a,a28292a,a28293a,a28297a,a28298a,a28299a,a28303a,a28304a,a28308a,a28309a,a28310a,a28314a,a28315a,a28319a,a28320a,a28321a,a28325a,a28326a,a28330a,a28331a,a28332a,a28336a,a28337a,a28341a,a28342a,a28343a,a28347a,a28348a,a28352a,a28353a,a28354a,a28358a,a28359a,a28363a,a28364a,a28365a,a28369a,a28370a,a28374a,a28375a,a28376a,a28380a,a28381a,a28385a,a28386a,a28387a,a28391a,a28392a,a28396a,a28397a,a28398a,a28402a,a28403a,a28407a,a28408a,a28409a,a28413a,a28414a,a28418a,a28419a,a28420a,a28424a,a28425a,a28429a,a28430a,a28431a,a28435a,a28436a,a28440a,a28441a,a28442a,a28446a,a28447a,a28451a,a28452a,a28453a,a28457a,a28458a,a28462a,a28463a,a28464a,a28468a,a28469a,a28473a,a28474a,a28475a,a28479a,a28480a,a28484a,a28485a,a28486a,a28490a,a28491a,a28495a,a28496a,a28497a,a28501a,a28502a,a28506a,a28507a,a28508a,a28512a,a28513a,a28517a,a28518a,a28519a,a28523a,a28524a,a28528a,a28529a,a28530a,a28534a,a28535a,a28539a,a28540a,a28541a,a28545a,a28546a,a28550a,a28551a,a28552a,a28556a,a28557a,a28561a,a28562a,a28563a,a28567a,a28568a,a28572a,a28573a,a28574a,a28578a,a28579a,a28583a,a28584a,a28585a,a28589a,a28590a,a28594a,a28595a,a28596a,a28600a,a28601a,a28605a,a28606a,a28607a,a28611a,a28612a,a28616a,a28617a,a28618a,a28622a,a28623a,a28627a,a28628a,a28629a,a28633a,a28634a,a28638a,a28639a,a28640a,a28644a,a28645a,a28649a,a28650a,a28651a,a28655a,a28656a,a28660a,a28661a,a28662a,a28666a,a28667a,a28671a,a28672a,a28673a,a28677a,a28678a,a28682a,a28683a,a28684a,a28688a,a28689a,a28693a,a28694a,a28695a,a28699a,a28700a,a28704a,a28705a,a28706a,a28710a,a28711a,a28715a,a28716a,a28717a,a28721a,a28722a,a28726a,a28727a,a28728a,a28732a,a28733a,a28737a,a28738a,a28739a,a28743a,a28744a,a28748a,a28749a,a28750a,a28754a,a28755a,a28759a,a28760a,a28761a,a28765a,a28766a,a28770a,a28771a,a28772a,a28776a,a28777a,a28781a,a28782a,a28783a,a28787a,a28788a,a28792a,a28793a,a28794a,a28798a,a28799a,a28803a,a28804a,a28805a,a28809a,a28810a,a28814a,a28815a,a28816a,a28820a,a28821a,a28825a,a28826a,a28827a,a28831a,a28832a,a28836a,a28837a,a28838a,a28842a,a28843a,a28847a,a28848a,a28849a,a28853a,a28854a,a28858a,a28859a,a28860a,a28864a,a28865a,a28869a,a28870a,a28871a,a28875a,a28876a,a28880a,a28881a,a28882a,a28886a,a28887a,a28891a,a28892a,a28893a,a28897a,a28898a,a28902a,a28903a,a28904a,a28908a,a28909a,a28913a,a28914a,a28915a,a28919a,a28920a,a28924a,a28925a,a28926a,a28930a,a28931a,a28935a,a28936a,a28937a,a28941a,a28942a,a28946a,a28947a,a28948a,a28952a,a28953a,a28957a,a28958a,a28959a,a28963a,a28964a,a28968a,a28969a,a28970a,a28974a,a28975a,a28979a,a28980a,a28981a,a28985a,a28986a,a28990a,a28991a,a28992a,a28996a,a28997a,a29001a,a29002a,a29003a,a29007a,a29008a,a29012a,a29013a,a29014a,a29018a,a29019a,a29023a,a29024a,a29025a,a29029a,a29030a,a29034a,a29035a,a29036a,a29040a,a29041a,a29045a,a29046a,a29047a,a29051a,a29052a,a29056a,a29057a,a29058a,a29062a,a29063a,a29067a,a29068a,a29069a,a29073a,a29074a,a29078a,a29079a,a29080a,a29084a,a29085a,a29089a,a29090a,a29091a,a29095a,a29096a,a29100a,a29101a,a29102a,a29106a,a29107a,a29111a,a29112a,a29113a,a29117a,a29118a,a29122a,a29123a,a29124a,a29128a,a29129a,a29133a,a29134a,a29135a,a29139a,a29140a,a29144a,a29145a,a29146a,a29150a,a29151a,a29155a,a29156a,a29157a,a29161a,a29162a,a29166a,a29167a,a29168a,a29172a,a29173a,a29177a,a29178a,a29179a,a29183a,a29184a,a29188a,a29189a,a29190a,a29194a,a29195a,a29199a,a29200a,a29201a,a29205a,a29206a,a29210a,a29211a,a29212a,a29216a,a29217a,a29221a,a29222a,a29223a,a29227a,a29228a,a29232a,a29233a,a29234a,a29238a,a29239a,a29243a,a29244a,a29245a,a29249a,a29250a,a29254a,a29255a,a29256a,a29260a,a29261a,a29265a,a29266a,a29267a,a29271a,a29272a,a29276a,a29277a,a29278a,a29282a,a29283a,a29287a,a29288a,a29289a,a29293a,a29294a,a29298a,a29299a,a29300a,a29304a,a29305a,a29309a,a29310a,a29311a,a29315a,a29316a,a29320a,a29321a,a29322a,a29326a,a29327a,a29331a,a29332a,a29333a,a29337a,a29338a,a29342a,a29343a,a29344a,a29348a,a29349a,a29353a,a29354a,a29355a,a29359a,a29360a,a29364a,a29365a,a29366a,a29370a,a29371a,a29375a,a29376a,a29377a,a29381a,a29382a,a29386a,a29387a,a29388a,a29392a,a29393a,a29397a,a29398a,a29399a,a29403a,a29404a,a29408a,a29409a,a29410a,a29414a,a29415a,a29419a,a29420a,a29421a,a29425a,a29426a,a29430a,a29431a,a29432a,a29436a,a29437a,a29441a,a29442a,a29443a,a29447a,a29448a,a29452a,a29453a,a29454a,a29458a,a29459a,a29463a,a29464a,a29465a,a29469a,a29470a,a29474a,a29475a,a29476a,a29480a,a29481a,a29485a,a29486a,a29487a,a29491a,a29492a,a29496a,a29497a,a29498a,a29502a,a29503a,a29507a,a29508a,a29509a,a29513a,a29514a,a29518a,a29519a,a29520a,a29524a,a29525a,a29529a,a29530a,a29531a,a29535a,a29536a,a29540a,a29541a,a29542a,a29546a,a29547a,a29551a,a29552a,a29553a,a29557a,a29558a,a29562a,a29563a,a29564a,a29568a,a29569a,a29573a,a29574a,a29575a,a29579a,a29580a,a29584a,a29585a,a29586a,a29590a,a29591a,a29595a,a29596a,a29597a,a29601a,a29602a,a29606a,a29607a,a29608a,a29612a,a29613a,a29617a,a29618a,a29619a,a29623a,a29624a,a29628a,a29629a,a29630a,a29634a,a29635a,a29639a,a29640a,a29641a,a29645a,a29646a,a29650a,a29651a,a29652a,a29656a,a29657a,a29661a,a29662a,a29663a,a29667a,a29668a,a29672a,a29673a,a29674a,a29678a,a29679a,a29683a,a29684a,a29685a,a29689a,a29690a,a29694a,a29695a,a29696a,a29700a,a29701a,a29705a,a29706a,a29707a,a29711a,a29712a,a29716a,a29717a,a29718a,a29722a,a29723a,a29727a,a29728a,a29729a,a29733a,a29734a,a29738a,a29739a,a29740a,a29744a,a29745a,a29749a,a29750a,a29751a,a29755a,a29756a,a29760a,a29761a,a29762a,a29766a,a29767a,a29771a,a29772a,a29773a,a29777a,a29778a,a29782a,a29783a,a29784a,a29788a,a29789a,a29793a,a29794a,a29795a,a29799a,a29800a,a29804a,a29805a,a29806a,a29810a,a29811a,a29815a,a29816a,a29817a,a29821a,a29822a,a29826a,a29827a,a29828a,a29832a,a29833a,a29837a,a29838a,a29839a,a29843a,a29844a,a29848a,a29849a,a29850a,a29854a,a29855a,a29859a,a29860a,a29861a,a29865a,a29866a,a29870a,a29871a,a29872a,a29876a,a29877a,a29881a,a29882a,a29883a,a29887a,a29888a,a29892a,a29893a,a29894a,a29898a,a29899a,a29903a,a29904a,a29905a,a29909a,a29910a,a29914a,a29915a,a29916a,a29920a,a29921a,a29925a,a29926a,a29927a,a29931a,a29932a,a29936a,a29937a,a29938a,a29942a,a29943a,a29947a,a29948a,a29949a,a29953a,a29954a,a29958a,a29959a,a29960a,a29964a,a29965a,a29969a,a29970a,a29971a,a29975a,a29976a,a29980a,a29981a,a29982a,a29986a,a29987a,a29991a,a29992a,a29993a,a29997a,a29998a,a30002a,a30003a,a30004a,a30008a,a30009a,a30013a,a30014a,a30015a,a30019a,a30020a,a30024a,a30025a,a30026a,a30030a,a30031a,a30035a,a30036a,a30037a,a30041a,a30042a,a30046a,a30047a,a30048a,a30052a,a30053a,a30057a,a30058a,a30059a,a30063a,a30064a,a30068a,a30069a,a30070a,a30074a,a30075a,a30079a,a30080a,a30081a,a30085a,a30086a,a30090a,a30091a,a30092a,a30096a,a30097a,a30101a,a30102a,a30103a,a30107a,a30108a,a30112a,a30113a,a30114a,a30118a,a30119a,a30123a,a30124a,a30125a,a30129a,a30130a,a30134a,a30135a,a30136a,a30140a,a30141a,a30145a,a30146a,a30147a,a30151a,a30152a,a30156a,a30157a,a30158a,a30162a,a30163a,a30167a,a30168a,a30169a,a30173a,a30174a,a30178a,a30179a,a30180a,a30184a,a30185a,a30189a,a30190a,a30191a,a30195a,a30196a,a30200a,a30201a,a30202a,a30206a,a30207a,a30211a,a30212a,a30213a,a30217a,a30218a,a30222a,a30223a,a30224a,a30228a,a30229a,a30233a,a30234a,a30235a,a30239a,a30240a,a30244a,a30245a,a30246a,a30250a,a30251a,a30255a,a30256a,a30257a,a30261a,a30262a,a30266a,a30267a,a30268a,a30272a,a30273a,a30277a,a30278a,a30279a,a30283a,a30284a,a30288a,a30289a,a30290a,a30294a,a30295a,a30299a,a30300a,a30301a,a30305a,a30306a,a30310a,a30311a,a30312a,a30316a,a30317a,a30321a,a30322a,a30323a,a30327a,a30328a,a30332a,a30333a,a30334a,a30338a,a30339a,a30343a,a30344a,a30345a,a30349a,a30350a,a30354a,a30355a,a30356a,a30360a,a30361a,a30365a,a30366a,a30367a,a30371a,a30372a,a30376a,a30377a,a30378a,a30382a,a30383a,a30387a,a30388a,a30389a,a30393a,a30394a,a30398a,a30399a,a30400a,a30404a,a30405a,a30409a,a30410a,a30411a,a30415a,a30416a,a30420a,a30421a,a30422a,a30426a,a30427a,a30431a,a30432a,a30433a,a30437a,a30438a,a30442a,a30443a,a30444a,a30448a,a30449a,a30453a,a30454a,a30455a,a30459a,a30460a,a30464a,a30465a,a30466a,a30470a,a30471a,a30475a,a30476a,a30477a,a30481a,a30482a,a30486a,a30487a,a30488a,a30492a,a30493a,a30497a,a30498a,a30499a,a30503a,a30504a,a30508a,a30509a,a30510a,a30514a,a30515a,a30519a,a30520a,a30521a,a30525a,a30526a,a30530a,a30531a,a30532a,a30536a,a30537a,a30541a,a30542a,a30543a,a30547a,a30548a,a30552a,a30553a,a30554a,a30558a,a30559a,a30563a,a30564a,a30565a,a30569a,a30570a,a30574a,a30575a,a30576a,a30580a,a30581a,a30585a,a30586a,a30587a,a30591a,a30592a,a30596a,a30597a,a30598a,a30602a,a30603a,a30607a,a30608a,a30609a,a30613a,a30614a,a30618a,a30619a,a30620a,a30624a,a30625a,a30629a,a30630a,a30631a,a30635a,a30636a,a30639a,a30642a,a30643a,a30644a,a30648a,a30649a,a30653a,a30654a,a30655a,a30659a,a30660a,a30663a,a30666a,a30667a,a30668a,a30672a,a30673a,a30677a,a30678a,a30679a,a30683a,a30684a,a30687a,a30690a,a30691a,a30692a,a30696a,a30697a,a30701a,a30702a,a30703a,a30707a,a30708a,a30711a,a30714a,a30715a,a30716a,a30720a,a30721a,a30725a,a30726a,a30727a,a30731a,a30732a,a30735a,a30738a,a30739a,a30740a,a30744a,a30745a,a30749a,a30750a,a30751a,a30755a,a30756a,a30759a,a30762a,a30763a,a30764a,a30768a,a30769a,a30773a,a30774a,a30775a,a30779a,a30780a,a30783a,a30786a,a30787a,a30788a,a30792a,a30793a,a30797a,a30798a,a30799a,a30803a,a30804a,a30807a,a30810a,a30811a,a30812a,a30816a,a30817a,a30821a,a30822a,a30823a,a30827a,a30828a,a30831a,a30834a,a30835a,a30836a,a30840a,a30841a,a30845a,a30846a,a30847a,a30851a,a30852a,a30855a,a30858a,a30859a,a30860a,a30864a,a30865a,a30869a,a30870a,a30871a,a30875a,a30876a,a30879a,a30882a,a30883a,a30884a,a30888a,a30889a,a30893a,a30894a,a30895a,a30899a,a30900a,a30903a,a30906a,a30907a,a30908a,a30912a,a30913a,a30917a,a30918a,a30919a,a30923a,a30924a,a30927a,a30930a,a30931a,a30932a,a30936a,a30937a,a30941a,a30942a,a30943a,a30947a,a30948a,a30951a,a30954a,a30955a,a30956a,a30960a,a30961a,a30965a,a30966a,a30967a,a30971a,a30972a,a30975a,a30978a,a30979a,a30980a,a30984a,a30985a,a30989a,a30990a,a30991a,a30995a,a30996a,a30999a,a31002a,a31003a,a31004a,a31008a,a31009a,a31013a,a31014a,a31015a,a31019a,a31020a,a31023a,a31026a,a31027a,a31028a,a31032a,a31033a,a31037a,a31038a,a31039a,a31043a,a31044a,a31047a,a31050a,a31051a,a31052a,a31056a,a31057a,a31061a,a31062a,a31063a,a31067a,a31068a,a31071a,a31074a,a31075a,a31076a,a31080a,a31081a,a31085a,a31086a,a31087a,a31091a,a31092a,a31095a,a31098a,a31099a,a31100a,a31104a,a31105a,a31109a,a31110a,a31111a,a31115a,a31116a,a31119a,a31122a,a31123a,a31124a,a31128a,a31129a,a31133a,a31134a,a31135a,a31139a,a31140a,a31143a,a31146a,a31147a,a31148a,a31152a,a31153a,a31157a,a31158a,a31159a,a31163a,a31164a,a31167a,a31170a,a31171a,a31172a,a31176a,a31177a,a31181a,a31182a,a31183a,a31187a,a31188a,a31191a,a31194a,a31195a,a31196a,a31200a,a31201a,a31205a,a31206a,a31207a,a31211a,a31212a,a31215a,a31218a,a31219a,a31220a,a31224a,a31225a,a31229a,a31230a,a31231a,a31235a,a31236a,a31239a,a31242a,a31243a,a31244a,a31248a,a31249a,a31253a,a31254a,a31255a,a31259a,a31260a,a31263a,a31266a,a31267a,a31268a,a31272a,a31273a,a31277a,a31278a,a31279a,a31283a,a31284a,a31287a,a31290a,a31291a,a31292a,a31296a,a31297a,a31301a,a31302a,a31303a,a31307a,a31308a,a31311a,a31314a,a31315a,a31316a,a31320a,a31321a,a31325a,a31326a,a31327a,a31331a,a31332a,a31335a,a31338a,a31339a,a31340a,a31344a,a31345a,a31349a,a31350a,a31351a,a31355a,a31356a,a31359a,a31362a,a31363a,a31364a,a31368a,a31369a,a31373a,a31374a,a31375a,a31379a,a31380a,a31383a,a31386a,a31387a,a31388a,a31392a,a31393a,a31397a,a31398a,a31399a,a31403a,a31404a,a31407a,a31410a,a31411a,a31412a,a31416a,a31417a,a31421a,a31422a,a31423a,a31427a,a31428a,a31431a,a31434a,a31435a,a31436a,a31440a,a31441a,a31445a,a31446a,a31447a,a31451a,a31452a,a31455a,a31458a,a31459a,a31460a,a31464a,a31465a,a31469a,a31470a,a31471a,a31475a,a31476a,a31479a,a31482a,a31483a,a31484a,a31488a,a31489a,a31493a,a31494a,a31495a,a31499a,a31500a,a31503a,a31506a,a31507a,a31508a,a31512a,a31513a,a31517a,a31518a,a31519a,a31523a,a31524a,a31527a,a31530a,a31531a,a31532a,a31536a,a31537a,a31541a,a31542a,a31543a,a31547a,a31548a,a31551a,a31554a,a31555a,a31556a,a31560a,a31561a,a31565a,a31566a,a31567a,a31571a,a31572a,a31575a,a31578a,a31579a,a31580a,a31584a,a31585a,a31589a,a31590a,a31591a,a31595a,a31596a,a31599a,a31602a,a31603a,a31604a,a31608a,a31609a,a31613a,a31614a,a31615a,a31619a,a31620a,a31623a,a31626a,a31627a,a31628a,a31632a,a31633a,a31637a,a31638a,a31639a,a31643a,a31644a,a31647a,a31650a,a31651a,a31652a,a31656a,a31657a,a31661a,a31662a,a31663a,a31667a,a31668a,a31671a,a31674a,a31675a,a31676a,a31680a,a31681a,a31685a,a31686a,a31687a,a31691a,a31692a,a31695a,a31698a,a31699a,a31700a,a31704a,a31705a,a31709a,a31710a,a31711a,a31715a,a31716a,a31719a,a31722a,a31723a,a31724a,a31728a,a31729a,a31733a,a31734a,a31735a,a31739a,a31740a,a31743a,a31746a,a31747a,a31748a,a31752a,a31753a,a31757a,a31758a,a31759a,a31763a,a31764a,a31767a,a31770a,a31771a,a31772a,a31776a,a31777a,a31781a,a31782a,a31783a,a31787a,a31788a,a31791a,a31794a,a31795a,a31796a,a31800a,a31801a,a31805a,a31806a,a31807a,a31811a,a31812a,a31815a,a31818a,a31819a,a31820a,a31824a,a31825a,a31829a,a31830a,a31831a,a31835a,a31836a,a31839a,a31842a,a31843a,a31844a,a31848a,a31849a,a31853a,a31854a,a31855a,a31859a,a31860a,a31863a,a31866a,a31867a,a31868a,a31872a,a31873a,a31877a,a31878a,a31879a,a31883a,a31884a,a31887a,a31890a,a31891a,a31892a,a31896a,a31897a,a31901a,a31902a,a31903a,a31907a,a31908a,a31911a,a31914a,a31915a,a31916a,a31920a,a31921a,a31925a,a31926a,a31927a,a31931a,a31932a,a31935a,a31938a,a31939a,a31940a,a31944a,a31945a,a31949a,a31950a,a31951a,a31955a,a31956a,a31959a,a31962a,a31963a,a31964a,a31968a,a31969a,a31973a,a31974a,a31975a,a31979a,a31980a,a31983a,a31986a,a31987a,a31988a,a31992a,a31993a,a31997a,a31998a,a31999a,a32003a,a32004a,a32007a,a32010a,a32011a,a32012a,a32016a,a32017a,a32021a,a32022a,a32023a,a32027a,a32028a,a32031a,a32034a,a32035a,a32036a,a32040a,a32041a,a32045a,a32046a,a32047a,a32051a,a32052a,a32055a,a32058a,a32059a,a32060a,a32064a,a32065a,a32069a,a32070a,a32071a,a32075a,a32076a,a32079a,a32082a,a32083a,a32084a,a32088a,a32089a,a32093a,a32094a,a32095a,a32099a,a32100a,a32103a,a32106a,a32107a,a32108a,a32112a,a32113a,a32117a,a32118a,a32119a,a32123a,a32124a,a32127a,a32130a,a32131a,a32132a,a32136a,a32137a,a32141a,a32142a,a32143a,a32147a,a32148a,a32151a,a32154a,a32155a,a32156a,a32160a,a32161a,a32165a,a32166a,a32167a,a32171a,a32172a,a32175a,a32178a,a32179a,a32180a,a32184a,a32185a,a32189a,a32190a,a32191a,a32195a,a32196a,a32199a,a32202a,a32203a,a32204a,a32208a,a32209a,a32213a,a32214a,a32215a,a32219a,a32220a,a32223a,a32226a,a32227a,a32228a,a32232a,a32233a,a32237a,a32238a,a32239a,a32243a,a32244a,a32247a,a32250a,a32251a,a32252a,a32256a,a32257a,a32261a,a32262a,a32263a,a32267a,a32268a,a32271a,a32274a,a32275a,a32276a,a32280a,a32281a,a32285a,a32286a,a32287a,a32291a,a32292a,a32295a,a32298a,a32299a,a32300a,a32304a,a32305a,a32309a,a32310a,a32311a,a32315a,a32316a,a32319a,a32322a,a32323a,a32324a,a32328a,a32329a,a32333a,a32334a,a32335a,a32339a,a32340a,a32343a,a32346a,a32347a,a32348a,a32352a,a32353a,a32357a,a32358a,a32359a,a32363a,a32364a,a32367a,a32370a,a32371a,a32372a,a32376a,a32377a,a32381a,a32382a,a32383a,a32387a,a32388a,a32391a,a32394a,a32395a,a32396a,a32400a,a32401a,a32405a,a32406a,a32407a,a32411a,a32412a,a32415a,a32418a,a32419a,a32420a,a32424a,a32425a,a32429a,a32430a,a32431a,a32435a,a32436a,a32439a,a32442a,a32443a,a32444a,a32448a,a32449a,a32453a,a32454a,a32455a,a32459a,a32460a,a32463a,a32466a,a32467a,a32468a,a32472a,a32473a,a32477a,a32478a,a32479a,a32483a,a32484a,a32487a,a32490a,a32491a,a32492a,a32496a,a32497a,a32501a,a32502a,a32503a,a32507a,a32508a,a32511a,a32514a,a32515a,a32516a,a32520a,a32521a,a32525a,a32526a,a32527a,a32531a,a32532a,a32535a,a32538a,a32539a,a32540a,a32544a,a32545a,a32549a,a32550a,a32551a,a32555a,a32556a,a32559a,a32562a,a32563a,a32564a,a32568a,a32569a,a32573a,a32574a,a32575a,a32579a,a32580a,a32583a,a32586a,a32587a,a32588a,a32592a,a32593a,a32597a,a32598a,a32599a,a32603a,a32604a,a32607a,a32610a,a32611a,a32612a,a32616a,a32617a,a32621a,a32622a,a32623a,a32627a,a32628a,a32631a,a32634a,a32635a,a32636a,a32640a,a32641a,a32645a,a32646a,a32647a,a32651a,a32652a,a32655a,a32658a,a32659a,a32660a,a32664a,a32665a,a32669a,a32670a,a32671a,a32675a,a32676a,a32679a,a32682a,a32683a,a32684a,a32688a,a32689a,a32693a,a32694a,a32695a,a32699a,a32700a,a32703a,a32706a,a32707a,a32708a,a32712a,a32713a,a32717a,a32718a,a32719a,a32723a,a32724a,a32727a,a32730a,a32731a,a32732a,a32736a,a32737a,a32741a,a32742a,a32743a,a32747a,a32748a,a32751a,a32754a,a32755a,a32756a,a32760a,a32761a,a32765a,a32766a,a32767a,a32771a,a32772a,a32775a,a32778a,a32779a,a32780a,a32784a,a32785a,a32789a,a32790a,a32791a,a32795a,a32796a,a32799a,a32802a,a32803a,a32804a,a32808a,a32809a,a32813a,a32814a,a32815a,a32819a,a32820a,a32823a,a32826a,a32827a,a32828a,a32832a,a32833a,a32837a,a32838a,a32839a,a32843a,a32844a,a32847a,a32850a,a32851a,a32852a,a32856a,a32857a,a32861a,a32862a,a32863a,a32867a,a32868a,a32871a,a32874a,a32875a,a32876a,a32880a,a32881a,a32885a,a32886a,a32887a,a32891a,a32892a,a32895a,a32898a,a32899a,a32900a,a32904a,a32905a,a32909a,a32910a,a32911a,a32915a,a32916a,a32919a,a32922a,a32923a,a32924a,a32928a,a32929a,a32933a,a32934a,a32935a,a32939a,a32940a,a32943a,a32946a,a32947a,a32948a,a32952a,a32953a,a32957a,a32958a,a32959a,a32963a,a32964a,a32967a,a32970a,a32971a,a32972a,a32976a,a32977a,a32981a,a32982a,a32983a,a32987a,a32988a,a32991a,a32994a,a32995a,a32996a,a33000a,a33001a,a33005a,a33006a,a33007a,a33011a,a33012a,a33015a,a33018a,a33019a,a33020a,a33024a,a33025a,a33029a,a33030a,a33031a,a33035a,a33036a,a33039a,a33042a,a33043a,a33044a,a33048a,a33049a,a33053a,a33054a,a33055a,a33059a,a33060a,a33063a,a33066a,a33067a,a33068a,a33072a,a33073a,a33077a,a33078a,a33079a,a33083a,a33084a,a33087a,a33090a,a33091a,a33092a,a33096a,a33097a,a33101a,a33102a,a33103a,a33107a,a33108a,a33111a,a33114a,a33115a,a33116a,a33120a,a33121a,a33125a,a33126a,a33127a,a33131a,a33132a,a33135a,a33138a,a33139a,a33140a,a33144a,a33145a,a33149a,a33150a,a33151a,a33155a,a33156a,a33159a,a33162a,a33163a,a33164a,a33168a,a33169a,a33173a,a33174a,a33175a,a33179a,a33180a,a33183a,a33186a,a33187a,a33188a,a33192a,a33193a,a33197a,a33198a,a33199a,a33203a,a33204a,a33207a,a33210a,a33211a,a33212a,a33216a,a33217a,a33221a,a33222a,a33223a,a33227a,a33228a,a33231a,a33234a,a33235a,a33236a,a33240a,a33241a,a33245a,a33246a,a33247a,a33251a,a33252a,a33255a,a33258a,a33259a,a33260a,a33264a,a33265a,a33269a,a33270a,a33271a,a33275a,a33276a,a33279a,a33282a,a33283a,a33284a,a33288a,a33289a,a33293a,a33294a,a33295a,a33299a,a33300a,a33303a,a33306a,a33307a,a33308a,a33312a,a33313a,a33317a,a33318a,a33319a,a33323a,a33324a,a33327a,a33330a,a33331a,a33332a,a33336a,a33337a,a33341a,a33342a,a33343a,a33347a,a33348a,a33351a,a33354a,a33355a,a33356a,a33360a,a33361a,a33365a,a33366a,a33367a,a33371a,a33372a,a33375a,a33378a,a33379a,a33380a,a33384a,a33385a,a33389a,a33390a,a33391a,a33395a,a33396a,a33399a,a33402a,a33403a,a33404a,a33408a,a33409a,a33413a,a33414a,a33415a,a33419a,a33420a,a33423a,a33426a,a33427a,a33428a,a33432a,a33433a,a33437a,a33438a,a33439a,a33443a,a33444a,a33447a,a33450a,a33451a,a33452a,a33456a,a33457a,a33461a,a33462a,a33463a,a33467a,a33468a,a33471a,a33474a,a33475a,a33476a,a33480a,a33481a,a33485a,a33486a,a33487a,a33491a,a33492a,a33495a,a33498a,a33499a,a33500a,a33504a,a33505a,a33509a,a33510a,a33511a,a33515a,a33516a,a33519a,a33522a,a33523a,a33524a,a33528a,a33529a,a33533a,a33534a,a33535a,a33539a,a33540a,a33543a,a33546a,a33547a,a33548a,a33552a,a33553a,a33557a,a33558a,a33559a,a33563a,a33564a,a33567a,a33570a,a33571a,a33572a,a33576a,a33577a,a33581a,a33582a,a33583a,a33587a,a33588a,a33591a,a33594a,a33595a,a33596a,a33600a,a33601a,a33605a,a33606a,a33607a,a33611a,a33612a,a33615a,a33618a,a33619a,a33620a,a33624a,a33625a,a33629a,a33630a,a33631a,a33635a,a33636a,a33639a,a33642a,a33643a,a33644a,a33648a,a33649a,a33653a,a33654a,a33655a,a33659a,a33660a,a33663a,a33666a,a33667a,a33668a,a33672a,a33673a,a33677a,a33678a,a33679a,a33683a,a33684a,a33687a,a33690a,a33691a,a33692a,a33696a,a33697a,a33701a,a33702a,a33703a,a33707a,a33708a,a33711a,a33714a,a33715a,a33716a,a33720a,a33721a,a33725a,a33726a,a33727a,a33731a,a33732a,a33735a,a33738a,a33739a,a33740a,a33744a,a33745a,a33749a,a33750a,a33751a,a33755a,a33756a,a33759a,a33762a,a33763a,a33764a,a33768a,a33769a,a33773a,a33774a,a33775a,a33779a,a33780a,a33783a,a33786a,a33787a,a33788a,a33792a,a33793a,a33797a,a33798a,a33799a,a33803a,a33804a,a33807a,a33810a,a33811a,a33812a,a33816a,a33817a,a33821a,a33822a,a33823a,a33827a,a33828a,a33831a,a33834a,a33835a,a33836a,a33840a,a33841a,a33845a,a33846a,a33847a,a33851a,a33852a,a33855a,a33858a,a33859a,a33860a,a33864a,a33865a,a33869a,a33870a,a33871a,a33875a,a33876a,a33879a,a33882a,a33883a,a33884a,a33888a,a33889a,a33893a,a33894a,a33895a,a33899a,a33900a,a33903a,a33906a,a33907a,a33908a,a33912a,a33913a,a33917a,a33918a,a33919a,a33923a,a33924a,a33927a,a33930a,a33931a,a33932a,a33936a,a33937a,a33941a,a33942a,a33943a,a33947a,a33948a,a33951a,a33954a,a33955a,a33956a,a33960a,a33961a,a33965a,a33966a,a33967a,a33971a,a33972a,a33975a,a33978a,a33979a,a33980a,a33984a,a33985a,a33989a,a33990a,a33991a,a33995a,a33996a,a33999a,a34002a,a34003a,a34004a,a34008a,a34009a,a34013a,a34014a,a34015a,a34019a,a34020a,a34023a,a34026a,a34027a,a34028a,a34032a,a34033a,a34037a,a34038a,a34039a,a34043a,a34044a,a34047a,a34050a,a34051a,a34052a,a34056a,a34057a,a34061a,a34062a,a34063a,a34067a,a34068a,a34071a,a34074a,a34075a,a34076a,a34080a,a34081a,a34085a,a34086a,a34087a,a34091a,a34092a,a34095a,a34098a,a34099a,a34100a,a34104a,a34105a,a34109a,a34110a,a34111a,a34115a,a34116a,a34119a,a34122a,a34123a,a34124a,a34128a,a34129a,a34133a,a34134a,a34135a,a34139a,a34140a,a34143a,a34146a,a34147a,a34148a,a34152a,a34153a,a34157a,a34158a,a34159a,a34163a,a34164a,a34167a,a34170a,a34171a,a34172a,a34176a,a34177a,a34181a,a34182a,a34183a,a34187a,a34188a,a34191a,a34194a,a34195a,a34196a,a34200a,a34201a,a34205a,a34206a,a34207a,a34211a,a34212a,a34215a,a34218a,a34219a,a34220a,a34224a,a34225a,a34229a,a34230a,a34231a,a34235a,a34236a,a34239a,a34242a,a34243a,a34244a,a34248a,a34249a,a34253a,a34254a,a34255a,a34259a,a34260a,a34263a,a34266a,a34267a,a34268a,a34272a,a34273a,a34277a,a34278a,a34279a,a34283a,a34284a,a34287a,a34290a,a34291a,a34292a,a34296a,a34297a,a34301a,a34302a,a34303a,a34307a,a34308a,a34311a,a34314a,a34315a,a34316a,a34320a,a34321a,a34325a,a34326a,a34327a,a34331a,a34332a,a34335a,a34338a,a34339a,a34340a,a34344a,a34345a,a34349a,a34350a,a34351a,a34355a,a34356a,a34359a,a34362a,a34363a,a34364a,a34368a,a34369a,a34373a,a34374a,a34375a,a34379a,a34380a,a34383a,a34386a,a34387a,a34388a,a34392a,a34393a,a34397a,a34398a,a34399a,a34403a,a34404a,a34407a,a34410a,a34411a,a34412a,a34416a,a34417a,a34421a,a34422a,a34423a,a34427a,a34428a,a34431a,a34434a,a34435a,a34436a,a34440a,a34441a,a34445a,a34446a,a34447a,a34451a,a34452a,a34455a,a34458a,a34459a,a34460a,a34464a,a34465a,a34469a,a34470a,a34471a,a34475a,a34476a,a34479a,a34482a,a34483a,a34484a,a34488a,a34489a,a34493a,a34494a,a34495a,a34499a,a34500a,a34503a,a34506a,a34507a,a34508a,a34512a,a34513a,a34517a,a34518a,a34519a,a34523a,a34524a,a34527a,a34530a,a34531a,a34532a,a34536a,a34537a,a34541a,a34542a,a34543a,a34547a,a34548a,a34551a,a34554a,a34555a,a34556a,a34560a,a34561a,a34565a,a34566a,a34567a,a34571a,a34572a,a34575a,a34578a,a34579a,a34580a,a34584a,a34585a,a34589a,a34590a,a34591a,a34595a,a34596a,a34599a,a34602a,a34603a,a34604a,a34608a,a34609a,a34613a,a34614a,a34615a,a34619a,a34620a,a34623a,a34626a,a34627a,a34628a,a34632a,a34633a,a34637a,a34638a,a34639a,a34643a,a34644a,a34647a,a34650a,a34651a,a34652a,a34656a,a34657a,a34661a,a34662a,a34663a,a34667a,a34668a,a34671a,a34674a,a34675a,a34676a,a34680a,a34681a,a34685a,a34686a,a34687a,a34691a,a34692a,a34695a,a34698a,a34699a,a34700a,a34704a,a34705a,a34709a,a34710a,a34711a,a34715a,a34716a,a34719a,a34722a,a34723a,a34724a,a34728a,a34729a,a34733a,a34734a,a34735a,a34739a,a34740a,a34743a,a34746a,a34747a,a34748a,a34752a,a34753a,a34757a,a34758a,a34759a,a34763a,a34764a,a34767a,a34770a,a34771a,a34772a,a34776a,a34777a,a34781a,a34782a,a34783a,a34787a,a34788a,a34791a,a34794a,a34795a,a34796a,a34800a,a34801a,a34805a,a34806a,a34807a,a34811a,a34812a,a34815a,a34818a,a34819a,a34820a,a34824a,a34825a,a34829a,a34830a,a34831a,a34835a,a34836a,a34839a,a34842a,a34843a,a34844a,a34848a,a34849a,a34853a,a34854a,a34855a,a34859a,a34860a,a34863a,a34866a,a34867a,a34868a,a34872a,a34873a,a34877a,a34878a,a34879a,a34883a,a34884a,a34887a,a34890a,a34891a,a34892a,a34896a,a34897a,a34901a,a34902a,a34903a,a34907a,a34908a,a34911a,a34914a,a34915a,a34916a,a34920a,a34921a,a34925a,a34926a,a34927a,a34931a,a34932a,a34935a,a34938a,a34939a,a34940a,a34944a,a34945a,a34949a,a34950a,a34951a,a34955a,a34956a,a34959a,a34962a,a34963a,a34964a,a34968a,a34969a,a34973a,a34974a,a34975a,a34979a,a34980a,a34983a,a34986a,a34987a,a34988a,a34992a,a34993a,a34997a,a34998a,a34999a,a35003a,a35004a,a35007a,a35010a,a35011a,a35012a,a35016a,a35017a,a35021a,a35022a,a35023a,a35027a,a35028a,a35031a,a35034a,a35035a,a35036a,a35040a,a35041a,a35045a,a35046a,a35047a,a35051a,a35052a,a35055a,a35058a,a35059a,a35060a,a35064a,a35065a,a35069a,a35070a,a35071a,a35075a,a35076a,a35079a,a35082a,a35083a,a35084a,a35088a,a35089a,a35093a,a35094a,a35095a,a35099a,a35100a,a35103a,a35106a,a35107a,a35108a,a35112a,a35113a,a35117a,a35118a,a35119a,a35123a,a35124a,a35127a,a35130a,a35131a,a35132a,a35136a,a35137a,a35141a,a35142a,a35143a,a35147a,a35148a,a35151a,a35154a,a35155a,a35156a,a35160a,a35161a,a35165a,a35166a,a35167a,a35171a,a35172a,a35175a,a35178a,a35179a,a35180a,a35184a,a35185a,a35189a,a35190a,a35191a,a35195a,a35196a,a35199a,a35202a,a35203a,a35204a,a35208a,a35209a,a35213a,a35214a,a35215a,a35219a,a35220a,a35223a,a35226a,a35227a,a35228a,a35232a,a35233a,a35237a,a35238a,a35239a,a35243a,a35244a,a35247a,a35250a,a35251a,a35252a,a35256a,a35257a,a35261a,a35262a,a35263a,a35267a,a35268a,a35271a,a35274a,a35275a,a35276a,a35280a,a35281a,a35285a,a35286a,a35287a,a35291a,a35292a,a35295a,a35298a,a35299a,a35300a,a35304a,a35305a,a35309a,a35310a,a35311a,a35315a,a35316a,a35319a,a35322a,a35323a,a35324a,a35328a,a35329a,a35333a,a35334a,a35335a,a35339a,a35340a,a35343a,a35346a,a35347a,a35348a,a35352a,a35353a,a35357a,a35358a,a35359a,a35363a,a35364a,a35367a,a35370a,a35371a,a35372a,a35376a,a35377a,a35381a,a35382a,a35383a,a35387a,a35388a,a35391a,a35394a,a35395a,a35396a,a35400a,a35401a,a35405a,a35406a,a35407a,a35411a,a35412a,a35415a,a35418a,a35419a,a35420a,a35424a,a35425a,a35429a,a35430a,a35431a,a35435a,a35436a,a35439a,a35442a,a35443a,a35444a,a35448a,a35449a,a35453a,a35454a,a35455a,a35459a,a35460a,a35463a,a35466a,a35467a,a35468a,a35472a,a35473a,a35477a,a35478a,a35479a,a35483a,a35484a,a35487a,a35490a,a35491a,a35492a,a35496a,a35497a,a35501a,a35502a,a35503a,a35507a,a35508a,a35511a,a35514a,a35515a,a35516a,a35520a,a35521a,a35525a,a35526a,a35527a,a35531a,a35532a,a35535a,a35538a,a35539a,a35540a,a35544a,a35545a,a35549a,a35550a,a35551a,a35555a,a35556a,a35559a,a35562a,a35563a,a35564a,a35568a,a35569a,a35573a,a35574a,a35575a,a35579a,a35580a,a35583a,a35586a,a35587a,a35588a,a35592a,a35593a,a35597a,a35598a,a35599a,a35603a,a35604a,a35607a,a35610a,a35611a,a35612a,a35616a,a35617a,a35621a,a35622a,a35623a,a35627a,a35628a,a35631a,a35634a,a35635a,a35636a,a35640a,a35641a,a35645a,a35646a,a35647a,a35651a,a35652a,a35655a,a35658a,a35659a,a35660a,a35664a,a35665a,a35669a,a35670a,a35671a,a35675a,a35676a,a35679a,a35682a,a35683a,a35684a,a35688a,a35689a,a35693a,a35694a,a35695a,a35699a,a35700a,a35703a,a35706a,a35707a,a35708a,a35712a,a35713a,a35717a,a35718a,a35719a,a35723a,a35724a,a35727a,a35730a,a35731a,a35732a,a35736a,a35737a,a35741a,a35742a,a35743a,a35747a,a35748a,a35751a,a35754a,a35755a,a35756a,a35760a,a35761a,a35765a,a35766a,a35767a,a35771a,a35772a,a35775a,a35778a,a35779a,a35780a,a35784a,a35785a,a35789a,a35790a,a35791a,a35795a,a35796a,a35799a,a35802a,a35803a,a35804a,a35808a,a35809a,a35813a,a35814a,a35815a,a35819a,a35820a,a35823a,a35826a,a35827a,a35828a,a35832a,a35833a,a35837a,a35838a,a35839a,a35843a,a35844a,a35847a,a35850a,a35851a,a35852a,a35856a,a35857a,a35861a,a35862a,a35863a,a35867a,a35868a,a35871a,a35874a,a35875a,a35876a,a35880a,a35881a,a35885a,a35886a,a35887a,a35891a,a35892a,a35895a,a35898a,a35899a,a35900a,a35904a,a35905a,a35909a,a35910a,a35911a,a35915a,a35916a,a35919a,a35922a,a35923a,a35924a,a35928a,a35929a,a35933a,a35934a,a35935a,a35939a,a35940a,a35943a,a35946a,a35947a,a35948a,a35952a,a35953a,a35957a,a35958a,a35959a,a35963a,a35964a,a35967a,a35970a,a35971a,a35972a,a35976a,a35977a,a35981a,a35982a,a35983a,a35987a,a35988a,a35991a,a35994a,a35995a,a35996a,a36000a,a36001a,a36005a,a36006a,a36007a,a36011a,a36012a,a36015a,a36018a,a36019a,a36020a,a36024a,a36025a,a36029a,a36030a,a36031a,a36035a,a36036a,a36039a,a36042a,a36043a,a36044a,a36048a,a36049a,a36053a,a36054a,a36055a,a36059a,a36060a,a36063a,a36066a,a36067a,a36068a,a36072a,a36073a,a36077a,a36078a,a36079a,a36083a,a36084a,a36087a,a36090a,a36091a,a36092a,a36096a,a36097a,a36101a,a36102a,a36103a,a36107a,a36108a,a36111a,a36114a,a36115a,a36116a,a36120a,a36121a,a36125a,a36126a,a36127a,a36131a,a36132a,a36135a,a36138a,a36139a,a36140a,a36144a,a36145a,a36149a,a36150a,a36151a,a36155a,a36156a,a36159a,a36162a,a36163a,a36164a,a36168a,a36169a,a36173a,a36174a,a36175a,a36179a,a36180a,a36183a,a36186a,a36187a,a36188a,a36192a,a36193a,a36197a,a36198a,a36199a,a36203a,a36204a,a36207a,a36210a,a36211a,a36212a,a36216a,a36217a,a36221a,a36222a,a36223a,a36227a,a36228a,a36231a,a36234a,a36235a,a36236a,a36240a,a36241a,a36245a,a36246a,a36247a,a36251a,a36252a,a36255a,a36258a,a36259a,a36260a,a36264a,a36265a,a36269a,a36270a,a36271a,a36275a,a36276a,a36279a,a36282a,a36283a,a36284a,a36288a,a36289a,a36293a,a36294a,a36295a,a36299a,a36300a,a36303a,a36306a,a36307a,a36308a,a36312a,a36313a,a36317a,a36318a,a36319a,a36323a,a36324a,a36327a,a36330a,a36331a,a36332a,a36336a,a36337a,a36341a,a36342a,a36343a,a36347a,a36348a,a36351a,a36354a,a36355a,a36356a,a36360a,a36361a,a36365a,a36366a,a36367a,a36371a,a36372a,a36375a,a36378a,a36379a,a36380a,a36384a,a36385a,a36389a,a36390a,a36391a,a36395a,a36396a,a36399a,a36402a,a36403a,a36404a,a36408a,a36409a,a36413a,a36414a,a36415a,a36419a,a36420a,a36423a,a36426a,a36427a,a36428a,a36432a,a36433a,a36437a,a36438a,a36439a,a36443a,a36444a,a36447a,a36450a,a36451a,a36452a,a36456a,a36457a,a36461a,a36462a,a36463a,a36467a,a36468a,a36471a,a36474a,a36475a,a36476a,a36480a,a36481a,a36485a,a36486a,a36487a,a36491a,a36492a,a36495a,a36498a,a36499a,a36500a,a36504a,a36505a,a36509a,a36510a,a36511a,a36515a,a36516a,a36519a,a36522a,a36523a,a36524a,a36528a,a36529a,a36533a,a36534a,a36535a,a36539a,a36540a,a36543a,a36546a,a36547a,a36548a,a36552a,a36553a,a36557a,a36558a,a36559a,a36563a,a36564a,a36567a,a36570a,a36571a,a36572a,a36576a,a36577a,a36581a,a36582a,a36583a,a36587a,a36588a,a36591a,a36594a,a36595a,a36596a,a36600a,a36601a,a36605a,a36606a,a36607a,a36611a,a36612a,a36615a,a36618a,a36619a,a36620a,a36624a,a36625a,a36629a,a36630a,a36631a,a36635a,a36636a,a36639a,a36642a,a36643a,a36644a,a36648a,a36649a,a36653a,a36654a,a36655a,a36659a,a36660a,a36663a,a36666a,a36667a,a36668a,a36672a,a36673a,a36677a,a36678a,a36679a,a36683a,a36684a,a36687a,a36690a,a36691a,a36692a,a36696a,a36697a,a36701a,a36702a,a36703a,a36707a,a36708a,a36711a,a36714a,a36715a,a36716a,a36720a,a36721a,a36725a,a36726a,a36727a,a36731a,a36732a,a36735a,a36738a,a36739a,a36740a,a36744a,a36745a,a36749a,a36750a,a36751a,a36755a,a36756a,a36759a,a36762a,a36763a,a36764a,a36768a,a36769a,a36773a,a36774a,a36775a,a36779a,a36780a,a36783a,a36786a,a36787a,a36788a,a36792a,a36793a,a36797a,a36798a,a36799a,a36803a,a36804a,a36807a,a36810a,a36811a,a36812a,a36816a,a36817a,a36821a,a36822a,a36823a,a36827a,a36828a,a36831a,a36834a,a36835a,a36836a,a36840a,a36841a,a36845a,a36846a,a36847a,a36851a,a36852a,a36855a,a36858a,a36859a,a36860a,a36864a,a36865a,a36869a,a36870a,a36871a,a36875a,a36876a,a36879a,a36882a,a36883a,a36884a,a36888a,a36889a,a36893a,a36894a,a36895a,a36899a,a36900a,a36903a,a36906a,a36907a,a36908a,a36912a,a36913a,a36917a,a36918a,a36919a,a36923a,a36924a,a36927a,a36930a,a36931a,a36932a,a36936a,a36937a,a36941a,a36942a,a36943a,a36947a,a36948a,a36951a,a36954a,a36955a,a36956a,a36960a,a36961a,a36965a,a36966a,a36967a,a36971a,a36972a,a36975a,a36978a,a36979a,a36980a,a36984a,a36985a,a36989a,a36990a,a36991a,a36995a,a36996a,a36999a,a37002a,a37003a,a37004a,a37008a,a37009a,a37013a,a37014a,a37015a,a37019a,a37020a,a37023a,a37026a,a37027a,a37028a,a37032a,a37033a,a37037a,a37038a,a37039a,a37043a,a37044a,a37047a,a37050a,a37051a,a37052a,a37056a,a37057a,a37061a,a37062a,a37063a,a37067a,a37068a,a37071a,a37074a,a37075a,a37076a,a37080a,a37081a,a37085a,a37086a,a37087a,a37091a,a37092a,a37095a,a37098a,a37099a,a37100a,a37104a,a37105a,a37109a,a37110a,a37111a,a37115a,a37116a,a37119a,a37122a,a37123a,a37124a,a37128a,a37129a,a37133a,a37134a,a37135a,a37139a,a37140a,a37143a,a37146a,a37147a,a37148a,a37152a,a37153a,a37157a,a37158a,a37159a,a37163a,a37164a,a37167a,a37170a,a37171a,a37172a,a37176a,a37177a,a37181a,a37182a,a37183a,a37187a,a37188a,a37191a,a37194a,a37195a,a37196a,a37200a,a37201a,a37205a,a37206a,a37207a,a37211a,a37212a,a37215a,a37218a,a37219a,a37220a,a37224a,a37225a,a37229a,a37230a,a37231a,a37235a,a37236a,a37239a,a37242a,a37243a,a37244a,a37248a,a37249a,a37253a,a37254a,a37255a,a37259a,a37260a,a37263a,a37266a,a37267a,a37268a,a37272a,a37273a,a37277a,a37278a,a37279a,a37283a,a37284a,a37287a,a37290a,a37291a,a37292a,a37296a,a37297a,a37301a,a37302a,a37303a,a37307a,a37308a,a37311a,a37314a,a37315a,a37316a,a37320a,a37321a,a37325a,a37326a,a37327a,a37331a,a37332a,a37335a,a37338a,a37339a,a37340a,a37344a,a37345a,a37349a,a37350a,a37351a,a37355a,a37356a,a37359a,a37362a,a37363a,a37364a,a37368a,a37369a,a37373a,a37374a,a37375a,a37379a,a37380a,a37383a,a37386a,a37387a,a37388a,a37392a,a37393a,a37397a,a37398a,a37399a,a37403a,a37404a,a37407a,a37410a,a37411a,a37412a,a37416a,a37417a,a37421a,a37422a,a37423a,a37427a,a37428a,a37431a,a37434a,a37435a,a37436a,a37440a,a37441a,a37445a,a37446a,a37447a,a37451a,a37452a,a37455a,a37458a,a37459a,a37460a,a37464a,a37465a,a37469a,a37470a,a37471a,a37475a,a37476a,a37479a,a37482a,a37483a,a37484a,a37488a,a37489a,a37493a,a37494a,a37495a,a37499a,a37500a,a37503a,a37506a,a37507a,a37508a,a37512a,a37513a,a37517a,a37518a,a37519a,a37523a,a37524a,a37527a,a37530a,a37531a,a37532a,a37536a,a37537a,a37541a,a37542a,a37543a,a37547a,a37548a,a37551a,a37554a,a37555a,a37556a,a37560a,a37561a,a37565a,a37566a,a37567a,a37571a,a37572a,a37575a,a37578a,a37579a,a37580a,a37584a,a37585a,a37589a,a37590a,a37591a,a37595a,a37596a,a37599a,a37602a,a37603a,a37604a,a37608a,a37609a,a37613a,a37614a,a37615a,a37619a,a37620a,a37623a,a37626a,a37627a,a37628a,a37632a,a37633a,a37637a,a37638a,a37639a,a37643a,a37644a,a37647a,a37650a,a37651a,a37652a,a37656a,a37657a,a37661a,a37662a,a37663a,a37667a,a37668a,a37671a,a37674a,a37675a,a37676a,a37680a,a37681a,a37685a,a37686a,a37687a,a37691a,a37692a,a37695a,a37698a,a37699a,a37700a,a37704a,a37705a,a37709a,a37710a,a37711a,a37715a,a37716a,a37719a,a37722a,a37723a,a37724a,a37728a,a37729a,a37733a,a37734a,a37735a,a37739a,a37740a,a37743a,a37746a,a37747a,a37748a,a37752a,a37753a,a37757a,a37758a,a37759a,a37763a,a37764a,a37767a,a37770a,a37771a,a37772a,a37776a,a37777a,a37781a,a37782a,a37783a,a37787a,a37788a,a37791a,a37794a,a37795a,a37796a,a37800a,a37801a,a37805a,a37806a,a37807a,a37811a,a37812a,a37815a,a37818a,a37819a,a37820a,a37824a,a37825a,a37828a,a37831a,a37832a,a37833a,a37837a,a37838a,a37841a,a37844a,a37845a,a37846a,a37850a,a37851a,a37854a,a37857a,a37858a,a37859a,a37863a,a37864a,a37867a,a37870a,a37871a,a37872a,a37876a,a37877a,a37880a,a37883a,a37884a,a37885a,a37889a,a37890a,a37893a,a37896a,a37897a,a37898a,a37902a,a37903a,a37906a,a37909a,a37910a,a37911a,a37915a,a37916a,a37919a,a37922a,a37923a,a37924a,a37928a,a37929a,a37932a,a37935a,a37936a,a37937a,a37941a,a37942a,a37945a,a37948a,a37949a,a37950a,a37954a,a37955a,a37958a,a37961a,a37962a,a37963a,a37967a,a37968a,a37971a,a37974a,a37975a,a37976a,a37980a,a37981a,a37984a,a37987a,a37988a,a37989a,a37993a,a37994a,a37997a,a38000a,a38001a,a38002a,a38006a,a38007a,a38010a,a38013a,a38014a,a38015a,a38019a,a38020a,a38023a,a38026a,a38027a,a38028a,a38032a,a38033a,a38036a,a38039a,a38040a,a38041a,a38045a,a38046a,a38049a,a38052a,a38053a,a38054a,a38058a,a38059a,a38062a,a38065a,a38066a,a38067a,a38071a,a38072a,a38075a,a38078a,a38079a,a38080a,a38084a,a38085a,a38088a,a38091a,a38092a,a38093a,a38097a,a38098a,a38101a,a38104a,a38105a,a38106a,a38110a,a38111a,a38114a,a38117a,a38118a,a38119a,a38123a,a38124a,a38127a,a38130a,a38131a,a38132a,a38136a,a38137a,a38140a,a38143a,a38144a,a38145a,a38149a,a38150a,a38153a,a38156a,a38157a,a38158a,a38162a,a38163a,a38166a,a38169a,a38170a,a38171a,a38175a,a38176a,a38179a,a38182a,a38183a,a38184a,a38188a,a38189a,a38192a,a38195a,a38196a,a38197a,a38201a,a38202a,a38205a,a38208a,a38209a,a38210a,a38214a,a38215a,a38218a,a38221a,a38222a,a38223a,a38227a,a38228a,a38231a,a38234a,a38235a,a38236a,a38240a,a38241a,a38244a,a38247a,a38248a,a38249a,a38253a,a38254a,a38257a,a38260a,a38261a,a38262a,a38266a,a38267a,a38270a,a38273a,a38274a,a38275a,a38279a,a38280a,a38283a,a38286a,a38287a,a38288a,a38292a,a38293a,a38296a,a38299a,a38300a,a38301a,a38305a,a38306a,a38309a,a38312a,a38313a,a38314a,a38318a,a38319a,a38322a,a38325a,a38326a,a38327a,a38331a,a38332a,a38335a,a38338a,a38339a,a38340a,a38344a,a38345a,a38348a,a38351a,a38352a,a38353a,a38357a,a38358a,a38361a,a38364a,a38365a,a38366a,a38370a,a38371a,a38374a,a38377a,a38378a,a38379a,a38383a,a38384a,a38387a,a38390a,a38391a,a38392a,a38396a,a38397a,a38400a,a38403a,a38404a,a38405a,a38409a,a38410a,a38413a,a38416a,a38417a,a38418a,a38422a,a38423a,a38426a,a38429a,a38430a,a38431a,a38435a,a38436a,a38439a,a38442a,a38443a,a38444a,a38448a,a38449a,a38452a,a38455a,a38456a,a38457a,a38461a,a38462a,a38465a,a38468a,a38469a,a38470a,a38474a,a38475a,a38478a,a38481a,a38482a,a38483a,a38487a,a38488a,a38491a,a38494a,a38495a,a38496a,a38500a,a38501a,a38504a,a38507a,a38508a,a38509a,a38513a,a38514a,a38517a,a38520a,a38521a,a38522a,a38526a,a38527a,a38530a,a38533a,a38534a,a38535a,a38539a,a38540a,a38543a,a38546a,a38547a,a38548a,a38552a,a38553a,a38556a,a38559a,a38560a,a38561a,a38565a,a38566a,a38569a,a38572a,a38573a,a38574a,a38578a,a38579a,a38582a,a38585a,a38586a,a38587a,a38591a,a38592a,a38595a,a38598a,a38599a,a38600a,a38604a,a38605a,a38608a,a38611a,a38612a,a38613a,a38617a,a38618a,a38621a,a38624a,a38625a,a38626a,a38630a,a38631a,a38634a,a38637a,a38638a,a38639a,a38643a,a38644a,a38647a,a38650a,a38651a,a38652a,a38656a,a38657a,a38660a,a38663a,a38664a,a38665a,a38669a,a38670a,a38673a,a38676a,a38677a,a38678a,a38682a,a38683a,a38686a,a38689a,a38690a,a38691a,a38695a,a38696a,a38699a,a38702a,a38703a,a38704a,a38708a,a38709a,a38712a,a38715a,a38716a,a38717a,a38721a,a38722a,a38725a,a38728a,a38729a,a38730a,a38734a,a38735a,a38738a,a38741a,a38742a,a38743a,a38747a,a38748a,a38751a,a38754a,a38755a,a38756a,a38760a,a38761a,a38764a,a38767a,a38768a,a38769a,a38773a,a38774a,a38777a,a38780a,a38781a,a38782a,a38786a,a38787a,a38790a,a38793a,a38794a,a38795a,a38799a,a38800a,a38803a,a38806a,a38807a,a38808a,a38812a,a38813a,a38816a,a38819a,a38820a,a38821a,a38825a,a38826a,a38829a,a38832a,a38833a,a38834a,a38838a,a38839a,a38842a,a38845a,a38846a,a38847a,a38851a,a38852a,a38855a,a38858a,a38859a,a38860a,a38864a,a38865a,a38868a,a38871a,a38872a,a38873a,a38877a,a38878a,a38881a,a38884a,a38885a,a38886a,a38890a,a38891a,a38894a,a38897a,a38898a,a38899a,a38903a,a38904a,a38907a,a38910a,a38911a,a38912a,a38916a,a38917a,a38920a,a38923a,a38924a,a38925a,a38929a,a38930a,a38933a,a38936a,a38937a,a38938a,a38942a,a38943a,a38946a,a38949a,a38950a,a38951a,a38955a,a38956a,a38959a,a38962a,a38963a,a38964a,a38968a,a38969a,a38972a,a38975a,a38976a,a38977a,a38981a,a38982a,a38985a,a38988a,a38989a,a38990a,a38994a,a38995a,a38998a,a39001a,a39002a,a39003a,a39007a,a39008a,a39011a,a39014a,a39015a,a39016a,a39020a,a39021a,a39024a,a39027a,a39028a,a39029a,a39033a,a39034a,a39037a,a39040a,a39041a,a39042a,a39046a,a39047a,a39050a,a39053a,a39054a,a39055a,a39059a,a39060a,a39063a,a39066a,a39067a,a39068a,a39072a,a39073a,a39076a,a39079a,a39080a,a39081a,a39085a,a39086a,a39089a,a39092a,a39093a,a39094a,a39098a,a39099a,a39102a,a39105a,a39106a,a39107a,a39111a,a39112a,a39115a,a39118a,a39119a,a39120a,a39124a,a39125a,a39128a,a39131a,a39132a,a39133a,a39137a,a39138a,a39141a,a39144a,a39145a,a39146a,a39150a,a39151a,a39154a,a39157a,a39158a,a39159a,a39163a,a39164a,a39167a,a39170a,a39171a,a39172a,a39176a,a39177a,a39180a,a39183a,a39184a,a39185a,a39189a,a39190a,a39193a,a39196a,a39197a,a39198a,a39202a,a39203a,a39206a,a39209a,a39210a,a39211a,a39215a,a39216a,a39219a,a39222a,a39223a,a39224a,a39228a,a39229a,a39232a,a39235a,a39236a,a39237a,a39241a,a39242a,a39245a,a39248a,a39249a,a39250a,a39254a,a39255a,a39258a,a39261a,a39262a,a39263a,a39267a,a39268a,a39271a,a39274a,a39275a,a39276a,a39280a,a39281a,a39284a,a39287a,a39288a,a39289a,a39293a,a39294a,a39297a,a39300a,a39301a,a39302a,a39306a,a39307a,a39310a,a39313a,a39314a,a39315a,a39319a,a39320a,a39323a,a39326a,a39327a,a39328a,a39332a,a39333a,a39336a,a39339a,a39340a,a39341a,a39345a,a39346a,a39349a,a39352a,a39353a,a39354a,a39358a,a39359a,a39362a,a39365a,a39366a,a39367a,a39371a,a39372a,a39375a,a39378a,a39379a,a39380a,a39384a,a39385a,a39388a,a39391a,a39392a,a39393a,a39397a,a39398a,a39401a,a39404a,a39405a,a39406a,a39410a,a39411a,a39414a,a39417a,a39418a,a39419a,a39423a,a39424a,a39427a,a39430a,a39431a,a39432a,a39436a,a39437a,a39440a,a39443a,a39444a,a39445a,a39449a,a39450a,a39453a,a39456a,a39457a,a39458a,a39462a,a39463a,a39466a,a39469a,a39470a,a39471a,a39475a,a39476a,a39479a,a39482a,a39483a,a39484a,a39488a,a39489a,a39492a,a39495a,a39496a,a39497a,a39501a,a39502a,a39505a,a39508a,a39509a,a39510a,a39514a,a39515a,a39518a,a39521a,a39522a,a39523a,a39527a,a39528a,a39531a,a39534a,a39535a,a39536a,a39540a,a39541a,a39544a,a39547a,a39548a,a39549a,a39553a,a39554a,a39557a,a39560a,a39561a,a39562a,a39566a,a39567a,a39570a,a39573a,a39574a,a39575a,a39579a,a39580a,a39583a,a39586a,a39587a,a39588a,a39592a,a39593a,a39596a,a39599a,a39600a,a39601a,a39605a,a39606a,a39609a,a39612a,a39613a,a39614a,a39618a,a39619a,a39622a,a39625a,a39626a,a39627a,a39631a,a39632a,a39635a,a39638a,a39639a,a39640a,a39644a,a39645a,a39648a,a39651a,a39652a,a39653a,a39657a,a39658a,a39661a,a39664a,a39665a,a39666a,a39670a,a39671a,a39674a,a39677a,a39678a,a39679a,a39683a,a39684a,a39687a,a39690a,a39691a,a39692a,a39696a,a39697a,a39700a,a39703a,a39704a,a39705a,a39709a,a39710a,a39713a,a39716a,a39717a,a39718a,a39722a,a39723a,a39726a,a39729a,a39730a,a39731a,a39735a,a39736a,a39739a,a39742a,a39743a,a39744a,a39748a,a39749a,a39752a,a39755a,a39756a,a39757a,a39761a,a39762a,a39765a,a39768a,a39769a,a39770a,a39774a,a39775a,a39778a,a39781a,a39782a,a39783a,a39787a,a39788a,a39791a,a39794a,a39795a,a39796a,a39800a,a39801a,a39804a,a39807a,a39808a,a39809a,a39813a,a39814a,a39817a,a39820a,a39821a,a39822a,a39826a,a39827a,a39830a,a39833a,a39834a,a39835a,a39839a,a39840a,a39843a,a39846a,a39847a,a39848a,a39852a,a39853a,a39856a,a39859a,a39860a,a39861a,a39865a,a39866a,a39869a,a39872a,a39873a,a39874a,a39878a,a39879a,a39882a,a39885a,a39886a,a39887a,a39891a,a39892a,a39895a,a39898a,a39899a,a39900a,a39904a,a39905a,a39908a,a39911a,a39912a,a39913a,a39917a,a39918a,a39921a,a39924a,a39925a,a39926a,a39930a,a39931a,a39934a,a39937a,a39938a,a39939a,a39943a,a39944a,a39947a,a39950a,a39951a,a39952a,a39956a,a39957a,a39960a,a39963a,a39964a,a39965a,a39969a,a39970a,a39973a,a39976a,a39977a,a39978a,a39982a,a39983a,a39986a,a39989a,a39990a,a39991a,a39995a,a39996a,a39999a,a40002a,a40003a,a40004a,a40008a,a40009a,a40012a,a40015a,a40016a,a40017a,a40021a,a40022a,a40025a,a40028a,a40029a,a40030a,a40034a,a40035a,a40038a,a40041a,a40042a,a40043a,a40047a,a40048a,a40051a,a40054a,a40055a,a40056a,a40060a,a40061a,a40064a,a40067a,a40068a,a40069a,a40073a,a40074a,a40077a,a40080a,a40081a,a40082a,a40086a,a40087a,a40090a,a40093a,a40094a,a40095a,a40099a,a40100a,a40103a,a40106a,a40107a,a40108a,a40112a,a40113a,a40116a,a40119a,a40120a,a40121a,a40125a,a40126a,a40129a,a40132a,a40133a,a40134a,a40138a,a40139a,a40142a,a40145a,a40146a,a40147a,a40151a,a40152a,a40155a,a40158a,a40159a,a40160a,a40164a,a40165a,a40168a,a40171a,a40172a,a40173a,a40177a,a40178a,a40181a,a40184a,a40185a,a40186a,a40190a,a40191a,a40194a,a40197a,a40198a,a40199a,a40203a,a40204a,a40207a,a40210a,a40211a,a40212a,a40216a,a40217a,a40220a,a40223a,a40224a,a40225a,a40229a,a40230a,a40233a,a40236a,a40237a,a40238a,a40242a,a40243a,a40246a,a40249a,a40250a,a40251a,a40255a,a40256a,a40259a,a40262a,a40263a,a40264a,a40268a,a40269a,a40272a,a40275a,a40276a,a40277a,a40281a,a40282a,a40285a,a40288a,a40289a,a40290a,a40294a,a40295a,a40298a,a40301a,a40302a,a40303a,a40307a,a40308a,a40311a,a40314a,a40315a,a40316a,a40320a,a40321a,a40324a,a40327a,a40328a,a40329a,a40333a,a40334a,a40337a,a40340a,a40341a,a40342a,a40346a,a40347a,a40350a,a40353a,a40354a,a40355a,a40359a,a40360a,a40363a,a40366a,a40367a,a40368a,a40372a,a40373a,a40376a,a40379a,a40380a,a40381a,a40385a,a40386a,a40389a,a40392a,a40393a,a40394a,a40398a,a40399a,a40402a,a40405a,a40406a,a40407a,a40411a,a40412a,a40415a,a40418a,a40419a,a40420a,a40424a,a40425a,a40428a,a40431a,a40432a,a40433a,a40437a,a40438a,a40441a,a40444a,a40445a,a40446a,a40450a,a40451a,a40454a,a40457a,a40458a,a40459a,a40463a,a40464a,a40467a,a40470a,a40471a,a40472a,a40476a,a40477a,a40480a,a40483a,a40484a,a40485a,a40489a,a40490a,a40493a,a40496a,a40497a,a40498a,a40502a,a40503a,a40506a,a40509a,a40510a,a40511a,a40515a,a40516a,a40519a,a40522a,a40523a,a40524a,a40528a,a40529a,a40532a,a40535a,a40536a,a40537a,a40541a,a40542a,a40545a,a40548a,a40549a,a40550a,a40554a,a40555a,a40558a,a40561a,a40562a,a40563a,a40567a,a40568a,a40571a,a40574a,a40575a,a40576a,a40580a,a40581a,a40584a,a40587a,a40588a,a40589a,a40593a,a40594a,a40597a,a40600a,a40601a,a40602a,a40606a,a40607a,a40610a,a40613a,a40614a,a40615a,a40619a,a40620a,a40623a,a40626a,a40627a,a40628a,a40632a,a40633a,a40636a,a40639a,a40640a,a40641a,a40645a,a40646a,a40649a,a40652a,a40653a,a40654a,a40658a,a40659a,a40662a,a40665a,a40666a,a40667a,a40671a,a40672a,a40675a,a40678a,a40679a,a40680a,a40684a,a40685a,a40688a,a40691a,a40692a,a40693a,a40697a,a40698a,a40701a,a40704a,a40705a,a40706a,a40710a,a40711a,a40714a,a40717a,a40718a,a40719a,a40723a,a40724a,a40727a,a40730a,a40731a,a40732a,a40736a,a40737a,a40740a,a40743a,a40744a,a40745a,a40749a,a40750a,a40753a,a40756a,a40757a,a40758a,a40762a,a40763a,a40766a,a40769a,a40770a,a40771a,a40775a,a40776a,a40779a,a40782a,a40783a,a40784a,a40788a,a40789a,a40792a,a40795a,a40796a,a40797a,a40801a,a40802a,a40805a,a40808a,a40809a,a40810a,a40814a,a40815a,a40818a,a40821a,a40822a,a40823a,a40827a,a40828a,a40831a,a40834a,a40835a,a40836a,a40840a,a40841a,a40844a,a40847a,a40848a,a40849a,a40853a,a40854a,a40857a,a40860a,a40861a,a40862a,a40866a,a40867a,a40870a,a40873a,a40874a,a40875a,a40879a,a40880a,a40883a,a40886a,a40887a,a40888a,a40892a,a40893a,a40896a,a40899a,a40900a,a40901a,a40905a,a40906a,a40909a,a40912a,a40913a,a40914a,a40918a,a40919a,a40922a,a40925a,a40926a,a40927a,a40931a,a40932a,a40935a,a40938a,a40939a,a40940a,a40944a,a40945a,a40948a,a40951a,a40952a,a40953a,a40957a,a40958a,a40961a,a40964a,a40965a,a40966a,a40970a,a40971a,a40974a,a40977a,a40978a,a40979a,a40983a,a40984a,a40987a,a40990a,a40991a,a40992a,a40996a,a40997a,a41000a,a41003a,a41004a,a41005a,a41009a,a41010a,a41013a,a41016a,a41017a,a41018a,a41022a,a41023a,a41026a,a41029a,a41030a,a41031a,a41035a,a41036a,a41039a,a41042a,a41043a,a41044a,a41048a,a41049a,a41052a,a41055a,a41056a,a41057a,a41061a,a41062a,a41065a,a41068a,a41069a,a41070a,a41074a,a41075a,a41078a,a41081a,a41082a,a41083a,a41087a,a41088a,a41091a,a41094a,a41095a,a41096a,a41100a,a41101a,a41104a,a41107a,a41108a,a41109a,a41113a,a41114a,a41117a,a41120a,a41121a,a41122a,a41126a,a41127a,a41130a,a41133a,a41134a,a41135a,a41139a,a41140a,a41143a,a41146a,a41147a,a41148a,a41152a,a41153a,a41156a,a41159a,a41160a,a41161a,a41165a,a41166a,a41169a,a41172a,a41173a,a41174a,a41178a,a41179a,a41182a,a41185a,a41186a,a41187a,a41191a,a41192a,a41195a,a41198a,a41199a,a41200a,a41204a,a41205a,a41208a,a41211a,a41212a,a41213a,a41217a,a41218a,a41221a,a41224a,a41225a,a41226a,a41230a,a41231a,a41234a,a41237a,a41238a,a41239a,a41243a,a41244a,a41247a,a41250a,a41251a,a41252a,a41256a,a41257a,a41260a,a41263a,a41264a,a41265a,a41269a,a41270a,a41273a,a41276a,a41277a,a41278a,a41282a,a41283a,a41286a,a41289a,a41290a,a41291a,a41295a,a41296a,a41299a,a41302a,a41303a,a41304a,a41308a,a41309a,a41312a,a41315a,a41316a,a41317a,a41321a,a41322a,a41325a,a41328a,a41329a,a41330a,a41334a,a41335a,a41338a,a41341a,a41342a,a41343a,a41347a,a41348a,a41351a,a41354a,a41355a,a41356a,a41360a,a41361a,a41364a,a41367a,a41368a,a41369a,a41373a,a41374a,a41377a,a41380a,a41381a,a41382a,a41386a,a41387a,a41390a,a41393a,a41394a,a41395a,a41399a,a41400a,a41403a,a41406a,a41407a,a41408a,a41412a,a41413a,a41416a,a41419a,a41420a,a41421a,a41425a,a41426a,a41429a,a41432a,a41433a,a41434a,a41438a,a41439a,a41442a,a41445a,a41446a,a41447a,a41451a,a41452a,a41455a,a41458a,a41459a,a41460a,a41464a,a41465a,a41468a,a41471a,a41472a,a41473a,a41477a,a41478a,a41481a,a41484a,a41485a,a41486a,a41490a,a41491a,a41494a,a41497a,a41498a,a41499a,a41503a,a41504a,a41507a,a41510a,a41511a,a41512a,a41516a,a41517a,a41520a,a41523a,a41524a,a41525a,a41529a,a41530a,a41533a,a41536a,a41537a,a41538a,a41542a,a41543a,a41546a,a41549a,a41550a,a41551a,a41555a,a41556a,a41559a,a41562a,a41563a,a41564a,a41568a,a41569a,a41572a,a41575a,a41576a,a41577a,a41581a,a41582a,a41585a,a41588a,a41589a,a41590a,a41594a,a41595a,a41598a,a41601a,a41602a,a41603a,a41607a,a41608a,a41611a,a41614a,a41615a,a41616a,a41620a,a41621a,a41624a,a41627a,a41628a,a41629a,a41633a,a41634a,a41637a,a41640a,a41641a,a41642a,a41646a,a41647a,a41650a,a41653a,a41654a,a41655a,a41659a,a41660a,a41663a,a41666a,a41667a,a41668a,a41672a,a41673a,a41676a,a41679a,a41680a,a41681a,a41685a,a41686a,a41689a,a41692a,a41693a,a41694a,a41698a,a41699a,a41702a,a41705a,a41706a,a41707a,a41711a,a41712a,a41715a,a41718a,a41719a,a41720a,a41724a,a41725a,a41728a,a41731a,a41732a,a41733a,a41737a,a41738a,a41741a,a41744a,a41745a,a41746a,a41750a,a41751a,a41754a,a41757a,a41758a,a41759a,a41763a,a41764a,a41767a,a41770a,a41771a,a41772a,a41776a,a41777a,a41780a,a41783a,a41784a,a41785a,a41789a,a41790a,a41793a,a41796a,a41797a,a41798a,a41802a,a41803a,a41806a,a41809a,a41810a,a41811a,a41815a,a41816a,a41819a,a41822a,a41823a,a41824a,a41828a,a41829a,a41832a,a41835a,a41836a,a41837a,a41841a,a41842a,a41845a,a41848a,a41849a,a41850a,a41854a,a41855a,a41858a,a41861a,a41862a,a41863a,a41867a,a41868a,a41871a,a41874a,a41875a,a41876a,a41880a,a41881a,a41884a,a41887a,a41888a,a41889a,a41893a,a41894a,a41897a,a41900a,a41901a,a41902a,a41906a,a41907a,a41910a,a41913a,a41914a,a41915a,a41919a,a41920a,a41923a,a41926a,a41927a,a41928a,a41932a,a41933a,a41936a,a41939a,a41940a,a41941a,a41945a,a41946a,a41949a,a41952a,a41953a,a41954a,a41958a,a41959a,a41962a,a41965a,a41966a,a41967a,a41971a,a41972a,a41975a,a41978a,a41979a,a41980a,a41984a,a41985a,a41988a,a41991a,a41992a,a41993a,a41997a,a41998a,a42001a,a42004a,a42005a,a42006a,a42010a,a42011a,a42014a,a42017a,a42018a,a42019a,a42023a,a42024a,a42027a,a42030a,a42031a,a42032a,a42036a,a42037a,a42040a,a42043a,a42044a,a42045a,a42049a,a42050a,a42053a,a42056a,a42057a,a42058a,a42062a,a42063a,a42066a,a42069a,a42070a,a42071a,a42075a,a42076a,a42079a,a42082a,a42083a,a42084a,a42088a,a42089a,a42092a,a42095a,a42096a,a42097a,a42101a,a42102a,a42105a,a42108a,a42109a,a42110a,a42114a,a42115a,a42118a,a42121a,a42122a,a42123a,a42127a,a42128a,a42131a,a42134a,a42135a,a42136a,a42140a,a42141a,a42144a,a42147a,a42148a,a42149a,a42153a,a42154a,a42157a,a42160a,a42161a,a42162a,a42166a,a42167a,a42170a,a42173a,a42174a,a42175a,a42179a,a42180a,a42183a,a42186a,a42187a,a42188a,a42192a,a42193a,a42196a,a42199a,a42200a,a42201a,a42205a,a42206a,a42209a,a42212a,a42213a,a42214a,a42218a,a42219a,a42222a,a42225a,a42226a,a42227a,a42231a,a42232a,a42235a,a42238a,a42239a,a42240a,a42244a,a42245a,a42248a,a42251a,a42252a,a42253a,a42257a,a42258a,a42261a,a42264a,a42265a,a42266a,a42270a,a42271a,a42274a,a42277a,a42278a,a42279a,a42283a,a42284a,a42287a,a42290a,a42291a,a42292a,a42296a,a42297a,a42300a,a42303a,a42304a,a42305a,a42309a,a42310a,a42313a,a42316a,a42317a,a42318a,a42322a,a42323a,a42326a,a42329a,a42330a,a42331a,a42335a,a42336a,a42339a,a42342a,a42343a,a42344a,a42348a,a42349a,a42352a,a42355a,a42356a,a42357a,a42361a,a42362a,a42365a,a42368a,a42369a,a42370a,a42374a,a42375a,a42378a,a42381a,a42382a,a42383a,a42387a,a42388a,a42391a,a42394a,a42395a,a42396a,a42400a,a42401a,a42404a,a42407a,a42408a,a42409a,a42413a,a42414a,a42417a,a42420a,a42421a,a42422a,a42426a,a42427a,a42430a,a42433a,a42434a,a42435a,a42439a,a42440a,a42443a,a42446a,a42447a,a42448a,a42452a,a42453a,a42456a,a42459a,a42460a,a42461a,a42465a,a42466a,a42469a,a42472a,a42473a,a42474a,a42478a,a42479a,a42482a,a42485a,a42486a,a42487a,a42491a,a42492a,a42495a,a42498a,a42499a,a42500a,a42504a,a42505a,a42508a,a42511a,a42512a,a42513a,a42517a,a42518a,a42521a,a42524a,a42525a,a42526a,a42530a,a42531a,a42534a,a42537a,a42538a,a42539a,a42543a,a42544a,a42547a,a42550a,a42551a,a42552a,a42556a,a42557a,a42560a,a42563a,a42564a,a42565a,a42569a,a42570a,a42573a,a42576a,a42577a,a42578a,a42582a,a42583a,a42586a,a42589a,a42590a,a42591a,a42595a,a42596a,a42599a,a42602a,a42603a,a42604a,a42608a,a42609a,a42612a,a42615a,a42616a,a42617a,a42621a,a42622a,a42625a,a42628a,a42629a,a42630a,a42634a,a42635a,a42638a,a42641a,a42642a,a42643a,a42647a,a42648a,a42651a,a42654a,a42655a,a42656a,a42660a,a42661a,a42664a,a42667a,a42668a,a42669a,a42673a,a42674a,a42677a,a42680a,a42681a,a42682a,a42686a,a42687a,a42690a,a42693a,a42694a,a42695a,a42699a,a42700a,a42703a,a42706a,a42707a,a42708a,a42712a,a42713a,a42716a,a42719a,a42720a,a42721a,a42725a,a42726a,a42729a,a42732a,a42733a,a42734a,a42738a,a42739a,a42742a,a42745a,a42746a,a42747a,a42751a,a42752a,a42755a,a42758a,a42759a,a42760a,a42764a,a42765a,a42768a,a42771a,a42772a,a42773a,a42777a,a42778a,a42781a,a42784a,a42785a,a42786a,a42790a,a42791a,a42794a,a42797a,a42798a,a42799a,a42803a,a42804a,a42807a,a42810a,a42811a,a42812a,a42816a,a42817a,a42820a,a42823a,a42824a,a42825a,a42829a,a42830a,a42833a,a42836a,a42837a,a42838a,a42842a,a42843a,a42846a,a42849a,a42850a,a42851a,a42855a,a42856a,a42859a,a42862a,a42863a,a42864a,a42868a,a42869a,a42872a,a42875a,a42876a,a42877a,a42881a,a42882a,a42885a,a42888a,a42889a,a42890a,a42894a,a42895a,a42898a,a42901a,a42902a,a42903a,a42907a,a42908a,a42911a,a42914a,a42915a,a42916a,a42920a,a42921a,a42924a,a42927a,a42928a,a42929a,a42933a,a42934a,a42937a,a42940a,a42941a,a42942a,a42946a,a42947a,a42950a,a42953a,a42954a,a42955a,a42959a,a42960a,a42963a,a42966a,a42967a,a42968a,a42972a,a42973a,a42976a,a42979a,a42980a,a42981a,a42985a,a42986a,a42989a,a42992a,a42993a,a42994a,a42998a,a42999a,a43002a,a43005a,a43006a,a43007a,a43011a,a43012a,a43015a,a43018a,a43019a,a43020a,a43024a,a43025a,a43028a,a43031a,a43032a,a43033a,a43037a,a43038a,a43041a,a43044a,a43045a,a43046a,a43050a,a43051a,a43054a,a43057a,a43058a,a43059a,a43063a,a43064a,a43067a,a43070a,a43071a,a43072a,a43076a,a43077a,a43080a,a43083a,a43084a,a43085a,a43089a,a43090a,a43093a,a43096a,a43097a,a43098a,a43102a,a43103a,a43106a,a43109a,a43110a,a43111a,a43115a,a43116a,a43119a,a43122a,a43123a,a43124a,a43128a,a43129a,a43132a,a43135a,a43136a,a43137a,a43141a,a43142a,a43145a,a43148a,a43149a,a43150a,a43154a,a43155a,a43158a,a43161a,a43162a,a43163a,a43167a,a43168a,a43171a,a43174a,a43175a,a43176a,a43180a,a43181a,a43184a,a43187a,a43188a,a43189a,a43193a,a43194a,a43197a,a43200a,a43201a,a43202a,a43206a,a43207a,a43210a,a43213a,a43214a,a43215a,a43219a,a43220a,a43223a,a43226a,a43227a,a43228a,a43232a,a43233a,a43236a,a43239a,a43240a,a43241a,a43245a,a43246a,a43249a,a43252a,a43253a,a43254a,a43258a,a43259a,a43262a,a43265a,a43266a,a43267a,a43271a,a43272a,a43275a,a43278a,a43279a,a43280a,a43284a,a43285a,a43288a,a43291a,a43292a,a43293a,a43297a,a43298a,a43301a,a43304a,a43305a,a43306a,a43310a,a43311a,a43314a,a43317a,a43318a,a43319a,a43323a,a43324a,a43327a,a43330a,a43331a,a43332a,a43336a,a43337a,a43340a,a43343a,a43344a,a43345a,a43349a,a43350a,a43353a,a43356a,a43357a,a43358a,a43362a,a43363a,a43366a,a43369a,a43370a,a43371a,a43375a,a43376a,a43379a,a43382a,a43383a,a43384a,a43388a,a43389a,a43392a,a43395a,a43396a,a43397a,a43401a,a43402a,a43405a,a43408a,a43409a,a43410a,a43414a,a43415a,a43418a,a43421a,a43422a,a43423a,a43427a,a43428a,a43431a,a43434a,a43435a,a43436a,a43440a,a43441a,a43444a,a43447a,a43448a,a43449a,a43453a,a43454a,a43457a,a43460a,a43461a,a43462a,a43466a,a43467a,a43470a,a43473a,a43474a,a43475a,a43479a,a43480a,a43483a,a43486a,a43487a,a43488a,a43492a,a43493a,a43496a,a43499a,a43500a,a43501a,a43505a,a43506a,a43509a,a43512a,a43513a,a43514a,a43518a,a43519a,a43522a,a43525a,a43526a,a43527a,a43531a,a43532a,a43535a,a43538a,a43539a,a43540a,a43544a,a43545a,a43548a,a43551a,a43552a,a43553a,a43557a,a43558a,a43561a,a43564a,a43565a,a43566a,a43570a,a43571a,a43574a,a43577a,a43578a,a43579a,a43583a,a43584a,a43587a,a43590a,a43591a,a43592a,a43596a,a43597a,a43600a,a43603a,a43604a,a43605a,a43609a,a43610a,a43613a,a43616a,a43617a,a43618a,a43622a,a43623a,a43626a,a43629a,a43630a,a43631a,a43635a,a43636a,a43639a,a43642a,a43643a,a43644a,a43648a,a43649a,a43652a,a43655a,a43656a,a43657a,a43661a,a43662a,a43665a,a43668a,a43669a,a43670a,a43674a,a43675a,a43678a,a43681a,a43682a,a43683a,a43687a,a43688a,a43691a,a43694a,a43695a,a43696a,a43700a,a43701a,a43704a,a43707a,a43708a,a43709a,a43713a,a43714a,a43717a,a43720a,a43721a,a43722a,a43726a,a43727a,a43730a,a43733a,a43734a,a43735a,a43739a,a43740a,a43743a,a43746a,a43747a,a43748a,a43752a,a43753a,a43756a,a43759a,a43760a,a43761a,a43765a,a43766a,a43769a,a43772a,a43773a,a43774a,a43778a,a43779a,a43782a,a43785a,a43786a,a43787a,a43791a,a43792a,a43795a,a43798a,a43799a,a43800a,a43804a,a43805a,a43808a,a43811a,a43812a,a43813a,a43817a,a43818a,a43821a,a43824a,a43825a,a43826a,a43830a,a43831a,a43834a,a43837a,a43838a,a43839a,a43843a,a43844a,a43847a,a43850a,a43851a,a43852a,a43856a,a43857a,a43860a,a43863a,a43864a,a43865a,a43869a,a43870a,a43873a,a43876a,a43877a,a43878a,a43882a,a43883a,a43886a,a43889a,a43890a,a43891a,a43895a,a43896a,a43899a,a43902a,a43903a,a43904a,a43908a,a43909a,a43912a,a43915a,a43916a,a43917a,a43921a,a43922a,a43925a,a43928a,a43929a,a43930a,a43934a,a43935a,a43938a,a43941a,a43942a,a43943a,a43947a,a43948a,a43951a,a43954a,a43955a,a43956a,a43960a,a43961a,a43964a,a43967a,a43968a,a43969a,a43973a,a43974a,a43977a,a43980a,a43981a,a43982a,a43986a,a43987a,a43990a,a43993a,a43994a,a43995a,a43999a,a44000a,a44003a,a44006a,a44007a,a44008a,a44012a,a44013a,a44016a,a44019a,a44020a,a44021a,a44025a,a44026a,a44029a,a44032a,a44033a,a44034a,a44038a,a44039a,a44042a,a44045a,a44046a,a44047a,a44051a,a44052a,a44055a,a44058a,a44059a,a44060a,a44064a,a44065a,a44068a,a44071a,a44072a,a44073a,a44077a,a44078a,a44081a,a44084a,a44085a,a44086a,a44090a,a44091a,a44094a,a44097a,a44098a,a44099a,a44103a,a44104a,a44107a,a44110a,a44111a,a44112a,a44116a,a44117a,a44120a,a44123a,a44124a,a44125a,a44129a,a44130a,a44133a,a44136a,a44137a,a44138a,a44142a,a44143a,a44146a,a44149a,a44150a,a44151a,a44155a,a44156a,a44159a,a44162a,a44163a,a44164a,a44168a,a44169a,a44172a,a44175a,a44176a,a44177a,a44181a,a44182a,a44185a,a44188a,a44189a,a44190a,a44194a,a44195a,a44198a,a44201a,a44202a,a44203a,a44207a,a44208a,a44211a,a44214a,a44215a,a44216a,a44220a,a44221a,a44224a,a44227a,a44228a,a44229a,a44233a,a44234a,a44237a,a44240a,a44241a,a44242a,a44246a,a44247a,a44250a,a44253a,a44254a,a44255a,a44259a,a44260a,a44263a,a44266a,a44267a,a44268a,a44272a,a44273a,a44276a,a44279a,a44280a,a44281a,a44285a,a44286a,a44289a,a44292a,a44293a,a44294a,a44298a,a44299a,a44302a,a44305a,a44306a,a44307a,a44311a,a44312a,a44315a,a44318a,a44319a,a44320a,a44324a,a44325a,a44328a,a44331a,a44332a,a44333a,a44337a,a44338a,a44341a,a44344a,a44345a,a44346a,a44350a,a44351a,a44354a,a44357a,a44358a,a44359a,a44363a,a44364a,a44367a,a44370a,a44371a,a44372a,a44376a,a44377a,a44380a,a44383a,a44384a,a44385a,a44389a,a44390a,a44393a,a44396a,a44397a,a44398a,a44402a,a44403a,a44406a,a44409a,a44410a,a44411a,a44415a,a44416a,a44419a,a44422a,a44423a,a44424a,a44428a,a44429a,a44432a,a44435a,a44436a,a44437a,a44441a,a44442a,a44445a,a44448a,a44449a,a44450a,a44454a,a44455a,a44458a,a44461a,a44462a,a44463a,a44467a,a44468a,a44471a,a44474a,a44475a,a44476a,a44480a,a44481a,a44484a,a44487a,a44488a,a44489a,a44493a,a44494a,a44497a,a44500a,a44501a,a44502a,a44506a,a44507a,a44510a,a44513a,a44514a,a44515a,a44519a,a44520a,a44523a,a44526a,a44527a,a44528a,a44532a,a44533a,a44536a,a44539a,a44540a,a44541a,a44545a,a44546a,a44549a,a44552a,a44553a,a44554a,a44558a,a44559a,a44562a,a44565a,a44566a,a44567a,a44571a,a44572a,a44575a,a44578a,a44579a,a44580a,a44584a,a44585a,a44588a,a44591a,a44592a,a44593a,a44597a,a44598a,a44601a,a44604a,a44605a,a44606a,a44610a,a44611a,a44614a,a44617a,a44618a,a44619a,a44623a,a44624a,a44627a,a44630a,a44631a,a44632a,a44636a,a44637a,a44640a,a44643a,a44644a,a44645a,a44649a,a44650a,a44653a,a44656a,a44657a,a44658a,a44662a,a44663a,a44666a,a44669a,a44670a,a44671a,a44675a,a44676a,a44679a,a44682a,a44683a,a44684a,a44688a,a44689a,a44692a,a44695a,a44696a,a44697a,a44701a,a44702a,a44705a,a44708a,a44709a,a44710a,a44714a,a44715a,a44718a,a44721a,a44722a,a44723a,a44727a,a44728a,a44731a,a44734a,a44735a,a44736a,a44740a,a44741a,a44744a,a44747a,a44748a,a44749a,a44753a,a44754a,a44757a,a44760a,a44761a,a44762a,a44766a,a44767a,a44770a,a44773a,a44774a,a44775a,a44779a,a44780a,a44783a,a44786a,a44787a,a44788a,a44792a,a44793a,a44796a,a44799a,a44800a,a44801a,a44805a,a44806a,a44809a,a44812a,a44813a,a44814a,a44818a,a44819a,a44822a,a44825a,a44826a,a44827a,a44831a,a44832a,a44835a,a44838a,a44839a,a44840a,a44844a,a44845a,a44848a,a44851a,a44852a,a44853a,a44857a,a44858a,a44861a,a44864a,a44865a,a44866a,a44870a,a44871a,a44874a,a44877a,a44878a,a44879a,a44883a,a44884a,a44887a,a44890a,a44891a,a44892a,a44896a,a44897a,a44900a,a44903a,a44904a,a44905a,a44909a,a44910a,a44913a,a44916a,a44917a,a44918a,a44922a,a44923a,a44926a,a44929a,a44930a,a44931a,a44935a,a44936a,a44939a,a44942a,a44943a,a44944a,a44948a,a44949a,a44952a,a44955a,a44956a,a44957a,a44961a,a44962a,a44965a,a44968a,a44969a,a44970a,a44974a,a44975a,a44978a,a44981a,a44982a,a44983a,a44987a,a44988a,a44991a,a44994a,a44995a,a44996a,a45000a,a45001a,a45004a,a45007a,a45008a,a45009a,a45013a,a45014a,a45017a,a45020a,a45021a,a45022a,a45026a,a45027a,a45030a,a45033a,a45034a,a45035a,a45039a,a45040a,a45043a,a45046a,a45047a,a45048a,a45052a,a45053a,a45056a,a45059a,a45060a,a45061a,a45065a,a45066a,a45069a,a45072a,a45073a,a45074a,a45078a,a45079a,a45082a,a45085a,a45086a,a45087a,a45091a,a45092a,a45095a,a45098a,a45099a,a45100a,a45104a,a45105a,a45108a,a45111a,a45112a,a45113a,a45117a,a45118a,a45121a,a45124a,a45125a,a45126a,a45130a,a45131a,a45134a,a45137a,a45138a,a45139a,a45143a,a45144a,a45147a,a45150a,a45151a,a45152a,a45156a,a45157a,a45160a,a45163a,a45164a,a45165a,a45169a,a45170a,a45173a,a45176a,a45177a,a45178a,a45182a,a45183a,a45186a,a45189a,a45190a,a45191a,a45195a,a45196a,a45199a,a45202a,a45203a,a45204a,a45208a,a45209a,a45212a,a45215a,a45216a,a45217a,a45221a,a45222a,a45225a,a45228a,a45229a,a45230a,a45234a,a45235a,a45238a,a45241a,a45242a,a45243a,a45247a,a45248a,a45251a,a45254a,a45255a,a45256a,a45260a,a45261a,a45264a,a45267a,a45268a,a45269a,a45273a,a45274a,a45277a,a45280a,a45281a,a45282a,a45286a,a45287a,a45290a,a45293a,a45294a,a45295a,a45299a,a45300a,a45303a,a45306a,a45307a,a45308a,a45312a,a45313a,a45316a,a45319a,a45320a,a45321a,a45325a,a45326a,a45329a,a45332a,a45333a,a45334a,a45338a,a45339a,a45342a,a45345a,a45346a,a45347a,a45351a,a45352a,a45355a,a45358a,a45359a,a45360a,a45364a,a45365a,a45368a,a45371a,a45372a,a45373a,a45377a,a45378a,a45381a,a45384a,a45385a,a45386a,a45390a,a45391a,a45394a,a45397a,a45398a,a45399a,a45403a,a45404a,a45407a,a45410a,a45411a,a45412a,a45416a,a45417a,a45420a,a45423a,a45424a,a45425a,a45429a,a45430a,a45433a,a45436a,a45437a,a45438a,a45442a,a45443a,a45446a,a45449a,a45450a,a45451a,a45455a,a45456a,a45459a,a45462a,a45463a,a45464a,a45468a,a45469a,a45472a,a45475a,a45476a,a45477a,a45481a,a45482a,a45485a,a45488a,a45489a,a45490a,a45494a,a45495a,a45498a,a45501a,a45502a,a45503a,a45507a,a45508a,a45511a,a45514a,a45515a,a45516a,a45520a,a45521a,a45524a,a45527a,a45528a,a45529a,a45533a,a45534a,a45537a,a45540a,a45541a,a45542a,a45546a,a45547a,a45550a,a45553a,a45554a,a45555a,a45559a,a45560a,a45563a,a45566a,a45567a,a45568a,a45572a,a45573a,a45576a,a45579a,a45580a,a45581a,a45585a,a45586a,a45589a,a45592a,a45593a,a45594a,a45598a,a45599a,a45602a,a45605a,a45606a,a45607a,a45611a,a45612a,a45615a,a45618a,a45619a,a45620a,a45624a,a45625a,a45628a,a45631a,a45632a,a45633a,a45637a,a45638a,a45641a,a45644a,a45645a,a45646a,a45650a,a45651a,a45654a,a45657a,a45658a,a45659a,a45663a,a45664a,a45667a,a45670a,a45671a,a45672a,a45676a,a45677a,a45680a,a45683a,a45684a,a45685a,a45689a,a45690a,a45693a,a45696a,a45697a,a45698a,a45702a,a45703a,a45706a,a45709a,a45710a,a45711a,a45715a,a45716a,a45719a,a45722a,a45723a,a45724a,a45728a,a45729a,a45732a,a45735a,a45736a,a45737a,a45741a,a45742a,a45745a,a45748a,a45749a,a45750a,a45754a,a45755a,a45758a,a45761a,a45762a,a45763a,a45767a,a45768a,a45771a,a45774a,a45775a,a45776a,a45780a,a45781a,a45784a,a45787a,a45788a,a45789a,a45793a,a45794a,a45797a,a45800a,a45801a,a45802a,a45806a,a45807a,a45810a,a45813a,a45814a,a45815a,a45819a,a45820a,a45823a,a45826a,a45827a,a45828a,a45832a,a45833a,a45836a,a45839a,a45840a,a45841a,a45845a,a45846a,a45849a,a45852a,a45853a,a45854a,a45858a,a45859a,a45862a,a45865a,a45866a,a45867a,a45871a,a45872a,a45875a,a45878a,a45879a,a45880a,a45884a,a45885a,a45888a,a45891a,a45892a,a45893a,a45897a,a45898a,a45901a,a45904a,a45905a,a45906a,a45910a,a45911a,a45914a,a45917a,a45918a,a45919a,a45923a,a45924a,a45927a,a45930a,a45931a,a45932a,a45936a,a45937a,a45940a,a45943a,a45944a,a45945a,a45949a,a45950a,a45953a,a45956a,a45957a,a45958a,a45962a,a45963a,a45966a,a45969a,a45970a,a45971a,a45975a,a45976a,a45979a,a45982a,a45983a,a45984a,a45988a,a45989a,a45992a,a45995a,a45996a,a45997a,a46001a,a46002a,a46005a,a46008a,a46009a,a46010a,a46014a,a46015a,a46018a,a46021a,a46022a,a46023a,a46027a,a46028a,a46031a,a46034a,a46035a,a46036a,a46040a,a46041a,a46044a,a46047a,a46048a,a46049a,a46053a,a46054a,a46057a,a46060a,a46061a,a46062a,a46066a,a46067a,a46070a,a46073a,a46074a,a46075a,a46079a,a46080a,a46083a,a46086a,a46087a,a46088a,a46092a,a46093a,a46096a,a46099a,a46100a,a46101a,a46105a,a46106a,a46109a,a46112a,a46113a,a46114a,a46118a,a46119a,a46122a,a46125a,a46126a,a46127a,a46131a,a46132a,a46135a,a46138a,a46139a,a46140a,a46144a,a46145a,a46148a,a46151a,a46152a,a46153a,a46157a,a46158a,a46161a,a46164a,a46165a,a46166a,a46170a,a46171a,a46174a,a46177a,a46178a,a46179a,a46183a,a46184a,a46187a,a46190a,a46191a,a46192a,a46196a,a46197a,a46200a,a46203a,a46204a,a46205a,a46209a,a46210a,a46213a,a46216a,a46217a,a46218a,a46222a,a46223a,a46226a,a46229a,a46230a,a46231a,a46235a,a46236a,a46239a,a46242a,a46243a,a46244a,a46248a,a46249a,a46252a,a46255a,a46256a,a46257a,a46261a,a46262a,a46265a,a46268a,a46269a,a46270a,a46274a,a46275a,a46278a,a46281a,a46282a,a46283a,a46287a,a46288a,a46291a,a46294a,a46295a,a46296a,a46300a,a46301a,a46304a,a46307a,a46308a,a46309a,a46313a,a46314a,a46317a,a46320a,a46321a,a46322a,a46326a,a46327a,a46330a,a46333a,a46334a,a46335a,a46339a,a46340a,a46343a,a46346a,a46347a,a46348a,a46352a,a46353a,a46356a,a46359a,a46360a,a46361a,a46365a,a46366a,a46369a,a46372a,a46373a,a46374a,a46378a,a46379a,a46382a,a46385a,a46386a,a46387a,a46391a,a46392a,a46395a,a46398a,a46399a,a46400a,a46404a,a46405a,a46408a,a46411a,a46412a,a46413a,a46417a,a46418a,a46421a,a46424a,a46425a,a46426a,a46430a,a46431a,a46434a,a46437a,a46438a,a46439a,a46443a,a46444a,a46447a,a46450a,a46451a,a46452a,a46456a,a46457a,a46460a,a46463a,a46464a,a46465a,a46469a,a46470a,a46473a,a46476a,a46477a,a46478a,a46482a,a46483a,a46486a,a46489a,a46490a,a46491a,a46495a,a46496a,a46499a,a46502a,a46503a,a46504a,a46508a,a46509a,a46512a,a46515a,a46516a,a46517a,a46521a,a46522a,a46525a,a46528a,a46529a,a46530a,a46534a,a46535a,a46538a,a46541a,a46542a,a46543a,a46547a,a46548a,a46551a,a46554a,a46555a,a46556a,a46560a,a46561a,a46564a,a46567a,a46568a,a46569a,a46573a,a46574a,a46577a,a46580a,a46581a,a46582a,a46586a,a46587a,a46590a,a46593a,a46594a,a46595a,a46599a,a46600a,a46603a,a46606a,a46607a,a46608a,a46612a,a46613a,a46616a,a46619a,a46620a,a46621a,a46625a,a46626a,a46629a,a46632a,a46633a,a46634a,a46638a,a46639a,a46642a,a46645a,a46646a,a46647a,a46651a,a46652a,a46655a,a46658a,a46659a,a46660a,a46664a,a46665a,a46668a,a46671a,a46672a,a46673a,a46677a,a46678a,a46681a,a46684a,a46685a,a46686a,a46690a,a46691a,a46694a,a46697a,a46698a,a46699a,a46703a,a46704a,a46707a,a46710a,a46711a,a46712a,a46716a,a46717a,a46720a,a46723a,a46724a,a46725a,a46729a,a46730a,a46733a,a46736a,a46737a,a46738a,a46742a,a46743a,a46746a,a46749a,a46750a,a46751a,a46755a,a46756a,a46759a,a46762a,a46763a,a46764a,a46768a,a46769a,a46772a,a46775a,a46776a,a46777a,a46781a,a46782a,a46785a,a46788a,a46789a,a46790a,a46794a,a46795a,a46798a,a46801a,a46802a,a46803a,a46807a,a46808a,a46811a,a46814a,a46815a,a46816a,a46820a,a46821a,a46824a,a46827a,a46828a,a46829a,a46833a,a46834a,a46837a,a46840a,a46841a,a46842a,a46846a,a46847a,a46850a,a46853a,a46854a,a46855a,a46859a,a46860a,a46863a,a46866a,a46867a,a46868a,a46872a,a46873a,a46876a,a46879a,a46880a,a46881a,a46885a,a46886a,a46889a,a46892a,a46893a,a46894a,a46898a,a46899a,a46902a,a46905a,a46906a,a46907a,a46911a,a46912a,a46915a,a46918a,a46919a,a46920a,a46924a,a46925a,a46928a,a46931a,a46932a,a46933a,a46937a,a46938a,a46941a,a46944a,a46945a,a46946a,a46950a,a46951a,a46954a,a46957a,a46958a,a46959a,a46963a,a46964a,a46967a,a46970a,a46971a,a46972a,a46976a,a46977a,a46980a,a46983a,a46984a,a46985a,a46989a,a46990a,a46993a,a46996a,a46997a,a46998a,a47002a,a47003a,a47006a,a47009a,a47010a,a47011a,a47015a,a47016a,a47019a,a47022a,a47023a,a47024a,a47028a,a47029a,a47032a,a47035a,a47036a,a47037a,a47041a,a47042a,a47045a,a47048a,a47049a,a47050a,a47054a,a47055a,a47058a,a47061a,a47062a,a47063a,a47067a,a47068a,a47071a,a47074a,a47075a,a47076a,a47080a,a47081a,a47084a,a47087a,a47088a,a47089a,a47093a,a47094a,a47097a,a47100a,a47101a,a47102a,a47106a,a47107a,a47110a,a47113a,a47114a,a47115a,a47119a,a47120a,a47123a,a47126a,a47127a,a47128a,a47132a,a47133a,a47136a,a47139a,a47140a,a47141a,a47145a,a47146a,a47149a,a47152a,a47153a,a47154a,a47158a,a47159a,a47162a,a47165a,a47166a,a47167a,a47171a,a47172a,a47175a,a47178a,a47179a,a47180a,a47184a,a47185a,a47188a,a47191a,a47192a,a47193a,a47197a,a47198a,a47201a,a47204a,a47205a,a47206a,a47210a,a47211a,a47214a,a47217a,a47218a,a47219a,a47223a,a47224a,a47227a,a47230a,a47231a,a47232a,a47236a,a47237a,a47240a,a47243a,a47244a,a47245a,a47249a,a47250a,a47253a,a47256a,a47257a,a47258a,a47262a,a47263a,a47266a,a47269a,a47270a,a47271a,a47275a,a47276a,a47279a,a47282a,a47283a,a47284a,a47288a,a47289a,a47292a,a47295a,a47296a,a47297a,a47301a,a47302a,a47305a,a47308a,a47309a,a47310a,a47314a,a47315a,a47318a,a47321a,a47322a,a47323a,a47327a,a47328a,a47331a,a47334a,a47335a,a47336a,a47340a,a47341a,a47344a,a47347a,a47348a,a47349a,a47353a,a47354a,a47357a,a47360a,a47361a,a47362a,a47366a,a47367a,a47370a,a47373a,a47374a,a47375a,a47379a,a47380a,a47383a,a47386a,a47387a,a47388a,a47392a,a47393a,a47396a,a47399a,a47400a,a47401a,a47405a,a47406a,a47409a,a47412a,a47413a,a47414a,a47418a,a47419a,a47422a,a47425a,a47426a,a47427a,a47431a,a47432a,a47435a,a47438a,a47439a,a47440a,a47444a,a47445a,a47448a,a47451a,a47452a,a47453a,a47457a,a47458a,a47461a,a47464a,a47465a,a47466a,a47470a,a47471a,a47474a,a47477a,a47478a,a47479a,a47483a,a47484a,a47487a,a47490a,a47491a,a47492a,a47496a,a47497a,a47500a,a47503a,a47504a,a47505a,a47509a,a47510a,a47513a,a47516a,a47517a,a47518a,a47522a,a47523a,a47526a,a47529a,a47530a,a47531a,a47535a,a47536a,a47539a,a47542a,a47543a,a47544a,a47548a,a47549a,a47552a,a47555a,a47556a,a47557a,a47561a,a47562a,a47565a,a47568a,a47569a,a47570a,a47574a,a47575a,a47578a,a47581a,a47582a,a47583a,a47587a,a47588a,a47591a,a47594a,a47595a,a47596a,a47600a,a47601a,a47604a,a47607a,a47608a,a47609a,a47613a,a47614a,a47617a,a47620a,a47621a,a47622a,a47626a,a47627a,a47630a,a47633a,a47634a,a47635a,a47639a,a47640a,a47643a,a47646a,a47647a,a47648a,a47652a,a47653a,a47656a,a47659a,a47660a,a47661a,a47664a,a47667a,a47668a,a47671a,a47674a,a47675a,a47676a,a47680a,a47681a,a47684a,a47687a,a47688a,a47689a,a47692a,a47695a,a47696a,a47699a,a47702a,a47703a,a47704a,a47708a,a47709a,a47712a,a47715a,a47716a,a47717a,a47720a,a47723a,a47724a,a47727a,a47730a,a47731a,a47732a,a47736a,a47737a,a47740a,a47743a,a47744a,a47745a,a47748a,a47751a,a47752a,a47755a,a47758a,a47759a,a47760a,a47764a,a47765a,a47768a,a47771a,a47772a,a47773a,a47776a,a47779a,a47780a,a47783a,a47786a,a47787a,a47788a,a47792a,a47793a,a47796a,a47799a,a47800a,a47801a,a47804a,a47807a,a47808a,a47811a,a47814a,a47815a,a47816a,a47820a,a47821a,a47824a,a47827a,a47828a,a47829a,a47832a,a47835a,a47836a,a47839a,a47842a,a47843a,a47844a,a47848a,a47849a,a47852a,a47855a,a47856a,a47857a,a47860a,a47863a,a47864a,a47867a,a47870a,a47871a,a47872a,a47876a,a47877a,a47880a,a47883a,a47884a,a47885a,a47888a,a47891a,a47892a,a47895a,a47898a,a47899a,a47900a,a47904a,a47905a,a47908a,a47911a,a47912a,a47913a,a47916a,a47919a,a47920a,a47923a,a47926a,a47927a,a47928a,a47932a,a47933a,a47936a,a47939a,a47940a,a47941a,a47944a,a47947a,a47948a,a47951a,a47954a,a47955a,a47956a,a47960a,a47961a,a47964a,a47967a,a47968a,a47969a,a47972a,a47975a,a47976a,a47979a,a47982a,a47983a,a47984a,a47988a,a47989a,a47992a,a47995a,a47996a,a47997a,a48000a,a48003a,a48004a,a48007a,a48010a,a48011a,a48012a,a48016a,a48017a,a48020a,a48023a,a48024a,a48025a,a48028a,a48031a,a48032a,a48035a,a48038a,a48039a,a48040a,a48044a,a48045a,a48048a,a48051a,a48052a,a48053a,a48056a,a48059a,a48060a,a48063a,a48066a,a48067a,a48068a,a48072a,a48073a,a48076a,a48079a,a48080a,a48081a,a48084a,a48087a,a48088a,a48091a,a48094a,a48095a,a48096a,a48100a,a48101a,a48104a,a48107a,a48108a,a48109a,a48112a,a48115a,a48116a,a48119a,a48122a,a48123a,a48124a,a48128a,a48129a,a48132a,a48135a,a48136a,a48137a,a48140a,a48143a,a48144a,a48147a,a48150a,a48151a,a48152a,a48156a,a48157a,a48160a,a48163a,a48164a,a48165a,a48168a,a48171a,a48172a,a48175a,a48178a,a48179a,a48180a,a48184a,a48185a,a48188a,a48191a,a48192a,a48193a,a48196a,a48199a,a48200a,a48203a,a48206a,a48207a,a48208a,a48212a,a48213a,a48216a,a48219a,a48220a,a48221a,a48224a,a48227a,a48228a,a48231a,a48234a,a48235a,a48236a,a48240a,a48241a,a48244a,a48247a,a48248a,a48249a,a48252a,a48255a,a48256a,a48259a,a48262a,a48263a,a48264a,a48268a,a48269a,a48272a,a48275a,a48276a,a48277a,a48280a,a48283a,a48284a,a48287a,a48290a,a48291a,a48292a,a48296a,a48297a,a48300a,a48303a,a48304a,a48305a,a48308a,a48311a,a48312a,a48315a,a48318a,a48319a,a48320a,a48324a,a48325a,a48328a,a48331a,a48332a,a48333a,a48336a,a48339a,a48340a,a48343a,a48346a,a48347a,a48348a,a48352a,a48353a,a48356a,a48359a,a48360a,a48361a,a48364a,a48367a,a48368a,a48371a,a48374a,a48375a,a48376a,a48380a,a48381a,a48384a,a48387a,a48388a,a48389a,a48392a,a48395a,a48396a,a48399a,a48402a,a48403a,a48404a,a48408a,a48409a,a48412a,a48415a,a48416a,a48417a,a48420a,a48423a,a48424a,a48427a,a48430a,a48431a,a48432a,a48436a,a48437a,a48440a,a48443a,a48444a,a48445a,a48448a,a48451a,a48452a,a48455a,a48458a,a48459a,a48460a,a48464a,a48465a,a48468a,a48471a,a48472a,a48473a,a48476a,a48479a,a48480a,a48483a,a48486a,a48487a,a48488a,a48492a,a48493a,a48496a,a48499a,a48500a,a48501a,a48504a,a48507a,a48508a,a48511a,a48514a,a48515a,a48516a,a48520a,a48521a,a48524a,a48527a,a48528a,a48529a,a48532a,a48535a,a48536a,a48539a,a48542a,a48543a,a48544a,a48548a,a48549a,a48552a,a48555a,a48556a,a48557a,a48560a,a48563a,a48564a,a48567a,a48570a,a48571a,a48572a,a48576a,a48577a,a48580a,a48583a,a48584a,a48585a,a48588a,a48591a,a48592a,a48595a,a48598a,a48599a,a48600a,a48604a,a48605a,a48608a,a48611a,a48612a,a48613a,a48616a,a48619a,a48620a,a48623a,a48626a,a48627a,a48628a,a48632a,a48633a,a48636a,a48639a,a48640a,a48641a,a48644a,a48647a,a48648a,a48651a,a48654a,a48655a,a48656a,a48660a,a48661a,a48664a,a48667a,a48668a,a48669a,a48672a,a48675a,a48676a,a48679a,a48682a,a48683a,a48684a,a48688a,a48689a,a48692a,a48695a,a48696a,a48697a,a48700a,a48703a,a48704a,a48707a,a48710a,a48711a,a48712a,a48716a,a48717a,a48720a,a48723a,a48724a,a48725a,a48728a,a48731a,a48732a,a48735a,a48738a,a48739a,a48740a,a48744a,a48745a,a48748a,a48751a,a48752a,a48753a,a48756a,a48759a,a48760a,a48763a,a48766a,a48767a,a48768a,a48772a,a48773a,a48776a,a48779a,a48780a,a48781a,a48784a,a48787a,a48788a,a48791a,a48794a,a48795a,a48796a,a48800a,a48801a,a48804a,a48807a,a48808a,a48809a,a48812a,a48815a,a48816a,a48819a,a48822a,a48823a,a48824a,a48828a,a48829a,a48832a,a48835a,a48836a,a48837a,a48840a,a48843a,a48844a,a48847a,a48850a,a48851a,a48852a,a48856a,a48857a,a48860a,a48863a,a48864a,a48865a,a48868a,a48871a,a48872a,a48875a,a48878a,a48879a,a48880a,a48884a,a48885a,a48888a,a48891a,a48892a,a48893a,a48896a,a48899a,a48900a,a48903a,a48906a,a48907a,a48908a,a48912a,a48913a,a48916a,a48919a,a48920a,a48921a,a48924a,a48927a,a48928a,a48931a,a48934a,a48935a,a48936a,a48940a,a48941a,a48944a,a48947a,a48948a,a48949a,a48952a,a48955a,a48956a,a48959a,a48962a,a48963a,a48964a,a48968a,a48969a,a48972a,a48975a,a48976a,a48977a,a48980a,a48983a,a48984a,a48987a,a48990a,a48991a,a48992a,a48996a,a48997a,a49000a,a49003a,a49004a,a49005a,a49008a,a49011a,a49012a,a49015a,a49018a,a49019a,a49020a,a49024a,a49025a,a49028a,a49031a,a49032a,a49033a,a49036a,a49039a,a49040a,a49043a,a49046a,a49047a,a49048a,a49052a,a49053a,a49056a,a49059a,a49060a,a49061a,a49064a,a49067a,a49068a,a49071a,a49074a,a49075a,a49076a,a49080a,a49081a,a49084a,a49087a,a49088a,a49089a,a49092a,a49095a,a49096a,a49099a,a49102a,a49103a,a49104a,a49108a,a49109a,a49112a,a49115a,a49116a,a49117a,a49120a,a49123a,a49124a,a49127a,a49130a,a49131a,a49132a,a49136a,a49137a,a49140a,a49143a,a49144a,a49145a,a49148a,a49151a,a49152a,a49155a,a49158a,a49159a,a49160a,a49164a,a49165a,a49168a,a49171a,a49172a,a49173a,a49176a,a49179a,a49180a,a49183a,a49186a,a49187a,a49188a,a49192a,a49193a,a49196a,a49199a,a49200a,a49201a,a49204a,a49207a,a49208a,a49211a,a49214a,a49215a,a49216a,a49220a,a49221a,a49224a,a49227a,a49228a,a49229a,a49232a,a49235a,a49236a,a49239a,a49242a,a49243a,a49244a,a49248a,a49249a,a49252a,a49255a,a49256a,a49257a,a49260a,a49263a,a49264a,a49267a,a49270a,a49271a,a49272a,a49276a,a49277a,a49280a,a49283a,a49284a,a49285a,a49288a,a49291a,a49292a,a49295a,a49298a,a49299a,a49300a,a49304a,a49305a,a49308a,a49311a,a49312a,a49313a,a49316a,a49319a,a49320a,a49323a,a49326a,a49327a,a49328a,a49332a,a49333a,a49336a,a49339a,a49340a,a49341a,a49344a,a49347a,a49348a,a49351a,a49354a,a49355a,a49356a,a49360a,a49361a,a49364a,a49367a,a49368a,a49369a,a49372a,a49375a,a49376a,a49379a,a49382a,a49383a,a49384a,a49388a,a49389a,a49392a,a49395a,a49396a,a49397a,a49400a,a49403a,a49404a,a49407a,a49410a,a49411a,a49412a,a49416a,a49417a,a49420a,a49423a,a49424a,a49425a,a49428a,a49431a,a49432a,a49435a,a49438a,a49439a,a49440a,a49444a,a49445a,a49448a,a49451a,a49452a,a49453a,a49456a,a49459a,a49460a,a49463a,a49466a,a49467a,a49468a,a49472a,a49473a,a49476a,a49479a,a49480a,a49481a,a49484a,a49487a,a49488a,a49491a,a49494a,a49495a,a49496a,a49500a,a49501a,a49504a,a49507a,a49508a,a49509a,a49512a,a49515a,a49516a,a49519a,a49522a,a49523a,a49524a,a49528a,a49529a,a49532a,a49535a,a49536a,a49537a,a49540a,a49543a,a49544a,a49547a,a49550a,a49551a,a49552a,a49556a,a49557a,a49560a,a49563a,a49564a,a49565a,a49568a,a49571a,a49572a,a49575a,a49578a,a49579a,a49580a,a49584a,a49585a,a49588a,a49591a,a49592a,a49593a,a49596a,a49599a,a49600a,a49603a,a49606a,a49607a,a49608a,a49612a,a49613a,a49616a,a49619a,a49620a,a49621a,a49624a,a49627a,a49628a,a49631a,a49634a,a49635a,a49636a,a49640a,a49641a,a49644a,a49647a,a49648a,a49649a,a49652a,a49655a,a49656a,a49659a,a49662a,a49663a,a49664a,a49668a,a49669a,a49672a,a49675a,a49676a,a49677a,a49680a,a49683a,a49684a,a49687a,a49690a,a49691a,a49692a,a49696a,a49697a,a49700a,a49703a,a49704a,a49705a,a49708a,a49711a,a49712a,a49715a,a49718a,a49719a,a49720a,a49724a,a49725a,a49728a,a49731a,a49732a,a49733a,a49736a,a49739a,a49740a,a49743a,a49746a,a49747a,a49748a,a49752a,a49753a,a49756a,a49759a,a49760a,a49761a,a49764a,a49767a,a49768a,a49771a,a49774a,a49775a,a49776a,a49780a,a49781a,a49784a,a49787a,a49788a,a49789a,a49792a,a49795a,a49796a,a49799a,a49802a,a49803a,a49804a,a49808a,a49809a,a49812a,a49815a,a49816a,a49817a,a49820a,a49823a,a49824a,a49827a,a49830a,a49831a,a49832a,a49836a,a49837a,a49840a,a49843a,a49844a,a49845a,a49848a,a49851a,a49852a,a49855a,a49858a,a49859a,a49860a,a49864a,a49865a,a49868a,a49871a,a49872a,a49873a,a49876a,a49879a,a49880a,a49883a,a49886a,a49887a,a49888a,a49892a,a49893a,a49896a,a49899a,a49900a,a49901a,a49904a,a49907a,a49908a,a49911a,a49914a,a49915a,a49916a,a49920a,a49921a,a49924a,a49927a,a49928a,a49929a,a49932a,a49935a,a49936a,a49939a,a49942a,a49943a,a49944a,a49948a,a49949a,a49952a,a49955a,a49956a,a49957a,a49960a,a49963a,a49964a,a49967a,a49970a,a49971a,a49972a,a49976a,a49977a,a49980a,a49983a,a49984a,a49985a,a49988a,a49991a,a49992a,a49995a,a49998a,a49999a,a50000a,a50004a,a50005a,a50008a,a50011a,a50012a,a50013a,a50016a,a50019a,a50020a,a50023a,a50026a,a50027a,a50028a,a50032a,a50033a,a50036a,a50039a,a50040a,a50041a,a50044a,a50047a,a50048a,a50051a,a50054a,a50055a,a50056a,a50060a,a50061a,a50064a,a50067a,a50068a,a50069a,a50072a,a50075a,a50076a,a50079a,a50082a,a50083a,a50084a,a50088a,a50089a,a50092a,a50095a,a50096a,a50097a,a50100a,a50103a,a50104a,a50107a,a50110a,a50111a,a50112a,a50116a,a50117a,a50120a,a50123a,a50124a,a50125a,a50128a,a50131a,a50132a,a50135a,a50138a,a50139a,a50140a,a50144a,a50145a,a50148a,a50151a,a50152a,a50153a,a50156a,a50159a,a50160a,a50163a,a50166a,a50167a,a50168a,a50172a,a50173a,a50176a,a50179a,a50180a,a50181a,a50184a,a50187a,a50188a,a50191a,a50194a,a50195a,a50196a,a50200a,a50201a,a50204a,a50207a,a50208a,a50209a,a50212a,a50215a,a50216a,a50219a,a50222a,a50223a,a50224a,a50228a,a50229a,a50232a,a50235a,a50236a,a50237a,a50240a,a50243a,a50244a,a50247a,a50250a,a50251a,a50252a,a50256a,a50257a,a50260a,a50263a,a50264a,a50265a,a50268a,a50271a,a50272a,a50275a,a50278a,a50279a,a50280a,a50284a,a50285a,a50288a,a50291a,a50292a,a50293a,a50296a,a50299a,a50300a,a50303a,a50306a,a50307a,a50308a,a50312a,a50313a,a50316a,a50319a,a50320a,a50321a,a50324a,a50327a,a50328a,a50331a,a50334a,a50335a,a50336a,a50340a,a50341a,a50344a,a50347a,a50348a,a50349a,a50352a,a50355a,a50356a,a50359a,a50362a,a50363a,a50364a,a50368a,a50369a,a50372a,a50375a,a50376a,a50377a,a50380a,a50383a,a50384a,a50387a,a50390a,a50391a,a50392a,a50396a,a50397a,a50400a,a50403a,a50404a,a50405a,a50408a,a50411a,a50412a,a50415a,a50418a,a50419a,a50420a,a50424a,a50425a,a50428a,a50431a,a50432a,a50433a,a50436a,a50439a,a50440a,a50443a,a50446a,a50447a,a50448a,a50452a,a50453a,a50456a,a50459a,a50460a,a50461a,a50464a,a50467a,a50468a,a50471a,a50474a,a50475a,a50476a,a50480a,a50481a,a50484a,a50487a,a50488a,a50489a,a50492a,a50495a,a50496a,a50499a,a50502a,a50503a,a50504a,a50508a,a50509a,a50512a,a50515a,a50516a,a50517a,a50520a,a50523a,a50524a,a50527a,a50530a,a50531a,a50532a,a50536a,a50537a,a50540a,a50543a,a50544a,a50545a,a50548a,a50551a,a50552a,a50555a,a50558a,a50559a,a50560a,a50564a,a50565a,a50568a,a50571a,a50572a,a50573a,a50576a,a50579a,a50580a,a50583a,a50586a,a50587a,a50588a,a50592a,a50593a,a50596a,a50599a,a50600a,a50601a,a50604a,a50607a,a50608a,a50611a,a50614a,a50615a,a50616a,a50620a,a50621a,a50624a,a50627a,a50628a,a50629a,a50632a,a50635a,a50636a,a50639a,a50642a,a50643a,a50644a,a50648a,a50649a,a50652a,a50655a,a50656a,a50657a,a50660a,a50663a,a50664a,a50667a,a50670a,a50671a,a50672a,a50676a,a50677a,a50680a,a50683a,a50684a,a50685a,a50688a,a50691a,a50692a,a50695a,a50698a,a50699a,a50700a,a50704a,a50705a,a50708a,a50711a,a50712a,a50713a,a50716a,a50719a,a50720a,a50723a,a50726a,a50727a,a50728a,a50732a,a50733a,a50736a,a50739a,a50740a,a50741a,a50744a,a50747a,a50748a,a50751a,a50754a,a50755a,a50756a,a50760a,a50761a,a50764a,a50767a,a50768a,a50769a,a50772a,a50775a,a50776a,a50779a,a50782a,a50783a,a50784a,a50788a,a50789a,a50792a,a50795a,a50796a,a50797a,a50800a,a50803a,a50804a,a50807a,a50810a,a50811a,a50812a,a50816a,a50817a,a50820a,a50823a,a50824a,a50825a,a50828a,a50831a,a50832a,a50835a,a50838a,a50839a,a50840a,a50844a,a50845a,a50848a,a50851a,a50852a,a50853a,a50856a,a50859a,a50860a,a50863a,a50866a,a50867a,a50868a,a50872a,a50873a,a50876a,a50879a,a50880a,a50881a,a50884a,a50887a,a50888a,a50891a,a50894a,a50895a,a50896a,a50900a,a50901a,a50904a,a50907a,a50908a,a50909a,a50912a,a50915a,a50916a,a50919a,a50922a,a50923a,a50924a,a50928a,a50929a,a50932a,a50935a,a50936a,a50937a,a50940a,a50943a,a50944a,a50947a,a50950a,a50951a,a50952a,a50956a,a50957a,a50960a,a50963a,a50964a,a50965a,a50968a,a50971a,a50972a,a50975a,a50978a,a50979a,a50980a,a50984a,a50985a,a50988a,a50991a,a50992a,a50993a,a50996a,a50999a,a51000a,a51003a,a51006a,a51007a,a51008a,a51012a,a51013a,a51016a,a51019a,a51020a,a51021a,a51024a,a51027a,a51028a,a51031a,a51034a,a51035a,a51036a,a51040a,a51041a,a51044a,a51047a,a51048a,a51049a,a51052a,a51055a,a51056a,a51059a,a51062a,a51063a,a51064a,a51068a,a51069a,a51072a,a51075a,a51076a,a51077a,a51080a,a51083a,a51084a,a51087a,a51090a,a51091a,a51092a,a51096a,a51097a,a51100a,a51103a,a51104a,a51105a,a51108a,a51111a,a51112a,a51115a,a51118a,a51119a,a51120a,a51124a,a51125a,a51128a,a51131a,a51132a,a51133a,a51136a,a51139a,a51140a,a51143a,a51146a,a51147a,a51148a,a51152a,a51153a,a51156a,a51159a,a51160a,a51161a,a51164a,a51167a,a51168a,a51171a,a51174a,a51175a,a51176a,a51180a,a51181a,a51184a,a51187a,a51188a,a51189a,a51192a,a51195a,a51196a,a51199a,a51202a,a51203a,a51204a,a51208a,a51209a,a51212a,a51215a,a51216a,a51217a,a51220a,a51223a,a51224a,a51227a,a51230a,a51231a,a51232a,a51236a,a51237a,a51240a,a51243a,a51244a,a51245a,a51248a,a51251a,a51252a,a51255a,a51258a,a51259a,a51260a,a51264a,a51265a,a51268a,a51271a,a51272a,a51273a,a51276a,a51279a,a51280a,a51283a,a51286a,a51287a,a51288a,a51292a,a51293a,a51296a,a51299a,a51300a,a51301a,a51304a,a51307a,a51308a,a51311a,a51314a,a51315a,a51316a,a51320a,a51321a,a51324a,a51327a,a51328a,a51329a,a51332a,a51335a,a51336a,a51339a,a51342a,a51343a,a51344a,a51348a,a51349a,a51352a,a51355a,a51356a,a51357a,a51360a,a51363a,a51364a,a51367a,a51370a,a51371a,a51372a,a51376a,a51377a,a51380a,a51383a,a51384a,a51385a,a51388a,a51391a,a51392a,a51395a,a51398a,a51399a,a51400a,a51404a,a51405a,a51408a,a51411a,a51412a,a51413a,a51416a,a51419a,a51420a,a51423a,a51426a,a51427a,a51428a,a51432a,a51433a,a51436a,a51439a,a51440a,a51441a,a51444a,a51447a,a51448a,a51451a,a51454a,a51455a,a51456a,a51460a,a51461a,a51464a,a51467a,a51468a,a51469a,a51472a,a51475a,a51476a,a51479a,a51482a,a51483a,a51484a,a51488a,a51489a,a51492a,a51495a,a51496a,a51497a,a51500a,a51503a,a51504a,a51507a,a51510a,a51511a,a51512a,a51516a,a51517a,a51520a,a51523a,a51524a,a51525a,a51528a,a51531a,a51532a,a51535a,a51538a,a51539a,a51540a,a51544a,a51545a,a51548a,a51551a,a51552a,a51553a,a51556a,a51559a,a51560a,a51563a,a51566a,a51567a,a51568a,a51572a,a51573a,a51576a,a51579a,a51580a,a51581a,a51584a,a51587a,a51588a,a51591a,a51594a,a51595a,a51596a,a51600a,a51601a,a51604a,a51607a,a51608a,a51609a,a51612a,a51615a,a51616a,a51619a,a51622a,a51623a,a51624a,a51628a,a51629a,a51632a,a51635a,a51636a,a51637a,a51640a,a51643a,a51644a,a51647a,a51650a,a51651a,a51652a,a51656a,a51657a,a51660a,a51663a,a51664a,a51665a,a51668a,a51671a,a51672a,a51675a,a51678a,a51679a,a51680a,a51684a,a51685a,a51688a,a51691a,a51692a,a51693a,a51696a,a51699a,a51700a,a51703a,a51706a,a51707a,a51708a,a51712a,a51713a,a51716a,a51719a,a51720a,a51721a,a51724a,a51727a,a51728a,a51731a,a51734a,a51735a,a51736a,a51740a,a51741a,a51744a,a51747a,a51748a,a51749a,a51752a,a51755a,a51756a,a51759a,a51762a,a51763a,a51764a,a51768a,a51769a,a51772a,a51775a,a51776a,a51777a,a51780a,a51783a,a51784a,a51787a,a51790a,a51791a,a51792a,a51796a,a51797a,a51800a,a51803a,a51804a,a51805a,a51808a,a51811a,a51812a,a51815a,a51818a,a51819a,a51820a,a51824a,a51825a,a51828a,a51831a,a51832a,a51833a,a51836a,a51839a,a51840a,a51843a,a51846a,a51847a,a51848a,a51852a,a51853a,a51856a,a51859a,a51860a,a51861a,a51864a,a51867a,a51868a,a51871a,a51874a,a51875a,a51876a,a51880a,a51881a,a51884a,a51887a,a51888a,a51889a,a51892a,a51895a,a51896a,a51899a,a51902a,a51903a,a51904a,a51908a,a51909a,a51912a,a51915a,a51916a,a51917a,a51920a,a51923a,a51924a,a51927a,a51930a,a51931a,a51932a,a51936a,a51937a,a51940a,a51943a,a51944a,a51945a,a51948a,a51951a,a51952a,a51955a,a51958a,a51959a,a51960a,a51964a,a51965a,a51968a,a51971a,a51972a,a51973a,a51976a,a51979a,a51980a,a51983a,a51986a,a51987a,a51988a,a51992a,a51993a,a51996a,a51999a,a52000a,a52001a,a52004a,a52007a,a52008a,a52011a,a52014a,a52015a,a52016a,a52020a,a52021a,a52024a,a52027a,a52028a,a52029a,a52032a,a52035a,a52036a,a52039a,a52042a,a52043a,a52044a,a52048a,a52049a,a52052a,a52055a,a52056a,a52057a,a52060a,a52063a,a52064a,a52067a,a52070a,a52071a,a52072a,a52076a,a52077a,a52080a,a52083a,a52084a,a52085a,a52088a,a52091a,a52092a,a52095a,a52098a,a52099a,a52100a,a52104a,a52105a,a52108a,a52111a,a52112a,a52113a,a52116a,a52119a,a52120a,a52123a,a52126a,a52127a,a52128a,a52132a,a52133a,a52136a,a52139a,a52140a,a52141a,a52144a,a52147a,a52148a,a52151a,a52154a,a52155a,a52156a,a52160a,a52161a,a52164a,a52167a,a52168a,a52169a,a52172a,a52175a,a52176a,a52179a,a52182a,a52183a,a52184a,a52188a,a52189a,a52192a,a52195a,a52196a,a52197a,a52200a,a52203a,a52204a,a52207a,a52210a,a52211a,a52212a,a52216a,a52217a,a52220a,a52223a,a52224a,a52225a,a52228a,a52231a,a52232a,a52235a,a52238a,a52239a,a52240a,a52244a,a52245a,a52248a,a52251a,a52252a,a52253a,a52256a,a52259a,a52260a,a52263a,a52266a,a52267a,a52268a,a52272a,a52273a,a52276a,a52279a,a52280a,a52281a,a52284a,a52287a,a52288a,a52291a,a52294a,a52295a,a52296a,a52300a,a52301a,a52304a,a52307a,a52308a,a52309a,a52312a,a52315a,a52316a,a52319a,a52322a,a52323a,a52324a,a52328a,a52329a,a52332a,a52335a,a52336a,a52337a,a52340a,a52343a,a52344a,a52347a,a52350a,a52351a,a52352a,a52356a,a52357a,a52360a,a52363a,a52364a,a52365a,a52368a,a52371a,a52372a,a52375a,a52378a,a52379a,a52380a,a52384a,a52385a,a52388a,a52391a,a52392a,a52393a,a52396a,a52399a,a52400a,a52403a,a52406a,a52407a,a52408a,a52412a,a52413a,a52416a,a52419a,a52420a,a52421a,a52424a,a52427a,a52428a,a52431a,a52434a,a52435a,a52436a,a52440a,a52441a,a52444a,a52447a,a52448a,a52449a,a52452a,a52455a,a52456a,a52459a,a52462a,a52463a,a52464a,a52468a,a52469a,a52472a,a52475a,a52476a,a52477a,a52480a,a52483a,a52484a,a52487a,a52490a,a52491a,a52492a,a52496a,a52497a,a52500a,a52503a,a52504a,a52505a,a52508a,a52511a,a52512a,a52515a,a52518a,a52519a,a52520a,a52524a,a52525a,a52528a,a52531a,a52532a,a52533a,a52536a,a52539a,a52540a,a52543a,a52546a,a52547a,a52548a,a52552a,a52553a,a52556a,a52559a,a52560a,a52561a,a52564a,a52567a,a52568a,a52571a,a52574a,a52575a,a52576a,a52580a,a52581a,a52584a,a52587a,a52588a,a52589a,a52592a,a52595a,a52596a,a52599a,a52602a,a52603a,a52604a,a52608a,a52609a,a52612a,a52615a,a52616a,a52617a,a52620a,a52623a,a52624a,a52627a,a52630a,a52631a,a52632a,a52636a,a52637a,a52640a,a52643a,a52644a,a52645a,a52648a,a52651a,a52652a,a52655a,a52658a,a52659a,a52660a,a52664a,a52665a,a52668a,a52671a,a52672a,a52673a,a52676a,a52679a,a52680a,a52683a,a52686a,a52687a,a52688a,a52692a,a52693a,a52696a,a52699a,a52700a,a52701a,a52704a,a52707a,a52708a,a52711a,a52714a,a52715a,a52716a,a52720a,a52721a,a52724a,a52727a,a52728a,a52729a,a52732a,a52735a,a52736a,a52739a,a52742a,a52743a,a52744a,a52748a,a52749a,a52752a,a52755a,a52756a,a52757a,a52760a,a52763a,a52764a,a52767a,a52770a,a52771a,a52772a,a52776a,a52777a,a52780a,a52783a,a52784a,a52785a,a52788a,a52791a,a52792a,a52795a,a52798a,a52799a,a52800a,a52804a,a52805a,a52808a,a52811a,a52812a,a52813a,a52816a,a52819a,a52820a,a52823a,a52826a,a52827a,a52828a,a52832a,a52833a,a52836a,a52839a,a52840a,a52841a,a52844a,a52847a,a52848a,a52851a,a52854a,a52855a,a52856a,a52860a,a52861a,a52864a,a52867a,a52868a,a52869a,a52872a,a52875a,a52876a,a52879a,a52882a,a52883a,a52884a,a52888a,a52889a,a52892a,a52895a,a52896a,a52897a,a52900a,a52903a,a52904a,a52907a,a52910a,a52911a,a52912a,a52916a,a52917a,a52920a,a52923a,a52924a,a52925a,a52928a,a52931a,a52932a,a52935a,a52938a,a52939a,a52940a,a52944a,a52945a,a52948a,a52951a,a52952a,a52953a,a52956a,a52959a,a52960a,a52963a,a52966a,a52967a,a52968a,a52972a,a52973a,a52976a,a52979a,a52980a,a52981a,a52984a,a52987a,a52988a,a52991a,a52994a,a52995a,a52996a,a53000a,a53001a,a53004a,a53007a,a53008a,a53009a,a53012a,a53015a,a53016a,a53019a,a53022a,a53023a,a53024a,a53028a,a53029a,a53032a,a53035a,a53036a,a53037a,a53040a,a53043a,a53044a,a53047a,a53050a,a53051a,a53052a,a53056a,a53057a,a53060a,a53063a,a53064a,a53065a,a53068a,a53071a,a53072a,a53075a,a53078a,a53079a,a53080a,a53084a,a53085a,a53088a,a53091a,a53092a,a53093a,a53096a,a53099a,a53100a,a53103a,a53106a,a53107a,a53108a,a53112a,a53113a,a53116a,a53119a,a53120a,a53121a,a53124a,a53127a,a53128a,a53131a,a53134a,a53135a,a53136a,a53140a,a53141a,a53144a,a53147a,a53148a,a53149a,a53152a,a53155a,a53156a,a53159a,a53162a,a53163a,a53164a,a53168a,a53169a,a53172a,a53175a,a53176a,a53177a,a53180a,a53183a,a53184a,a53187a,a53190a,a53191a,a53192a,a53196a,a53197a,a53200a,a53203a,a53204a,a53205a,a53208a,a53211a,a53212a,a53215a,a53218a,a53219a,a53220a,a53224a,a53225a,a53228a,a53231a,a53232a,a53233a,a53236a,a53239a,a53240a,a53243a,a53246a,a53247a,a53248a,a53252a,a53253a,a53256a,a53259a,a53260a,a53261a,a53264a,a53267a,a53268a,a53271a,a53274a,a53275a,a53276a,a53280a,a53281a,a53284a,a53287a,a53288a,a53289a,a53292a,a53295a,a53296a,a53299a,a53302a,a53303a,a53304a,a53308a,a53309a,a53312a,a53315a,a53316a,a53317a,a53320a,a53323a,a53324a,a53327a,a53330a,a53331a,a53332a,a53336a,a53337a,a53340a,a53343a,a53344a,a53345a,a53348a,a53351a,a53352a,a53355a,a53358a,a53359a,a53360a,a53364a,a53365a,a53368a,a53371a,a53372a,a53373a,a53376a,a53379a,a53380a,a53383a,a53386a,a53387a,a53388a,a53392a,a53393a,a53396a,a53399a,a53400a,a53401a,a53404a,a53407a,a53408a,a53411a,a53414a,a53415a,a53416a,a53420a,a53421a,a53424a,a53427a,a53428a,a53429a,a53432a,a53435a,a53436a,a53439a,a53442a,a53443a,a53444a,a53448a,a53449a,a53452a,a53455a,a53456a,a53457a,a53460a,a53463a,a53464a,a53467a,a53470a,a53471a,a53472a,a53476a,a53477a,a53480a,a53483a,a53484a,a53485a,a53488a,a53491a,a53492a,a53495a,a53498a,a53499a,a53500a,a53504a,a53505a,a53508a,a53511a,a53512a,a53513a,a53516a,a53519a,a53520a,a53523a,a53526a,a53527a,a53528a,a53532a,a53533a,a53536a,a53539a,a53540a,a53541a,a53544a,a53547a,a53548a,a53551a,a53554a,a53555a,a53556a,a53560a,a53561a,a53564a,a53567a,a53568a,a53569a,a53572a,a53575a,a53576a,a53579a,a53582a,a53583a,a53584a,a53588a,a53589a,a53592a,a53595a,a53596a,a53597a,a53600a,a53603a,a53604a,a53607a,a53610a,a53611a,a53612a,a53616a,a53617a,a53620a,a53623a,a53624a,a53625a,a53628a,a53631a,a53632a,a53635a,a53638a,a53639a,a53640a,a53644a,a53645a,a53648a,a53651a,a53652a,a53653a,a53656a,a53659a,a53660a,a53663a,a53666a,a53667a,a53668a,a53672a,a53673a,a53676a,a53679a,a53680a,a53681a,a53684a,a53687a,a53688a,a53691a,a53694a,a53695a,a53696a,a53700a,a53701a,a53704a,a53707a,a53708a,a53709a,a53712a,a53715a,a53716a,a53719a,a53722a,a53723a,a53724a,a53728a,a53729a,a53732a,a53735a,a53736a,a53737a,a53740a,a53743a,a53744a,a53747a,a53750a,a53751a,a53752a,a53756a,a53757a,a53760a,a53763a,a53764a,a53765a,a53768a,a53771a,a53772a,a53775a,a53778a,a53779a,a53780a,a53784a,a53785a,a53788a,a53791a,a53792a,a53793a,a53796a,a53799a,a53800a,a53803a,a53806a,a53807a,a53808a,a53812a,a53813a,a53816a,a53819a,a53820a,a53821a,a53824a,a53827a,a53828a,a53831a,a53834a,a53835a,a53836a,a53840a,a53841a,a53844a,a53847a,a53848a,a53849a,a53852a,a53855a,a53856a,a53859a,a53862a,a53863a,a53864a,a53868a,a53869a,a53872a,a53875a,a53876a,a53877a,a53880a,a53883a,a53884a,a53887a,a53890a,a53891a,a53892a,a53896a,a53897a,a53900a,a53903a,a53904a,a53905a,a53908a,a53911a,a53912a,a53915a,a53918a,a53919a,a53920a,a53924a,a53925a,a53928a,a53931a,a53932a,a53933a,a53936a,a53939a,a53940a,a53943a,a53946a,a53947a,a53948a,a53952a,a53953a,a53956a,a53959a,a53960a,a53961a,a53964a,a53967a,a53968a,a53971a,a53974a,a53975a,a53976a,a53980a,a53981a,a53984a,a53987a,a53988a,a53989a,a53992a,a53995a,a53996a,a53999a,a54002a,a54003a,a54004a,a54008a,a54009a,a54012a,a54015a,a54016a,a54017a,a54020a,a54023a,a54024a,a54027a,a54030a,a54031a,a54032a,a54036a,a54037a,a54040a,a54043a,a54044a,a54045a,a54048a,a54051a,a54052a,a54055a,a54058a,a54059a,a54060a,a54064a,a54065a,a54068a,a54071a,a54072a,a54073a,a54076a,a54079a,a54080a,a54083a,a54086a,a54087a,a54088a,a54092a,a54093a,a54096a,a54099a,a54100a,a54101a,a54104a,a54107a,a54108a,a54111a,a54114a,a54115a,a54116a,a54120a,a54121a,a54124a,a54127a,a54128a,a54129a,a54132a,a54135a,a54136a,a54139a,a54142a,a54143a,a54144a,a54148a,a54149a,a54152a,a54155a,a54156a,a54157a,a54160a,a54163a,a54164a,a54167a,a54170a,a54171a,a54172a,a54176a,a54177a,a54180a,a54183a,a54184a,a54185a,a54188a,a54191a,a54192a,a54195a,a54198a,a54199a,a54200a,a54204a,a54205a,a54208a,a54211a,a54212a,a54213a,a54216a,a54219a,a54220a,a54223a,a54226a,a54227a,a54228a,a54232a,a54233a,a54236a,a54239a,a54240a,a54241a,a54244a,a54247a,a54248a,a54251a,a54254a,a54255a,a54256a,a54260a,a54261a,a54264a,a54267a,a54268a,a54269a,a54272a,a54275a,a54276a,a54279a,a54282a,a54283a,a54284a,a54288a,a54289a,a54292a,a54295a,a54296a,a54297a,a54300a,a54303a,a54304a,a54307a,a54310a,a54311a,a54312a,a54316a,a54317a,a54320a,a54323a,a54324a,a54325a,a54328a,a54331a,a54332a,a54335a,a54338a,a54339a,a54340a,a54344a,a54345a,a54348a,a54351a,a54352a,a54353a,a54356a,a54359a,a54360a,a54363a,a54366a,a54367a,a54368a,a54372a,a54373a,a54376a,a54379a,a54380a,a54381a,a54384a,a54387a,a54388a,a54391a,a54394a,a54395a,a54396a,a54400a,a54401a,a54404a,a54407a,a54408a,a54409a,a54412a,a54415a,a54416a,a54419a,a54422a,a54423a,a54424a,a54428a,a54429a,a54432a,a54435a,a54436a,a54437a,a54440a,a54443a,a54444a,a54447a,a54450a,a54451a,a54452a,a54456a,a54457a,a54460a,a54463a,a54464a,a54465a,a54468a,a54471a,a54472a,a54475a,a54478a,a54479a,a54480a,a54484a,a54485a,a54488a,a54491a,a54492a,a54493a,a54496a,a54499a,a54500a,a54503a,a54506a,a54507a,a54508a,a54512a,a54513a,a54516a,a54519a,a54520a,a54521a,a54524a,a54527a,a54528a,a54531a,a54534a,a54535a,a54536a,a54540a,a54541a,a54544a,a54547a,a54548a,a54549a,a54552a,a54555a,a54556a,a54559a,a54562a,a54563a,a54564a,a54568a,a54569a,a54572a,a54575a,a54576a,a54577a,a54580a,a54583a,a54584a,a54587a,a54590a,a54591a,a54592a,a54596a,a54597a,a54600a,a54603a,a54604a,a54605a,a54608a,a54611a,a54612a,a54615a,a54618a,a54619a,a54620a,a54624a,a54625a,a54628a,a54631a,a54632a,a54633a,a54636a,a54639a,a54640a,a54643a,a54646a,a54647a,a54648a,a54652a,a54653a,a54656a,a54659a,a54660a,a54661a,a54664a,a54667a,a54668a,a54671a,a54674a,a54675a,a54676a,a54680a,a54681a,a54684a,a54687a,a54688a,a54689a,a54692a,a54695a,a54696a,a54699a,a54702a,a54703a,a54704a,a54708a,a54709a,a54712a,a54715a,a54716a,a54717a,a54720a,a54723a,a54724a,a54727a,a54730a,a54731a,a54732a,a54736a,a54737a,a54740a,a54743a,a54744a,a54745a,a54748a,a54751a,a54752a,a54755a,a54758a,a54759a,a54760a,a54764a,a54765a,a54768a,a54771a,a54772a,a54773a,a54776a,a54779a,a54780a,a54783a,a54786a,a54787a,a54788a,a54792a,a54793a,a54796a,a54799a,a54800a,a54801a,a54804a,a54807a,a54808a,a54811a,a54814a,a54815a,a54816a,a54820a,a54821a,a54824a,a54827a,a54828a,a54829a,a54832a,a54835a,a54836a,a54839a,a54842a,a54843a,a54844a,a54848a,a54849a,a54852a,a54855a,a54856a,a54857a,a54860a,a54863a,a54864a,a54867a,a54870a,a54871a,a54872a,a54876a,a54877a,a54880a,a54883a,a54884a,a54885a,a54888a,a54891a,a54892a,a54895a,a54898a,a54899a,a54900a,a54904a,a54905a,a54908a,a54911a,a54912a,a54913a,a54916a,a54919a,a54920a,a54923a,a54926a,a54927a,a54928a,a54932a,a54933a,a54936a,a54939a,a54940a,a54941a,a54944a,a54947a,a54948a,a54951a,a54954a,a54955a,a54956a,a54960a,a54961a,a54964a,a54967a,a54968a,a54969a,a54972a,a54975a,a54976a,a54979a,a54982a,a54983a,a54984a,a54988a,a54989a,a54992a,a54995a,a54996a,a54997a,a55000a,a55003a,a55004a,a55007a,a55010a,a55011a,a55012a,a55016a,a55017a,a55020a,a55023a,a55024a,a55025a,a55028a,a55031a,a55032a,a55035a,a55038a,a55039a,a55040a,a55044a,a55045a,a55048a,a55051a,a55052a,a55053a,a55056a,a55059a,a55060a,a55063a,a55066a,a55067a,a55068a,a55072a,a55073a,a55076a,a55079a,a55080a,a55081a,a55084a,a55087a,a55088a,a55091a,a55094a,a55095a,a55096a,a55100a,a55101a,a55104a,a55107a,a55108a,a55109a,a55112a,a55115a,a55116a,a55119a,a55122a,a55123a,a55124a,a55128a,a55129a,a55132a,a55135a,a55136a,a55137a,a55140a,a55143a,a55144a,a55147a,a55150a,a55151a,a55152a,a55156a,a55157a,a55160a,a55163a,a55164a,a55165a,a55168a,a55171a,a55172a,a55175a,a55178a,a55179a,a55180a,a55184a,a55185a,a55188a,a55191a,a55192a,a55193a,a55196a,a55199a,a55200a,a55203a,a55206a,a55207a,a55208a,a55212a,a55213a,a55216a,a55219a,a55220a,a55221a,a55224a,a55227a,a55228a,a55231a,a55234a,a55235a,a55236a,a55240a,a55241a,a55244a,a55247a,a55248a,a55249a,a55252a,a55255a,a55256a,a55259a,a55262a,a55263a,a55264a,a55268a,a55269a,a55272a,a55275a,a55276a,a55277a,a55280a,a55283a,a55284a,a55287a,a55290a,a55291a,a55292a,a55296a,a55297a,a55300a,a55303a,a55304a,a55305a,a55308a,a55311a,a55312a,a55315a,a55318a,a55319a,a55320a,a55324a,a55325a,a55328a,a55331a,a55332a,a55333a,a55336a,a55339a,a55340a,a55343a,a55346a,a55347a,a55348a,a55352a,a55353a,a55356a,a55359a,a55360a,a55361a,a55364a,a55367a,a55368a,a55371a,a55374a,a55375a,a55376a,a55380a,a55381a,a55384a,a55387a,a55388a,a55389a,a55392a,a55395a,a55396a,a55399a,a55402a,a55403a,a55404a,a55408a,a55409a,a55412a,a55415a,a55416a,a55417a,a55420a,a55423a,a55424a,a55427a,a55430a,a55431a,a55432a,a55436a,a55437a,a55440a,a55443a,a55444a,a55445a,a55448a,a55451a,a55452a,a55455a,a55458a,a55459a,a55460a,a55464a,a55465a,a55468a,a55471a,a55472a,a55473a,a55476a,a55479a,a55480a,a55483a,a55486a,a55487a,a55488a,a55492a,a55493a,a55496a,a55499a,a55500a,a55501a,a55504a,a55507a,a55508a,a55511a,a55514a,a55515a,a55516a,a55520a,a55521a,a55524a,a55527a,a55528a,a55529a,a55532a,a55535a,a55536a,a55539a,a55542a,a55543a,a55544a,a55548a,a55549a,a55552a,a55555a,a55556a,a55557a,a55560a,a55563a,a55564a,a55567a,a55570a,a55571a,a55572a,a55576a,a55577a,a55580a,a55583a,a55584a,a55585a,a55588a,a55591a,a55592a,a55595a,a55598a,a55599a,a55600a,a55604a,a55605a,a55608a,a55611a,a55612a,a55613a,a55616a,a55619a,a55620a,a55623a,a55626a,a55627a,a55628a,a55632a,a55633a,a55636a,a55639a,a55640a,a55641a,a55644a,a55647a,a55648a,a55651a,a55654a,a55655a,a55656a,a55660a,a55661a,a55664a,a55667a,a55668a,a55669a,a55672a,a55675a,a55676a,a55679a,a55682a,a55683a,a55684a,a55688a,a55689a,a55692a,a55695a,a55696a,a55697a,a55700a,a55703a,a55704a,a55707a,a55710a,a55711a,a55712a,a55716a,a55717a,a55720a,a55723a,a55724a,a55725a,a55728a,a55731a,a55732a,a55735a,a55738a,a55739a,a55740a,a55744a,a55745a,a55748a,a55751a,a55752a,a55753a,a55756a,a55759a,a55760a,a55763a,a55766a,a55767a,a55768a,a55772a,a55773a,a55776a,a55779a,a55780a,a55781a,a55784a,a55787a,a55788a,a55791a,a55794a,a55795a,a55796a,a55800a,a55801a,a55804a,a55807a,a55808a,a55809a,a55812a,a55815a,a55816a,a55819a,a55822a,a55823a,a55824a,a55828a,a55829a,a55832a,a55835a,a55836a,a55837a,a55840a,a55843a,a55844a,a55847a,a55850a,a55851a,a55852a,a55856a,a55857a,a55860a,a55863a,a55864a,a55865a,a55868a,a55871a,a55872a,a55875a,a55878a,a55879a,a55880a,a55884a,a55885a,a55888a,a55891a,a55892a,a55893a,a55896a,a55899a,a55900a,a55903a,a55906a,a55907a,a55908a,a55912a,a55913a,a55916a,a55919a,a55920a,a55921a,a55924a,a55927a,a55928a,a55931a,a55934a,a55935a,a55936a,a55940a,a55941a,a55944a,a55947a,a55948a,a55949a,a55952a,a55955a,a55956a,a55959a,a55962a,a55963a,a55964a,a55968a,a55969a,a55972a,a55975a,a55976a,a55977a,a55980a,a55983a,a55984a,a55987a,a55990a,a55991a,a55992a,a55996a,a55997a,a56000a,a56003a,a56004a,a56005a,a56008a,a56011a,a56012a,a56015a,a56018a,a56019a,a56020a,a56024a,a56025a,a56028a,a56031a,a56032a,a56033a,a56036a,a56039a,a56040a,a56043a,a56046a,a56047a,a56048a,a56052a,a56053a,a56056a,a56059a,a56060a,a56061a,a56064a,a56067a,a56068a,a56071a,a56074a,a56075a,a56076a,a56080a,a56081a,a56084a,a56087a,a56088a,a56089a,a56092a,a56095a,a56096a,a56099a,a56102a,a56103a,a56104a,a56108a,a56109a,a56112a,a56115a,a56116a,a56117a,a56120a,a56123a,a56124a,a56127a,a56130a,a56131a,a56132a,a56136a,a56137a,a56140a,a56143a,a56144a,a56145a,a56148a,a56151a,a56152a,a56155a,a56158a,a56159a,a56160a,a56164a,a56165a,a56168a,a56171a,a56172a,a56173a,a56176a,a56179a,a56180a,a56183a,a56186a,a56187a,a56188a,a56192a,a56193a,a56196a,a56199a,a56200a,a56201a,a56204a,a56207a,a56208a,a56211a,a56214a,a56215a,a56216a,a56220a,a56221a,a56224a,a56227a,a56228a,a56229a,a56232a,a56235a,a56236a,a56239a,a56242a,a56243a,a56244a,a56248a,a56249a,a56252a,a56255a,a56256a,a56257a,a56260a,a56263a,a56264a,a56267a,a56270a,a56271a,a56272a,a56276a,a56277a,a56280a,a56283a,a56284a,a56285a,a56288a,a56291a,a56292a,a56295a,a56298a,a56299a,a56300a,a56304a,a56305a,a56308a,a56311a,a56312a,a56313a,a56316a,a56319a,a56320a,a56323a,a56326a,a56327a,a56328a,a56332a,a56333a,a56336a,a56339a,a56340a,a56341a,a56344a,a56347a,a56348a,a56351a,a56354a,a56355a,a56356a,a56360a,a56361a,a56364a,a56367a,a56368a,a56369a,a56372a,a56375a,a56376a,a56379a,a56382a,a56383a,a56384a,a56388a,a56389a,a56392a,a56395a,a56396a,a56397a,a56400a,a56403a,a56404a,a56407a,a56410a,a56411a,a56412a,a56416a,a56417a,a56420a,a56423a,a56424a,a56425a,a56428a,a56431a,a56432a,a56435a,a56438a,a56439a,a56440a,a56444a,a56445a,a56448a,a56451a,a56452a,a56453a,a56456a,a56459a,a56460a,a56463a,a56466a,a56467a,a56468a,a56472a,a56473a,a56476a,a56479a,a56480a,a56481a,a56484a,a56487a,a56488a,a56491a,a56494a,a56495a,a56496a,a56500a,a56501a,a56504a,a56507a,a56508a,a56509a,a56512a,a56515a,a56516a,a56519a,a56522a,a56523a,a56524a,a56528a,a56529a,a56532a,a56535a,a56536a,a56537a,a56540a,a56543a,a56544a,a56547a,a56550a,a56551a,a56552a,a56556a,a56557a,a56560a,a56563a,a56564a,a56565a,a56568a,a56571a,a56572a,a56575a,a56578a,a56579a,a56580a,a56584a,a56585a,a56588a,a56591a,a56592a,a56593a,a56596a,a56599a,a56600a,a56603a,a56606a,a56607a,a56608a,a56612a,a56613a,a56616a,a56619a,a56620a,a56621a,a56624a,a56627a,a56628a,a56631a,a56634a,a56635a,a56636a,a56640a,a56641a,a56644a,a56647a,a56648a,a56649a,a56652a,a56655a,a56656a,a56659a,a56662a,a56663a,a56664a,a56668a,a56669a,a56672a,a56675a,a56676a,a56677a,a56680a,a56683a,a56684a,a56687a,a56690a,a56691a,a56692a,a56696a,a56697a,a56700a,a56703a,a56704a,a56705a,a56708a,a56711a,a56712a,a56715a,a56718a,a56719a,a56720a,a56724a,a56725a,a56728a,a56731a,a56732a,a56733a,a56736a,a56739a,a56740a,a56743a,a56746a,a56747a,a56748a,a56752a,a56753a,a56756a,a56759a,a56760a,a56761a,a56764a,a56767a,a56768a,a56771a,a56774a,a56775a,a56776a,a56780a,a56781a,a56784a,a56787a,a56788a,a56789a,a56792a,a56795a,a56796a,a56799a,a56802a,a56803a,a56804a,a56808a,a56809a,a56812a,a56815a,a56816a,a56817a,a56820a,a56823a,a56824a,a56827a,a56830a,a56831a,a56832a,a56836a,a56837a,a56840a,a56843a,a56844a,a56845a,a56848a,a56851a,a56852a,a56855a,a56858a,a56859a,a56860a,a56864a,a56865a,a56868a,a56871a,a56872a,a56873a,a56876a,a56879a,a56880a,a56883a,a56886a,a56887a,a56888a,a56892a,a56893a,a56896a,a56899a,a56900a,a56901a,a56904a,a56907a,a56908a,a56911a,a56914a,a56915a,a56916a,a56920a,a56921a,a56924a,a56927a,a56928a,a56929a,a56932a,a56935a,a56936a,a56939a,a56942a,a56943a,a56944a,a56948a,a56949a,a56952a,a56955a,a56956a,a56957a,a56960a,a56963a,a56964a,a56967a,a56970a,a56971a,a56972a,a56976a,a56977a,a56980a,a56983a,a56984a,a56985a,a56988a,a56991a,a56992a,a56995a,a56998a,a56999a,a57000a,a57004a,a57005a,a57008a,a57011a,a57012a,a57013a,a57016a,a57019a,a57020a,a57023a,a57026a,a57027a,a57028a,a57032a,a57033a,a57036a,a57039a,a57040a,a57041a,a57044a,a57047a,a57048a,a57051a,a57054a,a57055a,a57056a,a57060a,a57061a,a57064a,a57067a,a57068a,a57069a,a57072a,a57075a,a57076a,a57079a,a57082a,a57083a,a57084a,a57088a,a57089a,a57092a,a57095a,a57096a,a57097a,a57100a,a57103a,a57104a,a57107a,a57110a,a57111a,a57112a,a57116a,a57117a,a57120a,a57123a,a57124a,a57125a,a57128a,a57131a,a57132a,a57135a,a57138a,a57139a,a57140a,a57144a,a57145a,a57148a,a57151a,a57152a,a57153a,a57156a,a57159a,a57160a,a57163a,a57166a,a57167a,a57168a,a57172a,a57173a,a57176a,a57179a,a57180a,a57181a,a57184a,a57187a,a57188a,a57191a,a57194a,a57195a,a57196a,a57200a,a57201a,a57204a,a57207a,a57208a,a57209a,a57212a,a57215a,a57216a,a57219a,a57222a,a57223a,a57224a,a57228a,a57229a,a57232a,a57235a,a57236a,a57237a,a57240a,a57243a,a57244a,a57247a,a57250a,a57251a,a57252a,a57256a,a57257a,a57260a,a57263a,a57264a,a57265a,a57268a,a57271a,a57272a,a57275a,a57278a,a57279a,a57280a,a57284a,a57285a,a57288a,a57291a,a57292a,a57293a,a57296a,a57299a,a57300a,a57303a,a57306a,a57307a,a57308a,a57312a,a57313a,a57316a,a57319a,a57320a,a57321a,a57324a,a57327a,a57328a,a57331a,a57334a,a57335a,a57336a,a57340a,a57341a,a57344a,a57347a,a57348a,a57349a,a57352a,a57355a,a57356a,a57359a,a57362a,a57363a,a57364a,a57368a,a57369a,a57372a,a57375a,a57376a,a57377a,a57380a,a57383a,a57384a,a57387a,a57390a,a57391a,a57392a,a57396a,a57397a,a57400a,a57403a,a57404a,a57405a,a57408a,a57411a,a57412a,a57415a,a57418a,a57419a,a57420a,a57424a,a57425a,a57428a,a57431a,a57432a,a57433a,a57436a,a57439a,a57440a,a57443a,a57446a,a57447a,a57448a,a57452a,a57453a,a57456a,a57459a,a57460a,a57461a,a57464a,a57467a,a57468a,a57471a,a57474a,a57475a,a57476a,a57480a,a57481a,a57484a,a57487a,a57488a,a57489a,a57492a,a57495a,a57496a,a57499a,a57502a,a57503a,a57504a,a57508a,a57509a,a57512a,a57515a,a57516a,a57517a,a57520a,a57523a,a57524a,a57527a,a57530a,a57531a,a57532a,a57536a,a57537a,a57540a,a57543a,a57544a,a57545a,a57548a,a57551a,a57552a,a57555a,a57558a,a57559a,a57560a,a57564a,a57565a,a57568a,a57571a,a57572a,a57573a,a57576a,a57579a,a57580a,a57583a,a57586a,a57587a,a57588a,a57592a,a57593a,a57596a,a57599a,a57600a,a57601a,a57604a,a57607a,a57608a,a57611a,a57614a,a57615a,a57616a,a57620a,a57621a,a57624a,a57627a,a57628a,a57629a,a57632a,a57635a,a57636a,a57639a,a57642a,a57643a,a57644a,a57648a,a57649a,a57652a,a57655a,a57656a,a57657a,a57660a,a57663a,a57664a,a57667a,a57670a,a57671a,a57672a,a57676a,a57677a,a57680a,a57683a,a57684a,a57685a,a57688a,a57691a,a57692a,a57695a,a57698a,a57699a,a57700a,a57704a,a57705a,a57708a,a57711a,a57712a,a57713a,a57716a,a57719a,a57720a,a57723a,a57726a,a57727a,a57728a,a57731a,a57734a,a57735a,a57738a,a57741a,a57742a,a57743a,a57746a,a57749a,a57750a,a57753a,a57756a,a57757a,a57758a,a57761a,a57764a,a57765a,a57768a,a57771a,a57772a,a57773a,a57776a,a57779a,a57780a,a57783a,a57786a,a57787a,a57788a,a57791a,a57794a,a57795a,a57798a,a57801a,a57802a,a57803a,a57806a,a57809a,a57810a,a57813a,a57816a,a57817a,a57818a,a57821a,a57824a,a57825a,a57828a,a57831a,a57832a,a57833a,a57836a,a57839a,a57840a,a57843a,a57846a,a57847a,a57848a,a57851a,a57854a,a57855a,a57858a,a57861a,a57862a,a57863a,a57866a,a57869a,a57870a,a57873a,a57876a,a57877a,a57878a,a57881a,a57884a,a57885a,a57888a,a57891a,a57892a,a57893a,a57896a,a57899a,a57900a,a57903a,a57906a,a57907a,a57908a,a57911a,a57914a,a57915a,a57918a,a57921a,a57922a,a57923a,a57926a,a57929a,a57930a,a57933a,a57936a,a57937a,a57938a,a57941a,a57944a,a57945a,a57948a,a57951a,a57952a,a57953a,a57956a,a57959a,a57960a,a57963a,a57966a,a57967a,a57968a,a57971a,a57974a,a57975a,a57978a,a57981a,a57982a,a57983a,a57986a,a57989a,a57990a,a57993a,a57996a,a57997a,a57998a,a58001a,a58004a,a58005a,a58008a,a58011a,a58012a,a58013a,a58016a,a58019a,a58020a,a58023a,a58026a,a58027a,a58028a,a58031a,a58034a,a58035a,a58038a,a58041a,a58042a,a58043a,a58046a,a58049a,a58050a,a58053a,a58056a,a58057a,a58058a,a58061a,a58064a,a58065a,a58068a,a58071a,a58072a,a58073a,a58076a,a58079a,a58080a,a58083a,a58086a,a58087a,a58088a,a58091a,a58094a,a58095a,a58098a,a58101a,a58102a,a58103a,a58106a,a58109a,a58110a,a58113a,a58116a,a58117a,a58118a,a58121a,a58124a,a58125a,a58128a,a58131a,a58132a,a58133a,a58136a,a58139a,a58140a,a58143a,a58146a,a58147a,a58148a,a58151a,a58154a,a58155a,a58158a,a58161a,a58162a,a58163a,a58166a,a58169a,a58170a,a58173a,a58176a,a58177a,a58178a,a58181a,a58184a,a58185a,a58188a,a58191a,a58192a,a58193a,a58196a,a58199a,a58200a,a58203a,a58206a,a58207a,a58208a,a58211a,a58214a,a58215a,a58218a,a58221a,a58222a,a58223a,a58226a,a58229a,a58230a,a58233a,a58236a,a58237a,a58238a,a58241a,a58244a,a58245a,a58248a,a58251a,a58252a,a58253a,a58256a,a58259a,a58260a,a58263a,a58266a,a58267a,a58268a,a58271a,a58274a,a58275a,a58278a,a58281a,a58282a,a58283a,a58286a,a58289a,a58290a,a58293a,a58296a,a58297a,a58298a,a58301a,a58304a,a58305a,a58308a,a58311a,a58312a,a58313a,a58316a,a58319a,a58320a,a58323a,a58326a,a58327a,a58328a,a58331a,a58334a,a58335a,a58338a,a58341a,a58342a,a58343a,a58346a,a58349a,a58350a,a58353a,a58356a,a58357a,a58358a,a58361a,a58364a,a58365a,a58368a,a58371a,a58372a,a58373a,a58376a,a58379a,a58380a,a58383a,a58386a,a58387a,a58388a,a58391a,a58394a,a58395a,a58398a,a58401a,a58402a,a58403a,a58406a,a58409a,a58410a,a58413a,a58416a,a58417a,a58418a,a58421a,a58424a,a58425a,a58428a,a58431a,a58432a,a58433a,a58436a,a58439a,a58440a,a58443a,a58446a,a58447a,a58448a,a58451a,a58454a,a58455a,a58458a,a58461a,a58462a,a58463a,a58466a,a58469a,a58470a,a58473a,a58476a,a58477a,a58478a,a58481a,a58484a,a58485a,a58488a,a58491a,a58492a,a58493a,a58496a,a58499a,a58500a,a58503a,a58506a,a58507a,a58508a,a58511a,a58514a,a58515a,a58518a,a58521a,a58522a,a58523a,a58526a,a58529a,a58530a,a58533a,a58536a,a58537a,a58538a,a58541a,a58544a,a58545a,a58548a,a58551a,a58552a,a58553a,a58556a,a58559a,a58560a,a58563a,a58566a,a58567a,a58568a,a58571a,a58574a,a58575a,a58578a,a58581a,a58582a,a58583a,a58586a,a58589a,a58590a,a58593a,a58596a,a58597a,a58598a,a58601a,a58604a,a58605a,a58608a,a58611a,a58612a,a58613a,a58616a,a58619a,a58620a,a58623a,a58626a,a58627a,a58628a,a58631a,a58634a,a58635a,a58638a,a58641a,a58642a,a58643a,a58646a,a58649a,a58650a,a58653a,a58656a,a58657a,a58658a,a58661a,a58664a,a58665a,a58668a,a58671a,a58672a,a58673a,a58676a,a58679a,a58680a,a58683a,a58686a,a58687a,a58688a,a58691a,a58694a,a58695a,a58698a,a58701a,a58702a,a58703a,a58706a,a58709a,a58710a,a58713a,a58716a,a58717a,a58718a,a58721a,a58724a,a58725a,a58728a,a58731a,a58732a,a58733a,a58736a,a58739a,a58740a,a58743a,a58746a,a58747a,a58748a,a58751a,a58754a,a58755a,a58758a,a58761a,a58762a,a58763a,a58766a,a58769a,a58770a,a58773a,a58776a,a58777a,a58778a,a58781a,a58784a,a58785a,a58788a,a58791a,a58792a,a58793a,a58796a,a58799a,a58800a,a58803a,a58806a,a58807a,a58808a,a58811a,a58814a,a58815a,a58818a,a58821a,a58822a,a58823a,a58826a,a58829a,a58830a,a58833a,a58836a,a58837a,a58838a,a58841a,a58844a,a58845a,a58848a,a58851a,a58852a,a58853a,a58856a,a58859a,a58860a,a58863a,a58866a,a58867a,a58868a,a58871a,a58874a,a58875a,a58878a,a58881a,a58882a,a58883a,a58886a,a58889a,a58890a,a58893a,a58896a,a58897a,a58898a,a58901a,a58904a,a58905a,a58908a,a58911a,a58912a,a58913a,a58916a,a58919a,a58920a,a58923a,a58926a,a58927a,a58928a,a58931a,a58934a,a58935a,a58938a,a58941a,a58942a,a58943a,a58946a,a58949a,a58950a,a58953a,a58956a,a58957a,a58958a,a58961a,a58964a,a58965a,a58968a,a58971a,a58972a,a58973a,a58976a,a58979a,a58980a,a58983a,a58986a,a58987a,a58988a,a58991a,a58994a,a58995a,a58998a,a59001a,a59002a,a59003a,a59006a,a59009a,a59010a,a59013a,a59016a,a59017a,a59018a,a59021a,a59024a,a59025a,a59028a,a59031a,a59032a,a59033a,a59036a,a59039a,a59040a,a59043a,a59046a,a59047a,a59048a,a59051a,a59054a,a59055a,a59058a,a59061a,a59062a,a59063a,a59066a,a59069a,a59070a,a59073a,a59076a,a59077a,a59078a,a59081a,a59084a,a59085a,a59088a,a59091a,a59092a,a59093a,a59096a,a59099a,a59100a,a59103a,a59106a,a59107a,a59108a,a59111a,a59114a,a59115a,a59118a,a59121a,a59122a,a59123a,a59126a,a59129a,a59130a,a59133a,a59136a,a59137a,a59138a,a59141a,a59144a,a59145a,a59148a,a59151a,a59152a,a59153a,a59156a,a59159a,a59160a,a59163a,a59166a,a59167a,a59168a,a59171a,a59174a,a59175a,a59178a,a59181a,a59182a,a59183a,a59186a,a59189a,a59190a,a59193a,a59196a,a59197a,a59198a,a59201a,a59204a,a59205a,a59208a,a59211a,a59212a,a59213a,a59216a,a59219a,a59220a,a59223a,a59226a,a59227a,a59228a,a59231a,a59234a,a59235a,a59238a,a59241a,a59242a,a59243a,a59246a,a59249a,a59250a,a59253a,a59256a,a59257a,a59258a,a59261a,a59264a,a59265a,a59268a,a59271a,a59272a,a59273a,a59276a,a59279a,a59280a,a59283a,a59286a,a59287a,a59288a,a59291a,a59294a,a59295a,a59298a,a59301a,a59302a,a59303a,a59306a,a59309a,a59310a,a59313a,a59316a,a59317a,a59318a,a59321a,a59324a,a59325a,a59328a,a59331a,a59332a,a59333a,a59336a,a59339a,a59340a,a59343a,a59346a,a59347a,a59348a,a59351a,a59354a,a59355a,a59358a,a59361a,a59362a,a59363a,a59366a,a59369a,a59370a,a59373a,a59376a,a59377a,a59378a,a59381a,a59384a,a59385a,a59388a,a59391a,a59392a,a59393a,a59396a,a59399a,a59400a,a59403a,a59406a,a59407a,a59408a,a59411a,a59414a,a59415a,a59418a,a59421a,a59422a,a59423a,a59426a,a59429a,a59430a,a59433a,a59436a,a59437a,a59438a,a59441a,a59444a,a59445a,a59448a,a59451a,a59452a,a59453a,a59456a,a59459a,a59460a,a59463a,a59466a,a59467a,a59468a,a59471a,a59474a,a59475a,a59478a,a59481a,a59482a,a59483a,a59486a,a59489a,a59490a,a59493a,a59496a,a59497a,a59498a,a59501a,a59504a,a59505a,a59508a,a59511a,a59512a,a59513a,a59516a,a59519a,a59520a,a59523a,a59526a,a59527a,a59528a,a59531a,a59534a,a59535a,a59538a,a59541a,a59542a,a59543a,a59546a,a59549a,a59550a,a59553a,a59556a,a59557a,a59558a,a59561a,a59564a,a59565a,a59568a,a59571a,a59572a,a59573a,a59576a,a59579a,a59580a,a59583a,a59586a,a59587a,a59588a,a59591a,a59594a,a59595a,a59598a,a59601a,a59602a,a59603a,a59606a,a59609a,a59610a,a59613a,a59616a,a59617a,a59618a,a59621a,a59624a,a59625a,a59628a,a59631a,a59632a,a59633a,a59636a,a59639a,a59640a,a59643a,a59646a,a59647a,a59648a,a59651a,a59654a,a59655a,a59658a,a59661a,a59662a,a59663a,a59666a,a59669a,a59670a,a59673a,a59676a,a59677a,a59678a,a59681a,a59684a,a59685a,a59688a,a59691a,a59692a,a59693a,a59696a,a59699a,a59700a,a59703a,a59706a,a59707a,a59708a,a59711a,a59714a,a59715a,a59718a,a59721a,a59722a,a59723a,a59726a,a59729a,a59730a,a59733a,a59736a,a59737a,a59738a,a59741a,a59744a,a59745a,a59748a,a59751a,a59752a,a59753a,a59756a,a59759a,a59760a,a59763a,a59766a,a59767a,a59768a,a59771a,a59774a,a59775a,a59778a,a59781a,a59782a,a59783a,a59786a,a59789a,a59790a,a59793a,a59796a,a59797a,a59798a,a59801a,a59804a,a59805a,a59808a,a59811a,a59812a,a59813a,a59816a,a59819a,a59820a,a59823a,a59826a,a59827a,a59828a,a59831a,a59834a,a59835a,a59838a,a59841a,a59842a,a59843a,a59846a,a59849a,a59850a,a59853a,a59856a,a59857a,a59858a,a59861a,a59864a,a59865a,a59868a,a59871a,a59872a,a59873a,a59876a,a59879a,a59880a,a59883a,a59886a,a59887a,a59888a,a59891a,a59894a,a59895a,a59898a,a59901a,a59902a,a59903a,a59906a,a59909a,a59910a,a59913a,a59916a,a59917a,a59918a,a59921a,a59924a,a59925a,a59928a,a59931a,a59932a,a59933a,a59936a,a59939a,a59940a,a59943a,a59946a,a59947a,a59948a,a59951a,a59954a,a59955a,a59958a,a59961a,a59962a,a59963a,a59966a,a59969a,a59970a,a59973a,a59976a,a59977a,a59978a,a59981a,a59984a,a59985a,a59988a,a59991a,a59992a,a59993a,a59996a,a59999a,a60000a,a60003a,a60006a,a60007a,a60008a,a60011a,a60014a,a60015a,a60018a,a60021a,a60022a,a60023a,a60026a,a60029a,a60030a,a60033a,a60036a,a60037a,a60038a,a60041a,a60044a,a60045a,a60048a,a60051a,a60052a,a60053a,a60056a,a60059a,a60060a,a60063a,a60066a,a60067a,a60068a,a60071a,a60074a,a60075a,a60078a,a60081a,a60082a,a60083a,a60086a,a60089a,a60090a,a60093a,a60096a,a60097a,a60098a,a60101a,a60104a,a60105a,a60108a,a60111a,a60112a,a60113a,a60116a,a60119a,a60120a,a60123a,a60126a,a60127a,a60128a,a60131a,a60134a,a60135a,a60138a,a60141a,a60142a,a60143a,a60146a,a60149a,a60150a,a60153a,a60156a,a60157a,a60158a,a60161a,a60164a,a60165a,a60168a,a60171a,a60172a,a60173a,a60176a,a60179a,a60180a,a60183a,a60186a,a60187a,a60188a,a60191a,a60194a,a60195a,a60198a,a60201a,a60202a,a60203a,a60206a,a60209a,a60210a,a60213a,a60216a,a60217a,a60218a,a60221a,a60224a,a60225a,a60228a,a60231a,a60232a,a60233a,a60236a,a60239a,a60240a,a60243a,a60246a,a60247a,a60248a,a60251a,a60254a,a60255a,a60258a,a60261a,a60262a,a60263a,a60266a,a60269a,a60270a,a60273a,a60276a,a60277a,a60278a,a60281a,a60284a,a60285a,a60288a,a60291a,a60292a,a60293a,a60296a,a60299a,a60300a,a60303a,a60306a,a60307a,a60308a,a60311a,a60314a,a60315a,a60318a,a60321a,a60322a,a60323a,a60326a,a60329a,a60330a,a60333a,a60336a,a60337a,a60338a,a60341a,a60344a,a60345a,a60348a,a60351a,a60352a,a60353a,a60356a,a60359a,a60360a,a60363a,a60366a,a60367a,a60368a,a60371a,a60374a,a60375a,a60378a,a60381a,a60382a,a60383a,a60386a,a60389a,a60390a,a60393a,a60396a,a60397a,a60398a,a60401a,a60404a,a60405a,a60408a,a60411a,a60412a,a60413a,a60416a,a60419a,a60420a,a60423a,a60426a,a60427a,a60428a,a60431a,a60434a,a60435a,a60438a,a60441a,a60442a,a60443a,a60446a,a60449a,a60450a,a60453a,a60456a,a60457a,a60458a,a60461a,a60464a,a60465a,a60468a,a60471a,a60472a,a60473a,a60476a,a60479a,a60480a,a60483a,a60486a,a60487a,a60488a,a60491a,a60494a,a60495a,a60498a,a60501a,a60502a,a60503a,a60506a,a60509a,a60510a,a60513a,a60516a,a60517a,a60518a,a60521a,a60524a,a60525a,a60528a,a60531a,a60532a,a60533a,a60536a,a60539a,a60540a,a60543a,a60546a,a60547a,a60548a,a60551a,a60554a,a60555a,a60558a,a60561a,a60562a,a60563a,a60566a,a60569a,a60570a,a60573a,a60576a,a60577a,a60578a,a60581a,a60584a,a60585a,a60588a,a60591a,a60592a,a60593a,a60596a,a60599a,a60600a,a60603a,a60606a,a60607a,a60608a,a60611a,a60614a,a60615a,a60618a,a60621a,a60622a,a60623a,a60626a,a60629a,a60630a,a60633a,a60636a,a60637a,a60638a,a60641a,a60644a,a60645a,a60648a,a60651a,a60652a,a60653a,a60656a,a60659a,a60660a,a60663a,a60666a,a60667a,a60668a,a60671a,a60674a,a60675a,a60678a,a60681a,a60682a,a60683a,a60686a,a60689a,a60690a,a60693a,a60696a,a60697a,a60698a,a60701a,a60704a,a60705a,a60708a,a60711a,a60712a,a60713a,a60716a,a60719a,a60720a,a60723a,a60726a,a60727a,a60728a,a60731a,a60734a,a60735a,a60738a,a60741a,a60742a,a60743a,a60746a,a60749a,a60750a,a60753a,a60756a,a60757a,a60758a,a60761a,a60764a,a60765a,a60768a,a60771a,a60772a,a60773a,a60776a,a60779a,a60780a,a60783a,a60786a,a60787a,a60788a,a60791a,a60794a,a60795a,a60798a,a60801a,a60802a,a60803a,a60806a,a60809a,a60810a,a60813a,a60816a,a60817a,a60818a,a60821a,a60824a,a60825a,a60828a,a60831a,a60832a,a60833a,a60836a,a60839a,a60840a,a60843a,a60846a,a60847a,a60848a,a60851a,a60854a,a60855a,a60858a,a60861a,a60862a,a60863a,a60866a,a60869a,a60870a,a60873a,a60876a,a60877a,a60878a,a60881a,a60884a,a60885a,a60888a,a60891a,a60892a,a60893a,a60896a,a60899a,a60900a,a60903a,a60906a,a60907a,a60908a,a60911a,a60914a,a60915a,a60918a,a60921a,a60922a,a60923a,a60926a,a60929a,a60930a,a60933a,a60936a,a60937a,a60938a,a60941a,a60944a,a60945a,a60948a,a60951a,a60952a,a60953a,a60956a,a60959a,a60960a,a60963a,a60966a,a60967a,a60968a,a60971a,a60974a,a60975a,a60978a,a60981a,a60982a,a60983a,a60986a,a60989a,a60990a,a60993a,a60996a,a60997a,a60998a,a61001a,a61004a,a61005a,a61008a,a61011a,a61012a,a61013a,a61016a,a61019a,a61020a,a61023a,a61026a,a61027a,a61028a,a61031a,a61034a,a61035a,a61038a,a61041a,a61042a,a61043a,a61046a,a61049a,a61050a,a61053a,a61056a,a61057a,a61058a,a61061a,a61064a,a61065a,a61068a,a61071a,a61072a,a61073a,a61076a,a61079a,a61080a,a61083a,a61086a,a61087a,a61088a,a61091a,a61094a,a61095a,a61098a,a61101a,a61102a,a61103a,a61106a,a61109a,a61110a,a61113a,a61116a,a61117a,a61118a,a61121a,a61124a,a61125a,a61128a,a61131a,a61132a,a61133a,a61136a,a61139a,a61140a,a61143a,a61146a,a61147a,a61148a,a61151a,a61154a,a61155a,a61158a,a61161a,a61162a,a61163a,a61166a,a61169a,a61170a,a61173a,a61176a,a61177a,a61178a,a61181a,a61184a,a61185a,a61188a,a61191a,a61192a,a61193a,a61196a,a61199a,a61200a,a61203a,a61206a,a61207a,a61208a,a61211a,a61214a,a61215a,a61218a,a61221a,a61222a,a61223a,a61226a,a61229a,a61230a,a61233a,a61236a,a61237a,a61238a,a61241a,a61244a,a61245a,a61248a,a61251a,a61252a,a61253a,a61256a,a61259a,a61260a,a61263a,a61266a,a61267a,a61268a,a61271a,a61274a,a61275a,a61278a,a61281a,a61282a,a61283a,a61286a,a61289a,a61290a,a61293a,a61296a,a61297a,a61298a,a61301a,a61304a,a61305a,a61308a,a61311a,a61312a,a61313a,a61316a,a61319a,a61320a,a61323a,a61326a,a61327a,a61328a,a61331a,a61334a,a61335a,a61338a,a61341a,a61342a,a61343a,a61346a,a61349a,a61350a,a61353a,a61356a,a61357a,a61358a,a61361a,a61364a,a61365a,a61368a,a61371a,a61372a,a61373a,a61376a,a61379a,a61380a,a61383a,a61386a,a61387a,a61388a,a61391a,a61394a,a61395a,a61398a,a61401a,a61402a,a61403a,a61406a,a61409a,a61410a,a61413a,a61416a,a61417a,a61418a,a61421a,a61424a,a61425a,a61428a,a61431a,a61432a,a61433a,a61436a,a61439a,a61440a,a61443a,a61446a,a61447a,a61448a,a61451a,a61454a,a61455a,a61458a,a61461a,a61462a,a61463a,a61466a,a61469a,a61470a,a61473a,a61476a,a61477a,a61478a,a61481a,a61484a,a61485a,a61488a,a61491a,a61492a,a61493a,a61496a,a61499a,a61500a,a61503a,a61506a,a61507a,a61508a,a61511a,a61514a,a61515a,a61518a,a61521a,a61522a,a61523a,a61526a,a61529a,a61530a,a61533a,a61536a,a61537a,a61538a,a61541a,a61544a,a61545a,a61548a,a61551a,a61552a,a61553a,a61556a,a61559a,a61560a,a61563a,a61566a,a61567a,a61568a,a61571a,a61574a,a61575a,a61578a,a61581a,a61582a,a61583a,a61586a,a61589a,a61590a,a61593a,a61596a,a61597a,a61598a,a61601a,a61604a,a61605a,a61608a,a61611a,a61612a,a61613a,a61616a,a61619a,a61620a,a61623a,a61626a,a61627a,a61628a,a61631a,a61634a,a61635a,a61638a,a61641a,a61642a,a61643a,a61646a,a61649a,a61650a,a61653a,a61656a,a61657a,a61658a,a61661a,a61664a,a61665a,a61668a,a61671a,a61672a,a61673a,a61676a,a61679a,a61680a,a61683a,a61686a,a61687a,a61688a,a61691a,a61694a,a61695a,a61698a,a61701a,a61702a,a61703a,a61706a,a61709a,a61710a,a61713a,a61716a,a61717a,a61718a,a61721a,a61724a,a61725a,a61728a,a61731a,a61732a,a61733a,a61736a,a61739a,a61740a,a61743a,a61746a,a61747a,a61748a,a61751a,a61754a,a61755a,a61758a,a61761a,a61762a,a61763a,a61766a,a61769a,a61770a,a61773a,a61776a,a61777a,a61778a,a61781a,a61784a,a61785a,a61788a,a61791a,a61792a,a61793a,a61796a,a61799a,a61800a,a61803a,a61806a,a61807a,a61808a,a61811a,a61814a,a61815a,a61818a,a61821a,a61822a,a61823a,a61826a,a61829a,a61830a,a61833a,a61836a,a61837a,a61838a,a61841a,a61844a,a61845a,a61848a,a61851a,a61852a,a61853a,a61856a,a61859a,a61860a,a61863a,a61866a,a61867a,a61868a,a61871a,a61874a,a61875a,a61878a,a61881a,a61882a,a61883a,a61886a,a61889a,a61890a,a61893a,a61896a,a61897a,a61898a,a61901a,a61904a,a61905a,a61908a,a61911a,a61912a,a61913a,a61916a,a61919a,a61920a,a61923a,a61926a,a61927a,a61928a,a61931a,a61934a,a61935a,a61938a,a61941a,a61942a,a61943a,a61946a,a61949a,a61950a,a61953a,a61956a,a61957a,a61958a,a61961a,a61964a,a61965a,a61968a,a61971a,a61972a,a61973a,a61976a,a61979a,a61980a,a61983a,a61986a,a61987a,a61988a,a61991a,a61994a,a61995a,a61998a,a62001a,a62002a,a62003a,a62006a,a62009a,a62010a,a62013a,a62016a,a62017a,a62018a,a62021a,a62024a,a62025a,a62028a,a62031a,a62032a,a62033a,a62036a,a62039a,a62040a,a62043a,a62046a,a62047a,a62048a,a62051a,a62054a,a62055a,a62058a,a62061a,a62062a,a62063a,a62066a,a62069a,a62070a,a62073a,a62076a,a62077a,a62078a,a62081a,a62084a,a62085a,a62088a,a62091a,a62092a,a62093a,a62096a,a62099a,a62100a,a62103a,a62106a,a62107a,a62108a,a62111a,a62114a,a62115a,a62118a,a62121a,a62122a,a62123a,a62126a,a62129a,a62130a,a62133a,a62136a,a62137a,a62138a,a62141a,a62144a,a62145a,a62148a,a62151a,a62152a,a62153a,a62156a,a62159a,a62160a,a62163a,a62166a,a62167a,a62168a,a62171a,a62174a,a62175a,a62178a,a62181a,a62182a,a62183a,a62186a,a62189a,a62190a,a62193a,a62196a,a62197a,a62198a,a62201a,a62204a,a62205a,a62208a,a62211a,a62212a,a62213a,a62216a,a62219a,a62220a,a62223a,a62226a,a62227a,a62228a,a62231a,a62234a,a62235a,a62238a,a62241a,a62242a,a62243a,a62246a,a62249a,a62250a,a62253a,a62256a,a62257a,a62258a,a62261a,a62264a,a62265a,a62268a,a62271a,a62272a,a62273a,a62276a,a62279a,a62280a,a62283a,a62286a,a62287a,a62288a,a62291a,a62294a,a62295a,a62298a,a62301a,a62302a,a62303a,a62306a,a62309a,a62310a,a62313a,a62316a,a62317a,a62318a,a62321a,a62324a,a62325a,a62328a,a62331a,a62332a,a62333a,a62336a,a62339a,a62340a,a62343a,a62346a,a62347a,a62348a,a62351a,a62354a,a62355a,a62358a,a62361a,a62362a,a62363a,a62366a,a62369a,a62370a,a62373a,a62376a,a62377a,a62378a,a62381a,a62384a,a62385a,a62388a,a62391a,a62392a,a62393a,a62396a,a62399a,a62400a,a62403a,a62406a,a62407a,a62408a,a62411a,a62414a,a62415a,a62418a,a62421a,a62422a,a62423a,a62426a,a62429a,a62430a,a62433a,a62436a,a62437a,a62438a,a62441a,a62444a,a62445a,a62448a,a62451a,a62452a,a62453a,a62456a,a62459a,a62460a,a62463a,a62466a,a62467a,a62468a,a62471a,a62474a,a62475a,a62478a,a62481a,a62482a,a62483a,a62486a,a62489a,a62490a,a62493a,a62496a,a62497a,a62498a,a62501a,a62504a,a62505a,a62508a,a62511a,a62512a,a62513a,a62516a,a62519a,a62520a,a62523a,a62526a,a62527a,a62528a,a62531a,a62534a,a62535a,a62538a,a62541a,a62542a,a62543a,a62546a,a62549a,a62550a,a62553a,a62556a,a62557a,a62558a,a62561a,a62564a,a62565a,a62568a,a62571a,a62572a,a62573a,a62576a,a62579a,a62580a,a62583a,a62586a,a62587a,a62588a,a62591a,a62594a,a62595a,a62598a,a62601a,a62602a,a62603a,a62606a,a62609a,a62610a,a62613a,a62616a,a62617a,a62618a,a62621a,a62624a,a62625a,a62628a,a62631a,a62632a,a62633a,a62636a,a62639a,a62640a,a62643a,a62646a,a62647a,a62648a,a62651a,a62654a,a62655a,a62658a,a62661a,a62662a,a62663a,a62666a,a62669a,a62670a,a62673a,a62676a,a62677a,a62678a,a62681a,a62684a,a62685a,a62688a,a62691a,a62692a,a62693a,a62696a,a62699a,a62700a,a62703a,a62706a,a62707a,a62708a,a62711a,a62714a,a62715a,a62718a,a62721a,a62722a,a62723a,a62726a,a62729a,a62730a,a62733a,a62736a,a62737a,a62738a,a62741a,a62744a,a62745a,a62748a,a62751a,a62752a,a62753a,a62756a,a62759a,a62760a,a62763a,a62766a,a62767a,a62768a,a62771a,a62774a,a62775a,a62778a,a62781a,a62782a,a62783a,a62786a,a62789a,a62790a,a62793a,a62796a,a62797a,a62798a,a62801a,a62804a,a62805a,a62808a,a62811a,a62812a,a62813a,a62816a,a62819a,a62820a,a62823a,a62826a,a62827a,a62828a,a62831a,a62834a,a62835a,a62838a,a62841a,a62842a,a62843a,a62846a,a62849a,a62850a,a62853a,a62856a,a62857a,a62858a,a62861a,a62864a,a62865a,a62868a,a62871a,a62872a,a62873a,a62876a,a62879a,a62880a,a62883a,a62886a,a62887a,a62888a,a62891a,a62894a,a62895a,a62898a,a62901a,a62902a,a62903a,a62906a,a62909a,a62910a,a62913a,a62916a,a62917a,a62918a,a62921a,a62924a,a62925a,a62928a,a62931a,a62932a,a62933a,a62936a,a62939a,a62940a,a62943a,a62946a,a62947a,a62948a,a62951a,a62954a,a62955a,a62958a,a62961a,a62962a,a62963a,a62966a,a62969a,a62970a,a62973a,a62976a,a62977a,a62978a,a62981a,a62984a,a62985a,a62988a,a62991a,a62992a,a62993a,a62996a,a62999a,a63000a,a63003a,a63006a,a63007a,a63008a,a63011a,a63014a,a63015a,a63018a,a63021a,a63022a,a63023a,a63026a,a63029a,a63030a,a63033a,a63036a,a63037a,a63038a,a63041a,a63044a,a63045a,a63048a,a63051a,a63052a,a63053a,a63056a,a63059a,a63060a,a63063a,a63066a,a63067a,a63068a,a63071a,a63074a,a63075a,a63078a,a63081a,a63082a,a63083a,a63086a,a63089a,a63090a,a63093a,a63096a,a63097a,a63098a,a63101a,a63104a,a63105a,a63108a,a63111a,a63112a,a63113a,a63116a,a63119a,a63120a,a63123a,a63126a,a63127a,a63128a,a63131a,a63134a,a63135a,a63138a,a63141a,a63142a,a63143a,a63146a,a63149a,a63150a,a63153a,a63156a,a63157a,a63158a,a63161a,a63164a,a63165a,a63168a,a63171a,a63172a,a63173a,a63176a,a63179a,a63180a,a63183a,a63186a,a63187a,a63188a,a63191a,a63194a,a63195a,a63198a,a63201a,a63202a,a63203a,a63206a,a63209a,a63210a,a63213a,a63216a,a63217a,a63218a,a63221a,a63224a,a63225a,a63228a,a63231a,a63232a,a63233a,a63236a,a63239a,a63240a,a63243a,a63246a,a63247a,a63248a,a63251a,a63254a,a63255a,a63258a,a63261a,a63262a,a63263a,a63266a,a63269a,a63270a,a63273a,a63276a,a63277a,a63278a,a63281a,a63284a,a63285a,a63288a,a63291a,a63292a,a63293a,a63296a,a63299a,a63300a,a63303a,a63306a,a63307a,a63308a,a63311a,a63314a,a63315a,a63318a,a63321a,a63322a,a63323a,a63326a,a63329a,a63330a,a63333a,a63336a,a63337a,a63338a,a63341a,a63344a,a63345a,a63348a,a63351a,a63352a,a63353a,a63356a,a63359a,a63360a,a63363a,a63366a,a63367a,a63368a,a63371a,a63374a,a63375a,a63378a,a63381a,a63382a,a63383a,a63386a,a63389a,a63390a,a63393a,a63396a,a63397a,a63398a,a63401a,a63404a,a63405a,a63408a,a63411a,a63412a,a63413a,a63416a,a63419a,a63420a,a63423a,a63426a,a63427a,a63428a,a63431a,a63434a,a63435a,a63438a,a63441a,a63442a,a63443a,a63446a,a63449a,a63450a,a63453a,a63456a,a63457a,a63458a,a63461a,a63464a,a63465a,a63468a,a63471a,a63472a,a63473a,a63476a,a63479a,a63480a,a63483a,a63486a,a63487a,a63488a,a63491a,a63494a,a63495a,a63498a,a63501a,a63502a,a63503a,a63506a,a63509a,a63510a,a63513a,a63516a,a63517a,a63518a,a63521a,a63524a,a63525a,a63528a,a63531a,a63532a,a63533a,a63536a,a63539a,a63540a,a63543a,a63546a,a63547a,a63548a,a63551a,a63554a,a63555a,a63558a,a63561a,a63562a,a63563a,a63566a,a63569a,a63570a,a63573a,a63576a,a63577a,a63578a,a63581a,a63584a,a63585a,a63588a,a63591a,a63592a,a63593a,a63596a,a63599a,a63600a,a63603a,a63606a,a63607a,a63608a,a63611a,a63614a,a63615a,a63618a,a63621a,a63622a,a63623a,a63626a,a63629a,a63630a,a63633a,a63636a,a63637a,a63638a,a63641a,a63644a,a63645a,a63648a,a63651a,a63652a,a63653a,a63656a,a63659a,a63660a,a63663a,a63666a,a63667a,a63668a,a63671a,a63674a,a63675a,a63678a,a63681a,a63682a,a63683a,a63686a,a63689a,a63690a,a63693a,a63696a,a63697a,a63698a,a63701a,a63704a,a63705a,a63708a,a63711a,a63712a,a63713a,a63716a,a63719a,a63720a,a63723a,a63726a,a63727a,a63728a,a63731a,a63734a,a63735a,a63738a,a63741a,a63742a,a63743a,a63746a,a63749a,a63750a,a63753a,a63756a,a63757a,a63758a,a63761a,a63764a,a63765a,a63768a,a63771a,a63772a,a63773a,a63776a,a63779a,a63780a,a63783a,a63786a,a63787a,a63788a,a63791a,a63794a,a63795a,a63798a,a63801a,a63802a,a63803a,a63806a,a63809a,a63810a,a63813a,a63816a,a63817a,a63818a,a63821a,a63824a,a63825a,a63828a,a63831a,a63832a,a63833a,a63836a,a63839a,a63840a,a63843a,a63846a,a63847a,a63848a,a63851a,a63854a,a63855a,a63858a,a63861a,a63862a,a63863a,a63866a,a63869a,a63870a,a63873a,a63876a,a63877a,a63878a,a63881a,a63884a,a63885a,a63888a,a63891a,a63892a,a63893a,a63896a,a63899a,a63900a,a63903a,a63906a,a63907a,a63908a,a63911a,a63914a,a63915a,a63918a,a63921a,a63922a,a63923a,a63926a,a63929a,a63930a,a63933a,a63936a,a63937a,a63938a,a63941a,a63944a,a63945a,a63948a,a63951a,a63952a,a63953a,a63956a,a63959a,a63960a,a63963a,a63966a,a63967a,a63968a,a63971a,a63974a,a63975a,a63978a,a63981a,a63982a,a63983a,a63986a,a63989a,a63990a,a63993a,a63997a,a63998a,a63999a,a64000a,a64003a,a64006a,a64007a,a64010a,a64013a,a64014a,a64015a,a64018a,a64021a,a64022a,a64025a,a64029a,a64030a,a64031a,a64032a,a64035a,a64038a,a64039a,a64042a,a64045a,a64046a,a64047a,a64050a,a64053a,a64054a,a64057a,a64061a,a64062a,a64063a,a64064a,a64067a,a64070a,a64071a,a64074a,a64077a,a64078a,a64079a,a64082a,a64085a,a64086a,a64089a,a64093a,a64094a,a64095a,a64096a,a64099a,a64102a,a64103a,a64106a,a64109a,a64110a,a64111a,a64114a,a64117a,a64118a,a64121a,a64125a,a64126a,a64127a,a64128a,a64131a,a64134a,a64135a,a64138a,a64141a,a64142a,a64143a,a64146a,a64149a,a64150a,a64153a,a64157a,a64158a,a64159a,a64160a,a64163a,a64166a,a64167a,a64170a,a64173a,a64174a,a64175a,a64178a,a64181a,a64182a,a64185a,a64189a,a64190a,a64191a,a64192a,a64195a,a64198a,a64199a,a64202a,a64205a,a64206a,a64207a,a64210a,a64213a,a64214a,a64217a,a64221a,a64222a,a64223a,a64224a,a64227a,a64230a,a64231a,a64234a,a64237a,a64238a,a64239a,a64242a,a64245a,a64246a,a64249a,a64253a,a64254a,a64255a,a64256a,a64259a,a64262a,a64263a,a64266a,a64269a,a64270a,a64271a,a64274a,a64277a,a64278a,a64281a,a64285a,a64286a,a64287a,a64288a,a64291a,a64294a,a64295a,a64298a,a64301a,a64302a,a64303a,a64306a,a64309a,a64310a,a64313a,a64317a,a64318a,a64319a,a64320a,a64323a,a64326a,a64327a,a64330a,a64333a,a64334a,a64335a,a64338a,a64341a,a64342a,a64345a,a64349a,a64350a,a64351a,a64352a,a64355a,a64358a,a64359a,a64362a,a64365a,a64366a,a64367a,a64370a,a64373a,a64374a,a64377a,a64381a,a64382a,a64383a,a64384a,a64387a,a64390a,a64391a,a64394a,a64397a,a64398a,a64399a,a64402a,a64405a,a64406a,a64409a,a64413a,a64414a,a64415a,a64416a,a64419a,a64422a,a64423a,a64426a,a64429a,a64430a,a64431a,a64434a,a64437a,a64438a,a64441a,a64445a,a64446a,a64447a,a64448a,a64451a,a64454a,a64455a,a64458a,a64461a,a64462a,a64463a,a64466a,a64469a,a64470a,a64473a,a64477a,a64478a,a64479a,a64480a,a64483a,a64486a,a64487a,a64490a,a64493a,a64494a,a64495a,a64498a,a64501a,a64502a,a64505a,a64509a,a64510a,a64511a,a64512a,a64515a,a64518a,a64519a,a64522a,a64525a,a64526a,a64527a,a64530a,a64533a,a64534a,a64537a,a64541a,a64542a,a64543a,a64544a,a64547a,a64550a,a64551a,a64554a,a64557a,a64558a,a64559a,a64562a,a64565a,a64566a,a64569a,a64573a,a64574a,a64575a,a64576a,a64579a,a64582a,a64583a,a64586a,a64589a,a64590a,a64591a,a64594a,a64597a,a64598a,a64601a,a64605a,a64606a,a64607a,a64608a,a64611a,a64614a,a64615a,a64618a,a64621a,a64622a,a64623a,a64626a,a64629a,a64630a,a64633a,a64637a,a64638a,a64639a,a64640a,a64643a,a64646a,a64647a,a64650a,a64653a,a64654a,a64655a,a64658a,a64661a,a64662a,a64665a,a64669a,a64670a,a64671a,a64672a,a64675a,a64678a,a64679a,a64682a,a64685a,a64686a,a64687a,a64690a,a64693a,a64694a,a64697a,a64701a,a64702a,a64703a,a64704a,a64707a,a64710a,a64711a,a64714a,a64717a,a64718a,a64719a,a64722a,a64725a,a64726a,a64729a,a64733a,a64734a,a64735a,a64736a,a64739a,a64742a,a64743a,a64746a,a64749a,a64750a,a64751a,a64754a,a64757a,a64758a,a64761a,a64765a,a64766a,a64767a,a64768a,a64771a,a64774a,a64775a,a64778a,a64781a,a64782a,a64783a,a64786a,a64789a,a64790a,a64793a,a64797a,a64798a,a64799a,a64800a,a64803a,a64806a,a64807a,a64810a,a64813a,a64814a,a64815a,a64818a,a64821a,a64822a,a64825a,a64829a,a64830a,a64831a,a64832a,a64835a,a64838a,a64839a,a64842a,a64845a,a64846a,a64847a,a64850a,a64853a,a64854a,a64857a,a64861a,a64862a,a64863a,a64864a,a64867a,a64870a,a64871a,a64874a,a64877a,a64878a,a64879a,a64882a,a64885a,a64886a,a64889a,a64893a,a64894a,a64895a,a64896a,a64899a,a64902a,a64903a,a64906a,a64909a,a64910a,a64911a,a64914a,a64917a,a64918a,a64921a,a64925a,a64926a,a64927a,a64928a,a64931a,a64934a,a64935a,a64938a,a64941a,a64942a,a64943a,a64946a,a64949a,a64950a,a64953a,a64957a,a64958a,a64959a,a64960a,a64963a,a64966a,a64967a,a64970a,a64973a,a64974a,a64975a,a64978a,a64981a,a64982a,a64985a,a64989a,a64990a,a64991a,a64992a,a64995a,a64998a,a64999a,a65002a,a65005a,a65006a,a65007a,a65010a,a65013a,a65014a,a65017a,a65021a,a65022a,a65023a,a65024a,a65027a,a65030a,a65031a,a65034a,a65037a,a65038a,a65039a,a65042a,a65045a,a65046a,a65049a,a65053a,a65054a,a65055a,a65056a,a65059a,a65062a,a65063a,a65066a,a65069a,a65070a,a65071a,a65074a,a65077a,a65078a,a65081a,a65085a,a65086a,a65087a,a65088a,a65091a,a65094a,a65095a,a65098a,a65101a,a65102a,a65103a,a65106a,a65109a,a65110a,a65113a,a65117a,a65118a,a65119a,a65120a,a65123a,a65126a,a65127a,a65130a,a65133a,a65134a,a65135a,a65138a,a65141a,a65142a,a65145a,a65149a,a65150a,a65151a,a65152a,a65155a,a65158a,a65159a,a65162a,a65165a,a65166a,a65167a,a65170a,a65173a,a65174a,a65177a,a65181a,a65182a,a65183a,a65184a,a65187a,a65190a,a65191a,a65194a,a65197a,a65198a,a65199a,a65202a,a65205a,a65206a,a65209a,a65213a,a65214a,a65215a,a65216a,a65219a,a65222a,a65223a,a65226a,a65229a,a65230a,a65231a,a65234a,a65237a,a65238a,a65241a,a65245a,a65246a,a65247a,a65248a,a65251a,a65254a,a65255a,a65258a,a65261a,a65262a,a65263a,a65266a,a65269a,a65270a,a65273a,a65277a,a65278a,a65279a,a65280a,a65283a,a65286a,a65287a,a65290a,a65293a,a65294a,a65295a,a65298a,a65301a,a65302a,a65305a,a65309a,a65310a,a65311a,a65312a,a65315a,a65318a,a65319a,a65322a,a65325a,a65326a,a65327a,a65330a,a65333a,a65334a,a65337a,a65341a,a65342a,a65343a,a65344a,a65347a,a65350a,a65351a,a65354a,a65357a,a65358a,a65359a,a65362a,a65365a,a65366a,a65369a,a65373a,a65374a,a65375a,a65376a,a65379a,a65382a,a65383a,a65386a,a65389a,a65390a,a65391a,a65394a,a65397a,a65398a,a65401a,a65405a,a65406a,a65407a,a65408a,a65411a,a65414a,a65415a,a65418a,a65421a,a65422a,a65423a,a65426a,a65429a,a65430a,a65433a,a65437a,a65438a,a65439a,a65440a,a65443a,a65446a,a65447a,a65450a,a65453a,a65454a,a65455a,a65458a,a65461a,a65462a,a65465a,a65469a,a65470a,a65471a,a65472a,a65475a,a65478a,a65479a,a65482a,a65485a,a65486a,a65487a,a65490a,a65493a,a65494a,a65497a,a65501a,a65502a,a65503a,a65504a,a65507a,a65510a,a65511a,a65514a,a65517a,a65518a,a65519a,a65522a,a65525a,a65526a,a65529a,a65533a,a65534a,a65535a,a65536a,a65539a,a65542a,a65543a,a65546a,a65549a,a65550a,a65551a,a65554a,a65557a,a65558a,a65561a,a65565a,a65566a,a65567a,a65568a,a65571a,a65574a,a65575a,a65578a,a65581a,a65582a,a65583a,a65586a,a65589a,a65590a,a65593a,a65597a,a65598a,a65599a,a65600a,a65603a,a65606a,a65607a,a65610a,a65613a,a65614a,a65615a,a65618a,a65621a,a65622a,a65625a,a65629a,a65630a,a65631a,a65632a,a65635a,a65638a,a65639a,a65642a,a65645a,a65646a,a65647a,a65650a,a65653a,a65654a,a65657a,a65661a,a65662a,a65663a,a65664a,a65667a,a65670a,a65671a,a65674a,a65677a,a65678a,a65679a,a65682a,a65685a,a65686a,a65689a,a65693a,a65694a,a65695a,a65696a,a65699a,a65702a,a65703a,a65706a,a65709a,a65710a,a65711a,a65714a,a65717a,a65718a,a65721a,a65725a,a65726a,a65727a,a65728a,a65731a,a65734a,a65735a,a65738a,a65741a,a65742a,a65743a,a65746a,a65749a,a65750a,a65753a,a65757a,a65758a,a65759a,a65760a,a65763a,a65766a,a65767a,a65770a,a65773a,a65774a,a65775a,a65778a,a65781a,a65782a,a65785a,a65789a,a65790a,a65791a,a65792a,a65795a,a65798a,a65799a,a65802a,a65805a,a65806a,a65807a,a65810a,a65813a,a65814a,a65817a,a65821a,a65822a,a65823a,a65824a,a65827a,a65830a,a65831a,a65834a,a65837a,a65838a,a65839a,a65842a,a65845a,a65846a,a65849a,a65853a,a65854a,a65855a,a65856a,a65859a,a65862a,a65863a,a65866a,a65869a,a65870a,a65871a,a65874a,a65877a,a65878a,a65881a,a65885a,a65886a,a65887a,a65888a,a65891a,a65894a,a65895a,a65898a,a65901a,a65902a,a65903a,a65906a,a65909a,a65910a,a65913a,a65917a,a65918a,a65919a,a65920a,a65923a,a65926a,a65927a,a65930a,a65933a,a65934a,a65935a,a65938a,a65941a,a65942a,a65945a,a65949a,a65950a,a65951a,a65952a,a65955a,a65958a,a65959a,a65962a,a65965a,a65966a,a65967a,a65970a,a65973a,a65974a,a65977a,a65981a,a65982a,a65983a,a65984a,a65987a,a65990a,a65991a,a65994a,a65997a,a65998a,a65999a,a66002a,a66005a,a66006a,a66009a,a66013a,a66014a,a66015a,a66016a,a66019a,a66022a,a66023a,a66026a,a66030a,a66031a,a66032a,a66033a,a66036a,a66039a,a66040a,a66043a,a66047a,a66048a,a66049a,a66050a,a66053a,a66056a,a66057a,a66060a,a66064a,a66065a,a66066a,a66067a,a66070a,a66073a,a66074a,a66077a,a66081a,a66082a,a66083a,a66084a,a66087a,a66090a,a66091a,a66094a,a66098a,a66099a,a66100a,a66101a,a66104a,a66107a,a66108a,a66111a,a66115a,a66116a,a66117a,a66118a,a66121a,a66124a,a66125a,a66128a,a66132a,a66133a,a66134a,a66135a,a66138a,a66141a,a66142a,a66145a,a66149a,a66150a,a66151a,a66152a,a66155a,a66158a,a66159a,a66162a,a66166a,a66167a,a66168a,a66169a,a66172a,a66175a,a66176a,a66179a,a66183a,a66184a,a66185a,a66186a,a66189a,a66192a,a66193a,a66196a,a66200a,a66201a,a66202a,a66203a,a66206a,a66209a,a66210a,a66213a,a66217a,a66218a,a66219a,a66220a,a66223a,a66226a,a66227a,a66230a,a66234a,a66235a,a66236a,a66237a,a66240a,a66243a,a66244a,a66247a,a66251a,a66252a,a66253a,a66254a,a66257a,a66260a,a66261a,a66264a,a66268a,a66269a,a66270a,a66271a,a66274a,a66277a,a66278a,a66281a,a66285a,a66286a,a66287a,a66288a: std_logic;
begin

A72 <=( a7648a ) or ( a5099a );
 a1a <=( a66288a  and  a66271a );
 a2a <=( a66254a  and  a66237a );
 a3a <=( a66220a  and  a66203a );
 a4a <=( a66186a  and  a66169a );
 a5a <=( a66152a  and  a66135a );
 a6a <=( a66118a  and  a66101a );
 a7a <=( a66084a  and  a66067a );
 a8a <=( a66050a  and  a66033a );
 a9a <=( a66016a  and  a65999a );
 a10a <=( a65984a  and  a65967a );
 a11a <=( a65952a  and  a65935a );
 a12a <=( a65920a  and  a65903a );
 a13a <=( a65888a  and  a65871a );
 a14a <=( a65856a  and  a65839a );
 a15a <=( a65824a  and  a65807a );
 a16a <=( a65792a  and  a65775a );
 a17a <=( a65760a  and  a65743a );
 a18a <=( a65728a  and  a65711a );
 a19a <=( a65696a  and  a65679a );
 a20a <=( a65664a  and  a65647a );
 a21a <=( a65632a  and  a65615a );
 a22a <=( a65600a  and  a65583a );
 a23a <=( a65568a  and  a65551a );
 a24a <=( a65536a  and  a65519a );
 a25a <=( a65504a  and  a65487a );
 a26a <=( a65472a  and  a65455a );
 a27a <=( a65440a  and  a65423a );
 a28a <=( a65408a  and  a65391a );
 a29a <=( a65376a  and  a65359a );
 a30a <=( a65344a  and  a65327a );
 a31a <=( a65312a  and  a65295a );
 a32a <=( a65280a  and  a65263a );
 a33a <=( a65248a  and  a65231a );
 a34a <=( a65216a  and  a65199a );
 a35a <=( a65184a  and  a65167a );
 a36a <=( a65152a  and  a65135a );
 a37a <=( a65120a  and  a65103a );
 a38a <=( a65088a  and  a65071a );
 a39a <=( a65056a  and  a65039a );
 a40a <=( a65024a  and  a65007a );
 a41a <=( a64992a  and  a64975a );
 a42a <=( a64960a  and  a64943a );
 a43a <=( a64928a  and  a64911a );
 a44a <=( a64896a  and  a64879a );
 a45a <=( a64864a  and  a64847a );
 a46a <=( a64832a  and  a64815a );
 a47a <=( a64800a  and  a64783a );
 a48a <=( a64768a  and  a64751a );
 a49a <=( a64736a  and  a64719a );
 a50a <=( a64704a  and  a64687a );
 a51a <=( a64672a  and  a64655a );
 a52a <=( a64640a  and  a64623a );
 a53a <=( a64608a  and  a64591a );
 a54a <=( a64576a  and  a64559a );
 a55a <=( a64544a  and  a64527a );
 a56a <=( a64512a  and  a64495a );
 a57a <=( a64480a  and  a64463a );
 a58a <=( a64448a  and  a64431a );
 a59a <=( a64416a  and  a64399a );
 a60a <=( a64384a  and  a64367a );
 a61a <=( a64352a  and  a64335a );
 a62a <=( a64320a  and  a64303a );
 a63a <=( a64288a  and  a64271a );
 a64a <=( a64256a  and  a64239a );
 a65a <=( a64224a  and  a64207a );
 a66a <=( a64192a  and  a64175a );
 a67a <=( a64160a  and  a64143a );
 a68a <=( a64128a  and  a64111a );
 a69a <=( a64096a  and  a64079a );
 a70a <=( a64064a  and  a64047a );
 a71a <=( a64032a  and  a64015a );
 a72a <=( a64000a  and  a63983a );
 a73a <=( a63968a  and  a63953a );
 a74a <=( a63938a  and  a63923a );
 a75a <=( a63908a  and  a63893a );
 a76a <=( a63878a  and  a63863a );
 a77a <=( a63848a  and  a63833a );
 a78a <=( a63818a  and  a63803a );
 a79a <=( a63788a  and  a63773a );
 a80a <=( a63758a  and  a63743a );
 a81a <=( a63728a  and  a63713a );
 a82a <=( a63698a  and  a63683a );
 a83a <=( a63668a  and  a63653a );
 a84a <=( a63638a  and  a63623a );
 a85a <=( a63608a  and  a63593a );
 a86a <=( a63578a  and  a63563a );
 a87a <=( a63548a  and  a63533a );
 a88a <=( a63518a  and  a63503a );
 a89a <=( a63488a  and  a63473a );
 a90a <=( a63458a  and  a63443a );
 a91a <=( a63428a  and  a63413a );
 a92a <=( a63398a  and  a63383a );
 a93a <=( a63368a  and  a63353a );
 a94a <=( a63338a  and  a63323a );
 a95a <=( a63308a  and  a63293a );
 a96a <=( a63278a  and  a63263a );
 a97a <=( a63248a  and  a63233a );
 a98a <=( a63218a  and  a63203a );
 a99a <=( a63188a  and  a63173a );
 a100a <=( a63158a  and  a63143a );
 a101a <=( a63128a  and  a63113a );
 a102a <=( a63098a  and  a63083a );
 a103a <=( a63068a  and  a63053a );
 a104a <=( a63038a  and  a63023a );
 a105a <=( a63008a  and  a62993a );
 a106a <=( a62978a  and  a62963a );
 a107a <=( a62948a  and  a62933a );
 a108a <=( a62918a  and  a62903a );
 a109a <=( a62888a  and  a62873a );
 a110a <=( a62858a  and  a62843a );
 a111a <=( a62828a  and  a62813a );
 a112a <=( a62798a  and  a62783a );
 a113a <=( a62768a  and  a62753a );
 a114a <=( a62738a  and  a62723a );
 a115a <=( a62708a  and  a62693a );
 a116a <=( a62678a  and  a62663a );
 a117a <=( a62648a  and  a62633a );
 a118a <=( a62618a  and  a62603a );
 a119a <=( a62588a  and  a62573a );
 a120a <=( a62558a  and  a62543a );
 a121a <=( a62528a  and  a62513a );
 a122a <=( a62498a  and  a62483a );
 a123a <=( a62468a  and  a62453a );
 a124a <=( a62438a  and  a62423a );
 a125a <=( a62408a  and  a62393a );
 a126a <=( a62378a  and  a62363a );
 a127a <=( a62348a  and  a62333a );
 a128a <=( a62318a  and  a62303a );
 a129a <=( a62288a  and  a62273a );
 a130a <=( a62258a  and  a62243a );
 a131a <=( a62228a  and  a62213a );
 a132a <=( a62198a  and  a62183a );
 a133a <=( a62168a  and  a62153a );
 a134a <=( a62138a  and  a62123a );
 a135a <=( a62108a  and  a62093a );
 a136a <=( a62078a  and  a62063a );
 a137a <=( a62048a  and  a62033a );
 a138a <=( a62018a  and  a62003a );
 a139a <=( a61988a  and  a61973a );
 a140a <=( a61958a  and  a61943a );
 a141a <=( a61928a  and  a61913a );
 a142a <=( a61898a  and  a61883a );
 a143a <=( a61868a  and  a61853a );
 a144a <=( a61838a  and  a61823a );
 a145a <=( a61808a  and  a61793a );
 a146a <=( a61778a  and  a61763a );
 a147a <=( a61748a  and  a61733a );
 a148a <=( a61718a  and  a61703a );
 a149a <=( a61688a  and  a61673a );
 a150a <=( a61658a  and  a61643a );
 a151a <=( a61628a  and  a61613a );
 a152a <=( a61598a  and  a61583a );
 a153a <=( a61568a  and  a61553a );
 a154a <=( a61538a  and  a61523a );
 a155a <=( a61508a  and  a61493a );
 a156a <=( a61478a  and  a61463a );
 a157a <=( a61448a  and  a61433a );
 a158a <=( a61418a  and  a61403a );
 a159a <=( a61388a  and  a61373a );
 a160a <=( a61358a  and  a61343a );
 a161a <=( a61328a  and  a61313a );
 a162a <=( a61298a  and  a61283a );
 a163a <=( a61268a  and  a61253a );
 a164a <=( a61238a  and  a61223a );
 a165a <=( a61208a  and  a61193a );
 a166a <=( a61178a  and  a61163a );
 a167a <=( a61148a  and  a61133a );
 a168a <=( a61118a  and  a61103a );
 a169a <=( a61088a  and  a61073a );
 a170a <=( a61058a  and  a61043a );
 a171a <=( a61028a  and  a61013a );
 a172a <=( a60998a  and  a60983a );
 a173a <=( a60968a  and  a60953a );
 a174a <=( a60938a  and  a60923a );
 a175a <=( a60908a  and  a60893a );
 a176a <=( a60878a  and  a60863a );
 a177a <=( a60848a  and  a60833a );
 a178a <=( a60818a  and  a60803a );
 a179a <=( a60788a  and  a60773a );
 a180a <=( a60758a  and  a60743a );
 a181a <=( a60728a  and  a60713a );
 a182a <=( a60698a  and  a60683a );
 a183a <=( a60668a  and  a60653a );
 a184a <=( a60638a  and  a60623a );
 a185a <=( a60608a  and  a60593a );
 a186a <=( a60578a  and  a60563a );
 a187a <=( a60548a  and  a60533a );
 a188a <=( a60518a  and  a60503a );
 a189a <=( a60488a  and  a60473a );
 a190a <=( a60458a  and  a60443a );
 a191a <=( a60428a  and  a60413a );
 a192a <=( a60398a  and  a60383a );
 a193a <=( a60368a  and  a60353a );
 a194a <=( a60338a  and  a60323a );
 a195a <=( a60308a  and  a60293a );
 a196a <=( a60278a  and  a60263a );
 a197a <=( a60248a  and  a60233a );
 a198a <=( a60218a  and  a60203a );
 a199a <=( a60188a  and  a60173a );
 a200a <=( a60158a  and  a60143a );
 a201a <=( a60128a  and  a60113a );
 a202a <=( a60098a  and  a60083a );
 a203a <=( a60068a  and  a60053a );
 a204a <=( a60038a  and  a60023a );
 a205a <=( a60008a  and  a59993a );
 a206a <=( a59978a  and  a59963a );
 a207a <=( a59948a  and  a59933a );
 a208a <=( a59918a  and  a59903a );
 a209a <=( a59888a  and  a59873a );
 a210a <=( a59858a  and  a59843a );
 a211a <=( a59828a  and  a59813a );
 a212a <=( a59798a  and  a59783a );
 a213a <=( a59768a  and  a59753a );
 a214a <=( a59738a  and  a59723a );
 a215a <=( a59708a  and  a59693a );
 a216a <=( a59678a  and  a59663a );
 a217a <=( a59648a  and  a59633a );
 a218a <=( a59618a  and  a59603a );
 a219a <=( a59588a  and  a59573a );
 a220a <=( a59558a  and  a59543a );
 a221a <=( a59528a  and  a59513a );
 a222a <=( a59498a  and  a59483a );
 a223a <=( a59468a  and  a59453a );
 a224a <=( a59438a  and  a59423a );
 a225a <=( a59408a  and  a59393a );
 a226a <=( a59378a  and  a59363a );
 a227a <=( a59348a  and  a59333a );
 a228a <=( a59318a  and  a59303a );
 a229a <=( a59288a  and  a59273a );
 a230a <=( a59258a  and  a59243a );
 a231a <=( a59228a  and  a59213a );
 a232a <=( a59198a  and  a59183a );
 a233a <=( a59168a  and  a59153a );
 a234a <=( a59138a  and  a59123a );
 a235a <=( a59108a  and  a59093a );
 a236a <=( a59078a  and  a59063a );
 a237a <=( a59048a  and  a59033a );
 a238a <=( a59018a  and  a59003a );
 a239a <=( a58988a  and  a58973a );
 a240a <=( a58958a  and  a58943a );
 a241a <=( a58928a  and  a58913a );
 a242a <=( a58898a  and  a58883a );
 a243a <=( a58868a  and  a58853a );
 a244a <=( a58838a  and  a58823a );
 a245a <=( a58808a  and  a58793a );
 a246a <=( a58778a  and  a58763a );
 a247a <=( a58748a  and  a58733a );
 a248a <=( a58718a  and  a58703a );
 a249a <=( a58688a  and  a58673a );
 a250a <=( a58658a  and  a58643a );
 a251a <=( a58628a  and  a58613a );
 a252a <=( a58598a  and  a58583a );
 a253a <=( a58568a  and  a58553a );
 a254a <=( a58538a  and  a58523a );
 a255a <=( a58508a  and  a58493a );
 a256a <=( a58478a  and  a58463a );
 a257a <=( a58448a  and  a58433a );
 a258a <=( a58418a  and  a58403a );
 a259a <=( a58388a  and  a58373a );
 a260a <=( a58358a  and  a58343a );
 a261a <=( a58328a  and  a58313a );
 a262a <=( a58298a  and  a58283a );
 a263a <=( a58268a  and  a58253a );
 a264a <=( a58238a  and  a58223a );
 a265a <=( a58208a  and  a58193a );
 a266a <=( a58178a  and  a58163a );
 a267a <=( a58148a  and  a58133a );
 a268a <=( a58118a  and  a58103a );
 a269a <=( a58088a  and  a58073a );
 a270a <=( a58058a  and  a58043a );
 a271a <=( a58028a  and  a58013a );
 a272a <=( a57998a  and  a57983a );
 a273a <=( a57968a  and  a57953a );
 a274a <=( a57938a  and  a57923a );
 a275a <=( a57908a  and  a57893a );
 a276a <=( a57878a  and  a57863a );
 a277a <=( a57848a  and  a57833a );
 a278a <=( a57818a  and  a57803a );
 a279a <=( a57788a  and  a57773a );
 a280a <=( a57758a  and  a57743a );
 a281a <=( a57728a  and  a57713a );
 a282a <=( a57700a  and  a57685a );
 a283a <=( a57672a  and  a57657a );
 a284a <=( a57644a  and  a57629a );
 a285a <=( a57616a  and  a57601a );
 a286a <=( a57588a  and  a57573a );
 a287a <=( a57560a  and  a57545a );
 a288a <=( a57532a  and  a57517a );
 a289a <=( a57504a  and  a57489a );
 a290a <=( a57476a  and  a57461a );
 a291a <=( a57448a  and  a57433a );
 a292a <=( a57420a  and  a57405a );
 a293a <=( a57392a  and  a57377a );
 a294a <=( a57364a  and  a57349a );
 a295a <=( a57336a  and  a57321a );
 a296a <=( a57308a  and  a57293a );
 a297a <=( a57280a  and  a57265a );
 a298a <=( a57252a  and  a57237a );
 a299a <=( a57224a  and  a57209a );
 a300a <=( a57196a  and  a57181a );
 a301a <=( a57168a  and  a57153a );
 a302a <=( a57140a  and  a57125a );
 a303a <=( a57112a  and  a57097a );
 a304a <=( a57084a  and  a57069a );
 a305a <=( a57056a  and  a57041a );
 a306a <=( a57028a  and  a57013a );
 a307a <=( a57000a  and  a56985a );
 a308a <=( a56972a  and  a56957a );
 a309a <=( a56944a  and  a56929a );
 a310a <=( a56916a  and  a56901a );
 a311a <=( a56888a  and  a56873a );
 a312a <=( a56860a  and  a56845a );
 a313a <=( a56832a  and  a56817a );
 a314a <=( a56804a  and  a56789a );
 a315a <=( a56776a  and  a56761a );
 a316a <=( a56748a  and  a56733a );
 a317a <=( a56720a  and  a56705a );
 a318a <=( a56692a  and  a56677a );
 a319a <=( a56664a  and  a56649a );
 a320a <=( a56636a  and  a56621a );
 a321a <=( a56608a  and  a56593a );
 a322a <=( a56580a  and  a56565a );
 a323a <=( a56552a  and  a56537a );
 a324a <=( a56524a  and  a56509a );
 a325a <=( a56496a  and  a56481a );
 a326a <=( a56468a  and  a56453a );
 a327a <=( a56440a  and  a56425a );
 a328a <=( a56412a  and  a56397a );
 a329a <=( a56384a  and  a56369a );
 a330a <=( a56356a  and  a56341a );
 a331a <=( a56328a  and  a56313a );
 a332a <=( a56300a  and  a56285a );
 a333a <=( a56272a  and  a56257a );
 a334a <=( a56244a  and  a56229a );
 a335a <=( a56216a  and  a56201a );
 a336a <=( a56188a  and  a56173a );
 a337a <=( a56160a  and  a56145a );
 a338a <=( a56132a  and  a56117a );
 a339a <=( a56104a  and  a56089a );
 a340a <=( a56076a  and  a56061a );
 a341a <=( a56048a  and  a56033a );
 a342a <=( a56020a  and  a56005a );
 a343a <=( a55992a  and  a55977a );
 a344a <=( a55964a  and  a55949a );
 a345a <=( a55936a  and  a55921a );
 a346a <=( a55908a  and  a55893a );
 a347a <=( a55880a  and  a55865a );
 a348a <=( a55852a  and  a55837a );
 a349a <=( a55824a  and  a55809a );
 a350a <=( a55796a  and  a55781a );
 a351a <=( a55768a  and  a55753a );
 a352a <=( a55740a  and  a55725a );
 a353a <=( a55712a  and  a55697a );
 a354a <=( a55684a  and  a55669a );
 a355a <=( a55656a  and  a55641a );
 a356a <=( a55628a  and  a55613a );
 a357a <=( a55600a  and  a55585a );
 a358a <=( a55572a  and  a55557a );
 a359a <=( a55544a  and  a55529a );
 a360a <=( a55516a  and  a55501a );
 a361a <=( a55488a  and  a55473a );
 a362a <=( a55460a  and  a55445a );
 a363a <=( a55432a  and  a55417a );
 a364a <=( a55404a  and  a55389a );
 a365a <=( a55376a  and  a55361a );
 a366a <=( a55348a  and  a55333a );
 a367a <=( a55320a  and  a55305a );
 a368a <=( a55292a  and  a55277a );
 a369a <=( a55264a  and  a55249a );
 a370a <=( a55236a  and  a55221a );
 a371a <=( a55208a  and  a55193a );
 a372a <=( a55180a  and  a55165a );
 a373a <=( a55152a  and  a55137a );
 a374a <=( a55124a  and  a55109a );
 a375a <=( a55096a  and  a55081a );
 a376a <=( a55068a  and  a55053a );
 a377a <=( a55040a  and  a55025a );
 a378a <=( a55012a  and  a54997a );
 a379a <=( a54984a  and  a54969a );
 a380a <=( a54956a  and  a54941a );
 a381a <=( a54928a  and  a54913a );
 a382a <=( a54900a  and  a54885a );
 a383a <=( a54872a  and  a54857a );
 a384a <=( a54844a  and  a54829a );
 a385a <=( a54816a  and  a54801a );
 a386a <=( a54788a  and  a54773a );
 a387a <=( a54760a  and  a54745a );
 a388a <=( a54732a  and  a54717a );
 a389a <=( a54704a  and  a54689a );
 a390a <=( a54676a  and  a54661a );
 a391a <=( a54648a  and  a54633a );
 a392a <=( a54620a  and  a54605a );
 a393a <=( a54592a  and  a54577a );
 a394a <=( a54564a  and  a54549a );
 a395a <=( a54536a  and  a54521a );
 a396a <=( a54508a  and  a54493a );
 a397a <=( a54480a  and  a54465a );
 a398a <=( a54452a  and  a54437a );
 a399a <=( a54424a  and  a54409a );
 a400a <=( a54396a  and  a54381a );
 a401a <=( a54368a  and  a54353a );
 a402a <=( a54340a  and  a54325a );
 a403a <=( a54312a  and  a54297a );
 a404a <=( a54284a  and  a54269a );
 a405a <=( a54256a  and  a54241a );
 a406a <=( a54228a  and  a54213a );
 a407a <=( a54200a  and  a54185a );
 a408a <=( a54172a  and  a54157a );
 a409a <=( a54144a  and  a54129a );
 a410a <=( a54116a  and  a54101a );
 a411a <=( a54088a  and  a54073a );
 a412a <=( a54060a  and  a54045a );
 a413a <=( a54032a  and  a54017a );
 a414a <=( a54004a  and  a53989a );
 a415a <=( a53976a  and  a53961a );
 a416a <=( a53948a  and  a53933a );
 a417a <=( a53920a  and  a53905a );
 a418a <=( a53892a  and  a53877a );
 a419a <=( a53864a  and  a53849a );
 a420a <=( a53836a  and  a53821a );
 a421a <=( a53808a  and  a53793a );
 a422a <=( a53780a  and  a53765a );
 a423a <=( a53752a  and  a53737a );
 a424a <=( a53724a  and  a53709a );
 a425a <=( a53696a  and  a53681a );
 a426a <=( a53668a  and  a53653a );
 a427a <=( a53640a  and  a53625a );
 a428a <=( a53612a  and  a53597a );
 a429a <=( a53584a  and  a53569a );
 a430a <=( a53556a  and  a53541a );
 a431a <=( a53528a  and  a53513a );
 a432a <=( a53500a  and  a53485a );
 a433a <=( a53472a  and  a53457a );
 a434a <=( a53444a  and  a53429a );
 a435a <=( a53416a  and  a53401a );
 a436a <=( a53388a  and  a53373a );
 a437a <=( a53360a  and  a53345a );
 a438a <=( a53332a  and  a53317a );
 a439a <=( a53304a  and  a53289a );
 a440a <=( a53276a  and  a53261a );
 a441a <=( a53248a  and  a53233a );
 a442a <=( a53220a  and  a53205a );
 a443a <=( a53192a  and  a53177a );
 a444a <=( a53164a  and  a53149a );
 a445a <=( a53136a  and  a53121a );
 a446a <=( a53108a  and  a53093a );
 a447a <=( a53080a  and  a53065a );
 a448a <=( a53052a  and  a53037a );
 a449a <=( a53024a  and  a53009a );
 a450a <=( a52996a  and  a52981a );
 a451a <=( a52968a  and  a52953a );
 a452a <=( a52940a  and  a52925a );
 a453a <=( a52912a  and  a52897a );
 a454a <=( a52884a  and  a52869a );
 a455a <=( a52856a  and  a52841a );
 a456a <=( a52828a  and  a52813a );
 a457a <=( a52800a  and  a52785a );
 a458a <=( a52772a  and  a52757a );
 a459a <=( a52744a  and  a52729a );
 a460a <=( a52716a  and  a52701a );
 a461a <=( a52688a  and  a52673a );
 a462a <=( a52660a  and  a52645a );
 a463a <=( a52632a  and  a52617a );
 a464a <=( a52604a  and  a52589a );
 a465a <=( a52576a  and  a52561a );
 a466a <=( a52548a  and  a52533a );
 a467a <=( a52520a  and  a52505a );
 a468a <=( a52492a  and  a52477a );
 a469a <=( a52464a  and  a52449a );
 a470a <=( a52436a  and  a52421a );
 a471a <=( a52408a  and  a52393a );
 a472a <=( a52380a  and  a52365a );
 a473a <=( a52352a  and  a52337a );
 a474a <=( a52324a  and  a52309a );
 a475a <=( a52296a  and  a52281a );
 a476a <=( a52268a  and  a52253a );
 a477a <=( a52240a  and  a52225a );
 a478a <=( a52212a  and  a52197a );
 a479a <=( a52184a  and  a52169a );
 a480a <=( a52156a  and  a52141a );
 a481a <=( a52128a  and  a52113a );
 a482a <=( a52100a  and  a52085a );
 a483a <=( a52072a  and  a52057a );
 a484a <=( a52044a  and  a52029a );
 a485a <=( a52016a  and  a52001a );
 a486a <=( a51988a  and  a51973a );
 a487a <=( a51960a  and  a51945a );
 a488a <=( a51932a  and  a51917a );
 a489a <=( a51904a  and  a51889a );
 a490a <=( a51876a  and  a51861a );
 a491a <=( a51848a  and  a51833a );
 a492a <=( a51820a  and  a51805a );
 a493a <=( a51792a  and  a51777a );
 a494a <=( a51764a  and  a51749a );
 a495a <=( a51736a  and  a51721a );
 a496a <=( a51708a  and  a51693a );
 a497a <=( a51680a  and  a51665a );
 a498a <=( a51652a  and  a51637a );
 a499a <=( a51624a  and  a51609a );
 a500a <=( a51596a  and  a51581a );
 a501a <=( a51568a  and  a51553a );
 a502a <=( a51540a  and  a51525a );
 a503a <=( a51512a  and  a51497a );
 a504a <=( a51484a  and  a51469a );
 a505a <=( a51456a  and  a51441a );
 a506a <=( a51428a  and  a51413a );
 a507a <=( a51400a  and  a51385a );
 a508a <=( a51372a  and  a51357a );
 a509a <=( a51344a  and  a51329a );
 a510a <=( a51316a  and  a51301a );
 a511a <=( a51288a  and  a51273a );
 a512a <=( a51260a  and  a51245a );
 a513a <=( a51232a  and  a51217a );
 a514a <=( a51204a  and  a51189a );
 a515a <=( a51176a  and  a51161a );
 a516a <=( a51148a  and  a51133a );
 a517a <=( a51120a  and  a51105a );
 a518a <=( a51092a  and  a51077a );
 a519a <=( a51064a  and  a51049a );
 a520a <=( a51036a  and  a51021a );
 a521a <=( a51008a  and  a50993a );
 a522a <=( a50980a  and  a50965a );
 a523a <=( a50952a  and  a50937a );
 a524a <=( a50924a  and  a50909a );
 a525a <=( a50896a  and  a50881a );
 a526a <=( a50868a  and  a50853a );
 a527a <=( a50840a  and  a50825a );
 a528a <=( a50812a  and  a50797a );
 a529a <=( a50784a  and  a50769a );
 a530a <=( a50756a  and  a50741a );
 a531a <=( a50728a  and  a50713a );
 a532a <=( a50700a  and  a50685a );
 a533a <=( a50672a  and  a50657a );
 a534a <=( a50644a  and  a50629a );
 a535a <=( a50616a  and  a50601a );
 a536a <=( a50588a  and  a50573a );
 a537a <=( a50560a  and  a50545a );
 a538a <=( a50532a  and  a50517a );
 a539a <=( a50504a  and  a50489a );
 a540a <=( a50476a  and  a50461a );
 a541a <=( a50448a  and  a50433a );
 a542a <=( a50420a  and  a50405a );
 a543a <=( a50392a  and  a50377a );
 a544a <=( a50364a  and  a50349a );
 a545a <=( a50336a  and  a50321a );
 a546a <=( a50308a  and  a50293a );
 a547a <=( a50280a  and  a50265a );
 a548a <=( a50252a  and  a50237a );
 a549a <=( a50224a  and  a50209a );
 a550a <=( a50196a  and  a50181a );
 a551a <=( a50168a  and  a50153a );
 a552a <=( a50140a  and  a50125a );
 a553a <=( a50112a  and  a50097a );
 a554a <=( a50084a  and  a50069a );
 a555a <=( a50056a  and  a50041a );
 a556a <=( a50028a  and  a50013a );
 a557a <=( a50000a  and  a49985a );
 a558a <=( a49972a  and  a49957a );
 a559a <=( a49944a  and  a49929a );
 a560a <=( a49916a  and  a49901a );
 a561a <=( a49888a  and  a49873a );
 a562a <=( a49860a  and  a49845a );
 a563a <=( a49832a  and  a49817a );
 a564a <=( a49804a  and  a49789a );
 a565a <=( a49776a  and  a49761a );
 a566a <=( a49748a  and  a49733a );
 a567a <=( a49720a  and  a49705a );
 a568a <=( a49692a  and  a49677a );
 a569a <=( a49664a  and  a49649a );
 a570a <=( a49636a  and  a49621a );
 a571a <=( a49608a  and  a49593a );
 a572a <=( a49580a  and  a49565a );
 a573a <=( a49552a  and  a49537a );
 a574a <=( a49524a  and  a49509a );
 a575a <=( a49496a  and  a49481a );
 a576a <=( a49468a  and  a49453a );
 a577a <=( a49440a  and  a49425a );
 a578a <=( a49412a  and  a49397a );
 a579a <=( a49384a  and  a49369a );
 a580a <=( a49356a  and  a49341a );
 a581a <=( a49328a  and  a49313a );
 a582a <=( a49300a  and  a49285a );
 a583a <=( a49272a  and  a49257a );
 a584a <=( a49244a  and  a49229a );
 a585a <=( a49216a  and  a49201a );
 a586a <=( a49188a  and  a49173a );
 a587a <=( a49160a  and  a49145a );
 a588a <=( a49132a  and  a49117a );
 a589a <=( a49104a  and  a49089a );
 a590a <=( a49076a  and  a49061a );
 a591a <=( a49048a  and  a49033a );
 a592a <=( a49020a  and  a49005a );
 a593a <=( a48992a  and  a48977a );
 a594a <=( a48964a  and  a48949a );
 a595a <=( a48936a  and  a48921a );
 a596a <=( a48908a  and  a48893a );
 a597a <=( a48880a  and  a48865a );
 a598a <=( a48852a  and  a48837a );
 a599a <=( a48824a  and  a48809a );
 a600a <=( a48796a  and  a48781a );
 a601a <=( a48768a  and  a48753a );
 a602a <=( a48740a  and  a48725a );
 a603a <=( a48712a  and  a48697a );
 a604a <=( a48684a  and  a48669a );
 a605a <=( a48656a  and  a48641a );
 a606a <=( a48628a  and  a48613a );
 a607a <=( a48600a  and  a48585a );
 a608a <=( a48572a  and  a48557a );
 a609a <=( a48544a  and  a48529a );
 a610a <=( a48516a  and  a48501a );
 a611a <=( a48488a  and  a48473a );
 a612a <=( a48460a  and  a48445a );
 a613a <=( a48432a  and  a48417a );
 a614a <=( a48404a  and  a48389a );
 a615a <=( a48376a  and  a48361a );
 a616a <=( a48348a  and  a48333a );
 a617a <=( a48320a  and  a48305a );
 a618a <=( a48292a  and  a48277a );
 a619a <=( a48264a  and  a48249a );
 a620a <=( a48236a  and  a48221a );
 a621a <=( a48208a  and  a48193a );
 a622a <=( a48180a  and  a48165a );
 a623a <=( a48152a  and  a48137a );
 a624a <=( a48124a  and  a48109a );
 a625a <=( a48096a  and  a48081a );
 a626a <=( a48068a  and  a48053a );
 a627a <=( a48040a  and  a48025a );
 a628a <=( a48012a  and  a47997a );
 a629a <=( a47984a  and  a47969a );
 a630a <=( a47956a  and  a47941a );
 a631a <=( a47928a  and  a47913a );
 a632a <=( a47900a  and  a47885a );
 a633a <=( a47872a  and  a47857a );
 a634a <=( a47844a  and  a47829a );
 a635a <=( a47816a  and  a47801a );
 a636a <=( a47788a  and  a47773a );
 a637a <=( a47760a  and  a47745a );
 a638a <=( a47732a  and  a47717a );
 a639a <=( a47704a  and  a47689a );
 a640a <=( a47676a  and  a47661a );
 a641a <=( a47648a  and  a47635a );
 a642a <=( a47622a  and  a47609a );
 a643a <=( a47596a  and  a47583a );
 a644a <=( a47570a  and  a47557a );
 a645a <=( a47544a  and  a47531a );
 a646a <=( a47518a  and  a47505a );
 a647a <=( a47492a  and  a47479a );
 a648a <=( a47466a  and  a47453a );
 a649a <=( a47440a  and  a47427a );
 a650a <=( a47414a  and  a47401a );
 a651a <=( a47388a  and  a47375a );
 a652a <=( a47362a  and  a47349a );
 a653a <=( a47336a  and  a47323a );
 a654a <=( a47310a  and  a47297a );
 a655a <=( a47284a  and  a47271a );
 a656a <=( a47258a  and  a47245a );
 a657a <=( a47232a  and  a47219a );
 a658a <=( a47206a  and  a47193a );
 a659a <=( a47180a  and  a47167a );
 a660a <=( a47154a  and  a47141a );
 a661a <=( a47128a  and  a47115a );
 a662a <=( a47102a  and  a47089a );
 a663a <=( a47076a  and  a47063a );
 a664a <=( a47050a  and  a47037a );
 a665a <=( a47024a  and  a47011a );
 a666a <=( a46998a  and  a46985a );
 a667a <=( a46972a  and  a46959a );
 a668a <=( a46946a  and  a46933a );
 a669a <=( a46920a  and  a46907a );
 a670a <=( a46894a  and  a46881a );
 a671a <=( a46868a  and  a46855a );
 a672a <=( a46842a  and  a46829a );
 a673a <=( a46816a  and  a46803a );
 a674a <=( a46790a  and  a46777a );
 a675a <=( a46764a  and  a46751a );
 a676a <=( a46738a  and  a46725a );
 a677a <=( a46712a  and  a46699a );
 a678a <=( a46686a  and  a46673a );
 a679a <=( a46660a  and  a46647a );
 a680a <=( a46634a  and  a46621a );
 a681a <=( a46608a  and  a46595a );
 a682a <=( a46582a  and  a46569a );
 a683a <=( a46556a  and  a46543a );
 a684a <=( a46530a  and  a46517a );
 a685a <=( a46504a  and  a46491a );
 a686a <=( a46478a  and  a46465a );
 a687a <=( a46452a  and  a46439a );
 a688a <=( a46426a  and  a46413a );
 a689a <=( a46400a  and  a46387a );
 a690a <=( a46374a  and  a46361a );
 a691a <=( a46348a  and  a46335a );
 a692a <=( a46322a  and  a46309a );
 a693a <=( a46296a  and  a46283a );
 a694a <=( a46270a  and  a46257a );
 a695a <=( a46244a  and  a46231a );
 a696a <=( a46218a  and  a46205a );
 a697a <=( a46192a  and  a46179a );
 a698a <=( a46166a  and  a46153a );
 a699a <=( a46140a  and  a46127a );
 a700a <=( a46114a  and  a46101a );
 a701a <=( a46088a  and  a46075a );
 a702a <=( a46062a  and  a46049a );
 a703a <=( a46036a  and  a46023a );
 a704a <=( a46010a  and  a45997a );
 a705a <=( a45984a  and  a45971a );
 a706a <=( a45958a  and  a45945a );
 a707a <=( a45932a  and  a45919a );
 a708a <=( a45906a  and  a45893a );
 a709a <=( a45880a  and  a45867a );
 a710a <=( a45854a  and  a45841a );
 a711a <=( a45828a  and  a45815a );
 a712a <=( a45802a  and  a45789a );
 a713a <=( a45776a  and  a45763a );
 a714a <=( a45750a  and  a45737a );
 a715a <=( a45724a  and  a45711a );
 a716a <=( a45698a  and  a45685a );
 a717a <=( a45672a  and  a45659a );
 a718a <=( a45646a  and  a45633a );
 a719a <=( a45620a  and  a45607a );
 a720a <=( a45594a  and  a45581a );
 a721a <=( a45568a  and  a45555a );
 a722a <=( a45542a  and  a45529a );
 a723a <=( a45516a  and  a45503a );
 a724a <=( a45490a  and  a45477a );
 a725a <=( a45464a  and  a45451a );
 a726a <=( a45438a  and  a45425a );
 a727a <=( a45412a  and  a45399a );
 a728a <=( a45386a  and  a45373a );
 a729a <=( a45360a  and  a45347a );
 a730a <=( a45334a  and  a45321a );
 a731a <=( a45308a  and  a45295a );
 a732a <=( a45282a  and  a45269a );
 a733a <=( a45256a  and  a45243a );
 a734a <=( a45230a  and  a45217a );
 a735a <=( a45204a  and  a45191a );
 a736a <=( a45178a  and  a45165a );
 a737a <=( a45152a  and  a45139a );
 a738a <=( a45126a  and  a45113a );
 a739a <=( a45100a  and  a45087a );
 a740a <=( a45074a  and  a45061a );
 a741a <=( a45048a  and  a45035a );
 a742a <=( a45022a  and  a45009a );
 a743a <=( a44996a  and  a44983a );
 a744a <=( a44970a  and  a44957a );
 a745a <=( a44944a  and  a44931a );
 a746a <=( a44918a  and  a44905a );
 a747a <=( a44892a  and  a44879a );
 a748a <=( a44866a  and  a44853a );
 a749a <=( a44840a  and  a44827a );
 a750a <=( a44814a  and  a44801a );
 a751a <=( a44788a  and  a44775a );
 a752a <=( a44762a  and  a44749a );
 a753a <=( a44736a  and  a44723a );
 a754a <=( a44710a  and  a44697a );
 a755a <=( a44684a  and  a44671a );
 a756a <=( a44658a  and  a44645a );
 a757a <=( a44632a  and  a44619a );
 a758a <=( a44606a  and  a44593a );
 a759a <=( a44580a  and  a44567a );
 a760a <=( a44554a  and  a44541a );
 a761a <=( a44528a  and  a44515a );
 a762a <=( a44502a  and  a44489a );
 a763a <=( a44476a  and  a44463a );
 a764a <=( a44450a  and  a44437a );
 a765a <=( a44424a  and  a44411a );
 a766a <=( a44398a  and  a44385a );
 a767a <=( a44372a  and  a44359a );
 a768a <=( a44346a  and  a44333a );
 a769a <=( a44320a  and  a44307a );
 a770a <=( a44294a  and  a44281a );
 a771a <=( a44268a  and  a44255a );
 a772a <=( a44242a  and  a44229a );
 a773a <=( a44216a  and  a44203a );
 a774a <=( a44190a  and  a44177a );
 a775a <=( a44164a  and  a44151a );
 a776a <=( a44138a  and  a44125a );
 a777a <=( a44112a  and  a44099a );
 a778a <=( a44086a  and  a44073a );
 a779a <=( a44060a  and  a44047a );
 a780a <=( a44034a  and  a44021a );
 a781a <=( a44008a  and  a43995a );
 a782a <=( a43982a  and  a43969a );
 a783a <=( a43956a  and  a43943a );
 a784a <=( a43930a  and  a43917a );
 a785a <=( a43904a  and  a43891a );
 a786a <=( a43878a  and  a43865a );
 a787a <=( a43852a  and  a43839a );
 a788a <=( a43826a  and  a43813a );
 a789a <=( a43800a  and  a43787a );
 a790a <=( a43774a  and  a43761a );
 a791a <=( a43748a  and  a43735a );
 a792a <=( a43722a  and  a43709a );
 a793a <=( a43696a  and  a43683a );
 a794a <=( a43670a  and  a43657a );
 a795a <=( a43644a  and  a43631a );
 a796a <=( a43618a  and  a43605a );
 a797a <=( a43592a  and  a43579a );
 a798a <=( a43566a  and  a43553a );
 a799a <=( a43540a  and  a43527a );
 a800a <=( a43514a  and  a43501a );
 a801a <=( a43488a  and  a43475a );
 a802a <=( a43462a  and  a43449a );
 a803a <=( a43436a  and  a43423a );
 a804a <=( a43410a  and  a43397a );
 a805a <=( a43384a  and  a43371a );
 a806a <=( a43358a  and  a43345a );
 a807a <=( a43332a  and  a43319a );
 a808a <=( a43306a  and  a43293a );
 a809a <=( a43280a  and  a43267a );
 a810a <=( a43254a  and  a43241a );
 a811a <=( a43228a  and  a43215a );
 a812a <=( a43202a  and  a43189a );
 a813a <=( a43176a  and  a43163a );
 a814a <=( a43150a  and  a43137a );
 a815a <=( a43124a  and  a43111a );
 a816a <=( a43098a  and  a43085a );
 a817a <=( a43072a  and  a43059a );
 a818a <=( a43046a  and  a43033a );
 a819a <=( a43020a  and  a43007a );
 a820a <=( a42994a  and  a42981a );
 a821a <=( a42968a  and  a42955a );
 a822a <=( a42942a  and  a42929a );
 a823a <=( a42916a  and  a42903a );
 a824a <=( a42890a  and  a42877a );
 a825a <=( a42864a  and  a42851a );
 a826a <=( a42838a  and  a42825a );
 a827a <=( a42812a  and  a42799a );
 a828a <=( a42786a  and  a42773a );
 a829a <=( a42760a  and  a42747a );
 a830a <=( a42734a  and  a42721a );
 a831a <=( a42708a  and  a42695a );
 a832a <=( a42682a  and  a42669a );
 a833a <=( a42656a  and  a42643a );
 a834a <=( a42630a  and  a42617a );
 a835a <=( a42604a  and  a42591a );
 a836a <=( a42578a  and  a42565a );
 a837a <=( a42552a  and  a42539a );
 a838a <=( a42526a  and  a42513a );
 a839a <=( a42500a  and  a42487a );
 a840a <=( a42474a  and  a42461a );
 a841a <=( a42448a  and  a42435a );
 a842a <=( a42422a  and  a42409a );
 a843a <=( a42396a  and  a42383a );
 a844a <=( a42370a  and  a42357a );
 a845a <=( a42344a  and  a42331a );
 a846a <=( a42318a  and  a42305a );
 a847a <=( a42292a  and  a42279a );
 a848a <=( a42266a  and  a42253a );
 a849a <=( a42240a  and  a42227a );
 a850a <=( a42214a  and  a42201a );
 a851a <=( a42188a  and  a42175a );
 a852a <=( a42162a  and  a42149a );
 a853a <=( a42136a  and  a42123a );
 a854a <=( a42110a  and  a42097a );
 a855a <=( a42084a  and  a42071a );
 a856a <=( a42058a  and  a42045a );
 a857a <=( a42032a  and  a42019a );
 a858a <=( a42006a  and  a41993a );
 a859a <=( a41980a  and  a41967a );
 a860a <=( a41954a  and  a41941a );
 a861a <=( a41928a  and  a41915a );
 a862a <=( a41902a  and  a41889a );
 a863a <=( a41876a  and  a41863a );
 a864a <=( a41850a  and  a41837a );
 a865a <=( a41824a  and  a41811a );
 a866a <=( a41798a  and  a41785a );
 a867a <=( a41772a  and  a41759a );
 a868a <=( a41746a  and  a41733a );
 a869a <=( a41720a  and  a41707a );
 a870a <=( a41694a  and  a41681a );
 a871a <=( a41668a  and  a41655a );
 a872a <=( a41642a  and  a41629a );
 a873a <=( a41616a  and  a41603a );
 a874a <=( a41590a  and  a41577a );
 a875a <=( a41564a  and  a41551a );
 a876a <=( a41538a  and  a41525a );
 a877a <=( a41512a  and  a41499a );
 a878a <=( a41486a  and  a41473a );
 a879a <=( a41460a  and  a41447a );
 a880a <=( a41434a  and  a41421a );
 a881a <=( a41408a  and  a41395a );
 a882a <=( a41382a  and  a41369a );
 a883a <=( a41356a  and  a41343a );
 a884a <=( a41330a  and  a41317a );
 a885a <=( a41304a  and  a41291a );
 a886a <=( a41278a  and  a41265a );
 a887a <=( a41252a  and  a41239a );
 a888a <=( a41226a  and  a41213a );
 a889a <=( a41200a  and  a41187a );
 a890a <=( a41174a  and  a41161a );
 a891a <=( a41148a  and  a41135a );
 a892a <=( a41122a  and  a41109a );
 a893a <=( a41096a  and  a41083a );
 a894a <=( a41070a  and  a41057a );
 a895a <=( a41044a  and  a41031a );
 a896a <=( a41018a  and  a41005a );
 a897a <=( a40992a  and  a40979a );
 a898a <=( a40966a  and  a40953a );
 a899a <=( a40940a  and  a40927a );
 a900a <=( a40914a  and  a40901a );
 a901a <=( a40888a  and  a40875a );
 a902a <=( a40862a  and  a40849a );
 a903a <=( a40836a  and  a40823a );
 a904a <=( a40810a  and  a40797a );
 a905a <=( a40784a  and  a40771a );
 a906a <=( a40758a  and  a40745a );
 a907a <=( a40732a  and  a40719a );
 a908a <=( a40706a  and  a40693a );
 a909a <=( a40680a  and  a40667a );
 a910a <=( a40654a  and  a40641a );
 a911a <=( a40628a  and  a40615a );
 a912a <=( a40602a  and  a40589a );
 a913a <=( a40576a  and  a40563a );
 a914a <=( a40550a  and  a40537a );
 a915a <=( a40524a  and  a40511a );
 a916a <=( a40498a  and  a40485a );
 a917a <=( a40472a  and  a40459a );
 a918a <=( a40446a  and  a40433a );
 a919a <=( a40420a  and  a40407a );
 a920a <=( a40394a  and  a40381a );
 a921a <=( a40368a  and  a40355a );
 a922a <=( a40342a  and  a40329a );
 a923a <=( a40316a  and  a40303a );
 a924a <=( a40290a  and  a40277a );
 a925a <=( a40264a  and  a40251a );
 a926a <=( a40238a  and  a40225a );
 a927a <=( a40212a  and  a40199a );
 a928a <=( a40186a  and  a40173a );
 a929a <=( a40160a  and  a40147a );
 a930a <=( a40134a  and  a40121a );
 a931a <=( a40108a  and  a40095a );
 a932a <=( a40082a  and  a40069a );
 a933a <=( a40056a  and  a40043a );
 a934a <=( a40030a  and  a40017a );
 a935a <=( a40004a  and  a39991a );
 a936a <=( a39978a  and  a39965a );
 a937a <=( a39952a  and  a39939a );
 a938a <=( a39926a  and  a39913a );
 a939a <=( a39900a  and  a39887a );
 a940a <=( a39874a  and  a39861a );
 a941a <=( a39848a  and  a39835a );
 a942a <=( a39822a  and  a39809a );
 a943a <=( a39796a  and  a39783a );
 a944a <=( a39770a  and  a39757a );
 a945a <=( a39744a  and  a39731a );
 a946a <=( a39718a  and  a39705a );
 a947a <=( a39692a  and  a39679a );
 a948a <=( a39666a  and  a39653a );
 a949a <=( a39640a  and  a39627a );
 a950a <=( a39614a  and  a39601a );
 a951a <=( a39588a  and  a39575a );
 a952a <=( a39562a  and  a39549a );
 a953a <=( a39536a  and  a39523a );
 a954a <=( a39510a  and  a39497a );
 a955a <=( a39484a  and  a39471a );
 a956a <=( a39458a  and  a39445a );
 a957a <=( a39432a  and  a39419a );
 a958a <=( a39406a  and  a39393a );
 a959a <=( a39380a  and  a39367a );
 a960a <=( a39354a  and  a39341a );
 a961a <=( a39328a  and  a39315a );
 a962a <=( a39302a  and  a39289a );
 a963a <=( a39276a  and  a39263a );
 a964a <=( a39250a  and  a39237a );
 a965a <=( a39224a  and  a39211a );
 a966a <=( a39198a  and  a39185a );
 a967a <=( a39172a  and  a39159a );
 a968a <=( a39146a  and  a39133a );
 a969a <=( a39120a  and  a39107a );
 a970a <=( a39094a  and  a39081a );
 a971a <=( a39068a  and  a39055a );
 a972a <=( a39042a  and  a39029a );
 a973a <=( a39016a  and  a39003a );
 a974a <=( a38990a  and  a38977a );
 a975a <=( a38964a  and  a38951a );
 a976a <=( a38938a  and  a38925a );
 a977a <=( a38912a  and  a38899a );
 a978a <=( a38886a  and  a38873a );
 a979a <=( a38860a  and  a38847a );
 a980a <=( a38834a  and  a38821a );
 a981a <=( a38808a  and  a38795a );
 a982a <=( a38782a  and  a38769a );
 a983a <=( a38756a  and  a38743a );
 a984a <=( a38730a  and  a38717a );
 a985a <=( a38704a  and  a38691a );
 a986a <=( a38678a  and  a38665a );
 a987a <=( a38652a  and  a38639a );
 a988a <=( a38626a  and  a38613a );
 a989a <=( a38600a  and  a38587a );
 a990a <=( a38574a  and  a38561a );
 a991a <=( a38548a  and  a38535a );
 a992a <=( a38522a  and  a38509a );
 a993a <=( a38496a  and  a38483a );
 a994a <=( a38470a  and  a38457a );
 a995a <=( a38444a  and  a38431a );
 a996a <=( a38418a  and  a38405a );
 a997a <=( a38392a  and  a38379a );
 a998a <=( a38366a  and  a38353a );
 a999a <=( a38340a  and  a38327a );
 a1000a <=( a38314a  and  a38301a );
 a1001a <=( a38288a  and  a38275a );
 a1002a <=( a38262a  and  a38249a );
 a1003a <=( a38236a  and  a38223a );
 a1004a <=( a38210a  and  a38197a );
 a1005a <=( a38184a  and  a38171a );
 a1006a <=( a38158a  and  a38145a );
 a1007a <=( a38132a  and  a38119a );
 a1008a <=( a38106a  and  a38093a );
 a1009a <=( a38080a  and  a38067a );
 a1010a <=( a38054a  and  a38041a );
 a1011a <=( a38028a  and  a38015a );
 a1012a <=( a38002a  and  a37989a );
 a1013a <=( a37976a  and  a37963a );
 a1014a <=( a37950a  and  a37937a );
 a1015a <=( a37924a  and  a37911a );
 a1016a <=( a37898a  and  a37885a );
 a1017a <=( a37872a  and  a37859a );
 a1018a <=( a37846a  and  a37833a );
 a1019a <=( a37820a  and  a37807a );
 a1020a <=( a37796a  and  a37783a );
 a1021a <=( a37772a  and  a37759a );
 a1022a <=( a37748a  and  a37735a );
 a1023a <=( a37724a  and  a37711a );
 a1024a <=( a37700a  and  a37687a );
 a1025a <=( a37676a  and  a37663a );
 a1026a <=( a37652a  and  a37639a );
 a1027a <=( a37628a  and  a37615a );
 a1028a <=( a37604a  and  a37591a );
 a1029a <=( a37580a  and  a37567a );
 a1030a <=( a37556a  and  a37543a );
 a1031a <=( a37532a  and  a37519a );
 a1032a <=( a37508a  and  a37495a );
 a1033a <=( a37484a  and  a37471a );
 a1034a <=( a37460a  and  a37447a );
 a1035a <=( a37436a  and  a37423a );
 a1036a <=( a37412a  and  a37399a );
 a1037a <=( a37388a  and  a37375a );
 a1038a <=( a37364a  and  a37351a );
 a1039a <=( a37340a  and  a37327a );
 a1040a <=( a37316a  and  a37303a );
 a1041a <=( a37292a  and  a37279a );
 a1042a <=( a37268a  and  a37255a );
 a1043a <=( a37244a  and  a37231a );
 a1044a <=( a37220a  and  a37207a );
 a1045a <=( a37196a  and  a37183a );
 a1046a <=( a37172a  and  a37159a );
 a1047a <=( a37148a  and  a37135a );
 a1048a <=( a37124a  and  a37111a );
 a1049a <=( a37100a  and  a37087a );
 a1050a <=( a37076a  and  a37063a );
 a1051a <=( a37052a  and  a37039a );
 a1052a <=( a37028a  and  a37015a );
 a1053a <=( a37004a  and  a36991a );
 a1054a <=( a36980a  and  a36967a );
 a1055a <=( a36956a  and  a36943a );
 a1056a <=( a36932a  and  a36919a );
 a1057a <=( a36908a  and  a36895a );
 a1058a <=( a36884a  and  a36871a );
 a1059a <=( a36860a  and  a36847a );
 a1060a <=( a36836a  and  a36823a );
 a1061a <=( a36812a  and  a36799a );
 a1062a <=( a36788a  and  a36775a );
 a1063a <=( a36764a  and  a36751a );
 a1064a <=( a36740a  and  a36727a );
 a1065a <=( a36716a  and  a36703a );
 a1066a <=( a36692a  and  a36679a );
 a1067a <=( a36668a  and  a36655a );
 a1068a <=( a36644a  and  a36631a );
 a1069a <=( a36620a  and  a36607a );
 a1070a <=( a36596a  and  a36583a );
 a1071a <=( a36572a  and  a36559a );
 a1072a <=( a36548a  and  a36535a );
 a1073a <=( a36524a  and  a36511a );
 a1074a <=( a36500a  and  a36487a );
 a1075a <=( a36476a  and  a36463a );
 a1076a <=( a36452a  and  a36439a );
 a1077a <=( a36428a  and  a36415a );
 a1078a <=( a36404a  and  a36391a );
 a1079a <=( a36380a  and  a36367a );
 a1080a <=( a36356a  and  a36343a );
 a1081a <=( a36332a  and  a36319a );
 a1082a <=( a36308a  and  a36295a );
 a1083a <=( a36284a  and  a36271a );
 a1084a <=( a36260a  and  a36247a );
 a1085a <=( a36236a  and  a36223a );
 a1086a <=( a36212a  and  a36199a );
 a1087a <=( a36188a  and  a36175a );
 a1088a <=( a36164a  and  a36151a );
 a1089a <=( a36140a  and  a36127a );
 a1090a <=( a36116a  and  a36103a );
 a1091a <=( a36092a  and  a36079a );
 a1092a <=( a36068a  and  a36055a );
 a1093a <=( a36044a  and  a36031a );
 a1094a <=( a36020a  and  a36007a );
 a1095a <=( a35996a  and  a35983a );
 a1096a <=( a35972a  and  a35959a );
 a1097a <=( a35948a  and  a35935a );
 a1098a <=( a35924a  and  a35911a );
 a1099a <=( a35900a  and  a35887a );
 a1100a <=( a35876a  and  a35863a );
 a1101a <=( a35852a  and  a35839a );
 a1102a <=( a35828a  and  a35815a );
 a1103a <=( a35804a  and  a35791a );
 a1104a <=( a35780a  and  a35767a );
 a1105a <=( a35756a  and  a35743a );
 a1106a <=( a35732a  and  a35719a );
 a1107a <=( a35708a  and  a35695a );
 a1108a <=( a35684a  and  a35671a );
 a1109a <=( a35660a  and  a35647a );
 a1110a <=( a35636a  and  a35623a );
 a1111a <=( a35612a  and  a35599a );
 a1112a <=( a35588a  and  a35575a );
 a1113a <=( a35564a  and  a35551a );
 a1114a <=( a35540a  and  a35527a );
 a1115a <=( a35516a  and  a35503a );
 a1116a <=( a35492a  and  a35479a );
 a1117a <=( a35468a  and  a35455a );
 a1118a <=( a35444a  and  a35431a );
 a1119a <=( a35420a  and  a35407a );
 a1120a <=( a35396a  and  a35383a );
 a1121a <=( a35372a  and  a35359a );
 a1122a <=( a35348a  and  a35335a );
 a1123a <=( a35324a  and  a35311a );
 a1124a <=( a35300a  and  a35287a );
 a1125a <=( a35276a  and  a35263a );
 a1126a <=( a35252a  and  a35239a );
 a1127a <=( a35228a  and  a35215a );
 a1128a <=( a35204a  and  a35191a );
 a1129a <=( a35180a  and  a35167a );
 a1130a <=( a35156a  and  a35143a );
 a1131a <=( a35132a  and  a35119a );
 a1132a <=( a35108a  and  a35095a );
 a1133a <=( a35084a  and  a35071a );
 a1134a <=( a35060a  and  a35047a );
 a1135a <=( a35036a  and  a35023a );
 a1136a <=( a35012a  and  a34999a );
 a1137a <=( a34988a  and  a34975a );
 a1138a <=( a34964a  and  a34951a );
 a1139a <=( a34940a  and  a34927a );
 a1140a <=( a34916a  and  a34903a );
 a1141a <=( a34892a  and  a34879a );
 a1142a <=( a34868a  and  a34855a );
 a1143a <=( a34844a  and  a34831a );
 a1144a <=( a34820a  and  a34807a );
 a1145a <=( a34796a  and  a34783a );
 a1146a <=( a34772a  and  a34759a );
 a1147a <=( a34748a  and  a34735a );
 a1148a <=( a34724a  and  a34711a );
 a1149a <=( a34700a  and  a34687a );
 a1150a <=( a34676a  and  a34663a );
 a1151a <=( a34652a  and  a34639a );
 a1152a <=( a34628a  and  a34615a );
 a1153a <=( a34604a  and  a34591a );
 a1154a <=( a34580a  and  a34567a );
 a1155a <=( a34556a  and  a34543a );
 a1156a <=( a34532a  and  a34519a );
 a1157a <=( a34508a  and  a34495a );
 a1158a <=( a34484a  and  a34471a );
 a1159a <=( a34460a  and  a34447a );
 a1160a <=( a34436a  and  a34423a );
 a1161a <=( a34412a  and  a34399a );
 a1162a <=( a34388a  and  a34375a );
 a1163a <=( a34364a  and  a34351a );
 a1164a <=( a34340a  and  a34327a );
 a1165a <=( a34316a  and  a34303a );
 a1166a <=( a34292a  and  a34279a );
 a1167a <=( a34268a  and  a34255a );
 a1168a <=( a34244a  and  a34231a );
 a1169a <=( a34220a  and  a34207a );
 a1170a <=( a34196a  and  a34183a );
 a1171a <=( a34172a  and  a34159a );
 a1172a <=( a34148a  and  a34135a );
 a1173a <=( a34124a  and  a34111a );
 a1174a <=( a34100a  and  a34087a );
 a1175a <=( a34076a  and  a34063a );
 a1176a <=( a34052a  and  a34039a );
 a1177a <=( a34028a  and  a34015a );
 a1178a <=( a34004a  and  a33991a );
 a1179a <=( a33980a  and  a33967a );
 a1180a <=( a33956a  and  a33943a );
 a1181a <=( a33932a  and  a33919a );
 a1182a <=( a33908a  and  a33895a );
 a1183a <=( a33884a  and  a33871a );
 a1184a <=( a33860a  and  a33847a );
 a1185a <=( a33836a  and  a33823a );
 a1186a <=( a33812a  and  a33799a );
 a1187a <=( a33788a  and  a33775a );
 a1188a <=( a33764a  and  a33751a );
 a1189a <=( a33740a  and  a33727a );
 a1190a <=( a33716a  and  a33703a );
 a1191a <=( a33692a  and  a33679a );
 a1192a <=( a33668a  and  a33655a );
 a1193a <=( a33644a  and  a33631a );
 a1194a <=( a33620a  and  a33607a );
 a1195a <=( a33596a  and  a33583a );
 a1196a <=( a33572a  and  a33559a );
 a1197a <=( a33548a  and  a33535a );
 a1198a <=( a33524a  and  a33511a );
 a1199a <=( a33500a  and  a33487a );
 a1200a <=( a33476a  and  a33463a );
 a1201a <=( a33452a  and  a33439a );
 a1202a <=( a33428a  and  a33415a );
 a1203a <=( a33404a  and  a33391a );
 a1204a <=( a33380a  and  a33367a );
 a1205a <=( a33356a  and  a33343a );
 a1206a <=( a33332a  and  a33319a );
 a1207a <=( a33308a  and  a33295a );
 a1208a <=( a33284a  and  a33271a );
 a1209a <=( a33260a  and  a33247a );
 a1210a <=( a33236a  and  a33223a );
 a1211a <=( a33212a  and  a33199a );
 a1212a <=( a33188a  and  a33175a );
 a1213a <=( a33164a  and  a33151a );
 a1214a <=( a33140a  and  a33127a );
 a1215a <=( a33116a  and  a33103a );
 a1216a <=( a33092a  and  a33079a );
 a1217a <=( a33068a  and  a33055a );
 a1218a <=( a33044a  and  a33031a );
 a1219a <=( a33020a  and  a33007a );
 a1220a <=( a32996a  and  a32983a );
 a1221a <=( a32972a  and  a32959a );
 a1222a <=( a32948a  and  a32935a );
 a1223a <=( a32924a  and  a32911a );
 a1224a <=( a32900a  and  a32887a );
 a1225a <=( a32876a  and  a32863a );
 a1226a <=( a32852a  and  a32839a );
 a1227a <=( a32828a  and  a32815a );
 a1228a <=( a32804a  and  a32791a );
 a1229a <=( a32780a  and  a32767a );
 a1230a <=( a32756a  and  a32743a );
 a1231a <=( a32732a  and  a32719a );
 a1232a <=( a32708a  and  a32695a );
 a1233a <=( a32684a  and  a32671a );
 a1234a <=( a32660a  and  a32647a );
 a1235a <=( a32636a  and  a32623a );
 a1236a <=( a32612a  and  a32599a );
 a1237a <=( a32588a  and  a32575a );
 a1238a <=( a32564a  and  a32551a );
 a1239a <=( a32540a  and  a32527a );
 a1240a <=( a32516a  and  a32503a );
 a1241a <=( a32492a  and  a32479a );
 a1242a <=( a32468a  and  a32455a );
 a1243a <=( a32444a  and  a32431a );
 a1244a <=( a32420a  and  a32407a );
 a1245a <=( a32396a  and  a32383a );
 a1246a <=( a32372a  and  a32359a );
 a1247a <=( a32348a  and  a32335a );
 a1248a <=( a32324a  and  a32311a );
 a1249a <=( a32300a  and  a32287a );
 a1250a <=( a32276a  and  a32263a );
 a1251a <=( a32252a  and  a32239a );
 a1252a <=( a32228a  and  a32215a );
 a1253a <=( a32204a  and  a32191a );
 a1254a <=( a32180a  and  a32167a );
 a1255a <=( a32156a  and  a32143a );
 a1256a <=( a32132a  and  a32119a );
 a1257a <=( a32108a  and  a32095a );
 a1258a <=( a32084a  and  a32071a );
 a1259a <=( a32060a  and  a32047a );
 a1260a <=( a32036a  and  a32023a );
 a1261a <=( a32012a  and  a31999a );
 a1262a <=( a31988a  and  a31975a );
 a1263a <=( a31964a  and  a31951a );
 a1264a <=( a31940a  and  a31927a );
 a1265a <=( a31916a  and  a31903a );
 a1266a <=( a31892a  and  a31879a );
 a1267a <=( a31868a  and  a31855a );
 a1268a <=( a31844a  and  a31831a );
 a1269a <=( a31820a  and  a31807a );
 a1270a <=( a31796a  and  a31783a );
 a1271a <=( a31772a  and  a31759a );
 a1272a <=( a31748a  and  a31735a );
 a1273a <=( a31724a  and  a31711a );
 a1274a <=( a31700a  and  a31687a );
 a1275a <=( a31676a  and  a31663a );
 a1276a <=( a31652a  and  a31639a );
 a1277a <=( a31628a  and  a31615a );
 a1278a <=( a31604a  and  a31591a );
 a1279a <=( a31580a  and  a31567a );
 a1280a <=( a31556a  and  a31543a );
 a1281a <=( a31532a  and  a31519a );
 a1282a <=( a31508a  and  a31495a );
 a1283a <=( a31484a  and  a31471a );
 a1284a <=( a31460a  and  a31447a );
 a1285a <=( a31436a  and  a31423a );
 a1286a <=( a31412a  and  a31399a );
 a1287a <=( a31388a  and  a31375a );
 a1288a <=( a31364a  and  a31351a );
 a1289a <=( a31340a  and  a31327a );
 a1290a <=( a31316a  and  a31303a );
 a1291a <=( a31292a  and  a31279a );
 a1292a <=( a31268a  and  a31255a );
 a1293a <=( a31244a  and  a31231a );
 a1294a <=( a31220a  and  a31207a );
 a1295a <=( a31196a  and  a31183a );
 a1296a <=( a31172a  and  a31159a );
 a1297a <=( a31148a  and  a31135a );
 a1298a <=( a31124a  and  a31111a );
 a1299a <=( a31100a  and  a31087a );
 a1300a <=( a31076a  and  a31063a );
 a1301a <=( a31052a  and  a31039a );
 a1302a <=( a31028a  and  a31015a );
 a1303a <=( a31004a  and  a30991a );
 a1304a <=( a30980a  and  a30967a );
 a1305a <=( a30956a  and  a30943a );
 a1306a <=( a30932a  and  a30919a );
 a1307a <=( a30908a  and  a30895a );
 a1308a <=( a30884a  and  a30871a );
 a1309a <=( a30860a  and  a30847a );
 a1310a <=( a30836a  and  a30823a );
 a1311a <=( a30812a  and  a30799a );
 a1312a <=( a30788a  and  a30775a );
 a1313a <=( a30764a  and  a30751a );
 a1314a <=( a30740a  and  a30727a );
 a1315a <=( a30716a  and  a30703a );
 a1316a <=( a30692a  and  a30679a );
 a1317a <=( a30668a  and  a30655a );
 a1318a <=( a30644a  and  a30631a );
 a1319a <=( a30620a  and  a30609a );
 a1320a <=( a30598a  and  a30587a );
 a1321a <=( a30576a  and  a30565a );
 a1322a <=( a30554a  and  a30543a );
 a1323a <=( a30532a  and  a30521a );
 a1324a <=( a30510a  and  a30499a );
 a1325a <=( a30488a  and  a30477a );
 a1326a <=( a30466a  and  a30455a );
 a1327a <=( a30444a  and  a30433a );
 a1328a <=( a30422a  and  a30411a );
 a1329a <=( a30400a  and  a30389a );
 a1330a <=( a30378a  and  a30367a );
 a1331a <=( a30356a  and  a30345a );
 a1332a <=( a30334a  and  a30323a );
 a1333a <=( a30312a  and  a30301a );
 a1334a <=( a30290a  and  a30279a );
 a1335a <=( a30268a  and  a30257a );
 a1336a <=( a30246a  and  a30235a );
 a1337a <=( a30224a  and  a30213a );
 a1338a <=( a30202a  and  a30191a );
 a1339a <=( a30180a  and  a30169a );
 a1340a <=( a30158a  and  a30147a );
 a1341a <=( a30136a  and  a30125a );
 a1342a <=( a30114a  and  a30103a );
 a1343a <=( a30092a  and  a30081a );
 a1344a <=( a30070a  and  a30059a );
 a1345a <=( a30048a  and  a30037a );
 a1346a <=( a30026a  and  a30015a );
 a1347a <=( a30004a  and  a29993a );
 a1348a <=( a29982a  and  a29971a );
 a1349a <=( a29960a  and  a29949a );
 a1350a <=( a29938a  and  a29927a );
 a1351a <=( a29916a  and  a29905a );
 a1352a <=( a29894a  and  a29883a );
 a1353a <=( a29872a  and  a29861a );
 a1354a <=( a29850a  and  a29839a );
 a1355a <=( a29828a  and  a29817a );
 a1356a <=( a29806a  and  a29795a );
 a1357a <=( a29784a  and  a29773a );
 a1358a <=( a29762a  and  a29751a );
 a1359a <=( a29740a  and  a29729a );
 a1360a <=( a29718a  and  a29707a );
 a1361a <=( a29696a  and  a29685a );
 a1362a <=( a29674a  and  a29663a );
 a1363a <=( a29652a  and  a29641a );
 a1364a <=( a29630a  and  a29619a );
 a1365a <=( a29608a  and  a29597a );
 a1366a <=( a29586a  and  a29575a );
 a1367a <=( a29564a  and  a29553a );
 a1368a <=( a29542a  and  a29531a );
 a1369a <=( a29520a  and  a29509a );
 a1370a <=( a29498a  and  a29487a );
 a1371a <=( a29476a  and  a29465a );
 a1372a <=( a29454a  and  a29443a );
 a1373a <=( a29432a  and  a29421a );
 a1374a <=( a29410a  and  a29399a );
 a1375a <=( a29388a  and  a29377a );
 a1376a <=( a29366a  and  a29355a );
 a1377a <=( a29344a  and  a29333a );
 a1378a <=( a29322a  and  a29311a );
 a1379a <=( a29300a  and  a29289a );
 a1380a <=( a29278a  and  a29267a );
 a1381a <=( a29256a  and  a29245a );
 a1382a <=( a29234a  and  a29223a );
 a1383a <=( a29212a  and  a29201a );
 a1384a <=( a29190a  and  a29179a );
 a1385a <=( a29168a  and  a29157a );
 a1386a <=( a29146a  and  a29135a );
 a1387a <=( a29124a  and  a29113a );
 a1388a <=( a29102a  and  a29091a );
 a1389a <=( a29080a  and  a29069a );
 a1390a <=( a29058a  and  a29047a );
 a1391a <=( a29036a  and  a29025a );
 a1392a <=( a29014a  and  a29003a );
 a1393a <=( a28992a  and  a28981a );
 a1394a <=( a28970a  and  a28959a );
 a1395a <=( a28948a  and  a28937a );
 a1396a <=( a28926a  and  a28915a );
 a1397a <=( a28904a  and  a28893a );
 a1398a <=( a28882a  and  a28871a );
 a1399a <=( a28860a  and  a28849a );
 a1400a <=( a28838a  and  a28827a );
 a1401a <=( a28816a  and  a28805a );
 a1402a <=( a28794a  and  a28783a );
 a1403a <=( a28772a  and  a28761a );
 a1404a <=( a28750a  and  a28739a );
 a1405a <=( a28728a  and  a28717a );
 a1406a <=( a28706a  and  a28695a );
 a1407a <=( a28684a  and  a28673a );
 a1408a <=( a28662a  and  a28651a );
 a1409a <=( a28640a  and  a28629a );
 a1410a <=( a28618a  and  a28607a );
 a1411a <=( a28596a  and  a28585a );
 a1412a <=( a28574a  and  a28563a );
 a1413a <=( a28552a  and  a28541a );
 a1414a <=( a28530a  and  a28519a );
 a1415a <=( a28508a  and  a28497a );
 a1416a <=( a28486a  and  a28475a );
 a1417a <=( a28464a  and  a28453a );
 a1418a <=( a28442a  and  a28431a );
 a1419a <=( a28420a  and  a28409a );
 a1420a <=( a28398a  and  a28387a );
 a1421a <=( a28376a  and  a28365a );
 a1422a <=( a28354a  and  a28343a );
 a1423a <=( a28332a  and  a28321a );
 a1424a <=( a28310a  and  a28299a );
 a1425a <=( a28288a  and  a28277a );
 a1426a <=( a28266a  and  a28255a );
 a1427a <=( a28244a  and  a28233a );
 a1428a <=( a28222a  and  a28211a );
 a1429a <=( a28200a  and  a28189a );
 a1430a <=( a28178a  and  a28167a );
 a1431a <=( a28156a  and  a28145a );
 a1432a <=( a28134a  and  a28123a );
 a1433a <=( a28112a  and  a28101a );
 a1434a <=( a28090a  and  a28079a );
 a1435a <=( a28068a  and  a28057a );
 a1436a <=( a28046a  and  a28035a );
 a1437a <=( a28024a  and  a28013a );
 a1438a <=( a28002a  and  a27991a );
 a1439a <=( a27980a  and  a27969a );
 a1440a <=( a27958a  and  a27947a );
 a1441a <=( a27936a  and  a27925a );
 a1442a <=( a27914a  and  a27903a );
 a1443a <=( a27892a  and  a27881a );
 a1444a <=( a27870a  and  a27859a );
 a1445a <=( a27848a  and  a27837a );
 a1446a <=( a27826a  and  a27815a );
 a1447a <=( a27804a  and  a27793a );
 a1448a <=( a27782a  and  a27771a );
 a1449a <=( a27760a  and  a27749a );
 a1450a <=( a27738a  and  a27727a );
 a1451a <=( a27716a  and  a27705a );
 a1452a <=( a27694a  and  a27683a );
 a1453a <=( a27672a  and  a27661a );
 a1454a <=( a27650a  and  a27639a );
 a1455a <=( a27628a  and  a27617a );
 a1456a <=( a27606a  and  a27595a );
 a1457a <=( a27584a  and  a27573a );
 a1458a <=( a27562a  and  a27551a );
 a1459a <=( a27540a  and  a27529a );
 a1460a <=( a27518a  and  a27507a );
 a1461a <=( a27496a  and  a27485a );
 a1462a <=( a27474a  and  a27463a );
 a1463a <=( a27452a  and  a27441a );
 a1464a <=( a27430a  and  a27419a );
 a1465a <=( a27408a  and  a27397a );
 a1466a <=( a27386a  and  a27375a );
 a1467a <=( a27364a  and  a27353a );
 a1468a <=( a27342a  and  a27331a );
 a1469a <=( a27320a  and  a27309a );
 a1470a <=( a27298a  and  a27287a );
 a1471a <=( a27276a  and  a27265a );
 a1472a <=( a27254a  and  a27243a );
 a1473a <=( a27232a  and  a27221a );
 a1474a <=( a27210a  and  a27199a );
 a1475a <=( a27188a  and  a27177a );
 a1476a <=( a27166a  and  a27155a );
 a1477a <=( a27144a  and  a27133a );
 a1478a <=( a27122a  and  a27111a );
 a1479a <=( a27100a  and  a27089a );
 a1480a <=( a27078a  and  a27067a );
 a1481a <=( a27056a  and  a27045a );
 a1482a <=( a27034a  and  a27023a );
 a1483a <=( a27012a  and  a27001a );
 a1484a <=( a26990a  and  a26979a );
 a1485a <=( a26968a  and  a26957a );
 a1486a <=( a26946a  and  a26935a );
 a1487a <=( a26924a  and  a26913a );
 a1488a <=( a26902a  and  a26891a );
 a1489a <=( a26880a  and  a26869a );
 a1490a <=( a26858a  and  a26847a );
 a1491a <=( a26836a  and  a26825a );
 a1492a <=( a26814a  and  a26803a );
 a1493a <=( a26792a  and  a26781a );
 a1494a <=( a26770a  and  a26759a );
 a1495a <=( a26748a  and  a26737a );
 a1496a <=( a26726a  and  a26715a );
 a1497a <=( a26704a  and  a26693a );
 a1498a <=( a26682a  and  a26671a );
 a1499a <=( a26660a  and  a26649a );
 a1500a <=( a26638a  and  a26627a );
 a1501a <=( a26616a  and  a26605a );
 a1502a <=( a26594a  and  a26583a );
 a1503a <=( a26572a  and  a26561a );
 a1504a <=( a26550a  and  a26539a );
 a1505a <=( a26528a  and  a26517a );
 a1506a <=( a26506a  and  a26495a );
 a1507a <=( a26484a  and  a26473a );
 a1508a <=( a26462a  and  a26451a );
 a1509a <=( a26440a  and  a26429a );
 a1510a <=( a26418a  and  a26407a );
 a1511a <=( a26396a  and  a26385a );
 a1512a <=( a26374a  and  a26363a );
 a1513a <=( a26352a  and  a26341a );
 a1514a <=( a26330a  and  a26319a );
 a1515a <=( a26308a  and  a26297a );
 a1516a <=( a26286a  and  a26275a );
 a1517a <=( a26264a  and  a26253a );
 a1518a <=( a26242a  and  a26231a );
 a1519a <=( a26220a  and  a26209a );
 a1520a <=( a26198a  and  a26187a );
 a1521a <=( a26176a  and  a26165a );
 a1522a <=( a26154a  and  a26143a );
 a1523a <=( a26132a  and  a26121a );
 a1524a <=( a26110a  and  a26099a );
 a1525a <=( a26088a  and  a26077a );
 a1526a <=( a26066a  and  a26055a );
 a1527a <=( a26044a  and  a26033a );
 a1528a <=( a26022a  and  a26011a );
 a1529a <=( a26000a  and  a25989a );
 a1530a <=( a25978a  and  a25967a );
 a1531a <=( a25956a  and  a25945a );
 a1532a <=( a25934a  and  a25923a );
 a1533a <=( a25912a  and  a25901a );
 a1534a <=( a25890a  and  a25879a );
 a1535a <=( a25868a  and  a25857a );
 a1536a <=( a25846a  and  a25835a );
 a1537a <=( a25824a  and  a25813a );
 a1538a <=( a25802a  and  a25791a );
 a1539a <=( a25780a  and  a25769a );
 a1540a <=( a25758a  and  a25747a );
 a1541a <=( a25736a  and  a25725a );
 a1542a <=( a25714a  and  a25703a );
 a1543a <=( a25692a  and  a25681a );
 a1544a <=( a25670a  and  a25659a );
 a1545a <=( a25648a  and  a25637a );
 a1546a <=( a25626a  and  a25615a );
 a1547a <=( a25604a  and  a25593a );
 a1548a <=( a25582a  and  a25571a );
 a1549a <=( a25560a  and  a25549a );
 a1550a <=( a25538a  and  a25527a );
 a1551a <=( a25516a  and  a25505a );
 a1552a <=( a25494a  and  a25483a );
 a1553a <=( a25472a  and  a25461a );
 a1554a <=( a25450a  and  a25439a );
 a1555a <=( a25428a  and  a25417a );
 a1556a <=( a25406a  and  a25395a );
 a1557a <=( a25384a  and  a25373a );
 a1558a <=( a25362a  and  a25351a );
 a1559a <=( a25340a  and  a25329a );
 a1560a <=( a25318a  and  a25307a );
 a1561a <=( a25296a  and  a25285a );
 a1562a <=( a25274a  and  a25263a );
 a1563a <=( a25252a  and  a25241a );
 a1564a <=( a25230a  and  a25219a );
 a1565a <=( a25208a  and  a25197a );
 a1566a <=( a25186a  and  a25175a );
 a1567a <=( a25164a  and  a25153a );
 a1568a <=( a25142a  and  a25131a );
 a1569a <=( a25120a  and  a25109a );
 a1570a <=( a25098a  and  a25087a );
 a1571a <=( a25076a  and  a25065a );
 a1572a <=( a25054a  and  a25043a );
 a1573a <=( a25032a  and  a25021a );
 a1574a <=( a25010a  and  a24999a );
 a1575a <=( a24988a  and  a24977a );
 a1576a <=( a24966a  and  a24955a );
 a1577a <=( a24944a  and  a24933a );
 a1578a <=( a24922a  and  a24911a );
 a1579a <=( a24900a  and  a24889a );
 a1580a <=( a24878a  and  a24867a );
 a1581a <=( a24856a  and  a24845a );
 a1582a <=( a24834a  and  a24823a );
 a1583a <=( a24812a  and  a24801a );
 a1584a <=( a24790a  and  a24779a );
 a1585a <=( a24768a  and  a24757a );
 a1586a <=( a24746a  and  a24735a );
 a1587a <=( a24724a  and  a24713a );
 a1588a <=( a24702a  and  a24691a );
 a1589a <=( a24680a  and  a24669a );
 a1590a <=( a24658a  and  a24647a );
 a1591a <=( a24636a  and  a24625a );
 a1592a <=( a24614a  and  a24603a );
 a1593a <=( a24592a  and  a24581a );
 a1594a <=( a24570a  and  a24559a );
 a1595a <=( a24548a  and  a24537a );
 a1596a <=( a24526a  and  a24515a );
 a1597a <=( a24504a  and  a24493a );
 a1598a <=( a24482a  and  a24471a );
 a1599a <=( a24460a  and  a24449a );
 a1600a <=( a24440a  and  a24429a );
 a1601a <=( a24420a  and  a24409a );
 a1602a <=( a24400a  and  a24389a );
 a1603a <=( a24380a  and  a24369a );
 a1604a <=( a24360a  and  a24349a );
 a1605a <=( a24340a  and  a24329a );
 a1606a <=( a24320a  and  a24309a );
 a1607a <=( a24300a  and  a24289a );
 a1608a <=( a24280a  and  a24269a );
 a1609a <=( a24260a  and  a24249a );
 a1610a <=( a24240a  and  a24229a );
 a1611a <=( a24220a  and  a24209a );
 a1612a <=( a24200a  and  a24189a );
 a1613a <=( a24180a  and  a24169a );
 a1614a <=( a24160a  and  a24149a );
 a1615a <=( a24140a  and  a24129a );
 a1616a <=( a24120a  and  a24109a );
 a1617a <=( a24100a  and  a24089a );
 a1618a <=( a24080a  and  a24069a );
 a1619a <=( a24060a  and  a24049a );
 a1620a <=( a24040a  and  a24029a );
 a1621a <=( a24020a  and  a24009a );
 a1622a <=( a24000a  and  a23989a );
 a1623a <=( a23980a  and  a23969a );
 a1624a <=( a23960a  and  a23949a );
 a1625a <=( a23940a  and  a23929a );
 a1626a <=( a23920a  and  a23909a );
 a1627a <=( a23900a  and  a23889a );
 a1628a <=( a23880a  and  a23869a );
 a1629a <=( a23860a  and  a23849a );
 a1630a <=( a23840a  and  a23829a );
 a1631a <=( a23820a  and  a23809a );
 a1632a <=( a23800a  and  a23789a );
 a1633a <=( a23780a  and  a23769a );
 a1634a <=( a23760a  and  a23749a );
 a1635a <=( a23740a  and  a23729a );
 a1636a <=( a23720a  and  a23709a );
 a1637a <=( a23700a  and  a23689a );
 a1638a <=( a23680a  and  a23669a );
 a1639a <=( a23660a  and  a23649a );
 a1640a <=( a23640a  and  a23629a );
 a1641a <=( a23620a  and  a23609a );
 a1642a <=( a23600a  and  a23589a );
 a1643a <=( a23580a  and  a23569a );
 a1644a <=( a23560a  and  a23549a );
 a1645a <=( a23540a  and  a23529a );
 a1646a <=( a23520a  and  a23509a );
 a1647a <=( a23500a  and  a23489a );
 a1648a <=( a23480a  and  a23469a );
 a1649a <=( a23460a  and  a23449a );
 a1650a <=( a23440a  and  a23429a );
 a1651a <=( a23420a  and  a23409a );
 a1652a <=( a23400a  and  a23389a );
 a1653a <=( a23380a  and  a23369a );
 a1654a <=( a23360a  and  a23349a );
 a1655a <=( a23340a  and  a23329a );
 a1656a <=( a23320a  and  a23309a );
 a1657a <=( a23300a  and  a23289a );
 a1658a <=( a23280a  and  a23269a );
 a1659a <=( a23260a  and  a23249a );
 a1660a <=( a23240a  and  a23229a );
 a1661a <=( a23220a  and  a23209a );
 a1662a <=( a23200a  and  a23189a );
 a1663a <=( a23180a  and  a23169a );
 a1664a <=( a23160a  and  a23149a );
 a1665a <=( a23140a  and  a23129a );
 a1666a <=( a23120a  and  a23109a );
 a1667a <=( a23100a  and  a23089a );
 a1668a <=( a23080a  and  a23069a );
 a1669a <=( a23060a  and  a23049a );
 a1670a <=( a23040a  and  a23029a );
 a1671a <=( a23020a  and  a23009a );
 a1672a <=( a23000a  and  a22989a );
 a1673a <=( a22980a  and  a22969a );
 a1674a <=( a22960a  and  a22949a );
 a1675a <=( a22940a  and  a22929a );
 a1676a <=( a22920a  and  a22909a );
 a1677a <=( a22900a  and  a22889a );
 a1678a <=( a22880a  and  a22869a );
 a1679a <=( a22860a  and  a22849a );
 a1680a <=( a22840a  and  a22829a );
 a1681a <=( a22820a  and  a22809a );
 a1682a <=( a22800a  and  a22789a );
 a1683a <=( a22780a  and  a22769a );
 a1684a <=( a22760a  and  a22749a );
 a1685a <=( a22740a  and  a22729a );
 a1686a <=( a22720a  and  a22709a );
 a1687a <=( a22700a  and  a22689a );
 a1688a <=( a22680a  and  a22669a );
 a1689a <=( a22660a  and  a22649a );
 a1690a <=( a22640a  and  a22629a );
 a1691a <=( a22620a  and  a22609a );
 a1692a <=( a22600a  and  a22589a );
 a1693a <=( a22580a  and  a22569a );
 a1694a <=( a22560a  and  a22549a );
 a1695a <=( a22540a  and  a22529a );
 a1696a <=( a22520a  and  a22509a );
 a1697a <=( a22500a  and  a22489a );
 a1698a <=( a22480a  and  a22469a );
 a1699a <=( a22460a  and  a22449a );
 a1700a <=( a22440a  and  a22429a );
 a1701a <=( a22420a  and  a22409a );
 a1702a <=( a22400a  and  a22389a );
 a1703a <=( a22380a  and  a22369a );
 a1704a <=( a22360a  and  a22349a );
 a1705a <=( a22340a  and  a22329a );
 a1706a <=( a22320a  and  a22309a );
 a1707a <=( a22300a  and  a22289a );
 a1708a <=( a22280a  and  a22269a );
 a1709a <=( a22260a  and  a22249a );
 a1710a <=( a22240a  and  a22229a );
 a1711a <=( a22220a  and  a22209a );
 a1712a <=( a22200a  and  a22189a );
 a1713a <=( a22180a  and  a22169a );
 a1714a <=( a22160a  and  a22149a );
 a1715a <=( a22140a  and  a22129a );
 a1716a <=( a22120a  and  a22109a );
 a1717a <=( a22100a  and  a22089a );
 a1718a <=( a22080a  and  a22069a );
 a1719a <=( a22060a  and  a22049a );
 a1720a <=( a22040a  and  a22029a );
 a1721a <=( a22020a  and  a22009a );
 a1722a <=( a22000a  and  a21989a );
 a1723a <=( a21980a  and  a21969a );
 a1724a <=( a21960a  and  a21949a );
 a1725a <=( a21940a  and  a21929a );
 a1726a <=( a21920a  and  a21909a );
 a1727a <=( a21900a  and  a21889a );
 a1728a <=( a21880a  and  a21869a );
 a1729a <=( a21860a  and  a21849a );
 a1730a <=( a21840a  and  a21829a );
 a1731a <=( a21820a  and  a21809a );
 a1732a <=( a21800a  and  a21789a );
 a1733a <=( a21780a  and  a21769a );
 a1734a <=( a21760a  and  a21749a );
 a1735a <=( a21740a  and  a21729a );
 a1736a <=( a21720a  and  a21709a );
 a1737a <=( a21700a  and  a21689a );
 a1738a <=( a21680a  and  a21669a );
 a1739a <=( a21660a  and  a21649a );
 a1740a <=( a21640a  and  a21629a );
 a1741a <=( a21620a  and  a21609a );
 a1742a <=( a21600a  and  a21589a );
 a1743a <=( a21580a  and  a21569a );
 a1744a <=( a21560a  and  a21549a );
 a1745a <=( a21540a  and  a21529a );
 a1746a <=( a21520a  and  a21509a );
 a1747a <=( a21500a  and  a21489a );
 a1748a <=( a21480a  and  a21469a );
 a1749a <=( a21460a  and  a21449a );
 a1750a <=( a21440a  and  a21429a );
 a1751a <=( a21420a  and  a21409a );
 a1752a <=( a21400a  and  a21389a );
 a1753a <=( a21380a  and  a21369a );
 a1754a <=( a21360a  and  a21349a );
 a1755a <=( a21340a  and  a21329a );
 a1756a <=( a21320a  and  a21309a );
 a1757a <=( a21300a  and  a21289a );
 a1758a <=( a21280a  and  a21269a );
 a1759a <=( a21260a  and  a21249a );
 a1760a <=( a21240a  and  a21229a );
 a1761a <=( a21220a  and  a21209a );
 a1762a <=( a21200a  and  a21189a );
 a1763a <=( a21180a  and  a21169a );
 a1764a <=( a21160a  and  a21149a );
 a1765a <=( a21140a  and  a21129a );
 a1766a <=( a21120a  and  a21109a );
 a1767a <=( a21100a  and  a21089a );
 a1768a <=( a21080a  and  a21069a );
 a1769a <=( a21060a  and  a21049a );
 a1770a <=( a21040a  and  a21029a );
 a1771a <=( a21020a  and  a21009a );
 a1772a <=( a21000a  and  a20989a );
 a1773a <=( a20980a  and  a20969a );
 a1774a <=( a20960a  and  a20949a );
 a1775a <=( a20940a  and  a20929a );
 a1776a <=( a20920a  and  a20909a );
 a1777a <=( a20900a  and  a20889a );
 a1778a <=( a20880a  and  a20869a );
 a1779a <=( a20860a  and  a20849a );
 a1780a <=( a20840a  and  a20829a );
 a1781a <=( a20820a  and  a20809a );
 a1782a <=( a20800a  and  a20789a );
 a1783a <=( a20780a  and  a20769a );
 a1784a <=( a20760a  and  a20749a );
 a1785a <=( a20740a  and  a20729a );
 a1786a <=( a20720a  and  a20709a );
 a1787a <=( a20700a  and  a20689a );
 a1788a <=( a20680a  and  a20669a );
 a1789a <=( a20660a  and  a20649a );
 a1790a <=( a20640a  and  a20629a );
 a1791a <=( a20620a  and  a20609a );
 a1792a <=( a20600a  and  a20589a );
 a1793a <=( a20580a  and  a20569a );
 a1794a <=( a20560a  and  a20549a );
 a1795a <=( a20540a  and  a20529a );
 a1796a <=( a20520a  and  a20509a );
 a1797a <=( a20500a  and  a20489a );
 a1798a <=( a20480a  and  a20469a );
 a1799a <=( a20460a  and  a20449a );
 a1800a <=( a20440a  and  a20429a );
 a1801a <=( a20420a  and  a20409a );
 a1802a <=( a20400a  and  a20389a );
 a1803a <=( a20380a  and  a20369a );
 a1804a <=( a20360a  and  a20349a );
 a1805a <=( a20340a  and  a20329a );
 a1806a <=( a20320a  and  a20309a );
 a1807a <=( a20300a  and  a20289a );
 a1808a <=( a20280a  and  a20269a );
 a1809a <=( a20260a  and  a20249a );
 a1810a <=( a20240a  and  a20229a );
 a1811a <=( a20220a  and  a20209a );
 a1812a <=( a20200a  and  a20189a );
 a1813a <=( a20180a  and  a20169a );
 a1814a <=( a20160a  and  a20149a );
 a1815a <=( a20140a  and  a20129a );
 a1816a <=( a20120a  and  a20109a );
 a1817a <=( a20100a  and  a20089a );
 a1818a <=( a20080a  and  a20069a );
 a1819a <=( a20060a  and  a20049a );
 a1820a <=( a20040a  and  a20029a );
 a1821a <=( a20020a  and  a20009a );
 a1822a <=( a20000a  and  a19989a );
 a1823a <=( a19980a  and  a19969a );
 a1824a <=( a19960a  and  a19949a );
 a1825a <=( a19940a  and  a19929a );
 a1826a <=( a19920a  and  a19909a );
 a1827a <=( a19900a  and  a19889a );
 a1828a <=( a19880a  and  a19869a );
 a1829a <=( a19860a  and  a19849a );
 a1830a <=( a19840a  and  a19829a );
 a1831a <=( a19820a  and  a19809a );
 a1832a <=( a19800a  and  a19789a );
 a1833a <=( a19780a  and  a19769a );
 a1834a <=( a19760a  and  a19749a );
 a1835a <=( a19740a  and  a19729a );
 a1836a <=( a19720a  and  a19709a );
 a1837a <=( a19700a  and  a19689a );
 a1838a <=( a19680a  and  a19669a );
 a1839a <=( a19660a  and  a19649a );
 a1840a <=( a19640a  and  a19629a );
 a1841a <=( a19620a  and  a19609a );
 a1842a <=( a19600a  and  a19589a );
 a1843a <=( a19580a  and  a19569a );
 a1844a <=( a19560a  and  a19549a );
 a1845a <=( a19540a  and  a19529a );
 a1846a <=( a19520a  and  a19509a );
 a1847a <=( a19500a  and  a19489a );
 a1848a <=( a19480a  and  a19469a );
 a1849a <=( a19460a  and  a19449a );
 a1850a <=( a19440a  and  a19429a );
 a1851a <=( a19420a  and  a19409a );
 a1852a <=( a19400a  and  a19389a );
 a1853a <=( a19380a  and  a19369a );
 a1854a <=( a19360a  and  a19349a );
 a1855a <=( a19340a  and  a19329a );
 a1856a <=( a19320a  and  a19309a );
 a1857a <=( a19300a  and  a19289a );
 a1858a <=( a19280a  and  a19269a );
 a1859a <=( a19260a  and  a19249a );
 a1860a <=( a19240a  and  a19229a );
 a1861a <=( a19220a  and  a19209a );
 a1862a <=( a19200a  and  a19189a );
 a1863a <=( a19180a  and  a19169a );
 a1864a <=( a19160a  and  a19149a );
 a1865a <=( a19140a  and  a19129a );
 a1866a <=( a19120a  and  a19109a );
 a1867a <=( a19100a  and  a19089a );
 a1868a <=( a19080a  and  a19069a );
 a1869a <=( a19060a  and  a19049a );
 a1870a <=( a19040a  and  a19029a );
 a1871a <=( a19020a  and  a19009a );
 a1872a <=( a19000a  and  a18989a );
 a1873a <=( a18980a  and  a18969a );
 a1874a <=( a18960a  and  a18949a );
 a1875a <=( a18940a  and  a18929a );
 a1876a <=( a18920a  and  a18909a );
 a1877a <=( a18900a  and  a18889a );
 a1878a <=( a18880a  and  a18869a );
 a1879a <=( a18860a  and  a18849a );
 a1880a <=( a18840a  and  a18829a );
 a1881a <=( a18820a  and  a18809a );
 a1882a <=( a18800a  and  a18789a );
 a1883a <=( a18780a  and  a18769a );
 a1884a <=( a18760a  and  a18749a );
 a1885a <=( a18740a  and  a18729a );
 a1886a <=( a18720a  and  a18709a );
 a1887a <=( a18700a  and  a18689a );
 a1888a <=( a18680a  and  a18669a );
 a1889a <=( a18660a  and  a18649a );
 a1890a <=( a18640a  and  a18629a );
 a1891a <=( a18620a  and  a18609a );
 a1892a <=( a18600a  and  a18589a );
 a1893a <=( a18580a  and  a18569a );
 a1894a <=( a18560a  and  a18549a );
 a1895a <=( a18540a  and  a18529a );
 a1896a <=( a18520a  and  a18509a );
 a1897a <=( a18500a  and  a18489a );
 a1898a <=( a18480a  and  a18469a );
 a1899a <=( a18460a  and  a18449a );
 a1900a <=( a18440a  and  a18429a );
 a1901a <=( a18420a  and  a18409a );
 a1902a <=( a18400a  and  a18389a );
 a1903a <=( a18380a  and  a18369a );
 a1904a <=( a18360a  and  a18349a );
 a1905a <=( a18340a  and  a18329a );
 a1906a <=( a18320a  and  a18309a );
 a1907a <=( a18300a  and  a18289a );
 a1908a <=( a18280a  and  a18269a );
 a1909a <=( a18260a  and  a18249a );
 a1910a <=( a18240a  and  a18229a );
 a1911a <=( a18220a  and  a18209a );
 a1912a <=( a18200a  and  a18189a );
 a1913a <=( a18180a  and  a18169a );
 a1914a <=( a18160a  and  a18149a );
 a1915a <=( a18140a  and  a18129a );
 a1916a <=( a18120a  and  a18109a );
 a1917a <=( a18100a  and  a18089a );
 a1918a <=( a18080a  and  a18069a );
 a1919a <=( a18060a  and  a18051a );
 a1920a <=( a18042a  and  a18033a );
 a1921a <=( a18024a  and  a18015a );
 a1922a <=( a18006a  and  a17997a );
 a1923a <=( a17988a  and  a17979a );
 a1924a <=( a17970a  and  a17961a );
 a1925a <=( a17952a  and  a17943a );
 a1926a <=( a17934a  and  a17925a );
 a1927a <=( a17916a  and  a17907a );
 a1928a <=( a17898a  and  a17889a );
 a1929a <=( a17880a  and  a17871a );
 a1930a <=( a17862a  and  a17853a );
 a1931a <=( a17844a  and  a17835a );
 a1932a <=( a17826a  and  a17817a );
 a1933a <=( a17808a  and  a17799a );
 a1934a <=( a17790a  and  a17781a );
 a1935a <=( a17772a  and  a17763a );
 a1936a <=( a17754a  and  a17745a );
 a1937a <=( a17736a  and  a17727a );
 a1938a <=( a17718a  and  a17709a );
 a1939a <=( a17700a  and  a17691a );
 a1940a <=( a17682a  and  a17673a );
 a1941a <=( a17664a  and  a17655a );
 a1942a <=( a17646a  and  a17637a );
 a1943a <=( a17628a  and  a17619a );
 a1944a <=( a17610a  and  a17601a );
 a1945a <=( a17592a  and  a17583a );
 a1946a <=( a17574a  and  a17565a );
 a1947a <=( a17556a  and  a17547a );
 a1948a <=( a17538a  and  a17529a );
 a1949a <=( a17520a  and  a17511a );
 a1950a <=( a17502a  and  a17493a );
 a1951a <=( a17484a  and  a17475a );
 a1952a <=( a17466a  and  a17457a );
 a1953a <=( a17448a  and  a17439a );
 a1954a <=( a17430a  and  a17421a );
 a1955a <=( a17412a  and  a17403a );
 a1956a <=( a17394a  and  a17385a );
 a1957a <=( a17376a  and  a17367a );
 a1958a <=( a17358a  and  a17349a );
 a1959a <=( a17340a  and  a17331a );
 a1960a <=( a17322a  and  a17313a );
 a1961a <=( a17304a  and  a17295a );
 a1962a <=( a17286a  and  a17277a );
 a1963a <=( a17268a  and  a17259a );
 a1964a <=( a17250a  and  a17241a );
 a1965a <=( a17232a  and  a17223a );
 a1966a <=( a17214a  and  a17205a );
 a1967a <=( a17196a  and  a17187a );
 a1968a <=( a17178a  and  a17169a );
 a1969a <=( a17160a  and  a17151a );
 a1970a <=( a17142a  and  a17133a );
 a1971a <=( a17124a  and  a17115a );
 a1972a <=( a17106a  and  a17097a );
 a1973a <=( a17088a  and  a17079a );
 a1974a <=( a17070a  and  a17061a );
 a1975a <=( a17052a  and  a17043a );
 a1976a <=( a17034a  and  a17025a );
 a1977a <=( a17016a  and  a17007a );
 a1978a <=( a16998a  and  a16989a );
 a1979a <=( a16980a  and  a16971a );
 a1980a <=( a16962a  and  a16953a );
 a1981a <=( a16944a  and  a16935a );
 a1982a <=( a16926a  and  a16917a );
 a1983a <=( a16908a  and  a16899a );
 a1984a <=( a16890a  and  a16881a );
 a1985a <=( a16872a  and  a16863a );
 a1986a <=( a16854a  and  a16845a );
 a1987a <=( a16836a  and  a16827a );
 a1988a <=( a16818a  and  a16809a );
 a1989a <=( a16800a  and  a16791a );
 a1990a <=( a16782a  and  a16773a );
 a1991a <=( a16764a  and  a16755a );
 a1992a <=( a16746a  and  a16737a );
 a1993a <=( a16728a  and  a16719a );
 a1994a <=( a16710a  and  a16701a );
 a1995a <=( a16692a  and  a16683a );
 a1996a <=( a16674a  and  a16665a );
 a1997a <=( a16656a  and  a16647a );
 a1998a <=( a16638a  and  a16629a );
 a1999a <=( a16620a  and  a16611a );
 a2000a <=( a16602a  and  a16593a );
 a2001a <=( a16584a  and  a16575a );
 a2002a <=( a16566a  and  a16557a );
 a2003a <=( a16548a  and  a16539a );
 a2004a <=( a16530a  and  a16521a );
 a2005a <=( a16512a  and  a16503a );
 a2006a <=( a16494a  and  a16485a );
 a2007a <=( a16476a  and  a16467a );
 a2008a <=( a16458a  and  a16449a );
 a2009a <=( a16440a  and  a16431a );
 a2010a <=( a16422a  and  a16413a );
 a2011a <=( a16404a  and  a16395a );
 a2012a <=( a16386a  and  a16377a );
 a2013a <=( a16368a  and  a16359a );
 a2014a <=( a16350a  and  a16341a );
 a2015a <=( a16332a  and  a16323a );
 a2016a <=( a16314a  and  a16305a );
 a2017a <=( a16296a  and  a16287a );
 a2018a <=( a16278a  and  a16269a );
 a2019a <=( a16260a  and  a16251a );
 a2020a <=( a16242a  and  a16233a );
 a2021a <=( a16224a  and  a16215a );
 a2022a <=( a16206a  and  a16197a );
 a2023a <=( a16188a  and  a16179a );
 a2024a <=( a16170a  and  a16161a );
 a2025a <=( a16152a  and  a16143a );
 a2026a <=( a16134a  and  a16125a );
 a2027a <=( a16116a  and  a16107a );
 a2028a <=( a16098a  and  a16089a );
 a2029a <=( a16080a  and  a16071a );
 a2030a <=( a16062a  and  a16053a );
 a2031a <=( a16044a  and  a16035a );
 a2032a <=( a16026a  and  a16017a );
 a2033a <=( a16008a  and  a15999a );
 a2034a <=( a15990a  and  a15981a );
 a2035a <=( a15972a  and  a15963a );
 a2036a <=( a15954a  and  a15945a );
 a2037a <=( a15936a  and  a15927a );
 a2038a <=( a15918a  and  a15909a );
 a2039a <=( a15900a  and  a15891a );
 a2040a <=( a15882a  and  a15873a );
 a2041a <=( a15864a  and  a15855a );
 a2042a <=( a15846a  and  a15837a );
 a2043a <=( a15828a  and  a15819a );
 a2044a <=( a15810a  and  a15801a );
 a2045a <=( a15792a  and  a15783a );
 a2046a <=( a15774a  and  a15765a );
 a2047a <=( a15756a  and  a15747a );
 a2048a <=( a15738a  and  a15729a );
 a2049a <=( a15720a  and  a15711a );
 a2050a <=( a15702a  and  a15693a );
 a2051a <=( a15684a  and  a15675a );
 a2052a <=( a15666a  and  a15657a );
 a2053a <=( a15648a  and  a15639a );
 a2054a <=( a15630a  and  a15621a );
 a2055a <=( a15612a  and  a15603a );
 a2056a <=( a15594a  and  a15585a );
 a2057a <=( a15576a  and  a15567a );
 a2058a <=( a15558a  and  a15549a );
 a2059a <=( a15540a  and  a15531a );
 a2060a <=( a15522a  and  a15513a );
 a2061a <=( a15504a  and  a15495a );
 a2062a <=( a15486a  and  a15477a );
 a2063a <=( a15468a  and  a15459a );
 a2064a <=( a15450a  and  a15441a );
 a2065a <=( a15432a  and  a15423a );
 a2066a <=( a15414a  and  a15405a );
 a2067a <=( a15396a  and  a15387a );
 a2068a <=( a15378a  and  a15369a );
 a2069a <=( a15360a  and  a15351a );
 a2070a <=( a15342a  and  a15333a );
 a2071a <=( a15324a  and  a15315a );
 a2072a <=( a15306a  and  a15297a );
 a2073a <=( a15288a  and  a15279a );
 a2074a <=( a15270a  and  a15261a );
 a2075a <=( a15252a  and  a15243a );
 a2076a <=( a15234a  and  a15225a );
 a2077a <=( a15216a  and  a15207a );
 a2078a <=( a15198a  and  a15189a );
 a2079a <=( a15180a  and  a15171a );
 a2080a <=( a15162a  and  a15153a );
 a2081a <=( a15144a  and  a15135a );
 a2082a <=( a15126a  and  a15117a );
 a2083a <=( a15108a  and  a15099a );
 a2084a <=( a15090a  and  a15081a );
 a2085a <=( a15072a  and  a15063a );
 a2086a <=( a15054a  and  a15045a );
 a2087a <=( a15036a  and  a15027a );
 a2088a <=( a15018a  and  a15009a );
 a2089a <=( a15000a  and  a14991a );
 a2090a <=( a14982a  and  a14973a );
 a2091a <=( a14964a  and  a14955a );
 a2092a <=( a14946a  and  a14937a );
 a2093a <=( a14928a  and  a14919a );
 a2094a <=( a14910a  and  a14901a );
 a2095a <=( a14892a  and  a14883a );
 a2096a <=( a14874a  and  a14865a );
 a2097a <=( a14856a  and  a14847a );
 a2098a <=( a14838a  and  a14829a );
 a2099a <=( a14820a  and  a14811a );
 a2100a <=( a14802a  and  a14793a );
 a2101a <=( a14784a  and  a14775a );
 a2102a <=( a14766a  and  a14757a );
 a2103a <=( a14748a  and  a14739a );
 a2104a <=( a14730a  and  a14721a );
 a2105a <=( a14712a  and  a14703a );
 a2106a <=( a14694a  and  a14685a );
 a2107a <=( a14676a  and  a14667a );
 a2108a <=( a14658a  and  a14649a );
 a2109a <=( a14640a  and  a14631a );
 a2110a <=( a14622a  and  a14613a );
 a2111a <=( a14604a  and  a14595a );
 a2112a <=( a14586a  and  a14577a );
 a2113a <=( a14568a  and  a14559a );
 a2114a <=( a14550a  and  a14541a );
 a2115a <=( a14532a  and  a14523a );
 a2116a <=( a14514a  and  a14505a );
 a2117a <=( a14496a  and  a14487a );
 a2118a <=( a14478a  and  a14469a );
 a2119a <=( a14460a  and  a14451a );
 a2120a <=( a14442a  and  a14433a );
 a2121a <=( a14424a  and  a14415a );
 a2122a <=( a14406a  and  a14397a );
 a2123a <=( a14388a  and  a14379a );
 a2124a <=( a14370a  and  a14361a );
 a2125a <=( a14352a  and  a14343a );
 a2126a <=( a14334a  and  a14325a );
 a2127a <=( a14316a  and  a14307a );
 a2128a <=( a14298a  and  a14289a );
 a2129a <=( a14280a  and  a14271a );
 a2130a <=( a14262a  and  a14253a );
 a2131a <=( a14244a  and  a14235a );
 a2132a <=( a14226a  and  a14217a );
 a2133a <=( a14208a  and  a14199a );
 a2134a <=( a14190a  and  a14181a );
 a2135a <=( a14172a  and  a14163a );
 a2136a <=( a14154a  and  a14145a );
 a2137a <=( a14136a  and  a14127a );
 a2138a <=( a14118a  and  a14109a );
 a2139a <=( a14100a  and  a14091a );
 a2140a <=( a14082a  and  a14073a );
 a2141a <=( a14064a  and  a14055a );
 a2142a <=( a14046a  and  a14037a );
 a2143a <=( a14028a  and  a14019a );
 a2144a <=( a14010a  and  a14001a );
 a2145a <=( a13992a  and  a13983a );
 a2146a <=( a13974a  and  a13965a );
 a2147a <=( a13956a  and  a13947a );
 a2148a <=( a13938a  and  a13929a );
 a2149a <=( a13920a  and  a13911a );
 a2150a <=( a13902a  and  a13893a );
 a2151a <=( a13884a  and  a13875a );
 a2152a <=( a13866a  and  a13857a );
 a2153a <=( a13848a  and  a13839a );
 a2154a <=( a13830a  and  a13821a );
 a2155a <=( a13812a  and  a13803a );
 a2156a <=( a13794a  and  a13785a );
 a2157a <=( a13776a  and  a13767a );
 a2158a <=( a13758a  and  a13749a );
 a2159a <=( a13740a  and  a13731a );
 a2160a <=( a13722a  and  a13713a );
 a2161a <=( a13704a  and  a13695a );
 a2162a <=( a13686a  and  a13677a );
 a2163a <=( a13668a  and  a13659a );
 a2164a <=( a13650a  and  a13641a );
 a2165a <=( a13632a  and  a13623a );
 a2166a <=( a13614a  and  a13605a );
 a2167a <=( a13596a  and  a13587a );
 a2168a <=( a13578a  and  a13569a );
 a2169a <=( a13560a  and  a13551a );
 a2170a <=( a13542a  and  a13533a );
 a2171a <=( a13524a  and  a13515a );
 a2172a <=( a13506a  and  a13497a );
 a2173a <=( a13488a  and  a13479a );
 a2174a <=( a13470a  and  a13461a );
 a2175a <=( a13452a  and  a13443a );
 a2176a <=( a13434a  and  a13425a );
 a2177a <=( a13416a  and  a13407a );
 a2178a <=( a13398a  and  a13389a );
 a2179a <=( a13380a  and  a13371a );
 a2180a <=( a13362a  and  a13353a );
 a2181a <=( a13344a  and  a13335a );
 a2182a <=( a13326a  and  a13317a );
 a2183a <=( a13308a  and  a13299a );
 a2184a <=( a13290a  and  a13281a );
 a2185a <=( a13272a  and  a13263a );
 a2186a <=( a13254a  and  a13245a );
 a2187a <=( a13236a  and  a13227a );
 a2188a <=( a13218a  and  a13209a );
 a2189a <=( a13200a  and  a13191a );
 a2190a <=( a13182a  and  a13173a );
 a2191a <=( a13164a  and  a13155a );
 a2192a <=( a13146a  and  a13137a );
 a2193a <=( a13128a  and  a13119a );
 a2194a <=( a13110a  and  a13101a );
 a2195a <=( a13092a  and  a13083a );
 a2196a <=( a13074a  and  a13065a );
 a2197a <=( a13056a  and  a13047a );
 a2198a <=( a13038a  and  a13029a );
 a2199a <=( a13020a  and  a13011a );
 a2200a <=( a13002a  and  a12993a );
 a2201a <=( a12984a  and  a12975a );
 a2202a <=( a12966a  and  a12957a );
 a2203a <=( a12948a  and  a12939a );
 a2204a <=( a12930a  and  a12921a );
 a2205a <=( a12912a  and  a12903a );
 a2206a <=( a12894a  and  a12885a );
 a2207a <=( a12876a  and  a12867a );
 a2208a <=( a12858a  and  a12849a );
 a2209a <=( a12840a  and  a12831a );
 a2210a <=( a12822a  and  a12813a );
 a2211a <=( a12804a  and  a12795a );
 a2212a <=( a12786a  and  a12777a );
 a2213a <=( a12768a  and  a12759a );
 a2214a <=( a12750a  and  a12741a );
 a2215a <=( a12732a  and  a12723a );
 a2216a <=( a12714a  and  a12705a );
 a2217a <=( a12696a  and  a12687a );
 a2218a <=( a12678a  and  a12669a );
 a2219a <=( a12660a  and  a12651a );
 a2220a <=( a12642a  and  a12633a );
 a2221a <=( a12624a  and  a12615a );
 a2222a <=( a12606a  and  a12597a );
 a2223a <=( a12588a  and  a12579a );
 a2224a <=( a12570a  and  a12561a );
 a2225a <=( a12552a  and  a12543a );
 a2226a <=( a12536a  and  a12527a );
 a2227a <=( a12520a  and  a12511a );
 a2228a <=( a12504a  and  a12495a );
 a2229a <=( a12488a  and  a12479a );
 a2230a <=( a12472a  and  a12463a );
 a2231a <=( a12456a  and  a12447a );
 a2232a <=( a12440a  and  a12431a );
 a2233a <=( a12424a  and  a12415a );
 a2234a <=( a12408a  and  a12399a );
 a2235a <=( a12392a  and  a12383a );
 a2236a <=( a12376a  and  a12367a );
 a2237a <=( a12360a  and  a12351a );
 a2238a <=( a12344a  and  a12335a );
 a2239a <=( a12328a  and  a12319a );
 a2240a <=( a12312a  and  a12303a );
 a2241a <=( a12296a  and  a12287a );
 a2242a <=( a12280a  and  a12271a );
 a2243a <=( a12264a  and  a12255a );
 a2244a <=( a12248a  and  a12239a );
 a2245a <=( a12232a  and  a12223a );
 a2246a <=( a12216a  and  a12207a );
 a2247a <=( a12200a  and  a12191a );
 a2248a <=( a12184a  and  a12175a );
 a2249a <=( a12168a  and  a12159a );
 a2250a <=( a12152a  and  a12143a );
 a2251a <=( a12136a  and  a12127a );
 a2252a <=( a12120a  and  a12111a );
 a2253a <=( a12104a  and  a12095a );
 a2254a <=( a12088a  and  a12079a );
 a2255a <=( a12072a  and  a12063a );
 a2256a <=( a12056a  and  a12047a );
 a2257a <=( a12040a  and  a12031a );
 a2258a <=( a12024a  and  a12015a );
 a2259a <=( a12008a  and  a11999a );
 a2260a <=( a11992a  and  a11983a );
 a2261a <=( a11976a  and  a11967a );
 a2262a <=( a11960a  and  a11951a );
 a2263a <=( a11944a  and  a11935a );
 a2264a <=( a11928a  and  a11919a );
 a2265a <=( a11912a  and  a11903a );
 a2266a <=( a11896a  and  a11887a );
 a2267a <=( a11880a  and  a11871a );
 a2268a <=( a11864a  and  a11855a );
 a2269a <=( a11848a  and  a11839a );
 a2270a <=( a11832a  and  a11823a );
 a2271a <=( a11816a  and  a11807a );
 a2272a <=( a11800a  and  a11791a );
 a2273a <=( a11784a  and  a11775a );
 a2274a <=( a11768a  and  a11759a );
 a2275a <=( a11752a  and  a11743a );
 a2276a <=( a11736a  and  a11727a );
 a2277a <=( a11720a  and  a11711a );
 a2278a <=( a11704a  and  a11695a );
 a2279a <=( a11688a  and  a11679a );
 a2280a <=( a11672a  and  a11663a );
 a2281a <=( a11656a  and  a11647a );
 a2282a <=( a11640a  and  a11631a );
 a2283a <=( a11624a  and  a11615a );
 a2284a <=( a11608a  and  a11599a );
 a2285a <=( a11592a  and  a11583a );
 a2286a <=( a11576a  and  a11567a );
 a2287a <=( a11560a  and  a11551a );
 a2288a <=( a11544a  and  a11535a );
 a2289a <=( a11528a  and  a11519a );
 a2290a <=( a11512a  and  a11503a );
 a2291a <=( a11496a  and  a11487a );
 a2292a <=( a11480a  and  a11471a );
 a2293a <=( a11464a  and  a11455a );
 a2294a <=( a11448a  and  a11439a );
 a2295a <=( a11432a  and  a11423a );
 a2296a <=( a11416a  and  a11407a );
 a2297a <=( a11400a  and  a11391a );
 a2298a <=( a11384a  and  a11375a );
 a2299a <=( a11368a  and  a11359a );
 a2300a <=( a11352a  and  a11343a );
 a2301a <=( a11336a  and  a11327a );
 a2302a <=( a11320a  and  a11311a );
 a2303a <=( a11304a  and  a11295a );
 a2304a <=( a11288a  and  a11279a );
 a2305a <=( a11272a  and  a11263a );
 a2306a <=( a11256a  and  a11247a );
 a2307a <=( a11240a  and  a11231a );
 a2308a <=( a11224a  and  a11215a );
 a2309a <=( a11208a  and  a11199a );
 a2310a <=( a11192a  and  a11183a );
 a2311a <=( a11176a  and  a11167a );
 a2312a <=( a11160a  and  a11151a );
 a2313a <=( a11144a  and  a11135a );
 a2314a <=( a11128a  and  a11119a );
 a2315a <=( a11112a  and  a11103a );
 a2316a <=( a11096a  and  a11087a );
 a2317a <=( a11080a  and  a11071a );
 a2318a <=( a11064a  and  a11055a );
 a2319a <=( a11048a  and  a11039a );
 a2320a <=( a11032a  and  a11023a );
 a2321a <=( a11016a  and  a11007a );
 a2322a <=( a11000a  and  a10991a );
 a2323a <=( a10984a  and  a10975a );
 a2324a <=( a10968a  and  a10959a );
 a2325a <=( a10952a  and  a10943a );
 a2326a <=( a10936a  and  a10927a );
 a2327a <=( a10920a  and  a10911a );
 a2328a <=( a10904a  and  a10895a );
 a2329a <=( a10888a  and  a10879a );
 a2330a <=( a10872a  and  a10863a );
 a2331a <=( a10856a  and  a10847a );
 a2332a <=( a10840a  and  a10831a );
 a2333a <=( a10824a  and  a10815a );
 a2334a <=( a10808a  and  a10799a );
 a2335a <=( a10792a  and  a10783a );
 a2336a <=( a10776a  and  a10767a );
 a2337a <=( a10760a  and  a10751a );
 a2338a <=( a10744a  and  a10735a );
 a2339a <=( a10728a  and  a10719a );
 a2340a <=( a10712a  and  a10703a );
 a2341a <=( a10696a  and  a10687a );
 a2342a <=( a10680a  and  a10671a );
 a2343a <=( a10664a  and  a10655a );
 a2344a <=( a10648a  and  a10639a );
 a2345a <=( a10632a  and  a10623a );
 a2346a <=( a10616a  and  a10607a );
 a2347a <=( a10600a  and  a10591a );
 a2348a <=( a10584a  and  a10575a );
 a2349a <=( a10568a  and  a10559a );
 a2350a <=( a10552a  and  a10543a );
 a2351a <=( a10536a  and  a10527a );
 a2352a <=( a10520a  and  a10511a );
 a2353a <=( a10504a  and  a10495a );
 a2354a <=( a10488a  and  a10479a );
 a2355a <=( a10472a  and  a10463a );
 a2356a <=( a10456a  and  a10447a );
 a2357a <=( a10440a  and  a10431a );
 a2358a <=( a10424a  and  a10415a );
 a2359a <=( a10408a  and  a10399a );
 a2360a <=( a10392a  and  a10383a );
 a2361a <=( a10376a  and  a10367a );
 a2362a <=( a10360a  and  a10351a );
 a2363a <=( a10344a  and  a10335a );
 a2364a <=( a10328a  and  a10319a );
 a2365a <=( a10312a  and  a10303a );
 a2366a <=( a10296a  and  a10287a );
 a2367a <=( a10280a  and  a10271a );
 a2368a <=( a10264a  and  a10255a );
 a2369a <=( a10248a  and  a10239a );
 a2370a <=( a10232a  and  a10223a );
 a2371a <=( a10216a  and  a10207a );
 a2372a <=( a10200a  and  a10191a );
 a2373a <=( a10184a  and  a10175a );
 a2374a <=( a10168a  and  a10159a );
 a2375a <=( a10152a  and  a10143a );
 a2376a <=( a10136a  and  a10127a );
 a2377a <=( a10120a  and  a10111a );
 a2378a <=( a10104a  and  a10095a );
 a2379a <=( a10088a  and  a10079a );
 a2380a <=( a10072a  and  a10063a );
 a2381a <=( a10056a  and  a10047a );
 a2382a <=( a10040a  and  a10031a );
 a2383a <=( a10024a  and  a10015a );
 a2384a <=( a10008a  and  a9999a );
 a2385a <=( a9992a  and  a9983a );
 a2386a <=( a9976a  and  a9967a );
 a2387a <=( a9960a  and  a9951a );
 a2388a <=( a9944a  and  a9935a );
 a2389a <=( a9928a  and  a9919a );
 a2390a <=( a9912a  and  a9903a );
 a2391a <=( a9896a  and  a9887a );
 a2392a <=( a9880a  and  a9871a );
 a2393a <=( a9864a  and  a9855a );
 a2394a <=( a9848a  and  a9839a );
 a2395a <=( a9832a  and  a9823a );
 a2396a <=( a9816a  and  a9807a );
 a2397a <=( a9800a  and  a9791a );
 a2398a <=( a9784a  and  a9775a );
 a2399a <=( a9768a  and  a9759a );
 a2400a <=( a9752a  and  a9743a );
 a2401a <=( a9736a  and  a9727a );
 a2402a <=( a9720a  and  a9711a );
 a2403a <=( a9704a  and  a9695a );
 a2404a <=( a9688a  and  a9679a );
 a2405a <=( a9672a  and  a9663a );
 a2406a <=( a9656a  and  a9647a );
 a2407a <=( a9640a  and  a9631a );
 a2408a <=( a9624a  and  a9615a );
 a2409a <=( a9608a  and  a9599a );
 a2410a <=( a9592a  and  a9583a );
 a2411a <=( a9576a  and  a9567a );
 a2412a <=( a9560a  and  a9551a );
 a2413a <=( a9544a  and  a9535a );
 a2414a <=( a9528a  and  a9519a );
 a2415a <=( a9512a  and  a9503a );
 a2416a <=( a9496a  and  a9487a );
 a2417a <=( a9480a  and  a9471a );
 a2418a <=( a9464a  and  a9455a );
 a2419a <=( a9448a  and  a9439a );
 a2420a <=( a9432a  and  a9423a );
 a2421a <=( a9416a  and  a9407a );
 a2422a <=( a9400a  and  a9391a );
 a2423a <=( a9384a  and  a9375a );
 a2424a <=( a9368a  and  a9359a );
 a2425a <=( a9352a  and  a9343a );
 a2426a <=( a9336a  and  a9327a );
 a2427a <=( a9320a  and  a9311a );
 a2428a <=( a9304a  and  a9295a );
 a2429a <=( a9288a  and  a9281a );
 a2430a <=( a9274a  and  a9267a );
 a2431a <=( a9260a  and  a9253a );
 a2432a <=( a9246a  and  a9239a );
 a2433a <=( a9232a  and  a9225a );
 a2434a <=( a9218a  and  a9211a );
 a2435a <=( a9204a  and  a9197a );
 a2436a <=( a9190a  and  a9183a );
 a2437a <=( a9176a  and  a9169a );
 a2438a <=( a9162a  and  a9155a );
 a2439a <=( a9148a  and  a9141a );
 a2440a <=( a9134a  and  a9127a );
 a2441a <=( a9120a  and  a9113a );
 a2442a <=( a9106a  and  a9099a );
 a2443a <=( a9092a  and  a9085a );
 a2444a <=( a9078a  and  a9071a );
 a2445a <=( a9064a  and  a9057a );
 a2446a <=( a9050a  and  a9043a );
 a2447a <=( a9036a  and  a9029a );
 a2448a <=( a9022a  and  a9015a );
 a2449a <=( a9008a  and  a9001a );
 a2450a <=( a8994a  and  a8987a );
 a2451a <=( a8980a  and  a8973a );
 a2452a <=( a8966a  and  a8959a );
 a2453a <=( a8952a  and  a8945a );
 a2454a <=( a8938a  and  a8931a );
 a2455a <=( a8924a  and  a8917a );
 a2456a <=( a8910a  and  a8903a );
 a2457a <=( a8896a  and  a8889a );
 a2458a <=( a8882a  and  a8875a );
 a2459a <=( a8868a  and  a8861a );
 a2460a <=( a8854a  and  a8847a );
 a2461a <=( a8840a  and  a8833a );
 a2462a <=( a8826a  and  a8819a );
 a2463a <=( a8812a  and  a8805a );
 a2464a <=( a8798a  and  a8791a );
 a2465a <=( a8784a  and  a8777a );
 a2466a <=( a8770a  and  a8763a );
 a2467a <=( a8756a  and  a8749a );
 a2468a <=( a8742a  and  a8735a );
 a2469a <=( a8728a  and  a8721a );
 a2470a <=( a8714a  and  a8707a );
 a2471a <=( a8700a  and  a8693a );
 a2472a <=( a8686a  and  a8679a );
 a2473a <=( a8672a  and  a8665a );
 a2474a <=( a8658a  and  a8651a );
 a2475a <=( a8644a  and  a8637a );
 a2476a <=( a8630a  and  a8623a );
 a2477a <=( a8616a  and  a8609a );
 a2478a <=( a8602a  and  a8595a );
 a2479a <=( a8588a  and  a8581a );
 a2480a <=( a8574a  and  a8567a );
 a2481a <=( a8560a  and  a8553a );
 a2482a <=( a8546a  and  a8539a );
 a2483a <=( a8532a  and  a8525a );
 a2484a <=( a8518a  and  a8511a );
 a2485a <=( a8504a  and  a8497a );
 a2486a <=( a8490a  and  a8483a );
 a2487a <=( a8476a  and  a8469a );
 a2488a <=( a8462a  and  a8455a );
 a2489a <=( a8448a  and  a8441a );
 a2490a <=( a8434a  and  a8427a );
 a2491a <=( a8420a  and  a8413a );
 a2492a <=( a8406a  and  a8399a );
 a2493a <=( a8392a  and  a8385a );
 a2494a <=( a8378a  and  a8371a );
 a2495a <=( a8364a  and  a8357a );
 a2496a <=( a8350a  and  a8343a );
 a2497a <=( a8336a  and  a8329a );
 a2498a <=( a8322a  and  a8315a );
 a2499a <=( a8308a  and  a8301a );
 a2500a <=( a8294a  and  a8287a );
 a2501a <=( a8280a  and  a8273a );
 a2502a <=( a8266a  and  a8259a );
 a2503a <=( a8252a  and  a8245a );
 a2504a <=( a8238a  and  a8231a );
 a2505a <=( a8224a  and  a8217a );
 a2506a <=( a8210a  and  a8203a );
 a2507a <=( a8196a  and  a8189a );
 a2508a <=( a8182a  and  a8175a );
 a2509a <=( a8168a  and  a8161a );
 a2510a <=( a8154a  and  a8147a );
 a2511a <=( a8140a  and  a8133a );
 a2512a <=( a8126a  and  a8119a );
 a2513a <=( a8112a  and  a8105a );
 a2514a <=( a8098a  and  a8091a );
 a2515a <=( a8084a  and  a8077a );
 a2516a <=( a8070a  and  a8063a );
 a2517a <=( a8056a  and  a8049a );
 a2518a <=( a8042a  and  a8035a );
 a2519a <=( a8028a  and  a8021a );
 a2520a <=( a8014a  and  a8007a );
 a2521a <=( a8000a  and  a7993a );
 a2522a <=( a7988a  and  a7981a );
 a2523a <=( a7976a  and  a7969a );
 a2524a <=( a7964a  and  a7957a );
 a2525a <=( a7952a  and  a7945a );
 a2526a <=( a7940a  and  a7933a );
 a2527a <=( a7928a  and  a7921a );
 a2528a <=( a7916a  and  a7909a );
 a2529a <=( a7904a  and  a7897a );
 a2530a <=( a7892a  and  a7885a );
 a2531a <=( a7880a  and  a7873a );
 a2532a <=( a7868a  and  a7861a );
 a2533a <=( a7856a  and  a7849a );
 a2534a <=( a7844a  and  a7837a );
 a2535a <=( a7832a  and  a7825a );
 a2536a <=( a7820a  and  a7813a );
 a2537a <=( a7808a  and  a7801a );
 a2538a <=( a7796a  and  a7789a );
 a2539a <=( a7784a  and  a7777a );
 a2540a <=( a7772a  and  a7765a );
 a2541a <=( a7760a  and  a7753a );
 a2542a <=( a7748a  and  a7741a );
 a2543a <=( a7736a  and  a7729a );
 a2544a <=( a7724a  and  a7717a );
 a2545a <=( a7712a  and  a7705a );
 a2546a <=( a7700a  and  a7693a );
 a2547a <=( a7688a  and  a7683a );
 a2548a <=( a7678a  and  a7673a );
 a2549a <=( a7668a  and  a7663a );
 a2550a <=( a7658a  and  a7653a );
 a2553a <=( a2549a ) or ( a2550a );
 a2556a <=( a2547a ) or ( a2548a );
 a2557a <=( a2556a ) or ( a2553a );
 a2560a <=( a2545a ) or ( a2546a );
 a2564a <=( a2542a ) or ( a2543a );
 a2565a <=( a2544a ) or ( a2564a );
 a2566a <=( a2565a ) or ( a2560a );
 a2567a <=( a2566a ) or ( a2557a );
 a2570a <=( a2540a ) or ( a2541a );
 a2574a <=( a2537a ) or ( a2538a );
 a2575a <=( a2539a ) or ( a2574a );
 a2576a <=( a2575a ) or ( a2570a );
 a2579a <=( a2535a ) or ( a2536a );
 a2583a <=( a2532a ) or ( a2533a );
 a2584a <=( a2534a ) or ( a2583a );
 a2585a <=( a2584a ) or ( a2579a );
 a2586a <=( a2585a ) or ( a2576a );
 a2587a <=( a2586a ) or ( a2567a );
 a2590a <=( a2530a ) or ( a2531a );
 a2594a <=( a2527a ) or ( a2528a );
 a2595a <=( a2529a ) or ( a2594a );
 a2596a <=( a2595a ) or ( a2590a );
 a2599a <=( a2525a ) or ( a2526a );
 a2603a <=( a2522a ) or ( a2523a );
 a2604a <=( a2524a ) or ( a2603a );
 a2605a <=( a2604a ) or ( a2599a );
 a2606a <=( a2605a ) or ( a2596a );
 a2609a <=( a2520a ) or ( a2521a );
 a2613a <=( a2517a ) or ( a2518a );
 a2614a <=( a2519a ) or ( a2613a );
 a2615a <=( a2614a ) or ( a2609a );
 a2618a <=( a2515a ) or ( a2516a );
 a2622a <=( a2512a ) or ( a2513a );
 a2623a <=( a2514a ) or ( a2622a );
 a2624a <=( a2623a ) or ( a2618a );
 a2625a <=( a2624a ) or ( a2615a );
 a2626a <=( a2625a ) or ( a2606a );
 a2627a <=( a2626a ) or ( a2587a );
 a2630a <=( a2510a ) or ( a2511a );
 a2634a <=( a2507a ) or ( a2508a );
 a2635a <=( a2509a ) or ( a2634a );
 a2636a <=( a2635a ) or ( a2630a );
 a2639a <=( a2505a ) or ( a2506a );
 a2643a <=( a2502a ) or ( a2503a );
 a2644a <=( a2504a ) or ( a2643a );
 a2645a <=( a2644a ) or ( a2639a );
 a2646a <=( a2645a ) or ( a2636a );
 a2649a <=( a2500a ) or ( a2501a );
 a2653a <=( a2497a ) or ( a2498a );
 a2654a <=( a2499a ) or ( a2653a );
 a2655a <=( a2654a ) or ( a2649a );
 a2658a <=( a2495a ) or ( a2496a );
 a2662a <=( a2492a ) or ( a2493a );
 a2663a <=( a2494a ) or ( a2662a );
 a2664a <=( a2663a ) or ( a2658a );
 a2665a <=( a2664a ) or ( a2655a );
 a2666a <=( a2665a ) or ( a2646a );
 a2669a <=( a2490a ) or ( a2491a );
 a2673a <=( a2487a ) or ( a2488a );
 a2674a <=( a2489a ) or ( a2673a );
 a2675a <=( a2674a ) or ( a2669a );
 a2678a <=( a2485a ) or ( a2486a );
 a2682a <=( a2482a ) or ( a2483a );
 a2683a <=( a2484a ) or ( a2682a );
 a2684a <=( a2683a ) or ( a2678a );
 a2685a <=( a2684a ) or ( a2675a );
 a2688a <=( a2480a ) or ( a2481a );
 a2692a <=( a2477a ) or ( a2478a );
 a2693a <=( a2479a ) or ( a2692a );
 a2694a <=( a2693a ) or ( a2688a );
 a2697a <=( a2475a ) or ( a2476a );
 a2701a <=( a2472a ) or ( a2473a );
 a2702a <=( a2474a ) or ( a2701a );
 a2703a <=( a2702a ) or ( a2697a );
 a2704a <=( a2703a ) or ( a2694a );
 a2705a <=( a2704a ) or ( a2685a );
 a2706a <=( a2705a ) or ( a2666a );
 a2707a <=( a2706a ) or ( a2627a );
 a2710a <=( a2470a ) or ( a2471a );
 a2714a <=( a2467a ) or ( a2468a );
 a2715a <=( a2469a ) or ( a2714a );
 a2716a <=( a2715a ) or ( a2710a );
 a2719a <=( a2465a ) or ( a2466a );
 a2723a <=( a2462a ) or ( a2463a );
 a2724a <=( a2464a ) or ( a2723a );
 a2725a <=( a2724a ) or ( a2719a );
 a2726a <=( a2725a ) or ( a2716a );
 a2729a <=( a2460a ) or ( a2461a );
 a2733a <=( a2457a ) or ( a2458a );
 a2734a <=( a2459a ) or ( a2733a );
 a2735a <=( a2734a ) or ( a2729a );
 a2738a <=( a2455a ) or ( a2456a );
 a2742a <=( a2452a ) or ( a2453a );
 a2743a <=( a2454a ) or ( a2742a );
 a2744a <=( a2743a ) or ( a2738a );
 a2745a <=( a2744a ) or ( a2735a );
 a2746a <=( a2745a ) or ( a2726a );
 a2749a <=( a2450a ) or ( a2451a );
 a2753a <=( a2447a ) or ( a2448a );
 a2754a <=( a2449a ) or ( a2753a );
 a2755a <=( a2754a ) or ( a2749a );
 a2758a <=( a2445a ) or ( a2446a );
 a2762a <=( a2442a ) or ( a2443a );
 a2763a <=( a2444a ) or ( a2762a );
 a2764a <=( a2763a ) or ( a2758a );
 a2765a <=( a2764a ) or ( a2755a );
 a2768a <=( a2440a ) or ( a2441a );
 a2772a <=( a2437a ) or ( a2438a );
 a2773a <=( a2439a ) or ( a2772a );
 a2774a <=( a2773a ) or ( a2768a );
 a2777a <=( a2435a ) or ( a2436a );
 a2781a <=( a2432a ) or ( a2433a );
 a2782a <=( a2434a ) or ( a2781a );
 a2783a <=( a2782a ) or ( a2777a );
 a2784a <=( a2783a ) or ( a2774a );
 a2785a <=( a2784a ) or ( a2765a );
 a2786a <=( a2785a ) or ( a2746a );
 a2789a <=( a2430a ) or ( a2431a );
 a2793a <=( a2427a ) or ( a2428a );
 a2794a <=( a2429a ) or ( a2793a );
 a2795a <=( a2794a ) or ( a2789a );
 a2798a <=( a2425a ) or ( a2426a );
 a2802a <=( a2422a ) or ( a2423a );
 a2803a <=( a2424a ) or ( a2802a );
 a2804a <=( a2803a ) or ( a2798a );
 a2805a <=( a2804a ) or ( a2795a );
 a2808a <=( a2420a ) or ( a2421a );
 a2812a <=( a2417a ) or ( a2418a );
 a2813a <=( a2419a ) or ( a2812a );
 a2814a <=( a2813a ) or ( a2808a );
 a2817a <=( a2415a ) or ( a2416a );
 a2821a <=( a2412a ) or ( a2413a );
 a2822a <=( a2414a ) or ( a2821a );
 a2823a <=( a2822a ) or ( a2817a );
 a2824a <=( a2823a ) or ( a2814a );
 a2825a <=( a2824a ) or ( a2805a );
 a2828a <=( a2410a ) or ( a2411a );
 a2832a <=( a2407a ) or ( a2408a );
 a2833a <=( a2409a ) or ( a2832a );
 a2834a <=( a2833a ) or ( a2828a );
 a2837a <=( a2405a ) or ( a2406a );
 a2841a <=( a2402a ) or ( a2403a );
 a2842a <=( a2404a ) or ( a2841a );
 a2843a <=( a2842a ) or ( a2837a );
 a2844a <=( a2843a ) or ( a2834a );
 a2847a <=( a2400a ) or ( a2401a );
 a2851a <=( a2397a ) or ( a2398a );
 a2852a <=( a2399a ) or ( a2851a );
 a2853a <=( a2852a ) or ( a2847a );
 a2856a <=( a2395a ) or ( a2396a );
 a2860a <=( a2392a ) or ( a2393a );
 a2861a <=( a2394a ) or ( a2860a );
 a2862a <=( a2861a ) or ( a2856a );
 a2863a <=( a2862a ) or ( a2853a );
 a2864a <=( a2863a ) or ( a2844a );
 a2865a <=( a2864a ) or ( a2825a );
 a2866a <=( a2865a ) or ( a2786a );
 a2867a <=( a2866a ) or ( a2707a );
 a2870a <=( a2390a ) or ( a2391a );
 a2873a <=( a2388a ) or ( a2389a );
 a2874a <=( a2873a ) or ( a2870a );
 a2877a <=( a2386a ) or ( a2387a );
 a2881a <=( a2383a ) or ( a2384a );
 a2882a <=( a2385a ) or ( a2881a );
 a2883a <=( a2882a ) or ( a2877a );
 a2884a <=( a2883a ) or ( a2874a );
 a2887a <=( a2381a ) or ( a2382a );
 a2891a <=( a2378a ) or ( a2379a );
 a2892a <=( a2380a ) or ( a2891a );
 a2893a <=( a2892a ) or ( a2887a );
 a2896a <=( a2376a ) or ( a2377a );
 a2900a <=( a2373a ) or ( a2374a );
 a2901a <=( a2375a ) or ( a2900a );
 a2902a <=( a2901a ) or ( a2896a );
 a2903a <=( a2902a ) or ( a2893a );
 a2904a <=( a2903a ) or ( a2884a );
 a2907a <=( a2371a ) or ( a2372a );
 a2911a <=( a2368a ) or ( a2369a );
 a2912a <=( a2370a ) or ( a2911a );
 a2913a <=( a2912a ) or ( a2907a );
 a2916a <=( a2366a ) or ( a2367a );
 a2920a <=( a2363a ) or ( a2364a );
 a2921a <=( a2365a ) or ( a2920a );
 a2922a <=( a2921a ) or ( a2916a );
 a2923a <=( a2922a ) or ( a2913a );
 a2926a <=( a2361a ) or ( a2362a );
 a2930a <=( a2358a ) or ( a2359a );
 a2931a <=( a2360a ) or ( a2930a );
 a2932a <=( a2931a ) or ( a2926a );
 a2935a <=( a2356a ) or ( a2357a );
 a2939a <=( a2353a ) or ( a2354a );
 a2940a <=( a2355a ) or ( a2939a );
 a2941a <=( a2940a ) or ( a2935a );
 a2942a <=( a2941a ) or ( a2932a );
 a2943a <=( a2942a ) or ( a2923a );
 a2944a <=( a2943a ) or ( a2904a );
 a2947a <=( a2351a ) or ( a2352a );
 a2951a <=( a2348a ) or ( a2349a );
 a2952a <=( a2350a ) or ( a2951a );
 a2953a <=( a2952a ) or ( a2947a );
 a2956a <=( a2346a ) or ( a2347a );
 a2960a <=( a2343a ) or ( a2344a );
 a2961a <=( a2345a ) or ( a2960a );
 a2962a <=( a2961a ) or ( a2956a );
 a2963a <=( a2962a ) or ( a2953a );
 a2966a <=( a2341a ) or ( a2342a );
 a2970a <=( a2338a ) or ( a2339a );
 a2971a <=( a2340a ) or ( a2970a );
 a2972a <=( a2971a ) or ( a2966a );
 a2975a <=( a2336a ) or ( a2337a );
 a2979a <=( a2333a ) or ( a2334a );
 a2980a <=( a2335a ) or ( a2979a );
 a2981a <=( a2980a ) or ( a2975a );
 a2982a <=( a2981a ) or ( a2972a );
 a2983a <=( a2982a ) or ( a2963a );
 a2986a <=( a2331a ) or ( a2332a );
 a2990a <=( a2328a ) or ( a2329a );
 a2991a <=( a2330a ) or ( a2990a );
 a2992a <=( a2991a ) or ( a2986a );
 a2995a <=( a2326a ) or ( a2327a );
 a2999a <=( a2323a ) or ( a2324a );
 a3000a <=( a2325a ) or ( a2999a );
 a3001a <=( a3000a ) or ( a2995a );
 a3002a <=( a3001a ) or ( a2992a );
 a3005a <=( a2321a ) or ( a2322a );
 a3009a <=( a2318a ) or ( a2319a );
 a3010a <=( a2320a ) or ( a3009a );
 a3011a <=( a3010a ) or ( a3005a );
 a3014a <=( a2316a ) or ( a2317a );
 a3018a <=( a2313a ) or ( a2314a );
 a3019a <=( a2315a ) or ( a3018a );
 a3020a <=( a3019a ) or ( a3014a );
 a3021a <=( a3020a ) or ( a3011a );
 a3022a <=( a3021a ) or ( a3002a );
 a3023a <=( a3022a ) or ( a2983a );
 a3024a <=( a3023a ) or ( a2944a );
 a3027a <=( a2311a ) or ( a2312a );
 a3031a <=( a2308a ) or ( a2309a );
 a3032a <=( a2310a ) or ( a3031a );
 a3033a <=( a3032a ) or ( a3027a );
 a3036a <=( a2306a ) or ( a2307a );
 a3040a <=( a2303a ) or ( a2304a );
 a3041a <=( a2305a ) or ( a3040a );
 a3042a <=( a3041a ) or ( a3036a );
 a3043a <=( a3042a ) or ( a3033a );
 a3046a <=( a2301a ) or ( a2302a );
 a3050a <=( a2298a ) or ( a2299a );
 a3051a <=( a2300a ) or ( a3050a );
 a3052a <=( a3051a ) or ( a3046a );
 a3055a <=( a2296a ) or ( a2297a );
 a3059a <=( a2293a ) or ( a2294a );
 a3060a <=( a2295a ) or ( a3059a );
 a3061a <=( a3060a ) or ( a3055a );
 a3062a <=( a3061a ) or ( a3052a );
 a3063a <=( a3062a ) or ( a3043a );
 a3066a <=( a2291a ) or ( a2292a );
 a3070a <=( a2288a ) or ( a2289a );
 a3071a <=( a2290a ) or ( a3070a );
 a3072a <=( a3071a ) or ( a3066a );
 a3075a <=( a2286a ) or ( a2287a );
 a3079a <=( a2283a ) or ( a2284a );
 a3080a <=( a2285a ) or ( a3079a );
 a3081a <=( a3080a ) or ( a3075a );
 a3082a <=( a3081a ) or ( a3072a );
 a3085a <=( a2281a ) or ( a2282a );
 a3089a <=( a2278a ) or ( a2279a );
 a3090a <=( a2280a ) or ( a3089a );
 a3091a <=( a3090a ) or ( a3085a );
 a3094a <=( a2276a ) or ( a2277a );
 a3098a <=( a2273a ) or ( a2274a );
 a3099a <=( a2275a ) or ( a3098a );
 a3100a <=( a3099a ) or ( a3094a );
 a3101a <=( a3100a ) or ( a3091a );
 a3102a <=( a3101a ) or ( a3082a );
 a3103a <=( a3102a ) or ( a3063a );
 a3106a <=( a2271a ) or ( a2272a );
 a3110a <=( a2268a ) or ( a2269a );
 a3111a <=( a2270a ) or ( a3110a );
 a3112a <=( a3111a ) or ( a3106a );
 a3115a <=( a2266a ) or ( a2267a );
 a3119a <=( a2263a ) or ( a2264a );
 a3120a <=( a2265a ) or ( a3119a );
 a3121a <=( a3120a ) or ( a3115a );
 a3122a <=( a3121a ) or ( a3112a );
 a3125a <=( a2261a ) or ( a2262a );
 a3129a <=( a2258a ) or ( a2259a );
 a3130a <=( a2260a ) or ( a3129a );
 a3131a <=( a3130a ) or ( a3125a );
 a3134a <=( a2256a ) or ( a2257a );
 a3138a <=( a2253a ) or ( a2254a );
 a3139a <=( a2255a ) or ( a3138a );
 a3140a <=( a3139a ) or ( a3134a );
 a3141a <=( a3140a ) or ( a3131a );
 a3142a <=( a3141a ) or ( a3122a );
 a3145a <=( a2251a ) or ( a2252a );
 a3149a <=( a2248a ) or ( a2249a );
 a3150a <=( a2250a ) or ( a3149a );
 a3151a <=( a3150a ) or ( a3145a );
 a3154a <=( a2246a ) or ( a2247a );
 a3158a <=( a2243a ) or ( a2244a );
 a3159a <=( a2245a ) or ( a3158a );
 a3160a <=( a3159a ) or ( a3154a );
 a3161a <=( a3160a ) or ( a3151a );
 a3164a <=( a2241a ) or ( a2242a );
 a3168a <=( a2238a ) or ( a2239a );
 a3169a <=( a2240a ) or ( a3168a );
 a3170a <=( a3169a ) or ( a3164a );
 a3173a <=( a2236a ) or ( a2237a );
 a3177a <=( a2233a ) or ( a2234a );
 a3178a <=( a2235a ) or ( a3177a );
 a3179a <=( a3178a ) or ( a3173a );
 a3180a <=( a3179a ) or ( a3170a );
 a3181a <=( a3180a ) or ( a3161a );
 a3182a <=( a3181a ) or ( a3142a );
 a3183a <=( a3182a ) or ( a3103a );
 a3184a <=( a3183a ) or ( a3024a );
 a3185a <=( a3184a ) or ( a2867a );
 a3188a <=( a2231a ) or ( a2232a );
 a3191a <=( a2229a ) or ( a2230a );
 a3192a <=( a3191a ) or ( a3188a );
 a3195a <=( a2227a ) or ( a2228a );
 a3199a <=( a2224a ) or ( a2225a );
 a3200a <=( a2226a ) or ( a3199a );
 a3201a <=( a3200a ) or ( a3195a );
 a3202a <=( a3201a ) or ( a3192a );
 a3205a <=( a2222a ) or ( a2223a );
 a3209a <=( a2219a ) or ( a2220a );
 a3210a <=( a2221a ) or ( a3209a );
 a3211a <=( a3210a ) or ( a3205a );
 a3214a <=( a2217a ) or ( a2218a );
 a3218a <=( a2214a ) or ( a2215a );
 a3219a <=( a2216a ) or ( a3218a );
 a3220a <=( a3219a ) or ( a3214a );
 a3221a <=( a3220a ) or ( a3211a );
 a3222a <=( a3221a ) or ( a3202a );
 a3225a <=( a2212a ) or ( a2213a );
 a3229a <=( a2209a ) or ( a2210a );
 a3230a <=( a2211a ) or ( a3229a );
 a3231a <=( a3230a ) or ( a3225a );
 a3234a <=( a2207a ) or ( a2208a );
 a3238a <=( a2204a ) or ( a2205a );
 a3239a <=( a2206a ) or ( a3238a );
 a3240a <=( a3239a ) or ( a3234a );
 a3241a <=( a3240a ) or ( a3231a );
 a3244a <=( a2202a ) or ( a2203a );
 a3248a <=( a2199a ) or ( a2200a );
 a3249a <=( a2201a ) or ( a3248a );
 a3250a <=( a3249a ) or ( a3244a );
 a3253a <=( a2197a ) or ( a2198a );
 a3257a <=( a2194a ) or ( a2195a );
 a3258a <=( a2196a ) or ( a3257a );
 a3259a <=( a3258a ) or ( a3253a );
 a3260a <=( a3259a ) or ( a3250a );
 a3261a <=( a3260a ) or ( a3241a );
 a3262a <=( a3261a ) or ( a3222a );
 a3265a <=( a2192a ) or ( a2193a );
 a3269a <=( a2189a ) or ( a2190a );
 a3270a <=( a2191a ) or ( a3269a );
 a3271a <=( a3270a ) or ( a3265a );
 a3274a <=( a2187a ) or ( a2188a );
 a3278a <=( a2184a ) or ( a2185a );
 a3279a <=( a2186a ) or ( a3278a );
 a3280a <=( a3279a ) or ( a3274a );
 a3281a <=( a3280a ) or ( a3271a );
 a3284a <=( a2182a ) or ( a2183a );
 a3288a <=( a2179a ) or ( a2180a );
 a3289a <=( a2181a ) or ( a3288a );
 a3290a <=( a3289a ) or ( a3284a );
 a3293a <=( a2177a ) or ( a2178a );
 a3297a <=( a2174a ) or ( a2175a );
 a3298a <=( a2176a ) or ( a3297a );
 a3299a <=( a3298a ) or ( a3293a );
 a3300a <=( a3299a ) or ( a3290a );
 a3301a <=( a3300a ) or ( a3281a );
 a3304a <=( a2172a ) or ( a2173a );
 a3308a <=( a2169a ) or ( a2170a );
 a3309a <=( a2171a ) or ( a3308a );
 a3310a <=( a3309a ) or ( a3304a );
 a3313a <=( a2167a ) or ( a2168a );
 a3317a <=( a2164a ) or ( a2165a );
 a3318a <=( a2166a ) or ( a3317a );
 a3319a <=( a3318a ) or ( a3313a );
 a3320a <=( a3319a ) or ( a3310a );
 a3323a <=( a2162a ) or ( a2163a );
 a3327a <=( a2159a ) or ( a2160a );
 a3328a <=( a2161a ) or ( a3327a );
 a3329a <=( a3328a ) or ( a3323a );
 a3332a <=( a2157a ) or ( a2158a );
 a3336a <=( a2154a ) or ( a2155a );
 a3337a <=( a2156a ) or ( a3336a );
 a3338a <=( a3337a ) or ( a3332a );
 a3339a <=( a3338a ) or ( a3329a );
 a3340a <=( a3339a ) or ( a3320a );
 a3341a <=( a3340a ) or ( a3301a );
 a3342a <=( a3341a ) or ( a3262a );
 a3345a <=( a2152a ) or ( a2153a );
 a3349a <=( a2149a ) or ( a2150a );
 a3350a <=( a2151a ) or ( a3349a );
 a3351a <=( a3350a ) or ( a3345a );
 a3354a <=( a2147a ) or ( a2148a );
 a3358a <=( a2144a ) or ( a2145a );
 a3359a <=( a2146a ) or ( a3358a );
 a3360a <=( a3359a ) or ( a3354a );
 a3361a <=( a3360a ) or ( a3351a );
 a3364a <=( a2142a ) or ( a2143a );
 a3368a <=( a2139a ) or ( a2140a );
 a3369a <=( a2141a ) or ( a3368a );
 a3370a <=( a3369a ) or ( a3364a );
 a3373a <=( a2137a ) or ( a2138a );
 a3377a <=( a2134a ) or ( a2135a );
 a3378a <=( a2136a ) or ( a3377a );
 a3379a <=( a3378a ) or ( a3373a );
 a3380a <=( a3379a ) or ( a3370a );
 a3381a <=( a3380a ) or ( a3361a );
 a3384a <=( a2132a ) or ( a2133a );
 a3388a <=( a2129a ) or ( a2130a );
 a3389a <=( a2131a ) or ( a3388a );
 a3390a <=( a3389a ) or ( a3384a );
 a3393a <=( a2127a ) or ( a2128a );
 a3397a <=( a2124a ) or ( a2125a );
 a3398a <=( a2126a ) or ( a3397a );
 a3399a <=( a3398a ) or ( a3393a );
 a3400a <=( a3399a ) or ( a3390a );
 a3403a <=( a2122a ) or ( a2123a );
 a3407a <=( a2119a ) or ( a2120a );
 a3408a <=( a2121a ) or ( a3407a );
 a3409a <=( a3408a ) or ( a3403a );
 a3412a <=( a2117a ) or ( a2118a );
 a3416a <=( a2114a ) or ( a2115a );
 a3417a <=( a2116a ) or ( a3416a );
 a3418a <=( a3417a ) or ( a3412a );
 a3419a <=( a3418a ) or ( a3409a );
 a3420a <=( a3419a ) or ( a3400a );
 a3421a <=( a3420a ) or ( a3381a );
 a3424a <=( a2112a ) or ( a2113a );
 a3428a <=( a2109a ) or ( a2110a );
 a3429a <=( a2111a ) or ( a3428a );
 a3430a <=( a3429a ) or ( a3424a );
 a3433a <=( a2107a ) or ( a2108a );
 a3437a <=( a2104a ) or ( a2105a );
 a3438a <=( a2106a ) or ( a3437a );
 a3439a <=( a3438a ) or ( a3433a );
 a3440a <=( a3439a ) or ( a3430a );
 a3443a <=( a2102a ) or ( a2103a );
 a3447a <=( a2099a ) or ( a2100a );
 a3448a <=( a2101a ) or ( a3447a );
 a3449a <=( a3448a ) or ( a3443a );
 a3452a <=( a2097a ) or ( a2098a );
 a3456a <=( a2094a ) or ( a2095a );
 a3457a <=( a2096a ) or ( a3456a );
 a3458a <=( a3457a ) or ( a3452a );
 a3459a <=( a3458a ) or ( a3449a );
 a3460a <=( a3459a ) or ( a3440a );
 a3463a <=( a2092a ) or ( a2093a );
 a3467a <=( a2089a ) or ( a2090a );
 a3468a <=( a2091a ) or ( a3467a );
 a3469a <=( a3468a ) or ( a3463a );
 a3472a <=( a2087a ) or ( a2088a );
 a3476a <=( a2084a ) or ( a2085a );
 a3477a <=( a2086a ) or ( a3476a );
 a3478a <=( a3477a ) or ( a3472a );
 a3479a <=( a3478a ) or ( a3469a );
 a3482a <=( a2082a ) or ( a2083a );
 a3486a <=( a2079a ) or ( a2080a );
 a3487a <=( a2081a ) or ( a3486a );
 a3488a <=( a3487a ) or ( a3482a );
 a3491a <=( a2077a ) or ( a2078a );
 a3495a <=( a2074a ) or ( a2075a );
 a3496a <=( a2076a ) or ( a3495a );
 a3497a <=( a3496a ) or ( a3491a );
 a3498a <=( a3497a ) or ( a3488a );
 a3499a <=( a3498a ) or ( a3479a );
 a3500a <=( a3499a ) or ( a3460a );
 a3501a <=( a3500a ) or ( a3421a );
 a3502a <=( a3501a ) or ( a3342a );
 a3505a <=( a2072a ) or ( a2073a );
 a3509a <=( a2069a ) or ( a2070a );
 a3510a <=( a2071a ) or ( a3509a );
 a3511a <=( a3510a ) or ( a3505a );
 a3514a <=( a2067a ) or ( a2068a );
 a3518a <=( a2064a ) or ( a2065a );
 a3519a <=( a2066a ) or ( a3518a );
 a3520a <=( a3519a ) or ( a3514a );
 a3521a <=( a3520a ) or ( a3511a );
 a3524a <=( a2062a ) or ( a2063a );
 a3528a <=( a2059a ) or ( a2060a );
 a3529a <=( a2061a ) or ( a3528a );
 a3530a <=( a3529a ) or ( a3524a );
 a3533a <=( a2057a ) or ( a2058a );
 a3537a <=( a2054a ) or ( a2055a );
 a3538a <=( a2056a ) or ( a3537a );
 a3539a <=( a3538a ) or ( a3533a );
 a3540a <=( a3539a ) or ( a3530a );
 a3541a <=( a3540a ) or ( a3521a );
 a3544a <=( a2052a ) or ( a2053a );
 a3548a <=( a2049a ) or ( a2050a );
 a3549a <=( a2051a ) or ( a3548a );
 a3550a <=( a3549a ) or ( a3544a );
 a3553a <=( a2047a ) or ( a2048a );
 a3557a <=( a2044a ) or ( a2045a );
 a3558a <=( a2046a ) or ( a3557a );
 a3559a <=( a3558a ) or ( a3553a );
 a3560a <=( a3559a ) or ( a3550a );
 a3563a <=( a2042a ) or ( a2043a );
 a3567a <=( a2039a ) or ( a2040a );
 a3568a <=( a2041a ) or ( a3567a );
 a3569a <=( a3568a ) or ( a3563a );
 a3572a <=( a2037a ) or ( a2038a );
 a3576a <=( a2034a ) or ( a2035a );
 a3577a <=( a2036a ) or ( a3576a );
 a3578a <=( a3577a ) or ( a3572a );
 a3579a <=( a3578a ) or ( a3569a );
 a3580a <=( a3579a ) or ( a3560a );
 a3581a <=( a3580a ) or ( a3541a );
 a3584a <=( a2032a ) or ( a2033a );
 a3588a <=( a2029a ) or ( a2030a );
 a3589a <=( a2031a ) or ( a3588a );
 a3590a <=( a3589a ) or ( a3584a );
 a3593a <=( a2027a ) or ( a2028a );
 a3597a <=( a2024a ) or ( a2025a );
 a3598a <=( a2026a ) or ( a3597a );
 a3599a <=( a3598a ) or ( a3593a );
 a3600a <=( a3599a ) or ( a3590a );
 a3603a <=( a2022a ) or ( a2023a );
 a3607a <=( a2019a ) or ( a2020a );
 a3608a <=( a2021a ) or ( a3607a );
 a3609a <=( a3608a ) or ( a3603a );
 a3612a <=( a2017a ) or ( a2018a );
 a3616a <=( a2014a ) or ( a2015a );
 a3617a <=( a2016a ) or ( a3616a );
 a3618a <=( a3617a ) or ( a3612a );
 a3619a <=( a3618a ) or ( a3609a );
 a3620a <=( a3619a ) or ( a3600a );
 a3623a <=( a2012a ) or ( a2013a );
 a3627a <=( a2009a ) or ( a2010a );
 a3628a <=( a2011a ) or ( a3627a );
 a3629a <=( a3628a ) or ( a3623a );
 a3632a <=( a2007a ) or ( a2008a );
 a3636a <=( a2004a ) or ( a2005a );
 a3637a <=( a2006a ) or ( a3636a );
 a3638a <=( a3637a ) or ( a3632a );
 a3639a <=( a3638a ) or ( a3629a );
 a3642a <=( a2002a ) or ( a2003a );
 a3646a <=( a1999a ) or ( a2000a );
 a3647a <=( a2001a ) or ( a3646a );
 a3648a <=( a3647a ) or ( a3642a );
 a3651a <=( a1997a ) or ( a1998a );
 a3655a <=( a1994a ) or ( a1995a );
 a3656a <=( a1996a ) or ( a3655a );
 a3657a <=( a3656a ) or ( a3651a );
 a3658a <=( a3657a ) or ( a3648a );
 a3659a <=( a3658a ) or ( a3639a );
 a3660a <=( a3659a ) or ( a3620a );
 a3661a <=( a3660a ) or ( a3581a );
 a3664a <=( a1992a ) or ( a1993a );
 a3668a <=( a1989a ) or ( a1990a );
 a3669a <=( a1991a ) or ( a3668a );
 a3670a <=( a3669a ) or ( a3664a );
 a3673a <=( a1987a ) or ( a1988a );
 a3677a <=( a1984a ) or ( a1985a );
 a3678a <=( a1986a ) or ( a3677a );
 a3679a <=( a3678a ) or ( a3673a );
 a3680a <=( a3679a ) or ( a3670a );
 a3683a <=( a1982a ) or ( a1983a );
 a3687a <=( a1979a ) or ( a1980a );
 a3688a <=( a1981a ) or ( a3687a );
 a3689a <=( a3688a ) or ( a3683a );
 a3692a <=( a1977a ) or ( a1978a );
 a3696a <=( a1974a ) or ( a1975a );
 a3697a <=( a1976a ) or ( a3696a );
 a3698a <=( a3697a ) or ( a3692a );
 a3699a <=( a3698a ) or ( a3689a );
 a3700a <=( a3699a ) or ( a3680a );
 a3703a <=( a1972a ) or ( a1973a );
 a3707a <=( a1969a ) or ( a1970a );
 a3708a <=( a1971a ) or ( a3707a );
 a3709a <=( a3708a ) or ( a3703a );
 a3712a <=( a1967a ) or ( a1968a );
 a3716a <=( a1964a ) or ( a1965a );
 a3717a <=( a1966a ) or ( a3716a );
 a3718a <=( a3717a ) or ( a3712a );
 a3719a <=( a3718a ) or ( a3709a );
 a3722a <=( a1962a ) or ( a1963a );
 a3726a <=( a1959a ) or ( a1960a );
 a3727a <=( a1961a ) or ( a3726a );
 a3728a <=( a3727a ) or ( a3722a );
 a3731a <=( a1957a ) or ( a1958a );
 a3735a <=( a1954a ) or ( a1955a );
 a3736a <=( a1956a ) or ( a3735a );
 a3737a <=( a3736a ) or ( a3731a );
 a3738a <=( a3737a ) or ( a3728a );
 a3739a <=( a3738a ) or ( a3719a );
 a3740a <=( a3739a ) or ( a3700a );
 a3743a <=( a1952a ) or ( a1953a );
 a3747a <=( a1949a ) or ( a1950a );
 a3748a <=( a1951a ) or ( a3747a );
 a3749a <=( a3748a ) or ( a3743a );
 a3752a <=( a1947a ) or ( a1948a );
 a3756a <=( a1944a ) or ( a1945a );
 a3757a <=( a1946a ) or ( a3756a );
 a3758a <=( a3757a ) or ( a3752a );
 a3759a <=( a3758a ) or ( a3749a );
 a3762a <=( a1942a ) or ( a1943a );
 a3766a <=( a1939a ) or ( a1940a );
 a3767a <=( a1941a ) or ( a3766a );
 a3768a <=( a3767a ) or ( a3762a );
 a3771a <=( a1937a ) or ( a1938a );
 a3775a <=( a1934a ) or ( a1935a );
 a3776a <=( a1936a ) or ( a3775a );
 a3777a <=( a3776a ) or ( a3771a );
 a3778a <=( a3777a ) or ( a3768a );
 a3779a <=( a3778a ) or ( a3759a );
 a3782a <=( a1932a ) or ( a1933a );
 a3786a <=( a1929a ) or ( a1930a );
 a3787a <=( a1931a ) or ( a3786a );
 a3788a <=( a3787a ) or ( a3782a );
 a3791a <=( a1927a ) or ( a1928a );
 a3795a <=( a1924a ) or ( a1925a );
 a3796a <=( a1926a ) or ( a3795a );
 a3797a <=( a3796a ) or ( a3791a );
 a3798a <=( a3797a ) or ( a3788a );
 a3801a <=( a1922a ) or ( a1923a );
 a3805a <=( a1919a ) or ( a1920a );
 a3806a <=( a1921a ) or ( a3805a );
 a3807a <=( a3806a ) or ( a3801a );
 a3810a <=( a1917a ) or ( a1918a );
 a3814a <=( a1914a ) or ( a1915a );
 a3815a <=( a1916a ) or ( a3814a );
 a3816a <=( a3815a ) or ( a3810a );
 a3817a <=( a3816a ) or ( a3807a );
 a3818a <=( a3817a ) or ( a3798a );
 a3819a <=( a3818a ) or ( a3779a );
 a3820a <=( a3819a ) or ( a3740a );
 a3821a <=( a3820a ) or ( a3661a );
 a3822a <=( a3821a ) or ( a3502a );
 a3823a <=( a3822a ) or ( a3185a );
 a3826a <=( a1912a ) or ( a1913a );
 a3829a <=( a1910a ) or ( a1911a );
 a3830a <=( a3829a ) or ( a3826a );
 a3833a <=( a1908a ) or ( a1909a );
 a3837a <=( a1905a ) or ( a1906a );
 a3838a <=( a1907a ) or ( a3837a );
 a3839a <=( a3838a ) or ( a3833a );
 a3840a <=( a3839a ) or ( a3830a );
 a3843a <=( a1903a ) or ( a1904a );
 a3847a <=( a1900a ) or ( a1901a );
 a3848a <=( a1902a ) or ( a3847a );
 a3849a <=( a3848a ) or ( a3843a );
 a3852a <=( a1898a ) or ( a1899a );
 a3856a <=( a1895a ) or ( a1896a );
 a3857a <=( a1897a ) or ( a3856a );
 a3858a <=( a3857a ) or ( a3852a );
 a3859a <=( a3858a ) or ( a3849a );
 a3860a <=( a3859a ) or ( a3840a );
 a3863a <=( a1893a ) or ( a1894a );
 a3867a <=( a1890a ) or ( a1891a );
 a3868a <=( a1892a ) or ( a3867a );
 a3869a <=( a3868a ) or ( a3863a );
 a3872a <=( a1888a ) or ( a1889a );
 a3876a <=( a1885a ) or ( a1886a );
 a3877a <=( a1887a ) or ( a3876a );
 a3878a <=( a3877a ) or ( a3872a );
 a3879a <=( a3878a ) or ( a3869a );
 a3882a <=( a1883a ) or ( a1884a );
 a3886a <=( a1880a ) or ( a1881a );
 a3887a <=( a1882a ) or ( a3886a );
 a3888a <=( a3887a ) or ( a3882a );
 a3891a <=( a1878a ) or ( a1879a );
 a3895a <=( a1875a ) or ( a1876a );
 a3896a <=( a1877a ) or ( a3895a );
 a3897a <=( a3896a ) or ( a3891a );
 a3898a <=( a3897a ) or ( a3888a );
 a3899a <=( a3898a ) or ( a3879a );
 a3900a <=( a3899a ) or ( a3860a );
 a3903a <=( a1873a ) or ( a1874a );
 a3907a <=( a1870a ) or ( a1871a );
 a3908a <=( a1872a ) or ( a3907a );
 a3909a <=( a3908a ) or ( a3903a );
 a3912a <=( a1868a ) or ( a1869a );
 a3916a <=( a1865a ) or ( a1866a );
 a3917a <=( a1867a ) or ( a3916a );
 a3918a <=( a3917a ) or ( a3912a );
 a3919a <=( a3918a ) or ( a3909a );
 a3922a <=( a1863a ) or ( a1864a );
 a3926a <=( a1860a ) or ( a1861a );
 a3927a <=( a1862a ) or ( a3926a );
 a3928a <=( a3927a ) or ( a3922a );
 a3931a <=( a1858a ) or ( a1859a );
 a3935a <=( a1855a ) or ( a1856a );
 a3936a <=( a1857a ) or ( a3935a );
 a3937a <=( a3936a ) or ( a3931a );
 a3938a <=( a3937a ) or ( a3928a );
 a3939a <=( a3938a ) or ( a3919a );
 a3942a <=( a1853a ) or ( a1854a );
 a3946a <=( a1850a ) or ( a1851a );
 a3947a <=( a1852a ) or ( a3946a );
 a3948a <=( a3947a ) or ( a3942a );
 a3951a <=( a1848a ) or ( a1849a );
 a3955a <=( a1845a ) or ( a1846a );
 a3956a <=( a1847a ) or ( a3955a );
 a3957a <=( a3956a ) or ( a3951a );
 a3958a <=( a3957a ) or ( a3948a );
 a3961a <=( a1843a ) or ( a1844a );
 a3965a <=( a1840a ) or ( a1841a );
 a3966a <=( a1842a ) or ( a3965a );
 a3967a <=( a3966a ) or ( a3961a );
 a3970a <=( a1838a ) or ( a1839a );
 a3974a <=( a1835a ) or ( a1836a );
 a3975a <=( a1837a ) or ( a3974a );
 a3976a <=( a3975a ) or ( a3970a );
 a3977a <=( a3976a ) or ( a3967a );
 a3978a <=( a3977a ) or ( a3958a );
 a3979a <=( a3978a ) or ( a3939a );
 a3980a <=( a3979a ) or ( a3900a );
 a3983a <=( a1833a ) or ( a1834a );
 a3987a <=( a1830a ) or ( a1831a );
 a3988a <=( a1832a ) or ( a3987a );
 a3989a <=( a3988a ) or ( a3983a );
 a3992a <=( a1828a ) or ( a1829a );
 a3996a <=( a1825a ) or ( a1826a );
 a3997a <=( a1827a ) or ( a3996a );
 a3998a <=( a3997a ) or ( a3992a );
 a3999a <=( a3998a ) or ( a3989a );
 a4002a <=( a1823a ) or ( a1824a );
 a4006a <=( a1820a ) or ( a1821a );
 a4007a <=( a1822a ) or ( a4006a );
 a4008a <=( a4007a ) or ( a4002a );
 a4011a <=( a1818a ) or ( a1819a );
 a4015a <=( a1815a ) or ( a1816a );
 a4016a <=( a1817a ) or ( a4015a );
 a4017a <=( a4016a ) or ( a4011a );
 a4018a <=( a4017a ) or ( a4008a );
 a4019a <=( a4018a ) or ( a3999a );
 a4022a <=( a1813a ) or ( a1814a );
 a4026a <=( a1810a ) or ( a1811a );
 a4027a <=( a1812a ) or ( a4026a );
 a4028a <=( a4027a ) or ( a4022a );
 a4031a <=( a1808a ) or ( a1809a );
 a4035a <=( a1805a ) or ( a1806a );
 a4036a <=( a1807a ) or ( a4035a );
 a4037a <=( a4036a ) or ( a4031a );
 a4038a <=( a4037a ) or ( a4028a );
 a4041a <=( a1803a ) or ( a1804a );
 a4045a <=( a1800a ) or ( a1801a );
 a4046a <=( a1802a ) or ( a4045a );
 a4047a <=( a4046a ) or ( a4041a );
 a4050a <=( a1798a ) or ( a1799a );
 a4054a <=( a1795a ) or ( a1796a );
 a4055a <=( a1797a ) or ( a4054a );
 a4056a <=( a4055a ) or ( a4050a );
 a4057a <=( a4056a ) or ( a4047a );
 a4058a <=( a4057a ) or ( a4038a );
 a4059a <=( a4058a ) or ( a4019a );
 a4062a <=( a1793a ) or ( a1794a );
 a4066a <=( a1790a ) or ( a1791a );
 a4067a <=( a1792a ) or ( a4066a );
 a4068a <=( a4067a ) or ( a4062a );
 a4071a <=( a1788a ) or ( a1789a );
 a4075a <=( a1785a ) or ( a1786a );
 a4076a <=( a1787a ) or ( a4075a );
 a4077a <=( a4076a ) or ( a4071a );
 a4078a <=( a4077a ) or ( a4068a );
 a4081a <=( a1783a ) or ( a1784a );
 a4085a <=( a1780a ) or ( a1781a );
 a4086a <=( a1782a ) or ( a4085a );
 a4087a <=( a4086a ) or ( a4081a );
 a4090a <=( a1778a ) or ( a1779a );
 a4094a <=( a1775a ) or ( a1776a );
 a4095a <=( a1777a ) or ( a4094a );
 a4096a <=( a4095a ) or ( a4090a );
 a4097a <=( a4096a ) or ( a4087a );
 a4098a <=( a4097a ) or ( a4078a );
 a4101a <=( a1773a ) or ( a1774a );
 a4105a <=( a1770a ) or ( a1771a );
 a4106a <=( a1772a ) or ( a4105a );
 a4107a <=( a4106a ) or ( a4101a );
 a4110a <=( a1768a ) or ( a1769a );
 a4114a <=( a1765a ) or ( a1766a );
 a4115a <=( a1767a ) or ( a4114a );
 a4116a <=( a4115a ) or ( a4110a );
 a4117a <=( a4116a ) or ( a4107a );
 a4120a <=( a1763a ) or ( a1764a );
 a4124a <=( a1760a ) or ( a1761a );
 a4125a <=( a1762a ) or ( a4124a );
 a4126a <=( a4125a ) or ( a4120a );
 a4129a <=( a1758a ) or ( a1759a );
 a4133a <=( a1755a ) or ( a1756a );
 a4134a <=( a1757a ) or ( a4133a );
 a4135a <=( a4134a ) or ( a4129a );
 a4136a <=( a4135a ) or ( a4126a );
 a4137a <=( a4136a ) or ( a4117a );
 a4138a <=( a4137a ) or ( a4098a );
 a4139a <=( a4138a ) or ( a4059a );
 a4140a <=( a4139a ) or ( a3980a );
 a4143a <=( a1753a ) or ( a1754a );
 a4147a <=( a1750a ) or ( a1751a );
 a4148a <=( a1752a ) or ( a4147a );
 a4149a <=( a4148a ) or ( a4143a );
 a4152a <=( a1748a ) or ( a1749a );
 a4156a <=( a1745a ) or ( a1746a );
 a4157a <=( a1747a ) or ( a4156a );
 a4158a <=( a4157a ) or ( a4152a );
 a4159a <=( a4158a ) or ( a4149a );
 a4162a <=( a1743a ) or ( a1744a );
 a4166a <=( a1740a ) or ( a1741a );
 a4167a <=( a1742a ) or ( a4166a );
 a4168a <=( a4167a ) or ( a4162a );
 a4171a <=( a1738a ) or ( a1739a );
 a4175a <=( a1735a ) or ( a1736a );
 a4176a <=( a1737a ) or ( a4175a );
 a4177a <=( a4176a ) or ( a4171a );
 a4178a <=( a4177a ) or ( a4168a );
 a4179a <=( a4178a ) or ( a4159a );
 a4182a <=( a1733a ) or ( a1734a );
 a4186a <=( a1730a ) or ( a1731a );
 a4187a <=( a1732a ) or ( a4186a );
 a4188a <=( a4187a ) or ( a4182a );
 a4191a <=( a1728a ) or ( a1729a );
 a4195a <=( a1725a ) or ( a1726a );
 a4196a <=( a1727a ) or ( a4195a );
 a4197a <=( a4196a ) or ( a4191a );
 a4198a <=( a4197a ) or ( a4188a );
 a4201a <=( a1723a ) or ( a1724a );
 a4205a <=( a1720a ) or ( a1721a );
 a4206a <=( a1722a ) or ( a4205a );
 a4207a <=( a4206a ) or ( a4201a );
 a4210a <=( a1718a ) or ( a1719a );
 a4214a <=( a1715a ) or ( a1716a );
 a4215a <=( a1717a ) or ( a4214a );
 a4216a <=( a4215a ) or ( a4210a );
 a4217a <=( a4216a ) or ( a4207a );
 a4218a <=( a4217a ) or ( a4198a );
 a4219a <=( a4218a ) or ( a4179a );
 a4222a <=( a1713a ) or ( a1714a );
 a4226a <=( a1710a ) or ( a1711a );
 a4227a <=( a1712a ) or ( a4226a );
 a4228a <=( a4227a ) or ( a4222a );
 a4231a <=( a1708a ) or ( a1709a );
 a4235a <=( a1705a ) or ( a1706a );
 a4236a <=( a1707a ) or ( a4235a );
 a4237a <=( a4236a ) or ( a4231a );
 a4238a <=( a4237a ) or ( a4228a );
 a4241a <=( a1703a ) or ( a1704a );
 a4245a <=( a1700a ) or ( a1701a );
 a4246a <=( a1702a ) or ( a4245a );
 a4247a <=( a4246a ) or ( a4241a );
 a4250a <=( a1698a ) or ( a1699a );
 a4254a <=( a1695a ) or ( a1696a );
 a4255a <=( a1697a ) or ( a4254a );
 a4256a <=( a4255a ) or ( a4250a );
 a4257a <=( a4256a ) or ( a4247a );
 a4258a <=( a4257a ) or ( a4238a );
 a4261a <=( a1693a ) or ( a1694a );
 a4265a <=( a1690a ) or ( a1691a );
 a4266a <=( a1692a ) or ( a4265a );
 a4267a <=( a4266a ) or ( a4261a );
 a4270a <=( a1688a ) or ( a1689a );
 a4274a <=( a1685a ) or ( a1686a );
 a4275a <=( a1687a ) or ( a4274a );
 a4276a <=( a4275a ) or ( a4270a );
 a4277a <=( a4276a ) or ( a4267a );
 a4280a <=( a1683a ) or ( a1684a );
 a4284a <=( a1680a ) or ( a1681a );
 a4285a <=( a1682a ) or ( a4284a );
 a4286a <=( a4285a ) or ( a4280a );
 a4289a <=( a1678a ) or ( a1679a );
 a4293a <=( a1675a ) or ( a1676a );
 a4294a <=( a1677a ) or ( a4293a );
 a4295a <=( a4294a ) or ( a4289a );
 a4296a <=( a4295a ) or ( a4286a );
 a4297a <=( a4296a ) or ( a4277a );
 a4298a <=( a4297a ) or ( a4258a );
 a4299a <=( a4298a ) or ( a4219a );
 a4302a <=( a1673a ) or ( a1674a );
 a4306a <=( a1670a ) or ( a1671a );
 a4307a <=( a1672a ) or ( a4306a );
 a4308a <=( a4307a ) or ( a4302a );
 a4311a <=( a1668a ) or ( a1669a );
 a4315a <=( a1665a ) or ( a1666a );
 a4316a <=( a1667a ) or ( a4315a );
 a4317a <=( a4316a ) or ( a4311a );
 a4318a <=( a4317a ) or ( a4308a );
 a4321a <=( a1663a ) or ( a1664a );
 a4325a <=( a1660a ) or ( a1661a );
 a4326a <=( a1662a ) or ( a4325a );
 a4327a <=( a4326a ) or ( a4321a );
 a4330a <=( a1658a ) or ( a1659a );
 a4334a <=( a1655a ) or ( a1656a );
 a4335a <=( a1657a ) or ( a4334a );
 a4336a <=( a4335a ) or ( a4330a );
 a4337a <=( a4336a ) or ( a4327a );
 a4338a <=( a4337a ) or ( a4318a );
 a4341a <=( a1653a ) or ( a1654a );
 a4345a <=( a1650a ) or ( a1651a );
 a4346a <=( a1652a ) or ( a4345a );
 a4347a <=( a4346a ) or ( a4341a );
 a4350a <=( a1648a ) or ( a1649a );
 a4354a <=( a1645a ) or ( a1646a );
 a4355a <=( a1647a ) or ( a4354a );
 a4356a <=( a4355a ) or ( a4350a );
 a4357a <=( a4356a ) or ( a4347a );
 a4360a <=( a1643a ) or ( a1644a );
 a4364a <=( a1640a ) or ( a1641a );
 a4365a <=( a1642a ) or ( a4364a );
 a4366a <=( a4365a ) or ( a4360a );
 a4369a <=( a1638a ) or ( a1639a );
 a4373a <=( a1635a ) or ( a1636a );
 a4374a <=( a1637a ) or ( a4373a );
 a4375a <=( a4374a ) or ( a4369a );
 a4376a <=( a4375a ) or ( a4366a );
 a4377a <=( a4376a ) or ( a4357a );
 a4378a <=( a4377a ) or ( a4338a );
 a4381a <=( a1633a ) or ( a1634a );
 a4385a <=( a1630a ) or ( a1631a );
 a4386a <=( a1632a ) or ( a4385a );
 a4387a <=( a4386a ) or ( a4381a );
 a4390a <=( a1628a ) or ( a1629a );
 a4394a <=( a1625a ) or ( a1626a );
 a4395a <=( a1627a ) or ( a4394a );
 a4396a <=( a4395a ) or ( a4390a );
 a4397a <=( a4396a ) or ( a4387a );
 a4400a <=( a1623a ) or ( a1624a );
 a4404a <=( a1620a ) or ( a1621a );
 a4405a <=( a1622a ) or ( a4404a );
 a4406a <=( a4405a ) or ( a4400a );
 a4409a <=( a1618a ) or ( a1619a );
 a4413a <=( a1615a ) or ( a1616a );
 a4414a <=( a1617a ) or ( a4413a );
 a4415a <=( a4414a ) or ( a4409a );
 a4416a <=( a4415a ) or ( a4406a );
 a4417a <=( a4416a ) or ( a4397a );
 a4420a <=( a1613a ) or ( a1614a );
 a4424a <=( a1610a ) or ( a1611a );
 a4425a <=( a1612a ) or ( a4424a );
 a4426a <=( a4425a ) or ( a4420a );
 a4429a <=( a1608a ) or ( a1609a );
 a4433a <=( a1605a ) or ( a1606a );
 a4434a <=( a1607a ) or ( a4433a );
 a4435a <=( a4434a ) or ( a4429a );
 a4436a <=( a4435a ) or ( a4426a );
 a4439a <=( a1603a ) or ( a1604a );
 a4443a <=( a1600a ) or ( a1601a );
 a4444a <=( a1602a ) or ( a4443a );
 a4445a <=( a4444a ) or ( a4439a );
 a4448a <=( a1598a ) or ( a1599a );
 a4452a <=( a1595a ) or ( a1596a );
 a4453a <=( a1597a ) or ( a4452a );
 a4454a <=( a4453a ) or ( a4448a );
 a4455a <=( a4454a ) or ( a4445a );
 a4456a <=( a4455a ) or ( a4436a );
 a4457a <=( a4456a ) or ( a4417a );
 a4458a <=( a4457a ) or ( a4378a );
 a4459a <=( a4458a ) or ( a4299a );
 a4460a <=( a4459a ) or ( a4140a );
 a4463a <=( a1593a ) or ( a1594a );
 a4466a <=( a1591a ) or ( a1592a );
 a4467a <=( a4466a ) or ( a4463a );
 a4470a <=( a1589a ) or ( a1590a );
 a4474a <=( a1586a ) or ( a1587a );
 a4475a <=( a1588a ) or ( a4474a );
 a4476a <=( a4475a ) or ( a4470a );
 a4477a <=( a4476a ) or ( a4467a );
 a4480a <=( a1584a ) or ( a1585a );
 a4484a <=( a1581a ) or ( a1582a );
 a4485a <=( a1583a ) or ( a4484a );
 a4486a <=( a4485a ) or ( a4480a );
 a4489a <=( a1579a ) or ( a1580a );
 a4493a <=( a1576a ) or ( a1577a );
 a4494a <=( a1578a ) or ( a4493a );
 a4495a <=( a4494a ) or ( a4489a );
 a4496a <=( a4495a ) or ( a4486a );
 a4497a <=( a4496a ) or ( a4477a );
 a4500a <=( a1574a ) or ( a1575a );
 a4504a <=( a1571a ) or ( a1572a );
 a4505a <=( a1573a ) or ( a4504a );
 a4506a <=( a4505a ) or ( a4500a );
 a4509a <=( a1569a ) or ( a1570a );
 a4513a <=( a1566a ) or ( a1567a );
 a4514a <=( a1568a ) or ( a4513a );
 a4515a <=( a4514a ) or ( a4509a );
 a4516a <=( a4515a ) or ( a4506a );
 a4519a <=( a1564a ) or ( a1565a );
 a4523a <=( a1561a ) or ( a1562a );
 a4524a <=( a1563a ) or ( a4523a );
 a4525a <=( a4524a ) or ( a4519a );
 a4528a <=( a1559a ) or ( a1560a );
 a4532a <=( a1556a ) or ( a1557a );
 a4533a <=( a1558a ) or ( a4532a );
 a4534a <=( a4533a ) or ( a4528a );
 a4535a <=( a4534a ) or ( a4525a );
 a4536a <=( a4535a ) or ( a4516a );
 a4537a <=( a4536a ) or ( a4497a );
 a4540a <=( a1554a ) or ( a1555a );
 a4544a <=( a1551a ) or ( a1552a );
 a4545a <=( a1553a ) or ( a4544a );
 a4546a <=( a4545a ) or ( a4540a );
 a4549a <=( a1549a ) or ( a1550a );
 a4553a <=( a1546a ) or ( a1547a );
 a4554a <=( a1548a ) or ( a4553a );
 a4555a <=( a4554a ) or ( a4549a );
 a4556a <=( a4555a ) or ( a4546a );
 a4559a <=( a1544a ) or ( a1545a );
 a4563a <=( a1541a ) or ( a1542a );
 a4564a <=( a1543a ) or ( a4563a );
 a4565a <=( a4564a ) or ( a4559a );
 a4568a <=( a1539a ) or ( a1540a );
 a4572a <=( a1536a ) or ( a1537a );
 a4573a <=( a1538a ) or ( a4572a );
 a4574a <=( a4573a ) or ( a4568a );
 a4575a <=( a4574a ) or ( a4565a );
 a4576a <=( a4575a ) or ( a4556a );
 a4579a <=( a1534a ) or ( a1535a );
 a4583a <=( a1531a ) or ( a1532a );
 a4584a <=( a1533a ) or ( a4583a );
 a4585a <=( a4584a ) or ( a4579a );
 a4588a <=( a1529a ) or ( a1530a );
 a4592a <=( a1526a ) or ( a1527a );
 a4593a <=( a1528a ) or ( a4592a );
 a4594a <=( a4593a ) or ( a4588a );
 a4595a <=( a4594a ) or ( a4585a );
 a4598a <=( a1524a ) or ( a1525a );
 a4602a <=( a1521a ) or ( a1522a );
 a4603a <=( a1523a ) or ( a4602a );
 a4604a <=( a4603a ) or ( a4598a );
 a4607a <=( a1519a ) or ( a1520a );
 a4611a <=( a1516a ) or ( a1517a );
 a4612a <=( a1518a ) or ( a4611a );
 a4613a <=( a4612a ) or ( a4607a );
 a4614a <=( a4613a ) or ( a4604a );
 a4615a <=( a4614a ) or ( a4595a );
 a4616a <=( a4615a ) or ( a4576a );
 a4617a <=( a4616a ) or ( a4537a );
 a4620a <=( a1514a ) or ( a1515a );
 a4624a <=( a1511a ) or ( a1512a );
 a4625a <=( a1513a ) or ( a4624a );
 a4626a <=( a4625a ) or ( a4620a );
 a4629a <=( a1509a ) or ( a1510a );
 a4633a <=( a1506a ) or ( a1507a );
 a4634a <=( a1508a ) or ( a4633a );
 a4635a <=( a4634a ) or ( a4629a );
 a4636a <=( a4635a ) or ( a4626a );
 a4639a <=( a1504a ) or ( a1505a );
 a4643a <=( a1501a ) or ( a1502a );
 a4644a <=( a1503a ) or ( a4643a );
 a4645a <=( a4644a ) or ( a4639a );
 a4648a <=( a1499a ) or ( a1500a );
 a4652a <=( a1496a ) or ( a1497a );
 a4653a <=( a1498a ) or ( a4652a );
 a4654a <=( a4653a ) or ( a4648a );
 a4655a <=( a4654a ) or ( a4645a );
 a4656a <=( a4655a ) or ( a4636a );
 a4659a <=( a1494a ) or ( a1495a );
 a4663a <=( a1491a ) or ( a1492a );
 a4664a <=( a1493a ) or ( a4663a );
 a4665a <=( a4664a ) or ( a4659a );
 a4668a <=( a1489a ) or ( a1490a );
 a4672a <=( a1486a ) or ( a1487a );
 a4673a <=( a1488a ) or ( a4672a );
 a4674a <=( a4673a ) or ( a4668a );
 a4675a <=( a4674a ) or ( a4665a );
 a4678a <=( a1484a ) or ( a1485a );
 a4682a <=( a1481a ) or ( a1482a );
 a4683a <=( a1483a ) or ( a4682a );
 a4684a <=( a4683a ) or ( a4678a );
 a4687a <=( a1479a ) or ( a1480a );
 a4691a <=( a1476a ) or ( a1477a );
 a4692a <=( a1478a ) or ( a4691a );
 a4693a <=( a4692a ) or ( a4687a );
 a4694a <=( a4693a ) or ( a4684a );
 a4695a <=( a4694a ) or ( a4675a );
 a4696a <=( a4695a ) or ( a4656a );
 a4699a <=( a1474a ) or ( a1475a );
 a4703a <=( a1471a ) or ( a1472a );
 a4704a <=( a1473a ) or ( a4703a );
 a4705a <=( a4704a ) or ( a4699a );
 a4708a <=( a1469a ) or ( a1470a );
 a4712a <=( a1466a ) or ( a1467a );
 a4713a <=( a1468a ) or ( a4712a );
 a4714a <=( a4713a ) or ( a4708a );
 a4715a <=( a4714a ) or ( a4705a );
 a4718a <=( a1464a ) or ( a1465a );
 a4722a <=( a1461a ) or ( a1462a );
 a4723a <=( a1463a ) or ( a4722a );
 a4724a <=( a4723a ) or ( a4718a );
 a4727a <=( a1459a ) or ( a1460a );
 a4731a <=( a1456a ) or ( a1457a );
 a4732a <=( a1458a ) or ( a4731a );
 a4733a <=( a4732a ) or ( a4727a );
 a4734a <=( a4733a ) or ( a4724a );
 a4735a <=( a4734a ) or ( a4715a );
 a4738a <=( a1454a ) or ( a1455a );
 a4742a <=( a1451a ) or ( a1452a );
 a4743a <=( a1453a ) or ( a4742a );
 a4744a <=( a4743a ) or ( a4738a );
 a4747a <=( a1449a ) or ( a1450a );
 a4751a <=( a1446a ) or ( a1447a );
 a4752a <=( a1448a ) or ( a4751a );
 a4753a <=( a4752a ) or ( a4747a );
 a4754a <=( a4753a ) or ( a4744a );
 a4757a <=( a1444a ) or ( a1445a );
 a4761a <=( a1441a ) or ( a1442a );
 a4762a <=( a1443a ) or ( a4761a );
 a4763a <=( a4762a ) or ( a4757a );
 a4766a <=( a1439a ) or ( a1440a );
 a4770a <=( a1436a ) or ( a1437a );
 a4771a <=( a1438a ) or ( a4770a );
 a4772a <=( a4771a ) or ( a4766a );
 a4773a <=( a4772a ) or ( a4763a );
 a4774a <=( a4773a ) or ( a4754a );
 a4775a <=( a4774a ) or ( a4735a );
 a4776a <=( a4775a ) or ( a4696a );
 a4777a <=( a4776a ) or ( a4617a );
 a4780a <=( a1434a ) or ( a1435a );
 a4784a <=( a1431a ) or ( a1432a );
 a4785a <=( a1433a ) or ( a4784a );
 a4786a <=( a4785a ) or ( a4780a );
 a4789a <=( a1429a ) or ( a1430a );
 a4793a <=( a1426a ) or ( a1427a );
 a4794a <=( a1428a ) or ( a4793a );
 a4795a <=( a4794a ) or ( a4789a );
 a4796a <=( a4795a ) or ( a4786a );
 a4799a <=( a1424a ) or ( a1425a );
 a4803a <=( a1421a ) or ( a1422a );
 a4804a <=( a1423a ) or ( a4803a );
 a4805a <=( a4804a ) or ( a4799a );
 a4808a <=( a1419a ) or ( a1420a );
 a4812a <=( a1416a ) or ( a1417a );
 a4813a <=( a1418a ) or ( a4812a );
 a4814a <=( a4813a ) or ( a4808a );
 a4815a <=( a4814a ) or ( a4805a );
 a4816a <=( a4815a ) or ( a4796a );
 a4819a <=( a1414a ) or ( a1415a );
 a4823a <=( a1411a ) or ( a1412a );
 a4824a <=( a1413a ) or ( a4823a );
 a4825a <=( a4824a ) or ( a4819a );
 a4828a <=( a1409a ) or ( a1410a );
 a4832a <=( a1406a ) or ( a1407a );
 a4833a <=( a1408a ) or ( a4832a );
 a4834a <=( a4833a ) or ( a4828a );
 a4835a <=( a4834a ) or ( a4825a );
 a4838a <=( a1404a ) or ( a1405a );
 a4842a <=( a1401a ) or ( a1402a );
 a4843a <=( a1403a ) or ( a4842a );
 a4844a <=( a4843a ) or ( a4838a );
 a4847a <=( a1399a ) or ( a1400a );
 a4851a <=( a1396a ) or ( a1397a );
 a4852a <=( a1398a ) or ( a4851a );
 a4853a <=( a4852a ) or ( a4847a );
 a4854a <=( a4853a ) or ( a4844a );
 a4855a <=( a4854a ) or ( a4835a );
 a4856a <=( a4855a ) or ( a4816a );
 a4859a <=( a1394a ) or ( a1395a );
 a4863a <=( a1391a ) or ( a1392a );
 a4864a <=( a1393a ) or ( a4863a );
 a4865a <=( a4864a ) or ( a4859a );
 a4868a <=( a1389a ) or ( a1390a );
 a4872a <=( a1386a ) or ( a1387a );
 a4873a <=( a1388a ) or ( a4872a );
 a4874a <=( a4873a ) or ( a4868a );
 a4875a <=( a4874a ) or ( a4865a );
 a4878a <=( a1384a ) or ( a1385a );
 a4882a <=( a1381a ) or ( a1382a );
 a4883a <=( a1383a ) or ( a4882a );
 a4884a <=( a4883a ) or ( a4878a );
 a4887a <=( a1379a ) or ( a1380a );
 a4891a <=( a1376a ) or ( a1377a );
 a4892a <=( a1378a ) or ( a4891a );
 a4893a <=( a4892a ) or ( a4887a );
 a4894a <=( a4893a ) or ( a4884a );
 a4895a <=( a4894a ) or ( a4875a );
 a4898a <=( a1374a ) or ( a1375a );
 a4902a <=( a1371a ) or ( a1372a );
 a4903a <=( a1373a ) or ( a4902a );
 a4904a <=( a4903a ) or ( a4898a );
 a4907a <=( a1369a ) or ( a1370a );
 a4911a <=( a1366a ) or ( a1367a );
 a4912a <=( a1368a ) or ( a4911a );
 a4913a <=( a4912a ) or ( a4907a );
 a4914a <=( a4913a ) or ( a4904a );
 a4917a <=( a1364a ) or ( a1365a );
 a4921a <=( a1361a ) or ( a1362a );
 a4922a <=( a1363a ) or ( a4921a );
 a4923a <=( a4922a ) or ( a4917a );
 a4926a <=( a1359a ) or ( a1360a );
 a4930a <=( a1356a ) or ( a1357a );
 a4931a <=( a1358a ) or ( a4930a );
 a4932a <=( a4931a ) or ( a4926a );
 a4933a <=( a4932a ) or ( a4923a );
 a4934a <=( a4933a ) or ( a4914a );
 a4935a <=( a4934a ) or ( a4895a );
 a4936a <=( a4935a ) or ( a4856a );
 a4939a <=( a1354a ) or ( a1355a );
 a4943a <=( a1351a ) or ( a1352a );
 a4944a <=( a1353a ) or ( a4943a );
 a4945a <=( a4944a ) or ( a4939a );
 a4948a <=( a1349a ) or ( a1350a );
 a4952a <=( a1346a ) or ( a1347a );
 a4953a <=( a1348a ) or ( a4952a );
 a4954a <=( a4953a ) or ( a4948a );
 a4955a <=( a4954a ) or ( a4945a );
 a4958a <=( a1344a ) or ( a1345a );
 a4962a <=( a1341a ) or ( a1342a );
 a4963a <=( a1343a ) or ( a4962a );
 a4964a <=( a4963a ) or ( a4958a );
 a4967a <=( a1339a ) or ( a1340a );
 a4971a <=( a1336a ) or ( a1337a );
 a4972a <=( a1338a ) or ( a4971a );
 a4973a <=( a4972a ) or ( a4967a );
 a4974a <=( a4973a ) or ( a4964a );
 a4975a <=( a4974a ) or ( a4955a );
 a4978a <=( a1334a ) or ( a1335a );
 a4982a <=( a1331a ) or ( a1332a );
 a4983a <=( a1333a ) or ( a4982a );
 a4984a <=( a4983a ) or ( a4978a );
 a4987a <=( a1329a ) or ( a1330a );
 a4991a <=( a1326a ) or ( a1327a );
 a4992a <=( a1328a ) or ( a4991a );
 a4993a <=( a4992a ) or ( a4987a );
 a4994a <=( a4993a ) or ( a4984a );
 a4997a <=( a1324a ) or ( a1325a );
 a5001a <=( a1321a ) or ( a1322a );
 a5002a <=( a1323a ) or ( a5001a );
 a5003a <=( a5002a ) or ( a4997a );
 a5006a <=( a1319a ) or ( a1320a );
 a5010a <=( a1316a ) or ( a1317a );
 a5011a <=( a1318a ) or ( a5010a );
 a5012a <=( a5011a ) or ( a5006a );
 a5013a <=( a5012a ) or ( a5003a );
 a5014a <=( a5013a ) or ( a4994a );
 a5015a <=( a5014a ) or ( a4975a );
 a5018a <=( a1314a ) or ( a1315a );
 a5022a <=( a1311a ) or ( a1312a );
 a5023a <=( a1313a ) or ( a5022a );
 a5024a <=( a5023a ) or ( a5018a );
 a5027a <=( a1309a ) or ( a1310a );
 a5031a <=( a1306a ) or ( a1307a );
 a5032a <=( a1308a ) or ( a5031a );
 a5033a <=( a5032a ) or ( a5027a );
 a5034a <=( a5033a ) or ( a5024a );
 a5037a <=( a1304a ) or ( a1305a );
 a5041a <=( a1301a ) or ( a1302a );
 a5042a <=( a1303a ) or ( a5041a );
 a5043a <=( a5042a ) or ( a5037a );
 a5046a <=( a1299a ) or ( a1300a );
 a5050a <=( a1296a ) or ( a1297a );
 a5051a <=( a1298a ) or ( a5050a );
 a5052a <=( a5051a ) or ( a5046a );
 a5053a <=( a5052a ) or ( a5043a );
 a5054a <=( a5053a ) or ( a5034a );
 a5057a <=( a1294a ) or ( a1295a );
 a5061a <=( a1291a ) or ( a1292a );
 a5062a <=( a1293a ) or ( a5061a );
 a5063a <=( a5062a ) or ( a5057a );
 a5066a <=( a1289a ) or ( a1290a );
 a5070a <=( a1286a ) or ( a1287a );
 a5071a <=( a1288a ) or ( a5070a );
 a5072a <=( a5071a ) or ( a5066a );
 a5073a <=( a5072a ) or ( a5063a );
 a5076a <=( a1284a ) or ( a1285a );
 a5080a <=( a1281a ) or ( a1282a );
 a5081a <=( a1283a ) or ( a5080a );
 a5082a <=( a5081a ) or ( a5076a );
 a5085a <=( a1279a ) or ( a1280a );
 a5089a <=( a1276a ) or ( a1277a );
 a5090a <=( a1278a ) or ( a5089a );
 a5091a <=( a5090a ) or ( a5085a );
 a5092a <=( a5091a ) or ( a5082a );
 a5093a <=( a5092a ) or ( a5073a );
 a5094a <=( a5093a ) or ( a5054a );
 a5095a <=( a5094a ) or ( a5015a );
 a5096a <=( a5095a ) or ( a4936a );
 a5097a <=( a5096a ) or ( a4777a );
 a5098a <=( a5097a ) or ( a4460a );
 a5099a <=( a5098a ) or ( a3823a );
 a5102a <=( a1274a ) or ( a1275a );
 a5105a <=( a1272a ) or ( a1273a );
 a5106a <=( a5105a ) or ( a5102a );
 a5109a <=( a1270a ) or ( a1271a );
 a5113a <=( a1267a ) or ( a1268a );
 a5114a <=( a1269a ) or ( a5113a );
 a5115a <=( a5114a ) or ( a5109a );
 a5116a <=( a5115a ) or ( a5106a );
 a5119a <=( a1265a ) or ( a1266a );
 a5123a <=( a1262a ) or ( a1263a );
 a5124a <=( a1264a ) or ( a5123a );
 a5125a <=( a5124a ) or ( a5119a );
 a5128a <=( a1260a ) or ( a1261a );
 a5132a <=( a1257a ) or ( a1258a );
 a5133a <=( a1259a ) or ( a5132a );
 a5134a <=( a5133a ) or ( a5128a );
 a5135a <=( a5134a ) or ( a5125a );
 a5136a <=( a5135a ) or ( a5116a );
 a5139a <=( a1255a ) or ( a1256a );
 a5143a <=( a1252a ) or ( a1253a );
 a5144a <=( a1254a ) or ( a5143a );
 a5145a <=( a5144a ) or ( a5139a );
 a5148a <=( a1250a ) or ( a1251a );
 a5152a <=( a1247a ) or ( a1248a );
 a5153a <=( a1249a ) or ( a5152a );
 a5154a <=( a5153a ) or ( a5148a );
 a5155a <=( a5154a ) or ( a5145a );
 a5158a <=( a1245a ) or ( a1246a );
 a5162a <=( a1242a ) or ( a1243a );
 a5163a <=( a1244a ) or ( a5162a );
 a5164a <=( a5163a ) or ( a5158a );
 a5167a <=( a1240a ) or ( a1241a );
 a5171a <=( a1237a ) or ( a1238a );
 a5172a <=( a1239a ) or ( a5171a );
 a5173a <=( a5172a ) or ( a5167a );
 a5174a <=( a5173a ) or ( a5164a );
 a5175a <=( a5174a ) or ( a5155a );
 a5176a <=( a5175a ) or ( a5136a );
 a5179a <=( a1235a ) or ( a1236a );
 a5183a <=( a1232a ) or ( a1233a );
 a5184a <=( a1234a ) or ( a5183a );
 a5185a <=( a5184a ) or ( a5179a );
 a5188a <=( a1230a ) or ( a1231a );
 a5192a <=( a1227a ) or ( a1228a );
 a5193a <=( a1229a ) or ( a5192a );
 a5194a <=( a5193a ) or ( a5188a );
 a5195a <=( a5194a ) or ( a5185a );
 a5198a <=( a1225a ) or ( a1226a );
 a5202a <=( a1222a ) or ( a1223a );
 a5203a <=( a1224a ) or ( a5202a );
 a5204a <=( a5203a ) or ( a5198a );
 a5207a <=( a1220a ) or ( a1221a );
 a5211a <=( a1217a ) or ( a1218a );
 a5212a <=( a1219a ) or ( a5211a );
 a5213a <=( a5212a ) or ( a5207a );
 a5214a <=( a5213a ) or ( a5204a );
 a5215a <=( a5214a ) or ( a5195a );
 a5218a <=( a1215a ) or ( a1216a );
 a5222a <=( a1212a ) or ( a1213a );
 a5223a <=( a1214a ) or ( a5222a );
 a5224a <=( a5223a ) or ( a5218a );
 a5227a <=( a1210a ) or ( a1211a );
 a5231a <=( a1207a ) or ( a1208a );
 a5232a <=( a1209a ) or ( a5231a );
 a5233a <=( a5232a ) or ( a5227a );
 a5234a <=( a5233a ) or ( a5224a );
 a5237a <=( a1205a ) or ( a1206a );
 a5241a <=( a1202a ) or ( a1203a );
 a5242a <=( a1204a ) or ( a5241a );
 a5243a <=( a5242a ) or ( a5237a );
 a5246a <=( a1200a ) or ( a1201a );
 a5250a <=( a1197a ) or ( a1198a );
 a5251a <=( a1199a ) or ( a5250a );
 a5252a <=( a5251a ) or ( a5246a );
 a5253a <=( a5252a ) or ( a5243a );
 a5254a <=( a5253a ) or ( a5234a );
 a5255a <=( a5254a ) or ( a5215a );
 a5256a <=( a5255a ) or ( a5176a );
 a5259a <=( a1195a ) or ( a1196a );
 a5263a <=( a1192a ) or ( a1193a );
 a5264a <=( a1194a ) or ( a5263a );
 a5265a <=( a5264a ) or ( a5259a );
 a5268a <=( a1190a ) or ( a1191a );
 a5272a <=( a1187a ) or ( a1188a );
 a5273a <=( a1189a ) or ( a5272a );
 a5274a <=( a5273a ) or ( a5268a );
 a5275a <=( a5274a ) or ( a5265a );
 a5278a <=( a1185a ) or ( a1186a );
 a5282a <=( a1182a ) or ( a1183a );
 a5283a <=( a1184a ) or ( a5282a );
 a5284a <=( a5283a ) or ( a5278a );
 a5287a <=( a1180a ) or ( a1181a );
 a5291a <=( a1177a ) or ( a1178a );
 a5292a <=( a1179a ) or ( a5291a );
 a5293a <=( a5292a ) or ( a5287a );
 a5294a <=( a5293a ) or ( a5284a );
 a5295a <=( a5294a ) or ( a5275a );
 a5298a <=( a1175a ) or ( a1176a );
 a5302a <=( a1172a ) or ( a1173a );
 a5303a <=( a1174a ) or ( a5302a );
 a5304a <=( a5303a ) or ( a5298a );
 a5307a <=( a1170a ) or ( a1171a );
 a5311a <=( a1167a ) or ( a1168a );
 a5312a <=( a1169a ) or ( a5311a );
 a5313a <=( a5312a ) or ( a5307a );
 a5314a <=( a5313a ) or ( a5304a );
 a5317a <=( a1165a ) or ( a1166a );
 a5321a <=( a1162a ) or ( a1163a );
 a5322a <=( a1164a ) or ( a5321a );
 a5323a <=( a5322a ) or ( a5317a );
 a5326a <=( a1160a ) or ( a1161a );
 a5330a <=( a1157a ) or ( a1158a );
 a5331a <=( a1159a ) or ( a5330a );
 a5332a <=( a5331a ) or ( a5326a );
 a5333a <=( a5332a ) or ( a5323a );
 a5334a <=( a5333a ) or ( a5314a );
 a5335a <=( a5334a ) or ( a5295a );
 a5338a <=( a1155a ) or ( a1156a );
 a5342a <=( a1152a ) or ( a1153a );
 a5343a <=( a1154a ) or ( a5342a );
 a5344a <=( a5343a ) or ( a5338a );
 a5347a <=( a1150a ) or ( a1151a );
 a5351a <=( a1147a ) or ( a1148a );
 a5352a <=( a1149a ) or ( a5351a );
 a5353a <=( a5352a ) or ( a5347a );
 a5354a <=( a5353a ) or ( a5344a );
 a5357a <=( a1145a ) or ( a1146a );
 a5361a <=( a1142a ) or ( a1143a );
 a5362a <=( a1144a ) or ( a5361a );
 a5363a <=( a5362a ) or ( a5357a );
 a5366a <=( a1140a ) or ( a1141a );
 a5370a <=( a1137a ) or ( a1138a );
 a5371a <=( a1139a ) or ( a5370a );
 a5372a <=( a5371a ) or ( a5366a );
 a5373a <=( a5372a ) or ( a5363a );
 a5374a <=( a5373a ) or ( a5354a );
 a5377a <=( a1135a ) or ( a1136a );
 a5381a <=( a1132a ) or ( a1133a );
 a5382a <=( a1134a ) or ( a5381a );
 a5383a <=( a5382a ) or ( a5377a );
 a5386a <=( a1130a ) or ( a1131a );
 a5390a <=( a1127a ) or ( a1128a );
 a5391a <=( a1129a ) or ( a5390a );
 a5392a <=( a5391a ) or ( a5386a );
 a5393a <=( a5392a ) or ( a5383a );
 a5396a <=( a1125a ) or ( a1126a );
 a5400a <=( a1122a ) or ( a1123a );
 a5401a <=( a1124a ) or ( a5400a );
 a5402a <=( a5401a ) or ( a5396a );
 a5405a <=( a1120a ) or ( a1121a );
 a5409a <=( a1117a ) or ( a1118a );
 a5410a <=( a1119a ) or ( a5409a );
 a5411a <=( a5410a ) or ( a5405a );
 a5412a <=( a5411a ) or ( a5402a );
 a5413a <=( a5412a ) or ( a5393a );
 a5414a <=( a5413a ) or ( a5374a );
 a5415a <=( a5414a ) or ( a5335a );
 a5416a <=( a5415a ) or ( a5256a );
 a5419a <=( a1115a ) or ( a1116a );
 a5422a <=( a1113a ) or ( a1114a );
 a5423a <=( a5422a ) or ( a5419a );
 a5426a <=( a1111a ) or ( a1112a );
 a5430a <=( a1108a ) or ( a1109a );
 a5431a <=( a1110a ) or ( a5430a );
 a5432a <=( a5431a ) or ( a5426a );
 a5433a <=( a5432a ) or ( a5423a );
 a5436a <=( a1106a ) or ( a1107a );
 a5440a <=( a1103a ) or ( a1104a );
 a5441a <=( a1105a ) or ( a5440a );
 a5442a <=( a5441a ) or ( a5436a );
 a5445a <=( a1101a ) or ( a1102a );
 a5449a <=( a1098a ) or ( a1099a );
 a5450a <=( a1100a ) or ( a5449a );
 a5451a <=( a5450a ) or ( a5445a );
 a5452a <=( a5451a ) or ( a5442a );
 a5453a <=( a5452a ) or ( a5433a );
 a5456a <=( a1096a ) or ( a1097a );
 a5460a <=( a1093a ) or ( a1094a );
 a5461a <=( a1095a ) or ( a5460a );
 a5462a <=( a5461a ) or ( a5456a );
 a5465a <=( a1091a ) or ( a1092a );
 a5469a <=( a1088a ) or ( a1089a );
 a5470a <=( a1090a ) or ( a5469a );
 a5471a <=( a5470a ) or ( a5465a );
 a5472a <=( a5471a ) or ( a5462a );
 a5475a <=( a1086a ) or ( a1087a );
 a5479a <=( a1083a ) or ( a1084a );
 a5480a <=( a1085a ) or ( a5479a );
 a5481a <=( a5480a ) or ( a5475a );
 a5484a <=( a1081a ) or ( a1082a );
 a5488a <=( a1078a ) or ( a1079a );
 a5489a <=( a1080a ) or ( a5488a );
 a5490a <=( a5489a ) or ( a5484a );
 a5491a <=( a5490a ) or ( a5481a );
 a5492a <=( a5491a ) or ( a5472a );
 a5493a <=( a5492a ) or ( a5453a );
 a5496a <=( a1076a ) or ( a1077a );
 a5500a <=( a1073a ) or ( a1074a );
 a5501a <=( a1075a ) or ( a5500a );
 a5502a <=( a5501a ) or ( a5496a );
 a5505a <=( a1071a ) or ( a1072a );
 a5509a <=( a1068a ) or ( a1069a );
 a5510a <=( a1070a ) or ( a5509a );
 a5511a <=( a5510a ) or ( a5505a );
 a5512a <=( a5511a ) or ( a5502a );
 a5515a <=( a1066a ) or ( a1067a );
 a5519a <=( a1063a ) or ( a1064a );
 a5520a <=( a1065a ) or ( a5519a );
 a5521a <=( a5520a ) or ( a5515a );
 a5524a <=( a1061a ) or ( a1062a );
 a5528a <=( a1058a ) or ( a1059a );
 a5529a <=( a1060a ) or ( a5528a );
 a5530a <=( a5529a ) or ( a5524a );
 a5531a <=( a5530a ) or ( a5521a );
 a5532a <=( a5531a ) or ( a5512a );
 a5535a <=( a1056a ) or ( a1057a );
 a5539a <=( a1053a ) or ( a1054a );
 a5540a <=( a1055a ) or ( a5539a );
 a5541a <=( a5540a ) or ( a5535a );
 a5544a <=( a1051a ) or ( a1052a );
 a5548a <=( a1048a ) or ( a1049a );
 a5549a <=( a1050a ) or ( a5548a );
 a5550a <=( a5549a ) or ( a5544a );
 a5551a <=( a5550a ) or ( a5541a );
 a5554a <=( a1046a ) or ( a1047a );
 a5558a <=( a1043a ) or ( a1044a );
 a5559a <=( a1045a ) or ( a5558a );
 a5560a <=( a5559a ) or ( a5554a );
 a5563a <=( a1041a ) or ( a1042a );
 a5567a <=( a1038a ) or ( a1039a );
 a5568a <=( a1040a ) or ( a5567a );
 a5569a <=( a5568a ) or ( a5563a );
 a5570a <=( a5569a ) or ( a5560a );
 a5571a <=( a5570a ) or ( a5551a );
 a5572a <=( a5571a ) or ( a5532a );
 a5573a <=( a5572a ) or ( a5493a );
 a5576a <=( a1036a ) or ( a1037a );
 a5580a <=( a1033a ) or ( a1034a );
 a5581a <=( a1035a ) or ( a5580a );
 a5582a <=( a5581a ) or ( a5576a );
 a5585a <=( a1031a ) or ( a1032a );
 a5589a <=( a1028a ) or ( a1029a );
 a5590a <=( a1030a ) or ( a5589a );
 a5591a <=( a5590a ) or ( a5585a );
 a5592a <=( a5591a ) or ( a5582a );
 a5595a <=( a1026a ) or ( a1027a );
 a5599a <=( a1023a ) or ( a1024a );
 a5600a <=( a1025a ) or ( a5599a );
 a5601a <=( a5600a ) or ( a5595a );
 a5604a <=( a1021a ) or ( a1022a );
 a5608a <=( a1018a ) or ( a1019a );
 a5609a <=( a1020a ) or ( a5608a );
 a5610a <=( a5609a ) or ( a5604a );
 a5611a <=( a5610a ) or ( a5601a );
 a5612a <=( a5611a ) or ( a5592a );
 a5615a <=( a1016a ) or ( a1017a );
 a5619a <=( a1013a ) or ( a1014a );
 a5620a <=( a1015a ) or ( a5619a );
 a5621a <=( a5620a ) or ( a5615a );
 a5624a <=( a1011a ) or ( a1012a );
 a5628a <=( a1008a ) or ( a1009a );
 a5629a <=( a1010a ) or ( a5628a );
 a5630a <=( a5629a ) or ( a5624a );
 a5631a <=( a5630a ) or ( a5621a );
 a5634a <=( a1006a ) or ( a1007a );
 a5638a <=( a1003a ) or ( a1004a );
 a5639a <=( a1005a ) or ( a5638a );
 a5640a <=( a5639a ) or ( a5634a );
 a5643a <=( a1001a ) or ( a1002a );
 a5647a <=( a998a ) or ( a999a );
 a5648a <=( a1000a ) or ( a5647a );
 a5649a <=( a5648a ) or ( a5643a );
 a5650a <=( a5649a ) or ( a5640a );
 a5651a <=( a5650a ) or ( a5631a );
 a5652a <=( a5651a ) or ( a5612a );
 a5655a <=( a996a ) or ( a997a );
 a5659a <=( a993a ) or ( a994a );
 a5660a <=( a995a ) or ( a5659a );
 a5661a <=( a5660a ) or ( a5655a );
 a5664a <=( a991a ) or ( a992a );
 a5668a <=( a988a ) or ( a989a );
 a5669a <=( a990a ) or ( a5668a );
 a5670a <=( a5669a ) or ( a5664a );
 a5671a <=( a5670a ) or ( a5661a );
 a5674a <=( a986a ) or ( a987a );
 a5678a <=( a983a ) or ( a984a );
 a5679a <=( a985a ) or ( a5678a );
 a5680a <=( a5679a ) or ( a5674a );
 a5683a <=( a981a ) or ( a982a );
 a5687a <=( a978a ) or ( a979a );
 a5688a <=( a980a ) or ( a5687a );
 a5689a <=( a5688a ) or ( a5683a );
 a5690a <=( a5689a ) or ( a5680a );
 a5691a <=( a5690a ) or ( a5671a );
 a5694a <=( a976a ) or ( a977a );
 a5698a <=( a973a ) or ( a974a );
 a5699a <=( a975a ) or ( a5698a );
 a5700a <=( a5699a ) or ( a5694a );
 a5703a <=( a971a ) or ( a972a );
 a5707a <=( a968a ) or ( a969a );
 a5708a <=( a970a ) or ( a5707a );
 a5709a <=( a5708a ) or ( a5703a );
 a5710a <=( a5709a ) or ( a5700a );
 a5713a <=( a966a ) or ( a967a );
 a5717a <=( a963a ) or ( a964a );
 a5718a <=( a965a ) or ( a5717a );
 a5719a <=( a5718a ) or ( a5713a );
 a5722a <=( a961a ) or ( a962a );
 a5726a <=( a958a ) or ( a959a );
 a5727a <=( a960a ) or ( a5726a );
 a5728a <=( a5727a ) or ( a5722a );
 a5729a <=( a5728a ) or ( a5719a );
 a5730a <=( a5729a ) or ( a5710a );
 a5731a <=( a5730a ) or ( a5691a );
 a5732a <=( a5731a ) or ( a5652a );
 a5733a <=( a5732a ) or ( a5573a );
 a5734a <=( a5733a ) or ( a5416a );
 a5737a <=( a956a ) or ( a957a );
 a5740a <=( a954a ) or ( a955a );
 a5741a <=( a5740a ) or ( a5737a );
 a5744a <=( a952a ) or ( a953a );
 a5748a <=( a949a ) or ( a950a );
 a5749a <=( a951a ) or ( a5748a );
 a5750a <=( a5749a ) or ( a5744a );
 a5751a <=( a5750a ) or ( a5741a );
 a5754a <=( a947a ) or ( a948a );
 a5758a <=( a944a ) or ( a945a );
 a5759a <=( a946a ) or ( a5758a );
 a5760a <=( a5759a ) or ( a5754a );
 a5763a <=( a942a ) or ( a943a );
 a5767a <=( a939a ) or ( a940a );
 a5768a <=( a941a ) or ( a5767a );
 a5769a <=( a5768a ) or ( a5763a );
 a5770a <=( a5769a ) or ( a5760a );
 a5771a <=( a5770a ) or ( a5751a );
 a5774a <=( a937a ) or ( a938a );
 a5778a <=( a934a ) or ( a935a );
 a5779a <=( a936a ) or ( a5778a );
 a5780a <=( a5779a ) or ( a5774a );
 a5783a <=( a932a ) or ( a933a );
 a5787a <=( a929a ) or ( a930a );
 a5788a <=( a931a ) or ( a5787a );
 a5789a <=( a5788a ) or ( a5783a );
 a5790a <=( a5789a ) or ( a5780a );
 a5793a <=( a927a ) or ( a928a );
 a5797a <=( a924a ) or ( a925a );
 a5798a <=( a926a ) or ( a5797a );
 a5799a <=( a5798a ) or ( a5793a );
 a5802a <=( a922a ) or ( a923a );
 a5806a <=( a919a ) or ( a920a );
 a5807a <=( a921a ) or ( a5806a );
 a5808a <=( a5807a ) or ( a5802a );
 a5809a <=( a5808a ) or ( a5799a );
 a5810a <=( a5809a ) or ( a5790a );
 a5811a <=( a5810a ) or ( a5771a );
 a5814a <=( a917a ) or ( a918a );
 a5818a <=( a914a ) or ( a915a );
 a5819a <=( a916a ) or ( a5818a );
 a5820a <=( a5819a ) or ( a5814a );
 a5823a <=( a912a ) or ( a913a );
 a5827a <=( a909a ) or ( a910a );
 a5828a <=( a911a ) or ( a5827a );
 a5829a <=( a5828a ) or ( a5823a );
 a5830a <=( a5829a ) or ( a5820a );
 a5833a <=( a907a ) or ( a908a );
 a5837a <=( a904a ) or ( a905a );
 a5838a <=( a906a ) or ( a5837a );
 a5839a <=( a5838a ) or ( a5833a );
 a5842a <=( a902a ) or ( a903a );
 a5846a <=( a899a ) or ( a900a );
 a5847a <=( a901a ) or ( a5846a );
 a5848a <=( a5847a ) or ( a5842a );
 a5849a <=( a5848a ) or ( a5839a );
 a5850a <=( a5849a ) or ( a5830a );
 a5853a <=( a897a ) or ( a898a );
 a5857a <=( a894a ) or ( a895a );
 a5858a <=( a896a ) or ( a5857a );
 a5859a <=( a5858a ) or ( a5853a );
 a5862a <=( a892a ) or ( a893a );
 a5866a <=( a889a ) or ( a890a );
 a5867a <=( a891a ) or ( a5866a );
 a5868a <=( a5867a ) or ( a5862a );
 a5869a <=( a5868a ) or ( a5859a );
 a5872a <=( a887a ) or ( a888a );
 a5876a <=( a884a ) or ( a885a );
 a5877a <=( a886a ) or ( a5876a );
 a5878a <=( a5877a ) or ( a5872a );
 a5881a <=( a882a ) or ( a883a );
 a5885a <=( a879a ) or ( a880a );
 a5886a <=( a881a ) or ( a5885a );
 a5887a <=( a5886a ) or ( a5881a );
 a5888a <=( a5887a ) or ( a5878a );
 a5889a <=( a5888a ) or ( a5869a );
 a5890a <=( a5889a ) or ( a5850a );
 a5891a <=( a5890a ) or ( a5811a );
 a5894a <=( a877a ) or ( a878a );
 a5898a <=( a874a ) or ( a875a );
 a5899a <=( a876a ) or ( a5898a );
 a5900a <=( a5899a ) or ( a5894a );
 a5903a <=( a872a ) or ( a873a );
 a5907a <=( a869a ) or ( a870a );
 a5908a <=( a871a ) or ( a5907a );
 a5909a <=( a5908a ) or ( a5903a );
 a5910a <=( a5909a ) or ( a5900a );
 a5913a <=( a867a ) or ( a868a );
 a5917a <=( a864a ) or ( a865a );
 a5918a <=( a866a ) or ( a5917a );
 a5919a <=( a5918a ) or ( a5913a );
 a5922a <=( a862a ) or ( a863a );
 a5926a <=( a859a ) or ( a860a );
 a5927a <=( a861a ) or ( a5926a );
 a5928a <=( a5927a ) or ( a5922a );
 a5929a <=( a5928a ) or ( a5919a );
 a5930a <=( a5929a ) or ( a5910a );
 a5933a <=( a857a ) or ( a858a );
 a5937a <=( a854a ) or ( a855a );
 a5938a <=( a856a ) or ( a5937a );
 a5939a <=( a5938a ) or ( a5933a );
 a5942a <=( a852a ) or ( a853a );
 a5946a <=( a849a ) or ( a850a );
 a5947a <=( a851a ) or ( a5946a );
 a5948a <=( a5947a ) or ( a5942a );
 a5949a <=( a5948a ) or ( a5939a );
 a5952a <=( a847a ) or ( a848a );
 a5956a <=( a844a ) or ( a845a );
 a5957a <=( a846a ) or ( a5956a );
 a5958a <=( a5957a ) or ( a5952a );
 a5961a <=( a842a ) or ( a843a );
 a5965a <=( a839a ) or ( a840a );
 a5966a <=( a841a ) or ( a5965a );
 a5967a <=( a5966a ) or ( a5961a );
 a5968a <=( a5967a ) or ( a5958a );
 a5969a <=( a5968a ) or ( a5949a );
 a5970a <=( a5969a ) or ( a5930a );
 a5973a <=( a837a ) or ( a838a );
 a5977a <=( a834a ) or ( a835a );
 a5978a <=( a836a ) or ( a5977a );
 a5979a <=( a5978a ) or ( a5973a );
 a5982a <=( a832a ) or ( a833a );
 a5986a <=( a829a ) or ( a830a );
 a5987a <=( a831a ) or ( a5986a );
 a5988a <=( a5987a ) or ( a5982a );
 a5989a <=( a5988a ) or ( a5979a );
 a5992a <=( a827a ) or ( a828a );
 a5996a <=( a824a ) or ( a825a );
 a5997a <=( a826a ) or ( a5996a );
 a5998a <=( a5997a ) or ( a5992a );
 a6001a <=( a822a ) or ( a823a );
 a6005a <=( a819a ) or ( a820a );
 a6006a <=( a821a ) or ( a6005a );
 a6007a <=( a6006a ) or ( a6001a );
 a6008a <=( a6007a ) or ( a5998a );
 a6009a <=( a6008a ) or ( a5989a );
 a6012a <=( a817a ) or ( a818a );
 a6016a <=( a814a ) or ( a815a );
 a6017a <=( a816a ) or ( a6016a );
 a6018a <=( a6017a ) or ( a6012a );
 a6021a <=( a812a ) or ( a813a );
 a6025a <=( a809a ) or ( a810a );
 a6026a <=( a811a ) or ( a6025a );
 a6027a <=( a6026a ) or ( a6021a );
 a6028a <=( a6027a ) or ( a6018a );
 a6031a <=( a807a ) or ( a808a );
 a6035a <=( a804a ) or ( a805a );
 a6036a <=( a806a ) or ( a6035a );
 a6037a <=( a6036a ) or ( a6031a );
 a6040a <=( a802a ) or ( a803a );
 a6044a <=( a799a ) or ( a800a );
 a6045a <=( a801a ) or ( a6044a );
 a6046a <=( a6045a ) or ( a6040a );
 a6047a <=( a6046a ) or ( a6037a );
 a6048a <=( a6047a ) or ( a6028a );
 a6049a <=( a6048a ) or ( a6009a );
 a6050a <=( a6049a ) or ( a5970a );
 a6051a <=( a6050a ) or ( a5891a );
 a6054a <=( a797a ) or ( a798a );
 a6058a <=( a794a ) or ( a795a );
 a6059a <=( a796a ) or ( a6058a );
 a6060a <=( a6059a ) or ( a6054a );
 a6063a <=( a792a ) or ( a793a );
 a6067a <=( a789a ) or ( a790a );
 a6068a <=( a791a ) or ( a6067a );
 a6069a <=( a6068a ) or ( a6063a );
 a6070a <=( a6069a ) or ( a6060a );
 a6073a <=( a787a ) or ( a788a );
 a6077a <=( a784a ) or ( a785a );
 a6078a <=( a786a ) or ( a6077a );
 a6079a <=( a6078a ) or ( a6073a );
 a6082a <=( a782a ) or ( a783a );
 a6086a <=( a779a ) or ( a780a );
 a6087a <=( a781a ) or ( a6086a );
 a6088a <=( a6087a ) or ( a6082a );
 a6089a <=( a6088a ) or ( a6079a );
 a6090a <=( a6089a ) or ( a6070a );
 a6093a <=( a777a ) or ( a778a );
 a6097a <=( a774a ) or ( a775a );
 a6098a <=( a776a ) or ( a6097a );
 a6099a <=( a6098a ) or ( a6093a );
 a6102a <=( a772a ) or ( a773a );
 a6106a <=( a769a ) or ( a770a );
 a6107a <=( a771a ) or ( a6106a );
 a6108a <=( a6107a ) or ( a6102a );
 a6109a <=( a6108a ) or ( a6099a );
 a6112a <=( a767a ) or ( a768a );
 a6116a <=( a764a ) or ( a765a );
 a6117a <=( a766a ) or ( a6116a );
 a6118a <=( a6117a ) or ( a6112a );
 a6121a <=( a762a ) or ( a763a );
 a6125a <=( a759a ) or ( a760a );
 a6126a <=( a761a ) or ( a6125a );
 a6127a <=( a6126a ) or ( a6121a );
 a6128a <=( a6127a ) or ( a6118a );
 a6129a <=( a6128a ) or ( a6109a );
 a6130a <=( a6129a ) or ( a6090a );
 a6133a <=( a757a ) or ( a758a );
 a6137a <=( a754a ) or ( a755a );
 a6138a <=( a756a ) or ( a6137a );
 a6139a <=( a6138a ) or ( a6133a );
 a6142a <=( a752a ) or ( a753a );
 a6146a <=( a749a ) or ( a750a );
 a6147a <=( a751a ) or ( a6146a );
 a6148a <=( a6147a ) or ( a6142a );
 a6149a <=( a6148a ) or ( a6139a );
 a6152a <=( a747a ) or ( a748a );
 a6156a <=( a744a ) or ( a745a );
 a6157a <=( a746a ) or ( a6156a );
 a6158a <=( a6157a ) or ( a6152a );
 a6161a <=( a742a ) or ( a743a );
 a6165a <=( a739a ) or ( a740a );
 a6166a <=( a741a ) or ( a6165a );
 a6167a <=( a6166a ) or ( a6161a );
 a6168a <=( a6167a ) or ( a6158a );
 a6169a <=( a6168a ) or ( a6149a );
 a6172a <=( a737a ) or ( a738a );
 a6176a <=( a734a ) or ( a735a );
 a6177a <=( a736a ) or ( a6176a );
 a6178a <=( a6177a ) or ( a6172a );
 a6181a <=( a732a ) or ( a733a );
 a6185a <=( a729a ) or ( a730a );
 a6186a <=( a731a ) or ( a6185a );
 a6187a <=( a6186a ) or ( a6181a );
 a6188a <=( a6187a ) or ( a6178a );
 a6191a <=( a727a ) or ( a728a );
 a6195a <=( a724a ) or ( a725a );
 a6196a <=( a726a ) or ( a6195a );
 a6197a <=( a6196a ) or ( a6191a );
 a6200a <=( a722a ) or ( a723a );
 a6204a <=( a719a ) or ( a720a );
 a6205a <=( a721a ) or ( a6204a );
 a6206a <=( a6205a ) or ( a6200a );
 a6207a <=( a6206a ) or ( a6197a );
 a6208a <=( a6207a ) or ( a6188a );
 a6209a <=( a6208a ) or ( a6169a );
 a6210a <=( a6209a ) or ( a6130a );
 a6213a <=( a717a ) or ( a718a );
 a6217a <=( a714a ) or ( a715a );
 a6218a <=( a716a ) or ( a6217a );
 a6219a <=( a6218a ) or ( a6213a );
 a6222a <=( a712a ) or ( a713a );
 a6226a <=( a709a ) or ( a710a );
 a6227a <=( a711a ) or ( a6226a );
 a6228a <=( a6227a ) or ( a6222a );
 a6229a <=( a6228a ) or ( a6219a );
 a6232a <=( a707a ) or ( a708a );
 a6236a <=( a704a ) or ( a705a );
 a6237a <=( a706a ) or ( a6236a );
 a6238a <=( a6237a ) or ( a6232a );
 a6241a <=( a702a ) or ( a703a );
 a6245a <=( a699a ) or ( a700a );
 a6246a <=( a701a ) or ( a6245a );
 a6247a <=( a6246a ) or ( a6241a );
 a6248a <=( a6247a ) or ( a6238a );
 a6249a <=( a6248a ) or ( a6229a );
 a6252a <=( a697a ) or ( a698a );
 a6256a <=( a694a ) or ( a695a );
 a6257a <=( a696a ) or ( a6256a );
 a6258a <=( a6257a ) or ( a6252a );
 a6261a <=( a692a ) or ( a693a );
 a6265a <=( a689a ) or ( a690a );
 a6266a <=( a691a ) or ( a6265a );
 a6267a <=( a6266a ) or ( a6261a );
 a6268a <=( a6267a ) or ( a6258a );
 a6271a <=( a687a ) or ( a688a );
 a6275a <=( a684a ) or ( a685a );
 a6276a <=( a686a ) or ( a6275a );
 a6277a <=( a6276a ) or ( a6271a );
 a6280a <=( a682a ) or ( a683a );
 a6284a <=( a679a ) or ( a680a );
 a6285a <=( a681a ) or ( a6284a );
 a6286a <=( a6285a ) or ( a6280a );
 a6287a <=( a6286a ) or ( a6277a );
 a6288a <=( a6287a ) or ( a6268a );
 a6289a <=( a6288a ) or ( a6249a );
 a6292a <=( a677a ) or ( a678a );
 a6296a <=( a674a ) or ( a675a );
 a6297a <=( a676a ) or ( a6296a );
 a6298a <=( a6297a ) or ( a6292a );
 a6301a <=( a672a ) or ( a673a );
 a6305a <=( a669a ) or ( a670a );
 a6306a <=( a671a ) or ( a6305a );
 a6307a <=( a6306a ) or ( a6301a );
 a6308a <=( a6307a ) or ( a6298a );
 a6311a <=( a667a ) or ( a668a );
 a6315a <=( a664a ) or ( a665a );
 a6316a <=( a666a ) or ( a6315a );
 a6317a <=( a6316a ) or ( a6311a );
 a6320a <=( a662a ) or ( a663a );
 a6324a <=( a659a ) or ( a660a );
 a6325a <=( a661a ) or ( a6324a );
 a6326a <=( a6325a ) or ( a6320a );
 a6327a <=( a6326a ) or ( a6317a );
 a6328a <=( a6327a ) or ( a6308a );
 a6331a <=( a657a ) or ( a658a );
 a6335a <=( a654a ) or ( a655a );
 a6336a <=( a656a ) or ( a6335a );
 a6337a <=( a6336a ) or ( a6331a );
 a6340a <=( a652a ) or ( a653a );
 a6344a <=( a649a ) or ( a650a );
 a6345a <=( a651a ) or ( a6344a );
 a6346a <=( a6345a ) or ( a6340a );
 a6347a <=( a6346a ) or ( a6337a );
 a6350a <=( a647a ) or ( a648a );
 a6354a <=( a644a ) or ( a645a );
 a6355a <=( a646a ) or ( a6354a );
 a6356a <=( a6355a ) or ( a6350a );
 a6359a <=( a642a ) or ( a643a );
 a6363a <=( a639a ) or ( a640a );
 a6364a <=( a641a ) or ( a6363a );
 a6365a <=( a6364a ) or ( a6359a );
 a6366a <=( a6365a ) or ( a6356a );
 a6367a <=( a6366a ) or ( a6347a );
 a6368a <=( a6367a ) or ( a6328a );
 a6369a <=( a6368a ) or ( a6289a );
 a6370a <=( a6369a ) or ( a6210a );
 a6371a <=( a6370a ) or ( a6051a );
 a6372a <=( a6371a ) or ( a5734a );
 a6375a <=( a637a ) or ( a638a );
 a6378a <=( a635a ) or ( a636a );
 a6379a <=( a6378a ) or ( a6375a );
 a6382a <=( a633a ) or ( a634a );
 a6386a <=( a630a ) or ( a631a );
 a6387a <=( a632a ) or ( a6386a );
 a6388a <=( a6387a ) or ( a6382a );
 a6389a <=( a6388a ) or ( a6379a );
 a6392a <=( a628a ) or ( a629a );
 a6396a <=( a625a ) or ( a626a );
 a6397a <=( a627a ) or ( a6396a );
 a6398a <=( a6397a ) or ( a6392a );
 a6401a <=( a623a ) or ( a624a );
 a6405a <=( a620a ) or ( a621a );
 a6406a <=( a622a ) or ( a6405a );
 a6407a <=( a6406a ) or ( a6401a );
 a6408a <=( a6407a ) or ( a6398a );
 a6409a <=( a6408a ) or ( a6389a );
 a6412a <=( a618a ) or ( a619a );
 a6416a <=( a615a ) or ( a616a );
 a6417a <=( a617a ) or ( a6416a );
 a6418a <=( a6417a ) or ( a6412a );
 a6421a <=( a613a ) or ( a614a );
 a6425a <=( a610a ) or ( a611a );
 a6426a <=( a612a ) or ( a6425a );
 a6427a <=( a6426a ) or ( a6421a );
 a6428a <=( a6427a ) or ( a6418a );
 a6431a <=( a608a ) or ( a609a );
 a6435a <=( a605a ) or ( a606a );
 a6436a <=( a607a ) or ( a6435a );
 a6437a <=( a6436a ) or ( a6431a );
 a6440a <=( a603a ) or ( a604a );
 a6444a <=( a600a ) or ( a601a );
 a6445a <=( a602a ) or ( a6444a );
 a6446a <=( a6445a ) or ( a6440a );
 a6447a <=( a6446a ) or ( a6437a );
 a6448a <=( a6447a ) or ( a6428a );
 a6449a <=( a6448a ) or ( a6409a );
 a6452a <=( a598a ) or ( a599a );
 a6456a <=( a595a ) or ( a596a );
 a6457a <=( a597a ) or ( a6456a );
 a6458a <=( a6457a ) or ( a6452a );
 a6461a <=( a593a ) or ( a594a );
 a6465a <=( a590a ) or ( a591a );
 a6466a <=( a592a ) or ( a6465a );
 a6467a <=( a6466a ) or ( a6461a );
 a6468a <=( a6467a ) or ( a6458a );
 a6471a <=( a588a ) or ( a589a );
 a6475a <=( a585a ) or ( a586a );
 a6476a <=( a587a ) or ( a6475a );
 a6477a <=( a6476a ) or ( a6471a );
 a6480a <=( a583a ) or ( a584a );
 a6484a <=( a580a ) or ( a581a );
 a6485a <=( a582a ) or ( a6484a );
 a6486a <=( a6485a ) or ( a6480a );
 a6487a <=( a6486a ) or ( a6477a );
 a6488a <=( a6487a ) or ( a6468a );
 a6491a <=( a578a ) or ( a579a );
 a6495a <=( a575a ) or ( a576a );
 a6496a <=( a577a ) or ( a6495a );
 a6497a <=( a6496a ) or ( a6491a );
 a6500a <=( a573a ) or ( a574a );
 a6504a <=( a570a ) or ( a571a );
 a6505a <=( a572a ) or ( a6504a );
 a6506a <=( a6505a ) or ( a6500a );
 a6507a <=( a6506a ) or ( a6497a );
 a6510a <=( a568a ) or ( a569a );
 a6514a <=( a565a ) or ( a566a );
 a6515a <=( a567a ) or ( a6514a );
 a6516a <=( a6515a ) or ( a6510a );
 a6519a <=( a563a ) or ( a564a );
 a6523a <=( a560a ) or ( a561a );
 a6524a <=( a562a ) or ( a6523a );
 a6525a <=( a6524a ) or ( a6519a );
 a6526a <=( a6525a ) or ( a6516a );
 a6527a <=( a6526a ) or ( a6507a );
 a6528a <=( a6527a ) or ( a6488a );
 a6529a <=( a6528a ) or ( a6449a );
 a6532a <=( a558a ) or ( a559a );
 a6536a <=( a555a ) or ( a556a );
 a6537a <=( a557a ) or ( a6536a );
 a6538a <=( a6537a ) or ( a6532a );
 a6541a <=( a553a ) or ( a554a );
 a6545a <=( a550a ) or ( a551a );
 a6546a <=( a552a ) or ( a6545a );
 a6547a <=( a6546a ) or ( a6541a );
 a6548a <=( a6547a ) or ( a6538a );
 a6551a <=( a548a ) or ( a549a );
 a6555a <=( a545a ) or ( a546a );
 a6556a <=( a547a ) or ( a6555a );
 a6557a <=( a6556a ) or ( a6551a );
 a6560a <=( a543a ) or ( a544a );
 a6564a <=( a540a ) or ( a541a );
 a6565a <=( a542a ) or ( a6564a );
 a6566a <=( a6565a ) or ( a6560a );
 a6567a <=( a6566a ) or ( a6557a );
 a6568a <=( a6567a ) or ( a6548a );
 a6571a <=( a538a ) or ( a539a );
 a6575a <=( a535a ) or ( a536a );
 a6576a <=( a537a ) or ( a6575a );
 a6577a <=( a6576a ) or ( a6571a );
 a6580a <=( a533a ) or ( a534a );
 a6584a <=( a530a ) or ( a531a );
 a6585a <=( a532a ) or ( a6584a );
 a6586a <=( a6585a ) or ( a6580a );
 a6587a <=( a6586a ) or ( a6577a );
 a6590a <=( a528a ) or ( a529a );
 a6594a <=( a525a ) or ( a526a );
 a6595a <=( a527a ) or ( a6594a );
 a6596a <=( a6595a ) or ( a6590a );
 a6599a <=( a523a ) or ( a524a );
 a6603a <=( a520a ) or ( a521a );
 a6604a <=( a522a ) or ( a6603a );
 a6605a <=( a6604a ) or ( a6599a );
 a6606a <=( a6605a ) or ( a6596a );
 a6607a <=( a6606a ) or ( a6587a );
 a6608a <=( a6607a ) or ( a6568a );
 a6611a <=( a518a ) or ( a519a );
 a6615a <=( a515a ) or ( a516a );
 a6616a <=( a517a ) or ( a6615a );
 a6617a <=( a6616a ) or ( a6611a );
 a6620a <=( a513a ) or ( a514a );
 a6624a <=( a510a ) or ( a511a );
 a6625a <=( a512a ) or ( a6624a );
 a6626a <=( a6625a ) or ( a6620a );
 a6627a <=( a6626a ) or ( a6617a );
 a6630a <=( a508a ) or ( a509a );
 a6634a <=( a505a ) or ( a506a );
 a6635a <=( a507a ) or ( a6634a );
 a6636a <=( a6635a ) or ( a6630a );
 a6639a <=( a503a ) or ( a504a );
 a6643a <=( a500a ) or ( a501a );
 a6644a <=( a502a ) or ( a6643a );
 a6645a <=( a6644a ) or ( a6639a );
 a6646a <=( a6645a ) or ( a6636a );
 a6647a <=( a6646a ) or ( a6627a );
 a6650a <=( a498a ) or ( a499a );
 a6654a <=( a495a ) or ( a496a );
 a6655a <=( a497a ) or ( a6654a );
 a6656a <=( a6655a ) or ( a6650a );
 a6659a <=( a493a ) or ( a494a );
 a6663a <=( a490a ) or ( a491a );
 a6664a <=( a492a ) or ( a6663a );
 a6665a <=( a6664a ) or ( a6659a );
 a6666a <=( a6665a ) or ( a6656a );
 a6669a <=( a488a ) or ( a489a );
 a6673a <=( a485a ) or ( a486a );
 a6674a <=( a487a ) or ( a6673a );
 a6675a <=( a6674a ) or ( a6669a );
 a6678a <=( a483a ) or ( a484a );
 a6682a <=( a480a ) or ( a481a );
 a6683a <=( a482a ) or ( a6682a );
 a6684a <=( a6683a ) or ( a6678a );
 a6685a <=( a6684a ) or ( a6675a );
 a6686a <=( a6685a ) or ( a6666a );
 a6687a <=( a6686a ) or ( a6647a );
 a6688a <=( a6687a ) or ( a6608a );
 a6689a <=( a6688a ) or ( a6529a );
 a6692a <=( a478a ) or ( a479a );
 a6696a <=( a475a ) or ( a476a );
 a6697a <=( a477a ) or ( a6696a );
 a6698a <=( a6697a ) or ( a6692a );
 a6701a <=( a473a ) or ( a474a );
 a6705a <=( a470a ) or ( a471a );
 a6706a <=( a472a ) or ( a6705a );
 a6707a <=( a6706a ) or ( a6701a );
 a6708a <=( a6707a ) or ( a6698a );
 a6711a <=( a468a ) or ( a469a );
 a6715a <=( a465a ) or ( a466a );
 a6716a <=( a467a ) or ( a6715a );
 a6717a <=( a6716a ) or ( a6711a );
 a6720a <=( a463a ) or ( a464a );
 a6724a <=( a460a ) or ( a461a );
 a6725a <=( a462a ) or ( a6724a );
 a6726a <=( a6725a ) or ( a6720a );
 a6727a <=( a6726a ) or ( a6717a );
 a6728a <=( a6727a ) or ( a6708a );
 a6731a <=( a458a ) or ( a459a );
 a6735a <=( a455a ) or ( a456a );
 a6736a <=( a457a ) or ( a6735a );
 a6737a <=( a6736a ) or ( a6731a );
 a6740a <=( a453a ) or ( a454a );
 a6744a <=( a450a ) or ( a451a );
 a6745a <=( a452a ) or ( a6744a );
 a6746a <=( a6745a ) or ( a6740a );
 a6747a <=( a6746a ) or ( a6737a );
 a6750a <=( a448a ) or ( a449a );
 a6754a <=( a445a ) or ( a446a );
 a6755a <=( a447a ) or ( a6754a );
 a6756a <=( a6755a ) or ( a6750a );
 a6759a <=( a443a ) or ( a444a );
 a6763a <=( a440a ) or ( a441a );
 a6764a <=( a442a ) or ( a6763a );
 a6765a <=( a6764a ) or ( a6759a );
 a6766a <=( a6765a ) or ( a6756a );
 a6767a <=( a6766a ) or ( a6747a );
 a6768a <=( a6767a ) or ( a6728a );
 a6771a <=( a438a ) or ( a439a );
 a6775a <=( a435a ) or ( a436a );
 a6776a <=( a437a ) or ( a6775a );
 a6777a <=( a6776a ) or ( a6771a );
 a6780a <=( a433a ) or ( a434a );
 a6784a <=( a430a ) or ( a431a );
 a6785a <=( a432a ) or ( a6784a );
 a6786a <=( a6785a ) or ( a6780a );
 a6787a <=( a6786a ) or ( a6777a );
 a6790a <=( a428a ) or ( a429a );
 a6794a <=( a425a ) or ( a426a );
 a6795a <=( a427a ) or ( a6794a );
 a6796a <=( a6795a ) or ( a6790a );
 a6799a <=( a423a ) or ( a424a );
 a6803a <=( a420a ) or ( a421a );
 a6804a <=( a422a ) or ( a6803a );
 a6805a <=( a6804a ) or ( a6799a );
 a6806a <=( a6805a ) or ( a6796a );
 a6807a <=( a6806a ) or ( a6787a );
 a6810a <=( a418a ) or ( a419a );
 a6814a <=( a415a ) or ( a416a );
 a6815a <=( a417a ) or ( a6814a );
 a6816a <=( a6815a ) or ( a6810a );
 a6819a <=( a413a ) or ( a414a );
 a6823a <=( a410a ) or ( a411a );
 a6824a <=( a412a ) or ( a6823a );
 a6825a <=( a6824a ) or ( a6819a );
 a6826a <=( a6825a ) or ( a6816a );
 a6829a <=( a408a ) or ( a409a );
 a6833a <=( a405a ) or ( a406a );
 a6834a <=( a407a ) or ( a6833a );
 a6835a <=( a6834a ) or ( a6829a );
 a6838a <=( a403a ) or ( a404a );
 a6842a <=( a400a ) or ( a401a );
 a6843a <=( a402a ) or ( a6842a );
 a6844a <=( a6843a ) or ( a6838a );
 a6845a <=( a6844a ) or ( a6835a );
 a6846a <=( a6845a ) or ( a6826a );
 a6847a <=( a6846a ) or ( a6807a );
 a6848a <=( a6847a ) or ( a6768a );
 a6851a <=( a398a ) or ( a399a );
 a6855a <=( a395a ) or ( a396a );
 a6856a <=( a397a ) or ( a6855a );
 a6857a <=( a6856a ) or ( a6851a );
 a6860a <=( a393a ) or ( a394a );
 a6864a <=( a390a ) or ( a391a );
 a6865a <=( a392a ) or ( a6864a );
 a6866a <=( a6865a ) or ( a6860a );
 a6867a <=( a6866a ) or ( a6857a );
 a6870a <=( a388a ) or ( a389a );
 a6874a <=( a385a ) or ( a386a );
 a6875a <=( a387a ) or ( a6874a );
 a6876a <=( a6875a ) or ( a6870a );
 a6879a <=( a383a ) or ( a384a );
 a6883a <=( a380a ) or ( a381a );
 a6884a <=( a382a ) or ( a6883a );
 a6885a <=( a6884a ) or ( a6879a );
 a6886a <=( a6885a ) or ( a6876a );
 a6887a <=( a6886a ) or ( a6867a );
 a6890a <=( a378a ) or ( a379a );
 a6894a <=( a375a ) or ( a376a );
 a6895a <=( a377a ) or ( a6894a );
 a6896a <=( a6895a ) or ( a6890a );
 a6899a <=( a373a ) or ( a374a );
 a6903a <=( a370a ) or ( a371a );
 a6904a <=( a372a ) or ( a6903a );
 a6905a <=( a6904a ) or ( a6899a );
 a6906a <=( a6905a ) or ( a6896a );
 a6909a <=( a368a ) or ( a369a );
 a6913a <=( a365a ) or ( a366a );
 a6914a <=( a367a ) or ( a6913a );
 a6915a <=( a6914a ) or ( a6909a );
 a6918a <=( a363a ) or ( a364a );
 a6922a <=( a360a ) or ( a361a );
 a6923a <=( a362a ) or ( a6922a );
 a6924a <=( a6923a ) or ( a6918a );
 a6925a <=( a6924a ) or ( a6915a );
 a6926a <=( a6925a ) or ( a6906a );
 a6927a <=( a6926a ) or ( a6887a );
 a6930a <=( a358a ) or ( a359a );
 a6934a <=( a355a ) or ( a356a );
 a6935a <=( a357a ) or ( a6934a );
 a6936a <=( a6935a ) or ( a6930a );
 a6939a <=( a353a ) or ( a354a );
 a6943a <=( a350a ) or ( a351a );
 a6944a <=( a352a ) or ( a6943a );
 a6945a <=( a6944a ) or ( a6939a );
 a6946a <=( a6945a ) or ( a6936a );
 a6949a <=( a348a ) or ( a349a );
 a6953a <=( a345a ) or ( a346a );
 a6954a <=( a347a ) or ( a6953a );
 a6955a <=( a6954a ) or ( a6949a );
 a6958a <=( a343a ) or ( a344a );
 a6962a <=( a340a ) or ( a341a );
 a6963a <=( a342a ) or ( a6962a );
 a6964a <=( a6963a ) or ( a6958a );
 a6965a <=( a6964a ) or ( a6955a );
 a6966a <=( a6965a ) or ( a6946a );
 a6969a <=( a338a ) or ( a339a );
 a6973a <=( a335a ) or ( a336a );
 a6974a <=( a337a ) or ( a6973a );
 a6975a <=( a6974a ) or ( a6969a );
 a6978a <=( a333a ) or ( a334a );
 a6982a <=( a330a ) or ( a331a );
 a6983a <=( a332a ) or ( a6982a );
 a6984a <=( a6983a ) or ( a6978a );
 a6985a <=( a6984a ) or ( a6975a );
 a6988a <=( a328a ) or ( a329a );
 a6992a <=( a325a ) or ( a326a );
 a6993a <=( a327a ) or ( a6992a );
 a6994a <=( a6993a ) or ( a6988a );
 a6997a <=( a323a ) or ( a324a );
 a7001a <=( a320a ) or ( a321a );
 a7002a <=( a322a ) or ( a7001a );
 a7003a <=( a7002a ) or ( a6997a );
 a7004a <=( a7003a ) or ( a6994a );
 a7005a <=( a7004a ) or ( a6985a );
 a7006a <=( a7005a ) or ( a6966a );
 a7007a <=( a7006a ) or ( a6927a );
 a7008a <=( a7007a ) or ( a6848a );
 a7009a <=( a7008a ) or ( a6689a );
 a7012a <=( a318a ) or ( a319a );
 a7015a <=( a316a ) or ( a317a );
 a7016a <=( a7015a ) or ( a7012a );
 a7019a <=( a314a ) or ( a315a );
 a7023a <=( a311a ) or ( a312a );
 a7024a <=( a313a ) or ( a7023a );
 a7025a <=( a7024a ) or ( a7019a );
 a7026a <=( a7025a ) or ( a7016a );
 a7029a <=( a309a ) or ( a310a );
 a7033a <=( a306a ) or ( a307a );
 a7034a <=( a308a ) or ( a7033a );
 a7035a <=( a7034a ) or ( a7029a );
 a7038a <=( a304a ) or ( a305a );
 a7042a <=( a301a ) or ( a302a );
 a7043a <=( a303a ) or ( a7042a );
 a7044a <=( a7043a ) or ( a7038a );
 a7045a <=( a7044a ) or ( a7035a );
 a7046a <=( a7045a ) or ( a7026a );
 a7049a <=( a299a ) or ( a300a );
 a7053a <=( a296a ) or ( a297a );
 a7054a <=( a298a ) or ( a7053a );
 a7055a <=( a7054a ) or ( a7049a );
 a7058a <=( a294a ) or ( a295a );
 a7062a <=( a291a ) or ( a292a );
 a7063a <=( a293a ) or ( a7062a );
 a7064a <=( a7063a ) or ( a7058a );
 a7065a <=( a7064a ) or ( a7055a );
 a7068a <=( a289a ) or ( a290a );
 a7072a <=( a286a ) or ( a287a );
 a7073a <=( a288a ) or ( a7072a );
 a7074a <=( a7073a ) or ( a7068a );
 a7077a <=( a284a ) or ( a285a );
 a7081a <=( a281a ) or ( a282a );
 a7082a <=( a283a ) or ( a7081a );
 a7083a <=( a7082a ) or ( a7077a );
 a7084a <=( a7083a ) or ( a7074a );
 a7085a <=( a7084a ) or ( a7065a );
 a7086a <=( a7085a ) or ( a7046a );
 a7089a <=( a279a ) or ( a280a );
 a7093a <=( a276a ) or ( a277a );
 a7094a <=( a278a ) or ( a7093a );
 a7095a <=( a7094a ) or ( a7089a );
 a7098a <=( a274a ) or ( a275a );
 a7102a <=( a271a ) or ( a272a );
 a7103a <=( a273a ) or ( a7102a );
 a7104a <=( a7103a ) or ( a7098a );
 a7105a <=( a7104a ) or ( a7095a );
 a7108a <=( a269a ) or ( a270a );
 a7112a <=( a266a ) or ( a267a );
 a7113a <=( a268a ) or ( a7112a );
 a7114a <=( a7113a ) or ( a7108a );
 a7117a <=( a264a ) or ( a265a );
 a7121a <=( a261a ) or ( a262a );
 a7122a <=( a263a ) or ( a7121a );
 a7123a <=( a7122a ) or ( a7117a );
 a7124a <=( a7123a ) or ( a7114a );
 a7125a <=( a7124a ) or ( a7105a );
 a7128a <=( a259a ) or ( a260a );
 a7132a <=( a256a ) or ( a257a );
 a7133a <=( a258a ) or ( a7132a );
 a7134a <=( a7133a ) or ( a7128a );
 a7137a <=( a254a ) or ( a255a );
 a7141a <=( a251a ) or ( a252a );
 a7142a <=( a253a ) or ( a7141a );
 a7143a <=( a7142a ) or ( a7137a );
 a7144a <=( a7143a ) or ( a7134a );
 a7147a <=( a249a ) or ( a250a );
 a7151a <=( a246a ) or ( a247a );
 a7152a <=( a248a ) or ( a7151a );
 a7153a <=( a7152a ) or ( a7147a );
 a7156a <=( a244a ) or ( a245a );
 a7160a <=( a241a ) or ( a242a );
 a7161a <=( a243a ) or ( a7160a );
 a7162a <=( a7161a ) or ( a7156a );
 a7163a <=( a7162a ) or ( a7153a );
 a7164a <=( a7163a ) or ( a7144a );
 a7165a <=( a7164a ) or ( a7125a );
 a7166a <=( a7165a ) or ( a7086a );
 a7169a <=( a239a ) or ( a240a );
 a7173a <=( a236a ) or ( a237a );
 a7174a <=( a238a ) or ( a7173a );
 a7175a <=( a7174a ) or ( a7169a );
 a7178a <=( a234a ) or ( a235a );
 a7182a <=( a231a ) or ( a232a );
 a7183a <=( a233a ) or ( a7182a );
 a7184a <=( a7183a ) or ( a7178a );
 a7185a <=( a7184a ) or ( a7175a );
 a7188a <=( a229a ) or ( a230a );
 a7192a <=( a226a ) or ( a227a );
 a7193a <=( a228a ) or ( a7192a );
 a7194a <=( a7193a ) or ( a7188a );
 a7197a <=( a224a ) or ( a225a );
 a7201a <=( a221a ) or ( a222a );
 a7202a <=( a223a ) or ( a7201a );
 a7203a <=( a7202a ) or ( a7197a );
 a7204a <=( a7203a ) or ( a7194a );
 a7205a <=( a7204a ) or ( a7185a );
 a7208a <=( a219a ) or ( a220a );
 a7212a <=( a216a ) or ( a217a );
 a7213a <=( a218a ) or ( a7212a );
 a7214a <=( a7213a ) or ( a7208a );
 a7217a <=( a214a ) or ( a215a );
 a7221a <=( a211a ) or ( a212a );
 a7222a <=( a213a ) or ( a7221a );
 a7223a <=( a7222a ) or ( a7217a );
 a7224a <=( a7223a ) or ( a7214a );
 a7227a <=( a209a ) or ( a210a );
 a7231a <=( a206a ) or ( a207a );
 a7232a <=( a208a ) or ( a7231a );
 a7233a <=( a7232a ) or ( a7227a );
 a7236a <=( a204a ) or ( a205a );
 a7240a <=( a201a ) or ( a202a );
 a7241a <=( a203a ) or ( a7240a );
 a7242a <=( a7241a ) or ( a7236a );
 a7243a <=( a7242a ) or ( a7233a );
 a7244a <=( a7243a ) or ( a7224a );
 a7245a <=( a7244a ) or ( a7205a );
 a7248a <=( a199a ) or ( a200a );
 a7252a <=( a196a ) or ( a197a );
 a7253a <=( a198a ) or ( a7252a );
 a7254a <=( a7253a ) or ( a7248a );
 a7257a <=( a194a ) or ( a195a );
 a7261a <=( a191a ) or ( a192a );
 a7262a <=( a193a ) or ( a7261a );
 a7263a <=( a7262a ) or ( a7257a );
 a7264a <=( a7263a ) or ( a7254a );
 a7267a <=( a189a ) or ( a190a );
 a7271a <=( a186a ) or ( a187a );
 a7272a <=( a188a ) or ( a7271a );
 a7273a <=( a7272a ) or ( a7267a );
 a7276a <=( a184a ) or ( a185a );
 a7280a <=( a181a ) or ( a182a );
 a7281a <=( a183a ) or ( a7280a );
 a7282a <=( a7281a ) or ( a7276a );
 a7283a <=( a7282a ) or ( a7273a );
 a7284a <=( a7283a ) or ( a7264a );
 a7287a <=( a179a ) or ( a180a );
 a7291a <=( a176a ) or ( a177a );
 a7292a <=( a178a ) or ( a7291a );
 a7293a <=( a7292a ) or ( a7287a );
 a7296a <=( a174a ) or ( a175a );
 a7300a <=( a171a ) or ( a172a );
 a7301a <=( a173a ) or ( a7300a );
 a7302a <=( a7301a ) or ( a7296a );
 a7303a <=( a7302a ) or ( a7293a );
 a7306a <=( a169a ) or ( a170a );
 a7310a <=( a166a ) or ( a167a );
 a7311a <=( a168a ) or ( a7310a );
 a7312a <=( a7311a ) or ( a7306a );
 a7315a <=( a164a ) or ( a165a );
 a7319a <=( a161a ) or ( a162a );
 a7320a <=( a163a ) or ( a7319a );
 a7321a <=( a7320a ) or ( a7315a );
 a7322a <=( a7321a ) or ( a7312a );
 a7323a <=( a7322a ) or ( a7303a );
 a7324a <=( a7323a ) or ( a7284a );
 a7325a <=( a7324a ) or ( a7245a );
 a7326a <=( a7325a ) or ( a7166a );
 a7329a <=( a159a ) or ( a160a );
 a7333a <=( a156a ) or ( a157a );
 a7334a <=( a158a ) or ( a7333a );
 a7335a <=( a7334a ) or ( a7329a );
 a7338a <=( a154a ) or ( a155a );
 a7342a <=( a151a ) or ( a152a );
 a7343a <=( a153a ) or ( a7342a );
 a7344a <=( a7343a ) or ( a7338a );
 a7345a <=( a7344a ) or ( a7335a );
 a7348a <=( a149a ) or ( a150a );
 a7352a <=( a146a ) or ( a147a );
 a7353a <=( a148a ) or ( a7352a );
 a7354a <=( a7353a ) or ( a7348a );
 a7357a <=( a144a ) or ( a145a );
 a7361a <=( a141a ) or ( a142a );
 a7362a <=( a143a ) or ( a7361a );
 a7363a <=( a7362a ) or ( a7357a );
 a7364a <=( a7363a ) or ( a7354a );
 a7365a <=( a7364a ) or ( a7345a );
 a7368a <=( a139a ) or ( a140a );
 a7372a <=( a136a ) or ( a137a );
 a7373a <=( a138a ) or ( a7372a );
 a7374a <=( a7373a ) or ( a7368a );
 a7377a <=( a134a ) or ( a135a );
 a7381a <=( a131a ) or ( a132a );
 a7382a <=( a133a ) or ( a7381a );
 a7383a <=( a7382a ) or ( a7377a );
 a7384a <=( a7383a ) or ( a7374a );
 a7387a <=( a129a ) or ( a130a );
 a7391a <=( a126a ) or ( a127a );
 a7392a <=( a128a ) or ( a7391a );
 a7393a <=( a7392a ) or ( a7387a );
 a7396a <=( a124a ) or ( a125a );
 a7400a <=( a121a ) or ( a122a );
 a7401a <=( a123a ) or ( a7400a );
 a7402a <=( a7401a ) or ( a7396a );
 a7403a <=( a7402a ) or ( a7393a );
 a7404a <=( a7403a ) or ( a7384a );
 a7405a <=( a7404a ) or ( a7365a );
 a7408a <=( a119a ) or ( a120a );
 a7412a <=( a116a ) or ( a117a );
 a7413a <=( a118a ) or ( a7412a );
 a7414a <=( a7413a ) or ( a7408a );
 a7417a <=( a114a ) or ( a115a );
 a7421a <=( a111a ) or ( a112a );
 a7422a <=( a113a ) or ( a7421a );
 a7423a <=( a7422a ) or ( a7417a );
 a7424a <=( a7423a ) or ( a7414a );
 a7427a <=( a109a ) or ( a110a );
 a7431a <=( a106a ) or ( a107a );
 a7432a <=( a108a ) or ( a7431a );
 a7433a <=( a7432a ) or ( a7427a );
 a7436a <=( a104a ) or ( a105a );
 a7440a <=( a101a ) or ( a102a );
 a7441a <=( a103a ) or ( a7440a );
 a7442a <=( a7441a ) or ( a7436a );
 a7443a <=( a7442a ) or ( a7433a );
 a7444a <=( a7443a ) or ( a7424a );
 a7447a <=( a99a ) or ( a100a );
 a7451a <=( a96a ) or ( a97a );
 a7452a <=( a98a ) or ( a7451a );
 a7453a <=( a7452a ) or ( a7447a );
 a7456a <=( a94a ) or ( a95a );
 a7460a <=( a91a ) or ( a92a );
 a7461a <=( a93a ) or ( a7460a );
 a7462a <=( a7461a ) or ( a7456a );
 a7463a <=( a7462a ) or ( a7453a );
 a7466a <=( a89a ) or ( a90a );
 a7470a <=( a86a ) or ( a87a );
 a7471a <=( a88a ) or ( a7470a );
 a7472a <=( a7471a ) or ( a7466a );
 a7475a <=( a84a ) or ( a85a );
 a7479a <=( a81a ) or ( a82a );
 a7480a <=( a83a ) or ( a7479a );
 a7481a <=( a7480a ) or ( a7475a );
 a7482a <=( a7481a ) or ( a7472a );
 a7483a <=( a7482a ) or ( a7463a );
 a7484a <=( a7483a ) or ( a7444a );
 a7485a <=( a7484a ) or ( a7405a );
 a7488a <=( a79a ) or ( a80a );
 a7492a <=( a76a ) or ( a77a );
 a7493a <=( a78a ) or ( a7492a );
 a7494a <=( a7493a ) or ( a7488a );
 a7497a <=( a74a ) or ( a75a );
 a7501a <=( a71a ) or ( a72a );
 a7502a <=( a73a ) or ( a7501a );
 a7503a <=( a7502a ) or ( a7497a );
 a7504a <=( a7503a ) or ( a7494a );
 a7507a <=( a69a ) or ( a70a );
 a7511a <=( a66a ) or ( a67a );
 a7512a <=( a68a ) or ( a7511a );
 a7513a <=( a7512a ) or ( a7507a );
 a7516a <=( a64a ) or ( a65a );
 a7520a <=( a61a ) or ( a62a );
 a7521a <=( a63a ) or ( a7520a );
 a7522a <=( a7521a ) or ( a7516a );
 a7523a <=( a7522a ) or ( a7513a );
 a7524a <=( a7523a ) or ( a7504a );
 a7527a <=( a59a ) or ( a60a );
 a7531a <=( a56a ) or ( a57a );
 a7532a <=( a58a ) or ( a7531a );
 a7533a <=( a7532a ) or ( a7527a );
 a7536a <=( a54a ) or ( a55a );
 a7540a <=( a51a ) or ( a52a );
 a7541a <=( a53a ) or ( a7540a );
 a7542a <=( a7541a ) or ( a7536a );
 a7543a <=( a7542a ) or ( a7533a );
 a7546a <=( a49a ) or ( a50a );
 a7550a <=( a46a ) or ( a47a );
 a7551a <=( a48a ) or ( a7550a );
 a7552a <=( a7551a ) or ( a7546a );
 a7555a <=( a44a ) or ( a45a );
 a7559a <=( a41a ) or ( a42a );
 a7560a <=( a43a ) or ( a7559a );
 a7561a <=( a7560a ) or ( a7555a );
 a7562a <=( a7561a ) or ( a7552a );
 a7563a <=( a7562a ) or ( a7543a );
 a7564a <=( a7563a ) or ( a7524a );
 a7567a <=( a39a ) or ( a40a );
 a7571a <=( a36a ) or ( a37a );
 a7572a <=( a38a ) or ( a7571a );
 a7573a <=( a7572a ) or ( a7567a );
 a7576a <=( a34a ) or ( a35a );
 a7580a <=( a31a ) or ( a32a );
 a7581a <=( a33a ) or ( a7580a );
 a7582a <=( a7581a ) or ( a7576a );
 a7583a <=( a7582a ) or ( a7573a );
 a7586a <=( a29a ) or ( a30a );
 a7590a <=( a26a ) or ( a27a );
 a7591a <=( a28a ) or ( a7590a );
 a7592a <=( a7591a ) or ( a7586a );
 a7595a <=( a24a ) or ( a25a );
 a7599a <=( a21a ) or ( a22a );
 a7600a <=( a23a ) or ( a7599a );
 a7601a <=( a7600a ) or ( a7595a );
 a7602a <=( a7601a ) or ( a7592a );
 a7603a <=( a7602a ) or ( a7583a );
 a7606a <=( a19a ) or ( a20a );
 a7610a <=( a16a ) or ( a17a );
 a7611a <=( a18a ) or ( a7610a );
 a7612a <=( a7611a ) or ( a7606a );
 a7615a <=( a14a ) or ( a15a );
 a7619a <=( a11a ) or ( a12a );
 a7620a <=( a13a ) or ( a7619a );
 a7621a <=( a7620a ) or ( a7615a );
 a7622a <=( a7621a ) or ( a7612a );
 a7625a <=( a9a ) or ( a10a );
 a7629a <=( a6a ) or ( a7a );
 a7630a <=( a8a ) or ( a7629a );
 a7631a <=( a7630a ) or ( a7625a );
 a7634a <=( a4a ) or ( a5a );
 a7638a <=( a1a ) or ( a2a );
 a7639a <=( a3a ) or ( a7638a );
 a7640a <=( a7639a ) or ( a7634a );
 a7641a <=( a7640a ) or ( a7631a );
 a7642a <=( a7641a ) or ( a7622a );
 a7643a <=( a7642a ) or ( a7603a );
 a7644a <=( a7643a ) or ( a7564a );
 a7645a <=( a7644a ) or ( a7485a );
 a7646a <=( a7645a ) or ( a7326a );
 a7647a <=( a7646a ) or ( a7009a );
 a7648a <=( a7647a ) or ( a6372a );
 a7652a <=( (not A202)  and  (not A201) );
 a7653a <=( A169  and  a7652a );
 a7657a <=( A268  and  A235 );
 a7658a <=( (not A203)  and  a7657a );
 a7662a <=( (not A200)  and  (not A199) );
 a7663a <=( A169  and  a7662a );
 a7667a <=( A268  and  A235 );
 a7668a <=( (not A202)  and  a7667a );
 a7672a <=( (not A166)  and  (not A167) );
 a7673a <=( (not A169)  and  a7672a );
 a7677a <=( A268  and  A235 );
 a7678a <=( A202  and  a7677a );
 a7682a <=( (not A168)  and  (not A169) );
 a7683a <=( (not A170)  and  a7682a );
 a7687a <=( A268  and  A235 );
 a7688a <=( A202  and  a7687a );
 a7692a <=( (not A201)  and  A166 );
 a7693a <=( A168  and  a7692a );
 a7696a <=( (not A203)  and  (not A202) );
 a7699a <=( A268  and  A235 );
 a7700a <=( a7699a  and  a7696a );
 a7704a <=( (not A199)  and  A166 );
 a7705a <=( A168  and  a7704a );
 a7708a <=( (not A202)  and  (not A200) );
 a7711a <=( A268  and  A235 );
 a7712a <=( a7711a  and  a7708a );
 a7716a <=( (not A201)  and  A167 );
 a7717a <=( A168  and  a7716a );
 a7720a <=( (not A203)  and  (not A202) );
 a7723a <=( A268  and  A235 );
 a7724a <=( a7723a  and  a7720a );
 a7728a <=( (not A199)  and  A167 );
 a7729a <=( A168  and  a7728a );
 a7732a <=( (not A202)  and  (not A200) );
 a7735a <=( A268  and  A235 );
 a7736a <=( a7735a  and  a7732a );
 a7740a <=( (not A202)  and  (not A201) );
 a7741a <=( A169  and  a7740a );
 a7744a <=( A235  and  (not A203) );
 a7747a <=( A267  and  A265 );
 a7748a <=( a7747a  and  a7744a );
 a7752a <=( (not A202)  and  (not A201) );
 a7753a <=( A169  and  a7752a );
 a7756a <=( A235  and  (not A203) );
 a7759a <=( A267  and  A266 );
 a7760a <=( a7759a  and  a7756a );
 a7764a <=( (not A202)  and  (not A201) );
 a7765a <=( A169  and  a7764a );
 a7768a <=( A232  and  (not A203) );
 a7771a <=( A268  and  A234 );
 a7772a <=( a7771a  and  a7768a );
 a7776a <=( (not A202)  and  (not A201) );
 a7777a <=( A169  and  a7776a );
 a7780a <=( A233  and  (not A203) );
 a7783a <=( A268  and  A234 );
 a7784a <=( a7783a  and  a7780a );
 a7788a <=( A200  and  A199 );
 a7789a <=( A169  and  a7788a );
 a7792a <=( (not A202)  and  (not A201) );
 a7795a <=( A268  and  A235 );
 a7796a <=( a7795a  and  a7792a );
 a7800a <=( (not A200)  and  (not A199) );
 a7801a <=( A169  and  a7800a );
 a7804a <=( A235  and  (not A202) );
 a7807a <=( A267  and  A265 );
 a7808a <=( a7807a  and  a7804a );
 a7812a <=( (not A200)  and  (not A199) );
 a7813a <=( A169  and  a7812a );
 a7816a <=( A235  and  (not A202) );
 a7819a <=( A267  and  A266 );
 a7820a <=( a7819a  and  a7816a );
 a7824a <=( (not A200)  and  (not A199) );
 a7825a <=( A169  and  a7824a );
 a7828a <=( A232  and  (not A202) );
 a7831a <=( A268  and  A234 );
 a7832a <=( a7831a  and  a7828a );
 a7836a <=( (not A200)  and  (not A199) );
 a7837a <=( A169  and  a7836a );
 a7840a <=( A233  and  (not A202) );
 a7843a <=( A268  and  A234 );
 a7844a <=( a7843a  and  a7840a );
 a7848a <=( (not A166)  and  (not A167) );
 a7849a <=( (not A169)  and  a7848a );
 a7852a <=( A235  and  A202 );
 a7855a <=( A267  and  A265 );
 a7856a <=( a7855a  and  a7852a );
 a7860a <=( (not A166)  and  (not A167) );
 a7861a <=( (not A169)  and  a7860a );
 a7864a <=( A235  and  A202 );
 a7867a <=( A267  and  A266 );
 a7868a <=( a7867a  and  a7864a );
 a7872a <=( (not A166)  and  (not A167) );
 a7873a <=( (not A169)  and  a7872a );
 a7876a <=( A232  and  A202 );
 a7879a <=( A268  and  A234 );
 a7880a <=( a7879a  and  a7876a );
 a7884a <=( (not A166)  and  (not A167) );
 a7885a <=( (not A169)  and  a7884a );
 a7888a <=( A233  and  A202 );
 a7891a <=( A268  and  A234 );
 a7892a <=( a7891a  and  a7888a );
 a7896a <=( (not A166)  and  (not A167) );
 a7897a <=( (not A169)  and  a7896a );
 a7900a <=( A201  and  A199 );
 a7903a <=( A268  and  A235 );
 a7904a <=( a7903a  and  a7900a );
 a7908a <=( (not A166)  and  (not A167) );
 a7909a <=( (not A169)  and  a7908a );
 a7912a <=( A201  and  A200 );
 a7915a <=( A268  and  A235 );
 a7916a <=( a7915a  and  a7912a );
 a7920a <=( A167  and  (not A168) );
 a7921a <=( (not A169)  and  a7920a );
 a7924a <=( A202  and  A166 );
 a7927a <=( A268  and  A235 );
 a7928a <=( a7927a  and  a7924a );
 a7932a <=( (not A168)  and  (not A169) );
 a7933a <=( (not A170)  and  a7932a );
 a7936a <=( A235  and  A202 );
 a7939a <=( A267  and  A265 );
 a7940a <=( a7939a  and  a7936a );
 a7944a <=( (not A168)  and  (not A169) );
 a7945a <=( (not A170)  and  a7944a );
 a7948a <=( A235  and  A202 );
 a7951a <=( A267  and  A266 );
 a7952a <=( a7951a  and  a7948a );
 a7956a <=( (not A168)  and  (not A169) );
 a7957a <=( (not A170)  and  a7956a );
 a7960a <=( A232  and  A202 );
 a7963a <=( A268  and  A234 );
 a7964a <=( a7963a  and  a7960a );
 a7968a <=( (not A168)  and  (not A169) );
 a7969a <=( (not A170)  and  a7968a );
 a7972a <=( A233  and  A202 );
 a7975a <=( A268  and  A234 );
 a7976a <=( a7975a  and  a7972a );
 a7980a <=( (not A168)  and  (not A169) );
 a7981a <=( (not A170)  and  a7980a );
 a7984a <=( A201  and  A199 );
 a7987a <=( A268  and  A235 );
 a7988a <=( a7987a  and  a7984a );
 a7992a <=( (not A168)  and  (not A169) );
 a7993a <=( (not A170)  and  a7992a );
 a7996a <=( A201  and  A200 );
 a7999a <=( A268  and  A235 );
 a8000a <=( a7999a  and  a7996a );
 a8003a <=( A166  and  A168 );
 a8006a <=( (not A202)  and  (not A201) );
 a8007a <=( a8006a  and  a8003a );
 a8010a <=( A235  and  (not A203) );
 a8013a <=( A267  and  A265 );
 a8014a <=( a8013a  and  a8010a );
 a8017a <=( A166  and  A168 );
 a8020a <=( (not A202)  and  (not A201) );
 a8021a <=( a8020a  and  a8017a );
 a8024a <=( A235  and  (not A203) );
 a8027a <=( A267  and  A266 );
 a8028a <=( a8027a  and  a8024a );
 a8031a <=( A166  and  A168 );
 a8034a <=( (not A202)  and  (not A201) );
 a8035a <=( a8034a  and  a8031a );
 a8038a <=( A232  and  (not A203) );
 a8041a <=( A268  and  A234 );
 a8042a <=( a8041a  and  a8038a );
 a8045a <=( A166  and  A168 );
 a8048a <=( (not A202)  and  (not A201) );
 a8049a <=( a8048a  and  a8045a );
 a8052a <=( A233  and  (not A203) );
 a8055a <=( A268  and  A234 );
 a8056a <=( a8055a  and  a8052a );
 a8059a <=( A166  and  A168 );
 a8062a <=( A200  and  A199 );
 a8063a <=( a8062a  and  a8059a );
 a8066a <=( (not A202)  and  (not A201) );
 a8069a <=( A268  and  A235 );
 a8070a <=( a8069a  and  a8066a );
 a8073a <=( A166  and  A168 );
 a8076a <=( (not A200)  and  (not A199) );
 a8077a <=( a8076a  and  a8073a );
 a8080a <=( A235  and  (not A202) );
 a8083a <=( A267  and  A265 );
 a8084a <=( a8083a  and  a8080a );
 a8087a <=( A166  and  A168 );
 a8090a <=( (not A200)  and  (not A199) );
 a8091a <=( a8090a  and  a8087a );
 a8094a <=( A235  and  (not A202) );
 a8097a <=( A267  and  A266 );
 a8098a <=( a8097a  and  a8094a );
 a8101a <=( A166  and  A168 );
 a8104a <=( (not A200)  and  (not A199) );
 a8105a <=( a8104a  and  a8101a );
 a8108a <=( A232  and  (not A202) );
 a8111a <=( A268  and  A234 );
 a8112a <=( a8111a  and  a8108a );
 a8115a <=( A166  and  A168 );
 a8118a <=( (not A200)  and  (not A199) );
 a8119a <=( a8118a  and  a8115a );
 a8122a <=( A233  and  (not A202) );
 a8125a <=( A268  and  A234 );
 a8126a <=( a8125a  and  a8122a );
 a8129a <=( A167  and  A168 );
 a8132a <=( (not A202)  and  (not A201) );
 a8133a <=( a8132a  and  a8129a );
 a8136a <=( A235  and  (not A203) );
 a8139a <=( A267  and  A265 );
 a8140a <=( a8139a  and  a8136a );
 a8143a <=( A167  and  A168 );
 a8146a <=( (not A202)  and  (not A201) );
 a8147a <=( a8146a  and  a8143a );
 a8150a <=( A235  and  (not A203) );
 a8153a <=( A267  and  A266 );
 a8154a <=( a8153a  and  a8150a );
 a8157a <=( A167  and  A168 );
 a8160a <=( (not A202)  and  (not A201) );
 a8161a <=( a8160a  and  a8157a );
 a8164a <=( A232  and  (not A203) );
 a8167a <=( A268  and  A234 );
 a8168a <=( a8167a  and  a8164a );
 a8171a <=( A167  and  A168 );
 a8174a <=( (not A202)  and  (not A201) );
 a8175a <=( a8174a  and  a8171a );
 a8178a <=( A233  and  (not A203) );
 a8181a <=( A268  and  A234 );
 a8182a <=( a8181a  and  a8178a );
 a8185a <=( A167  and  A168 );
 a8188a <=( A200  and  A199 );
 a8189a <=( a8188a  and  a8185a );
 a8192a <=( (not A202)  and  (not A201) );
 a8195a <=( A268  and  A235 );
 a8196a <=( a8195a  and  a8192a );
 a8199a <=( A167  and  A168 );
 a8202a <=( (not A200)  and  (not A199) );
 a8203a <=( a8202a  and  a8199a );
 a8206a <=( A235  and  (not A202) );
 a8209a <=( A267  and  A265 );
 a8210a <=( a8209a  and  a8206a );
 a8213a <=( A167  and  A168 );
 a8216a <=( (not A200)  and  (not A199) );
 a8217a <=( a8216a  and  a8213a );
 a8220a <=( A235  and  (not A202) );
 a8223a <=( A267  and  A266 );
 a8224a <=( a8223a  and  a8220a );
 a8227a <=( A167  and  A168 );
 a8230a <=( (not A200)  and  (not A199) );
 a8231a <=( a8230a  and  a8227a );
 a8234a <=( A232  and  (not A202) );
 a8237a <=( A268  and  A234 );
 a8238a <=( a8237a  and  a8234a );
 a8241a <=( A167  and  A168 );
 a8244a <=( (not A200)  and  (not A199) );
 a8245a <=( a8244a  and  a8241a );
 a8248a <=( A233  and  (not A202) );
 a8251a <=( A268  and  A234 );
 a8252a <=( a8251a  and  a8248a );
 a8255a <=( A167  and  A170 );
 a8258a <=( (not A201)  and  (not A166) );
 a8259a <=( a8258a  and  a8255a );
 a8262a <=( (not A203)  and  (not A202) );
 a8265a <=( A268  and  A235 );
 a8266a <=( a8265a  and  a8262a );
 a8269a <=( A167  and  A170 );
 a8272a <=( (not A199)  and  (not A166) );
 a8273a <=( a8272a  and  a8269a );
 a8276a <=( (not A202)  and  (not A200) );
 a8279a <=( A268  and  A235 );
 a8280a <=( a8279a  and  a8276a );
 a8283a <=( (not A167)  and  A170 );
 a8286a <=( (not A201)  and  A166 );
 a8287a <=( a8286a  and  a8283a );
 a8290a <=( (not A203)  and  (not A202) );
 a8293a <=( A268  and  A235 );
 a8294a <=( a8293a  and  a8290a );
 a8297a <=( (not A167)  and  A170 );
 a8300a <=( (not A199)  and  A166 );
 a8301a <=( a8300a  and  a8297a );
 a8304a <=( (not A202)  and  (not A200) );
 a8307a <=( A268  and  A235 );
 a8308a <=( a8307a  and  a8304a );
 a8311a <=( (not A201)  and  A169 );
 a8314a <=( (not A203)  and  (not A202) );
 a8315a <=( a8314a  and  a8311a );
 a8318a <=( (not A300)  and  A235 );
 a8321a <=( (not A302)  and  (not A301) );
 a8322a <=( a8321a  and  a8318a );
 a8325a <=( (not A201)  and  A169 );
 a8328a <=( (not A203)  and  (not A202) );
 a8329a <=( a8328a  and  a8325a );
 a8332a <=( (not A298)  and  A235 );
 a8335a <=( (not A301)  and  (not A299) );
 a8336a <=( a8335a  and  a8332a );
 a8339a <=( (not A201)  and  A169 );
 a8342a <=( (not A203)  and  (not A202) );
 a8343a <=( a8342a  and  a8339a );
 a8346a <=( (not A265)  and  A235 );
 a8349a <=( A269  and  A266 );
 a8350a <=( a8349a  and  a8346a );
 a8353a <=( (not A201)  and  A169 );
 a8356a <=( (not A203)  and  (not A202) );
 a8357a <=( a8356a  and  a8353a );
 a8360a <=( A265  and  A235 );
 a8363a <=( A269  and  (not A266) );
 a8364a <=( a8363a  and  a8360a );
 a8367a <=( (not A201)  and  A169 );
 a8370a <=( (not A203)  and  (not A202) );
 a8371a <=( a8370a  and  a8367a );
 a8374a <=( A234  and  A232 );
 a8377a <=( A267  and  A265 );
 a8378a <=( a8377a  and  a8374a );
 a8381a <=( (not A201)  and  A169 );
 a8384a <=( (not A203)  and  (not A202) );
 a8385a <=( a8384a  and  a8381a );
 a8388a <=( A234  and  A232 );
 a8391a <=( A267  and  A266 );
 a8392a <=( a8391a  and  a8388a );
 a8395a <=( (not A201)  and  A169 );
 a8398a <=( (not A203)  and  (not A202) );
 a8399a <=( a8398a  and  a8395a );
 a8402a <=( A234  and  A233 );
 a8405a <=( A267  and  A265 );
 a8406a <=( a8405a  and  a8402a );
 a8409a <=( (not A201)  and  A169 );
 a8412a <=( (not A203)  and  (not A202) );
 a8413a <=( a8412a  and  a8409a );
 a8416a <=( A234  and  A233 );
 a8419a <=( A267  and  A266 );
 a8420a <=( a8419a  and  a8416a );
 a8423a <=( (not A201)  and  A169 );
 a8426a <=( (not A203)  and  (not A202) );
 a8427a <=( a8426a  and  a8423a );
 a8430a <=( A233  and  (not A232) );
 a8433a <=( A268  and  A236 );
 a8434a <=( a8433a  and  a8430a );
 a8437a <=( (not A201)  and  A169 );
 a8440a <=( (not A203)  and  (not A202) );
 a8441a <=( a8440a  and  a8437a );
 a8444a <=( (not A233)  and  A232 );
 a8447a <=( A268  and  A236 );
 a8448a <=( a8447a  and  a8444a );
 a8451a <=( A199  and  A169 );
 a8454a <=( (not A201)  and  A200 );
 a8455a <=( a8454a  and  a8451a );
 a8458a <=( A235  and  (not A202) );
 a8461a <=( A267  and  A265 );
 a8462a <=( a8461a  and  a8458a );
 a8465a <=( A199  and  A169 );
 a8468a <=( (not A201)  and  A200 );
 a8469a <=( a8468a  and  a8465a );
 a8472a <=( A235  and  (not A202) );
 a8475a <=( A267  and  A266 );
 a8476a <=( a8475a  and  a8472a );
 a8479a <=( A199  and  A169 );
 a8482a <=( (not A201)  and  A200 );
 a8483a <=( a8482a  and  a8479a );
 a8486a <=( A232  and  (not A202) );
 a8489a <=( A268  and  A234 );
 a8490a <=( a8489a  and  a8486a );
 a8493a <=( A199  and  A169 );
 a8496a <=( (not A201)  and  A200 );
 a8497a <=( a8496a  and  a8493a );
 a8500a <=( A233  and  (not A202) );
 a8503a <=( A268  and  A234 );
 a8504a <=( a8503a  and  a8500a );
 a8507a <=( (not A199)  and  A169 );
 a8510a <=( (not A202)  and  (not A200) );
 a8511a <=( a8510a  and  a8507a );
 a8514a <=( (not A300)  and  A235 );
 a8517a <=( (not A302)  and  (not A301) );
 a8518a <=( a8517a  and  a8514a );
 a8521a <=( (not A199)  and  A169 );
 a8524a <=( (not A202)  and  (not A200) );
 a8525a <=( a8524a  and  a8521a );
 a8528a <=( (not A298)  and  A235 );
 a8531a <=( (not A301)  and  (not A299) );
 a8532a <=( a8531a  and  a8528a );
 a8535a <=( (not A199)  and  A169 );
 a8538a <=( (not A202)  and  (not A200) );
 a8539a <=( a8538a  and  a8535a );
 a8542a <=( (not A265)  and  A235 );
 a8545a <=( A269  and  A266 );
 a8546a <=( a8545a  and  a8542a );
 a8549a <=( (not A199)  and  A169 );
 a8552a <=( (not A202)  and  (not A200) );
 a8553a <=( a8552a  and  a8549a );
 a8556a <=( A265  and  A235 );
 a8559a <=( A269  and  (not A266) );
 a8560a <=( a8559a  and  a8556a );
 a8563a <=( (not A199)  and  A169 );
 a8566a <=( (not A202)  and  (not A200) );
 a8567a <=( a8566a  and  a8563a );
 a8570a <=( A234  and  A232 );
 a8573a <=( A267  and  A265 );
 a8574a <=( a8573a  and  a8570a );
 a8577a <=( (not A199)  and  A169 );
 a8580a <=( (not A202)  and  (not A200) );
 a8581a <=( a8580a  and  a8577a );
 a8584a <=( A234  and  A232 );
 a8587a <=( A267  and  A266 );
 a8588a <=( a8587a  and  a8584a );
 a8591a <=( (not A199)  and  A169 );
 a8594a <=( (not A202)  and  (not A200) );
 a8595a <=( a8594a  and  a8591a );
 a8598a <=( A234  and  A233 );
 a8601a <=( A267  and  A265 );
 a8602a <=( a8601a  and  a8598a );
 a8605a <=( (not A199)  and  A169 );
 a8608a <=( (not A202)  and  (not A200) );
 a8609a <=( a8608a  and  a8605a );
 a8612a <=( A234  and  A233 );
 a8615a <=( A267  and  A266 );
 a8616a <=( a8615a  and  a8612a );
 a8619a <=( (not A199)  and  A169 );
 a8622a <=( (not A202)  and  (not A200) );
 a8623a <=( a8622a  and  a8619a );
 a8626a <=( A233  and  (not A232) );
 a8629a <=( A268  and  A236 );
 a8630a <=( a8629a  and  a8626a );
 a8633a <=( (not A199)  and  A169 );
 a8636a <=( (not A202)  and  (not A200) );
 a8637a <=( a8636a  and  a8633a );
 a8640a <=( (not A233)  and  A232 );
 a8643a <=( A268  and  A236 );
 a8644a <=( a8643a  and  a8640a );
 a8647a <=( (not A167)  and  (not A169) );
 a8650a <=( A202  and  (not A166) );
 a8651a <=( a8650a  and  a8647a );
 a8654a <=( (not A300)  and  A235 );
 a8657a <=( (not A302)  and  (not A301) );
 a8658a <=( a8657a  and  a8654a );
 a8661a <=( (not A167)  and  (not A169) );
 a8664a <=( A202  and  (not A166) );
 a8665a <=( a8664a  and  a8661a );
 a8668a <=( (not A298)  and  A235 );
 a8671a <=( (not A301)  and  (not A299) );
 a8672a <=( a8671a  and  a8668a );
 a8675a <=( (not A167)  and  (not A169) );
 a8678a <=( A202  and  (not A166) );
 a8679a <=( a8678a  and  a8675a );
 a8682a <=( (not A265)  and  A235 );
 a8685a <=( A269  and  A266 );
 a8686a <=( a8685a  and  a8682a );
 a8689a <=( (not A167)  and  (not A169) );
 a8692a <=( A202  and  (not A166) );
 a8693a <=( a8692a  and  a8689a );
 a8696a <=( A265  and  A235 );
 a8699a <=( A269  and  (not A266) );
 a8700a <=( a8699a  and  a8696a );
 a8703a <=( (not A167)  and  (not A169) );
 a8706a <=( A202  and  (not A166) );
 a8707a <=( a8706a  and  a8703a );
 a8710a <=( A234  and  A232 );
 a8713a <=( A267  and  A265 );
 a8714a <=( a8713a  and  a8710a );
 a8717a <=( (not A167)  and  (not A169) );
 a8720a <=( A202  and  (not A166) );
 a8721a <=( a8720a  and  a8717a );
 a8724a <=( A234  and  A232 );
 a8727a <=( A267  and  A266 );
 a8728a <=( a8727a  and  a8724a );
 a8731a <=( (not A167)  and  (not A169) );
 a8734a <=( A202  and  (not A166) );
 a8735a <=( a8734a  and  a8731a );
 a8738a <=( A234  and  A233 );
 a8741a <=( A267  and  A265 );
 a8742a <=( a8741a  and  a8738a );
 a8745a <=( (not A167)  and  (not A169) );
 a8748a <=( A202  and  (not A166) );
 a8749a <=( a8748a  and  a8745a );
 a8752a <=( A234  and  A233 );
 a8755a <=( A267  and  A266 );
 a8756a <=( a8755a  and  a8752a );
 a8759a <=( (not A167)  and  (not A169) );
 a8762a <=( A202  and  (not A166) );
 a8763a <=( a8762a  and  a8759a );
 a8766a <=( A233  and  (not A232) );
 a8769a <=( A268  and  A236 );
 a8770a <=( a8769a  and  a8766a );
 a8773a <=( (not A167)  and  (not A169) );
 a8776a <=( A202  and  (not A166) );
 a8777a <=( a8776a  and  a8773a );
 a8780a <=( (not A233)  and  A232 );
 a8783a <=( A268  and  A236 );
 a8784a <=( a8783a  and  a8780a );
 a8787a <=( (not A167)  and  (not A169) );
 a8790a <=( A199  and  (not A166) );
 a8791a <=( a8790a  and  a8787a );
 a8794a <=( A235  and  A201 );
 a8797a <=( A267  and  A265 );
 a8798a <=( a8797a  and  a8794a );
 a8801a <=( (not A167)  and  (not A169) );
 a8804a <=( A199  and  (not A166) );
 a8805a <=( a8804a  and  a8801a );
 a8808a <=( A235  and  A201 );
 a8811a <=( A267  and  A266 );
 a8812a <=( a8811a  and  a8808a );
 a8815a <=( (not A167)  and  (not A169) );
 a8818a <=( A199  and  (not A166) );
 a8819a <=( a8818a  and  a8815a );
 a8822a <=( A232  and  A201 );
 a8825a <=( A268  and  A234 );
 a8826a <=( a8825a  and  a8822a );
 a8829a <=( (not A167)  and  (not A169) );
 a8832a <=( A199  and  (not A166) );
 a8833a <=( a8832a  and  a8829a );
 a8836a <=( A233  and  A201 );
 a8839a <=( A268  and  A234 );
 a8840a <=( a8839a  and  a8836a );
 a8843a <=( (not A167)  and  (not A169) );
 a8846a <=( A200  and  (not A166) );
 a8847a <=( a8846a  and  a8843a );
 a8850a <=( A235  and  A201 );
 a8853a <=( A267  and  A265 );
 a8854a <=( a8853a  and  a8850a );
 a8857a <=( (not A167)  and  (not A169) );
 a8860a <=( A200  and  (not A166) );
 a8861a <=( a8860a  and  a8857a );
 a8864a <=( A235  and  A201 );
 a8867a <=( A267  and  A266 );
 a8868a <=( a8867a  and  a8864a );
 a8871a <=( (not A167)  and  (not A169) );
 a8874a <=( A200  and  (not A166) );
 a8875a <=( a8874a  and  a8871a );
 a8878a <=( A232  and  A201 );
 a8881a <=( A268  and  A234 );
 a8882a <=( a8881a  and  a8878a );
 a8885a <=( (not A167)  and  (not A169) );
 a8888a <=( A200  and  (not A166) );
 a8889a <=( a8888a  and  a8885a );
 a8892a <=( A233  and  A201 );
 a8895a <=( A268  and  A234 );
 a8896a <=( a8895a  and  a8892a );
 a8899a <=( (not A167)  and  (not A169) );
 a8902a <=( (not A199)  and  (not A166) );
 a8903a <=( a8902a  and  a8899a );
 a8906a <=( A203  and  A200 );
 a8909a <=( A268  and  A235 );
 a8910a <=( a8909a  and  a8906a );
 a8913a <=( (not A167)  and  (not A169) );
 a8916a <=( A199  and  (not A166) );
 a8917a <=( a8916a  and  a8913a );
 a8920a <=( A203  and  (not A200) );
 a8923a <=( A268  and  A235 );
 a8924a <=( a8923a  and  a8920a );
 a8927a <=( (not A168)  and  (not A169) );
 a8930a <=( A166  and  A167 );
 a8931a <=( a8930a  and  a8927a );
 a8934a <=( A235  and  A202 );
 a8937a <=( A267  and  A265 );
 a8938a <=( a8937a  and  a8934a );
 a8941a <=( (not A168)  and  (not A169) );
 a8944a <=( A166  and  A167 );
 a8945a <=( a8944a  and  a8941a );
 a8948a <=( A235  and  A202 );
 a8951a <=( A267  and  A266 );
 a8952a <=( a8951a  and  a8948a );
 a8955a <=( (not A168)  and  (not A169) );
 a8958a <=( A166  and  A167 );
 a8959a <=( a8958a  and  a8955a );
 a8962a <=( A232  and  A202 );
 a8965a <=( A268  and  A234 );
 a8966a <=( a8965a  and  a8962a );
 a8969a <=( (not A168)  and  (not A169) );
 a8972a <=( A166  and  A167 );
 a8973a <=( a8972a  and  a8969a );
 a8976a <=( A233  and  A202 );
 a8979a <=( A268  and  A234 );
 a8980a <=( a8979a  and  a8976a );
 a8983a <=( (not A168)  and  (not A169) );
 a8986a <=( A166  and  A167 );
 a8987a <=( a8986a  and  a8983a );
 a8990a <=( A201  and  A199 );
 a8993a <=( A268  and  A235 );
 a8994a <=( a8993a  and  a8990a );
 a8997a <=( (not A168)  and  (not A169) );
 a9000a <=( A166  and  A167 );
 a9001a <=( a9000a  and  a8997a );
 a9004a <=( A201  and  A200 );
 a9007a <=( A268  and  A235 );
 a9008a <=( a9007a  and  a9004a );
 a9011a <=( (not A169)  and  (not A170) );
 a9014a <=( A202  and  (not A168) );
 a9015a <=( a9014a  and  a9011a );
 a9018a <=( (not A300)  and  A235 );
 a9021a <=( (not A302)  and  (not A301) );
 a9022a <=( a9021a  and  a9018a );
 a9025a <=( (not A169)  and  (not A170) );
 a9028a <=( A202  and  (not A168) );
 a9029a <=( a9028a  and  a9025a );
 a9032a <=( (not A298)  and  A235 );
 a9035a <=( (not A301)  and  (not A299) );
 a9036a <=( a9035a  and  a9032a );
 a9039a <=( (not A169)  and  (not A170) );
 a9042a <=( A202  and  (not A168) );
 a9043a <=( a9042a  and  a9039a );
 a9046a <=( (not A265)  and  A235 );
 a9049a <=( A269  and  A266 );
 a9050a <=( a9049a  and  a9046a );
 a9053a <=( (not A169)  and  (not A170) );
 a9056a <=( A202  and  (not A168) );
 a9057a <=( a9056a  and  a9053a );
 a9060a <=( A265  and  A235 );
 a9063a <=( A269  and  (not A266) );
 a9064a <=( a9063a  and  a9060a );
 a9067a <=( (not A169)  and  (not A170) );
 a9070a <=( A202  and  (not A168) );
 a9071a <=( a9070a  and  a9067a );
 a9074a <=( A234  and  A232 );
 a9077a <=( A267  and  A265 );
 a9078a <=( a9077a  and  a9074a );
 a9081a <=( (not A169)  and  (not A170) );
 a9084a <=( A202  and  (not A168) );
 a9085a <=( a9084a  and  a9081a );
 a9088a <=( A234  and  A232 );
 a9091a <=( A267  and  A266 );
 a9092a <=( a9091a  and  a9088a );
 a9095a <=( (not A169)  and  (not A170) );
 a9098a <=( A202  and  (not A168) );
 a9099a <=( a9098a  and  a9095a );
 a9102a <=( A234  and  A233 );
 a9105a <=( A267  and  A265 );
 a9106a <=( a9105a  and  a9102a );
 a9109a <=( (not A169)  and  (not A170) );
 a9112a <=( A202  and  (not A168) );
 a9113a <=( a9112a  and  a9109a );
 a9116a <=( A234  and  A233 );
 a9119a <=( A267  and  A266 );
 a9120a <=( a9119a  and  a9116a );
 a9123a <=( (not A169)  and  (not A170) );
 a9126a <=( A202  and  (not A168) );
 a9127a <=( a9126a  and  a9123a );
 a9130a <=( A233  and  (not A232) );
 a9133a <=( A268  and  A236 );
 a9134a <=( a9133a  and  a9130a );
 a9137a <=( (not A169)  and  (not A170) );
 a9140a <=( A202  and  (not A168) );
 a9141a <=( a9140a  and  a9137a );
 a9144a <=( (not A233)  and  A232 );
 a9147a <=( A268  and  A236 );
 a9148a <=( a9147a  and  a9144a );
 a9151a <=( (not A169)  and  (not A170) );
 a9154a <=( A199  and  (not A168) );
 a9155a <=( a9154a  and  a9151a );
 a9158a <=( A235  and  A201 );
 a9161a <=( A267  and  A265 );
 a9162a <=( a9161a  and  a9158a );
 a9165a <=( (not A169)  and  (not A170) );
 a9168a <=( A199  and  (not A168) );
 a9169a <=( a9168a  and  a9165a );
 a9172a <=( A235  and  A201 );
 a9175a <=( A267  and  A266 );
 a9176a <=( a9175a  and  a9172a );
 a9179a <=( (not A169)  and  (not A170) );
 a9182a <=( A199  and  (not A168) );
 a9183a <=( a9182a  and  a9179a );
 a9186a <=( A232  and  A201 );
 a9189a <=( A268  and  A234 );
 a9190a <=( a9189a  and  a9186a );
 a9193a <=( (not A169)  and  (not A170) );
 a9196a <=( A199  and  (not A168) );
 a9197a <=( a9196a  and  a9193a );
 a9200a <=( A233  and  A201 );
 a9203a <=( A268  and  A234 );
 a9204a <=( a9203a  and  a9200a );
 a9207a <=( (not A169)  and  (not A170) );
 a9210a <=( A200  and  (not A168) );
 a9211a <=( a9210a  and  a9207a );
 a9214a <=( A235  and  A201 );
 a9217a <=( A267  and  A265 );
 a9218a <=( a9217a  and  a9214a );
 a9221a <=( (not A169)  and  (not A170) );
 a9224a <=( A200  and  (not A168) );
 a9225a <=( a9224a  and  a9221a );
 a9228a <=( A235  and  A201 );
 a9231a <=( A267  and  A266 );
 a9232a <=( a9231a  and  a9228a );
 a9235a <=( (not A169)  and  (not A170) );
 a9238a <=( A200  and  (not A168) );
 a9239a <=( a9238a  and  a9235a );
 a9242a <=( A232  and  A201 );
 a9245a <=( A268  and  A234 );
 a9246a <=( a9245a  and  a9242a );
 a9249a <=( (not A169)  and  (not A170) );
 a9252a <=( A200  and  (not A168) );
 a9253a <=( a9252a  and  a9249a );
 a9256a <=( A233  and  A201 );
 a9259a <=( A268  and  A234 );
 a9260a <=( a9259a  and  a9256a );
 a9263a <=( (not A169)  and  (not A170) );
 a9266a <=( (not A199)  and  (not A168) );
 a9267a <=( a9266a  and  a9263a );
 a9270a <=( A203  and  A200 );
 a9273a <=( A268  and  A235 );
 a9274a <=( a9273a  and  a9270a );
 a9277a <=( (not A169)  and  (not A170) );
 a9280a <=( A199  and  (not A168) );
 a9281a <=( a9280a  and  a9277a );
 a9284a <=( A203  and  (not A200) );
 a9287a <=( A268  and  A235 );
 a9288a <=( a9287a  and  a9284a );
 a9291a <=( A166  and  A168 );
 a9294a <=( (not A202)  and  (not A201) );
 a9295a <=( a9294a  and  a9291a );
 a9298a <=( A235  and  (not A203) );
 a9302a <=( (not A302)  and  (not A301) );
 a9303a <=( (not A300)  and  a9302a );
 a9304a <=( a9303a  and  a9298a );
 a9307a <=( A166  and  A168 );
 a9310a <=( (not A202)  and  (not A201) );
 a9311a <=( a9310a  and  a9307a );
 a9314a <=( A235  and  (not A203) );
 a9318a <=( (not A301)  and  (not A299) );
 a9319a <=( (not A298)  and  a9318a );
 a9320a <=( a9319a  and  a9314a );
 a9323a <=( A166  and  A168 );
 a9326a <=( (not A202)  and  (not A201) );
 a9327a <=( a9326a  and  a9323a );
 a9330a <=( A235  and  (not A203) );
 a9334a <=( A269  and  A266 );
 a9335a <=( (not A265)  and  a9334a );
 a9336a <=( a9335a  and  a9330a );
 a9339a <=( A166  and  A168 );
 a9342a <=( (not A202)  and  (not A201) );
 a9343a <=( a9342a  and  a9339a );
 a9346a <=( A235  and  (not A203) );
 a9350a <=( A269  and  (not A266) );
 a9351a <=( A265  and  a9350a );
 a9352a <=( a9351a  and  a9346a );
 a9355a <=( A166  and  A168 );
 a9358a <=( (not A202)  and  (not A201) );
 a9359a <=( a9358a  and  a9355a );
 a9362a <=( A232  and  (not A203) );
 a9366a <=( A267  and  A265 );
 a9367a <=( A234  and  a9366a );
 a9368a <=( a9367a  and  a9362a );
 a9371a <=( A166  and  A168 );
 a9374a <=( (not A202)  and  (not A201) );
 a9375a <=( a9374a  and  a9371a );
 a9378a <=( A232  and  (not A203) );
 a9382a <=( A267  and  A266 );
 a9383a <=( A234  and  a9382a );
 a9384a <=( a9383a  and  a9378a );
 a9387a <=( A166  and  A168 );
 a9390a <=( (not A202)  and  (not A201) );
 a9391a <=( a9390a  and  a9387a );
 a9394a <=( A233  and  (not A203) );
 a9398a <=( A267  and  A265 );
 a9399a <=( A234  and  a9398a );
 a9400a <=( a9399a  and  a9394a );
 a9403a <=( A166  and  A168 );
 a9406a <=( (not A202)  and  (not A201) );
 a9407a <=( a9406a  and  a9403a );
 a9410a <=( A233  and  (not A203) );
 a9414a <=( A267  and  A266 );
 a9415a <=( A234  and  a9414a );
 a9416a <=( a9415a  and  a9410a );
 a9419a <=( A166  and  A168 );
 a9422a <=( (not A202)  and  (not A201) );
 a9423a <=( a9422a  and  a9419a );
 a9426a <=( (not A232)  and  (not A203) );
 a9430a <=( A268  and  A236 );
 a9431a <=( A233  and  a9430a );
 a9432a <=( a9431a  and  a9426a );
 a9435a <=( A166  and  A168 );
 a9438a <=( (not A202)  and  (not A201) );
 a9439a <=( a9438a  and  a9435a );
 a9442a <=( A232  and  (not A203) );
 a9446a <=( A268  and  A236 );
 a9447a <=( (not A233)  and  a9446a );
 a9448a <=( a9447a  and  a9442a );
 a9451a <=( A166  and  A168 );
 a9454a <=( A200  and  A199 );
 a9455a <=( a9454a  and  a9451a );
 a9458a <=( (not A202)  and  (not A201) );
 a9462a <=( A267  and  A265 );
 a9463a <=( A235  and  a9462a );
 a9464a <=( a9463a  and  a9458a );
 a9467a <=( A166  and  A168 );
 a9470a <=( A200  and  A199 );
 a9471a <=( a9470a  and  a9467a );
 a9474a <=( (not A202)  and  (not A201) );
 a9478a <=( A267  and  A266 );
 a9479a <=( A235  and  a9478a );
 a9480a <=( a9479a  and  a9474a );
 a9483a <=( A166  and  A168 );
 a9486a <=( A200  and  A199 );
 a9487a <=( a9486a  and  a9483a );
 a9490a <=( (not A202)  and  (not A201) );
 a9494a <=( A268  and  A234 );
 a9495a <=( A232  and  a9494a );
 a9496a <=( a9495a  and  a9490a );
 a9499a <=( A166  and  A168 );
 a9502a <=( A200  and  A199 );
 a9503a <=( a9502a  and  a9499a );
 a9506a <=( (not A202)  and  (not A201) );
 a9510a <=( A268  and  A234 );
 a9511a <=( A233  and  a9510a );
 a9512a <=( a9511a  and  a9506a );
 a9515a <=( A166  and  A168 );
 a9518a <=( (not A200)  and  (not A199) );
 a9519a <=( a9518a  and  a9515a );
 a9522a <=( A235  and  (not A202) );
 a9526a <=( (not A302)  and  (not A301) );
 a9527a <=( (not A300)  and  a9526a );
 a9528a <=( a9527a  and  a9522a );
 a9531a <=( A166  and  A168 );
 a9534a <=( (not A200)  and  (not A199) );
 a9535a <=( a9534a  and  a9531a );
 a9538a <=( A235  and  (not A202) );
 a9542a <=( (not A301)  and  (not A299) );
 a9543a <=( (not A298)  and  a9542a );
 a9544a <=( a9543a  and  a9538a );
 a9547a <=( A166  and  A168 );
 a9550a <=( (not A200)  and  (not A199) );
 a9551a <=( a9550a  and  a9547a );
 a9554a <=( A235  and  (not A202) );
 a9558a <=( A269  and  A266 );
 a9559a <=( (not A265)  and  a9558a );
 a9560a <=( a9559a  and  a9554a );
 a9563a <=( A166  and  A168 );
 a9566a <=( (not A200)  and  (not A199) );
 a9567a <=( a9566a  and  a9563a );
 a9570a <=( A235  and  (not A202) );
 a9574a <=( A269  and  (not A266) );
 a9575a <=( A265  and  a9574a );
 a9576a <=( a9575a  and  a9570a );
 a9579a <=( A166  and  A168 );
 a9582a <=( (not A200)  and  (not A199) );
 a9583a <=( a9582a  and  a9579a );
 a9586a <=( A232  and  (not A202) );
 a9590a <=( A267  and  A265 );
 a9591a <=( A234  and  a9590a );
 a9592a <=( a9591a  and  a9586a );
 a9595a <=( A166  and  A168 );
 a9598a <=( (not A200)  and  (not A199) );
 a9599a <=( a9598a  and  a9595a );
 a9602a <=( A232  and  (not A202) );
 a9606a <=( A267  and  A266 );
 a9607a <=( A234  and  a9606a );
 a9608a <=( a9607a  and  a9602a );
 a9611a <=( A166  and  A168 );
 a9614a <=( (not A200)  and  (not A199) );
 a9615a <=( a9614a  and  a9611a );
 a9618a <=( A233  and  (not A202) );
 a9622a <=( A267  and  A265 );
 a9623a <=( A234  and  a9622a );
 a9624a <=( a9623a  and  a9618a );
 a9627a <=( A166  and  A168 );
 a9630a <=( (not A200)  and  (not A199) );
 a9631a <=( a9630a  and  a9627a );
 a9634a <=( A233  and  (not A202) );
 a9638a <=( A267  and  A266 );
 a9639a <=( A234  and  a9638a );
 a9640a <=( a9639a  and  a9634a );
 a9643a <=( A166  and  A168 );
 a9646a <=( (not A200)  and  (not A199) );
 a9647a <=( a9646a  and  a9643a );
 a9650a <=( (not A232)  and  (not A202) );
 a9654a <=( A268  and  A236 );
 a9655a <=( A233  and  a9654a );
 a9656a <=( a9655a  and  a9650a );
 a9659a <=( A166  and  A168 );
 a9662a <=( (not A200)  and  (not A199) );
 a9663a <=( a9662a  and  a9659a );
 a9666a <=( A232  and  (not A202) );
 a9670a <=( A268  and  A236 );
 a9671a <=( (not A233)  and  a9670a );
 a9672a <=( a9671a  and  a9666a );
 a9675a <=( A167  and  A168 );
 a9678a <=( (not A202)  and  (not A201) );
 a9679a <=( a9678a  and  a9675a );
 a9682a <=( A235  and  (not A203) );
 a9686a <=( (not A302)  and  (not A301) );
 a9687a <=( (not A300)  and  a9686a );
 a9688a <=( a9687a  and  a9682a );
 a9691a <=( A167  and  A168 );
 a9694a <=( (not A202)  and  (not A201) );
 a9695a <=( a9694a  and  a9691a );
 a9698a <=( A235  and  (not A203) );
 a9702a <=( (not A301)  and  (not A299) );
 a9703a <=( (not A298)  and  a9702a );
 a9704a <=( a9703a  and  a9698a );
 a9707a <=( A167  and  A168 );
 a9710a <=( (not A202)  and  (not A201) );
 a9711a <=( a9710a  and  a9707a );
 a9714a <=( A235  and  (not A203) );
 a9718a <=( A269  and  A266 );
 a9719a <=( (not A265)  and  a9718a );
 a9720a <=( a9719a  and  a9714a );
 a9723a <=( A167  and  A168 );
 a9726a <=( (not A202)  and  (not A201) );
 a9727a <=( a9726a  and  a9723a );
 a9730a <=( A235  and  (not A203) );
 a9734a <=( A269  and  (not A266) );
 a9735a <=( A265  and  a9734a );
 a9736a <=( a9735a  and  a9730a );
 a9739a <=( A167  and  A168 );
 a9742a <=( (not A202)  and  (not A201) );
 a9743a <=( a9742a  and  a9739a );
 a9746a <=( A232  and  (not A203) );
 a9750a <=( A267  and  A265 );
 a9751a <=( A234  and  a9750a );
 a9752a <=( a9751a  and  a9746a );
 a9755a <=( A167  and  A168 );
 a9758a <=( (not A202)  and  (not A201) );
 a9759a <=( a9758a  and  a9755a );
 a9762a <=( A232  and  (not A203) );
 a9766a <=( A267  and  A266 );
 a9767a <=( A234  and  a9766a );
 a9768a <=( a9767a  and  a9762a );
 a9771a <=( A167  and  A168 );
 a9774a <=( (not A202)  and  (not A201) );
 a9775a <=( a9774a  and  a9771a );
 a9778a <=( A233  and  (not A203) );
 a9782a <=( A267  and  A265 );
 a9783a <=( A234  and  a9782a );
 a9784a <=( a9783a  and  a9778a );
 a9787a <=( A167  and  A168 );
 a9790a <=( (not A202)  and  (not A201) );
 a9791a <=( a9790a  and  a9787a );
 a9794a <=( A233  and  (not A203) );
 a9798a <=( A267  and  A266 );
 a9799a <=( A234  and  a9798a );
 a9800a <=( a9799a  and  a9794a );
 a9803a <=( A167  and  A168 );
 a9806a <=( (not A202)  and  (not A201) );
 a9807a <=( a9806a  and  a9803a );
 a9810a <=( (not A232)  and  (not A203) );
 a9814a <=( A268  and  A236 );
 a9815a <=( A233  and  a9814a );
 a9816a <=( a9815a  and  a9810a );
 a9819a <=( A167  and  A168 );
 a9822a <=( (not A202)  and  (not A201) );
 a9823a <=( a9822a  and  a9819a );
 a9826a <=( A232  and  (not A203) );
 a9830a <=( A268  and  A236 );
 a9831a <=( (not A233)  and  a9830a );
 a9832a <=( a9831a  and  a9826a );
 a9835a <=( A167  and  A168 );
 a9838a <=( A200  and  A199 );
 a9839a <=( a9838a  and  a9835a );
 a9842a <=( (not A202)  and  (not A201) );
 a9846a <=( A267  and  A265 );
 a9847a <=( A235  and  a9846a );
 a9848a <=( a9847a  and  a9842a );
 a9851a <=( A167  and  A168 );
 a9854a <=( A200  and  A199 );
 a9855a <=( a9854a  and  a9851a );
 a9858a <=( (not A202)  and  (not A201) );
 a9862a <=( A267  and  A266 );
 a9863a <=( A235  and  a9862a );
 a9864a <=( a9863a  and  a9858a );
 a9867a <=( A167  and  A168 );
 a9870a <=( A200  and  A199 );
 a9871a <=( a9870a  and  a9867a );
 a9874a <=( (not A202)  and  (not A201) );
 a9878a <=( A268  and  A234 );
 a9879a <=( A232  and  a9878a );
 a9880a <=( a9879a  and  a9874a );
 a9883a <=( A167  and  A168 );
 a9886a <=( A200  and  A199 );
 a9887a <=( a9886a  and  a9883a );
 a9890a <=( (not A202)  and  (not A201) );
 a9894a <=( A268  and  A234 );
 a9895a <=( A233  and  a9894a );
 a9896a <=( a9895a  and  a9890a );
 a9899a <=( A167  and  A168 );
 a9902a <=( (not A200)  and  (not A199) );
 a9903a <=( a9902a  and  a9899a );
 a9906a <=( A235  and  (not A202) );
 a9910a <=( (not A302)  and  (not A301) );
 a9911a <=( (not A300)  and  a9910a );
 a9912a <=( a9911a  and  a9906a );
 a9915a <=( A167  and  A168 );
 a9918a <=( (not A200)  and  (not A199) );
 a9919a <=( a9918a  and  a9915a );
 a9922a <=( A235  and  (not A202) );
 a9926a <=( (not A301)  and  (not A299) );
 a9927a <=( (not A298)  and  a9926a );
 a9928a <=( a9927a  and  a9922a );
 a9931a <=( A167  and  A168 );
 a9934a <=( (not A200)  and  (not A199) );
 a9935a <=( a9934a  and  a9931a );
 a9938a <=( A235  and  (not A202) );
 a9942a <=( A269  and  A266 );
 a9943a <=( (not A265)  and  a9942a );
 a9944a <=( a9943a  and  a9938a );
 a9947a <=( A167  and  A168 );
 a9950a <=( (not A200)  and  (not A199) );
 a9951a <=( a9950a  and  a9947a );
 a9954a <=( A235  and  (not A202) );
 a9958a <=( A269  and  (not A266) );
 a9959a <=( A265  and  a9958a );
 a9960a <=( a9959a  and  a9954a );
 a9963a <=( A167  and  A168 );
 a9966a <=( (not A200)  and  (not A199) );
 a9967a <=( a9966a  and  a9963a );
 a9970a <=( A232  and  (not A202) );
 a9974a <=( A267  and  A265 );
 a9975a <=( A234  and  a9974a );
 a9976a <=( a9975a  and  a9970a );
 a9979a <=( A167  and  A168 );
 a9982a <=( (not A200)  and  (not A199) );
 a9983a <=( a9982a  and  a9979a );
 a9986a <=( A232  and  (not A202) );
 a9990a <=( A267  and  A266 );
 a9991a <=( A234  and  a9990a );
 a9992a <=( a9991a  and  a9986a );
 a9995a <=( A167  and  A168 );
 a9998a <=( (not A200)  and  (not A199) );
 a9999a <=( a9998a  and  a9995a );
 a10002a <=( A233  and  (not A202) );
 a10006a <=( A267  and  A265 );
 a10007a <=( A234  and  a10006a );
 a10008a <=( a10007a  and  a10002a );
 a10011a <=( A167  and  A168 );
 a10014a <=( (not A200)  and  (not A199) );
 a10015a <=( a10014a  and  a10011a );
 a10018a <=( A233  and  (not A202) );
 a10022a <=( A267  and  A266 );
 a10023a <=( A234  and  a10022a );
 a10024a <=( a10023a  and  a10018a );
 a10027a <=( A167  and  A168 );
 a10030a <=( (not A200)  and  (not A199) );
 a10031a <=( a10030a  and  a10027a );
 a10034a <=( (not A232)  and  (not A202) );
 a10038a <=( A268  and  A236 );
 a10039a <=( A233  and  a10038a );
 a10040a <=( a10039a  and  a10034a );
 a10043a <=( A167  and  A168 );
 a10046a <=( (not A200)  and  (not A199) );
 a10047a <=( a10046a  and  a10043a );
 a10050a <=( A232  and  (not A202) );
 a10054a <=( A268  and  A236 );
 a10055a <=( (not A233)  and  a10054a );
 a10056a <=( a10055a  and  a10050a );
 a10059a <=( A167  and  A170 );
 a10062a <=( (not A201)  and  (not A166) );
 a10063a <=( a10062a  and  a10059a );
 a10066a <=( (not A203)  and  (not A202) );
 a10070a <=( A267  and  A265 );
 a10071a <=( A235  and  a10070a );
 a10072a <=( a10071a  and  a10066a );
 a10075a <=( A167  and  A170 );
 a10078a <=( (not A201)  and  (not A166) );
 a10079a <=( a10078a  and  a10075a );
 a10082a <=( (not A203)  and  (not A202) );
 a10086a <=( A267  and  A266 );
 a10087a <=( A235  and  a10086a );
 a10088a <=( a10087a  and  a10082a );
 a10091a <=( A167  and  A170 );
 a10094a <=( (not A201)  and  (not A166) );
 a10095a <=( a10094a  and  a10091a );
 a10098a <=( (not A203)  and  (not A202) );
 a10102a <=( A268  and  A234 );
 a10103a <=( A232  and  a10102a );
 a10104a <=( a10103a  and  a10098a );
 a10107a <=( A167  and  A170 );
 a10110a <=( (not A201)  and  (not A166) );
 a10111a <=( a10110a  and  a10107a );
 a10114a <=( (not A203)  and  (not A202) );
 a10118a <=( A268  and  A234 );
 a10119a <=( A233  and  a10118a );
 a10120a <=( a10119a  and  a10114a );
 a10123a <=( A167  and  A170 );
 a10126a <=( A199  and  (not A166) );
 a10127a <=( a10126a  and  a10123a );
 a10130a <=( (not A201)  and  A200 );
 a10134a <=( A268  and  A235 );
 a10135a <=( (not A202)  and  a10134a );
 a10136a <=( a10135a  and  a10130a );
 a10139a <=( A167  and  A170 );
 a10142a <=( (not A199)  and  (not A166) );
 a10143a <=( a10142a  and  a10139a );
 a10146a <=( (not A202)  and  (not A200) );
 a10150a <=( A267  and  A265 );
 a10151a <=( A235  and  a10150a );
 a10152a <=( a10151a  and  a10146a );
 a10155a <=( A167  and  A170 );
 a10158a <=( (not A199)  and  (not A166) );
 a10159a <=( a10158a  and  a10155a );
 a10162a <=( (not A202)  and  (not A200) );
 a10166a <=( A267  and  A266 );
 a10167a <=( A235  and  a10166a );
 a10168a <=( a10167a  and  a10162a );
 a10171a <=( A167  and  A170 );
 a10174a <=( (not A199)  and  (not A166) );
 a10175a <=( a10174a  and  a10171a );
 a10178a <=( (not A202)  and  (not A200) );
 a10182a <=( A268  and  A234 );
 a10183a <=( A232  and  a10182a );
 a10184a <=( a10183a  and  a10178a );
 a10187a <=( A167  and  A170 );
 a10190a <=( (not A199)  and  (not A166) );
 a10191a <=( a10190a  and  a10187a );
 a10194a <=( (not A202)  and  (not A200) );
 a10198a <=( A268  and  A234 );
 a10199a <=( A233  and  a10198a );
 a10200a <=( a10199a  and  a10194a );
 a10203a <=( (not A167)  and  A170 );
 a10206a <=( (not A201)  and  A166 );
 a10207a <=( a10206a  and  a10203a );
 a10210a <=( (not A203)  and  (not A202) );
 a10214a <=( A267  and  A265 );
 a10215a <=( A235  and  a10214a );
 a10216a <=( a10215a  and  a10210a );
 a10219a <=( (not A167)  and  A170 );
 a10222a <=( (not A201)  and  A166 );
 a10223a <=( a10222a  and  a10219a );
 a10226a <=( (not A203)  and  (not A202) );
 a10230a <=( A267  and  A266 );
 a10231a <=( A235  and  a10230a );
 a10232a <=( a10231a  and  a10226a );
 a10235a <=( (not A167)  and  A170 );
 a10238a <=( (not A201)  and  A166 );
 a10239a <=( a10238a  and  a10235a );
 a10242a <=( (not A203)  and  (not A202) );
 a10246a <=( A268  and  A234 );
 a10247a <=( A232  and  a10246a );
 a10248a <=( a10247a  and  a10242a );
 a10251a <=( (not A167)  and  A170 );
 a10254a <=( (not A201)  and  A166 );
 a10255a <=( a10254a  and  a10251a );
 a10258a <=( (not A203)  and  (not A202) );
 a10262a <=( A268  and  A234 );
 a10263a <=( A233  and  a10262a );
 a10264a <=( a10263a  and  a10258a );
 a10267a <=( (not A167)  and  A170 );
 a10270a <=( A199  and  A166 );
 a10271a <=( a10270a  and  a10267a );
 a10274a <=( (not A201)  and  A200 );
 a10278a <=( A268  and  A235 );
 a10279a <=( (not A202)  and  a10278a );
 a10280a <=( a10279a  and  a10274a );
 a10283a <=( (not A167)  and  A170 );
 a10286a <=( (not A199)  and  A166 );
 a10287a <=( a10286a  and  a10283a );
 a10290a <=( (not A202)  and  (not A200) );
 a10294a <=( A267  and  A265 );
 a10295a <=( A235  and  a10294a );
 a10296a <=( a10295a  and  a10290a );
 a10299a <=( (not A167)  and  A170 );
 a10302a <=( (not A199)  and  A166 );
 a10303a <=( a10302a  and  a10299a );
 a10306a <=( (not A202)  and  (not A200) );
 a10310a <=( A267  and  A266 );
 a10311a <=( A235  and  a10310a );
 a10312a <=( a10311a  and  a10306a );
 a10315a <=( (not A167)  and  A170 );
 a10318a <=( (not A199)  and  A166 );
 a10319a <=( a10318a  and  a10315a );
 a10322a <=( (not A202)  and  (not A200) );
 a10326a <=( A268  and  A234 );
 a10327a <=( A232  and  a10326a );
 a10328a <=( a10327a  and  a10322a );
 a10331a <=( (not A167)  and  A170 );
 a10334a <=( (not A199)  and  A166 );
 a10335a <=( a10334a  and  a10331a );
 a10338a <=( (not A202)  and  (not A200) );
 a10342a <=( A268  and  A234 );
 a10343a <=( A233  and  a10342a );
 a10344a <=( a10343a  and  a10338a );
 a10347a <=( (not A201)  and  A169 );
 a10350a <=( (not A203)  and  (not A202) );
 a10351a <=( a10350a  and  a10347a );
 a10354a <=( A298  and  A235 );
 a10358a <=( (not A301)  and  (not A300) );
 a10359a <=( A299  and  a10358a );
 a10360a <=( a10359a  and  a10354a );
 a10363a <=( (not A201)  and  A169 );
 a10366a <=( (not A203)  and  (not A202) );
 a10367a <=( a10366a  and  a10363a );
 a10370a <=( A234  and  A232 );
 a10374a <=( (not A302)  and  (not A301) );
 a10375a <=( (not A300)  and  a10374a );
 a10376a <=( a10375a  and  a10370a );
 a10379a <=( (not A201)  and  A169 );
 a10382a <=( (not A203)  and  (not A202) );
 a10383a <=( a10382a  and  a10379a );
 a10386a <=( A234  and  A232 );
 a10390a <=( (not A301)  and  (not A299) );
 a10391a <=( (not A298)  and  a10390a );
 a10392a <=( a10391a  and  a10386a );
 a10395a <=( (not A201)  and  A169 );
 a10398a <=( (not A203)  and  (not A202) );
 a10399a <=( a10398a  and  a10395a );
 a10402a <=( A234  and  A232 );
 a10406a <=( A269  and  A266 );
 a10407a <=( (not A265)  and  a10406a );
 a10408a <=( a10407a  and  a10402a );
 a10411a <=( (not A201)  and  A169 );
 a10414a <=( (not A203)  and  (not A202) );
 a10415a <=( a10414a  and  a10411a );
 a10418a <=( A234  and  A232 );
 a10422a <=( A269  and  (not A266) );
 a10423a <=( A265  and  a10422a );
 a10424a <=( a10423a  and  a10418a );
 a10427a <=( (not A201)  and  A169 );
 a10430a <=( (not A203)  and  (not A202) );
 a10431a <=( a10430a  and  a10427a );
 a10434a <=( A234  and  A233 );
 a10438a <=( (not A302)  and  (not A301) );
 a10439a <=( (not A300)  and  a10438a );
 a10440a <=( a10439a  and  a10434a );
 a10443a <=( (not A201)  and  A169 );
 a10446a <=( (not A203)  and  (not A202) );
 a10447a <=( a10446a  and  a10443a );
 a10450a <=( A234  and  A233 );
 a10454a <=( (not A301)  and  (not A299) );
 a10455a <=( (not A298)  and  a10454a );
 a10456a <=( a10455a  and  a10450a );
 a10459a <=( (not A201)  and  A169 );
 a10462a <=( (not A203)  and  (not A202) );
 a10463a <=( a10462a  and  a10459a );
 a10466a <=( A234  and  A233 );
 a10470a <=( A269  and  A266 );
 a10471a <=( (not A265)  and  a10470a );
 a10472a <=( a10471a  and  a10466a );
 a10475a <=( (not A201)  and  A169 );
 a10478a <=( (not A203)  and  (not A202) );
 a10479a <=( a10478a  and  a10475a );
 a10482a <=( A234  and  A233 );
 a10486a <=( A269  and  (not A266) );
 a10487a <=( A265  and  a10486a );
 a10488a <=( a10487a  and  a10482a );
 a10491a <=( (not A201)  and  A169 );
 a10494a <=( (not A203)  and  (not A202) );
 a10495a <=( a10494a  and  a10491a );
 a10498a <=( A233  and  (not A232) );
 a10502a <=( A267  and  A265 );
 a10503a <=( A236  and  a10502a );
 a10504a <=( a10503a  and  a10498a );
 a10507a <=( (not A201)  and  A169 );
 a10510a <=( (not A203)  and  (not A202) );
 a10511a <=( a10510a  and  a10507a );
 a10514a <=( A233  and  (not A232) );
 a10518a <=( A267  and  A266 );
 a10519a <=( A236  and  a10518a );
 a10520a <=( a10519a  and  a10514a );
 a10523a <=( (not A201)  and  A169 );
 a10526a <=( (not A203)  and  (not A202) );
 a10527a <=( a10526a  and  a10523a );
 a10530a <=( (not A233)  and  A232 );
 a10534a <=( A267  and  A265 );
 a10535a <=( A236  and  a10534a );
 a10536a <=( a10535a  and  a10530a );
 a10539a <=( (not A201)  and  A169 );
 a10542a <=( (not A203)  and  (not A202) );
 a10543a <=( a10542a  and  a10539a );
 a10546a <=( (not A233)  and  A232 );
 a10550a <=( A267  and  A266 );
 a10551a <=( A236  and  a10550a );
 a10552a <=( a10551a  and  a10546a );
 a10555a <=( A199  and  A169 );
 a10558a <=( (not A201)  and  A200 );
 a10559a <=( a10558a  and  a10555a );
 a10562a <=( A235  and  (not A202) );
 a10566a <=( (not A302)  and  (not A301) );
 a10567a <=( (not A300)  and  a10566a );
 a10568a <=( a10567a  and  a10562a );
 a10571a <=( A199  and  A169 );
 a10574a <=( (not A201)  and  A200 );
 a10575a <=( a10574a  and  a10571a );
 a10578a <=( A235  and  (not A202) );
 a10582a <=( (not A301)  and  (not A299) );
 a10583a <=( (not A298)  and  a10582a );
 a10584a <=( a10583a  and  a10578a );
 a10587a <=( A199  and  A169 );
 a10590a <=( (not A201)  and  A200 );
 a10591a <=( a10590a  and  a10587a );
 a10594a <=( A235  and  (not A202) );
 a10598a <=( A269  and  A266 );
 a10599a <=( (not A265)  and  a10598a );
 a10600a <=( a10599a  and  a10594a );
 a10603a <=( A199  and  A169 );
 a10606a <=( (not A201)  and  A200 );
 a10607a <=( a10606a  and  a10603a );
 a10610a <=( A235  and  (not A202) );
 a10614a <=( A269  and  (not A266) );
 a10615a <=( A265  and  a10614a );
 a10616a <=( a10615a  and  a10610a );
 a10619a <=( A199  and  A169 );
 a10622a <=( (not A201)  and  A200 );
 a10623a <=( a10622a  and  a10619a );
 a10626a <=( A232  and  (not A202) );
 a10630a <=( A267  and  A265 );
 a10631a <=( A234  and  a10630a );
 a10632a <=( a10631a  and  a10626a );
 a10635a <=( A199  and  A169 );
 a10638a <=( (not A201)  and  A200 );
 a10639a <=( a10638a  and  a10635a );
 a10642a <=( A232  and  (not A202) );
 a10646a <=( A267  and  A266 );
 a10647a <=( A234  and  a10646a );
 a10648a <=( a10647a  and  a10642a );
 a10651a <=( A199  and  A169 );
 a10654a <=( (not A201)  and  A200 );
 a10655a <=( a10654a  and  a10651a );
 a10658a <=( A233  and  (not A202) );
 a10662a <=( A267  and  A265 );
 a10663a <=( A234  and  a10662a );
 a10664a <=( a10663a  and  a10658a );
 a10667a <=( A199  and  A169 );
 a10670a <=( (not A201)  and  A200 );
 a10671a <=( a10670a  and  a10667a );
 a10674a <=( A233  and  (not A202) );
 a10678a <=( A267  and  A266 );
 a10679a <=( A234  and  a10678a );
 a10680a <=( a10679a  and  a10674a );
 a10683a <=( A199  and  A169 );
 a10686a <=( (not A201)  and  A200 );
 a10687a <=( a10686a  and  a10683a );
 a10690a <=( (not A232)  and  (not A202) );
 a10694a <=( A268  and  A236 );
 a10695a <=( A233  and  a10694a );
 a10696a <=( a10695a  and  a10690a );
 a10699a <=( A199  and  A169 );
 a10702a <=( (not A201)  and  A200 );
 a10703a <=( a10702a  and  a10699a );
 a10706a <=( A232  and  (not A202) );
 a10710a <=( A268  and  A236 );
 a10711a <=( (not A233)  and  a10710a );
 a10712a <=( a10711a  and  a10706a );
 a10715a <=( (not A199)  and  A169 );
 a10718a <=( (not A202)  and  (not A200) );
 a10719a <=( a10718a  and  a10715a );
 a10722a <=( A298  and  A235 );
 a10726a <=( (not A301)  and  (not A300) );
 a10727a <=( A299  and  a10726a );
 a10728a <=( a10727a  and  a10722a );
 a10731a <=( (not A199)  and  A169 );
 a10734a <=( (not A202)  and  (not A200) );
 a10735a <=( a10734a  and  a10731a );
 a10738a <=( A234  and  A232 );
 a10742a <=( (not A302)  and  (not A301) );
 a10743a <=( (not A300)  and  a10742a );
 a10744a <=( a10743a  and  a10738a );
 a10747a <=( (not A199)  and  A169 );
 a10750a <=( (not A202)  and  (not A200) );
 a10751a <=( a10750a  and  a10747a );
 a10754a <=( A234  and  A232 );
 a10758a <=( (not A301)  and  (not A299) );
 a10759a <=( (not A298)  and  a10758a );
 a10760a <=( a10759a  and  a10754a );
 a10763a <=( (not A199)  and  A169 );
 a10766a <=( (not A202)  and  (not A200) );
 a10767a <=( a10766a  and  a10763a );
 a10770a <=( A234  and  A232 );
 a10774a <=( A269  and  A266 );
 a10775a <=( (not A265)  and  a10774a );
 a10776a <=( a10775a  and  a10770a );
 a10779a <=( (not A199)  and  A169 );
 a10782a <=( (not A202)  and  (not A200) );
 a10783a <=( a10782a  and  a10779a );
 a10786a <=( A234  and  A232 );
 a10790a <=( A269  and  (not A266) );
 a10791a <=( A265  and  a10790a );
 a10792a <=( a10791a  and  a10786a );
 a10795a <=( (not A199)  and  A169 );
 a10798a <=( (not A202)  and  (not A200) );
 a10799a <=( a10798a  and  a10795a );
 a10802a <=( A234  and  A233 );
 a10806a <=( (not A302)  and  (not A301) );
 a10807a <=( (not A300)  and  a10806a );
 a10808a <=( a10807a  and  a10802a );
 a10811a <=( (not A199)  and  A169 );
 a10814a <=( (not A202)  and  (not A200) );
 a10815a <=( a10814a  and  a10811a );
 a10818a <=( A234  and  A233 );
 a10822a <=( (not A301)  and  (not A299) );
 a10823a <=( (not A298)  and  a10822a );
 a10824a <=( a10823a  and  a10818a );
 a10827a <=( (not A199)  and  A169 );
 a10830a <=( (not A202)  and  (not A200) );
 a10831a <=( a10830a  and  a10827a );
 a10834a <=( A234  and  A233 );
 a10838a <=( A269  and  A266 );
 a10839a <=( (not A265)  and  a10838a );
 a10840a <=( a10839a  and  a10834a );
 a10843a <=( (not A199)  and  A169 );
 a10846a <=( (not A202)  and  (not A200) );
 a10847a <=( a10846a  and  a10843a );
 a10850a <=( A234  and  A233 );
 a10854a <=( A269  and  (not A266) );
 a10855a <=( A265  and  a10854a );
 a10856a <=( a10855a  and  a10850a );
 a10859a <=( (not A199)  and  A169 );
 a10862a <=( (not A202)  and  (not A200) );
 a10863a <=( a10862a  and  a10859a );
 a10866a <=( A233  and  (not A232) );
 a10870a <=( A267  and  A265 );
 a10871a <=( A236  and  a10870a );
 a10872a <=( a10871a  and  a10866a );
 a10875a <=( (not A199)  and  A169 );
 a10878a <=( (not A202)  and  (not A200) );
 a10879a <=( a10878a  and  a10875a );
 a10882a <=( A233  and  (not A232) );
 a10886a <=( A267  and  A266 );
 a10887a <=( A236  and  a10886a );
 a10888a <=( a10887a  and  a10882a );
 a10891a <=( (not A199)  and  A169 );
 a10894a <=( (not A202)  and  (not A200) );
 a10895a <=( a10894a  and  a10891a );
 a10898a <=( (not A233)  and  A232 );
 a10902a <=( A267  and  A265 );
 a10903a <=( A236  and  a10902a );
 a10904a <=( a10903a  and  a10898a );
 a10907a <=( (not A199)  and  A169 );
 a10910a <=( (not A202)  and  (not A200) );
 a10911a <=( a10910a  and  a10907a );
 a10914a <=( (not A233)  and  A232 );
 a10918a <=( A267  and  A266 );
 a10919a <=( A236  and  a10918a );
 a10920a <=( a10919a  and  a10914a );
 a10923a <=( (not A167)  and  (not A169) );
 a10926a <=( A202  and  (not A166) );
 a10927a <=( a10926a  and  a10923a );
 a10930a <=( A298  and  A235 );
 a10934a <=( (not A301)  and  (not A300) );
 a10935a <=( A299  and  a10934a );
 a10936a <=( a10935a  and  a10930a );
 a10939a <=( (not A167)  and  (not A169) );
 a10942a <=( A202  and  (not A166) );
 a10943a <=( a10942a  and  a10939a );
 a10946a <=( A234  and  A232 );
 a10950a <=( (not A302)  and  (not A301) );
 a10951a <=( (not A300)  and  a10950a );
 a10952a <=( a10951a  and  a10946a );
 a10955a <=( (not A167)  and  (not A169) );
 a10958a <=( A202  and  (not A166) );
 a10959a <=( a10958a  and  a10955a );
 a10962a <=( A234  and  A232 );
 a10966a <=( (not A301)  and  (not A299) );
 a10967a <=( (not A298)  and  a10966a );
 a10968a <=( a10967a  and  a10962a );
 a10971a <=( (not A167)  and  (not A169) );
 a10974a <=( A202  and  (not A166) );
 a10975a <=( a10974a  and  a10971a );
 a10978a <=( A234  and  A232 );
 a10982a <=( A269  and  A266 );
 a10983a <=( (not A265)  and  a10982a );
 a10984a <=( a10983a  and  a10978a );
 a10987a <=( (not A167)  and  (not A169) );
 a10990a <=( A202  and  (not A166) );
 a10991a <=( a10990a  and  a10987a );
 a10994a <=( A234  and  A232 );
 a10998a <=( A269  and  (not A266) );
 a10999a <=( A265  and  a10998a );
 a11000a <=( a10999a  and  a10994a );
 a11003a <=( (not A167)  and  (not A169) );
 a11006a <=( A202  and  (not A166) );
 a11007a <=( a11006a  and  a11003a );
 a11010a <=( A234  and  A233 );
 a11014a <=( (not A302)  and  (not A301) );
 a11015a <=( (not A300)  and  a11014a );
 a11016a <=( a11015a  and  a11010a );
 a11019a <=( (not A167)  and  (not A169) );
 a11022a <=( A202  and  (not A166) );
 a11023a <=( a11022a  and  a11019a );
 a11026a <=( A234  and  A233 );
 a11030a <=( (not A301)  and  (not A299) );
 a11031a <=( (not A298)  and  a11030a );
 a11032a <=( a11031a  and  a11026a );
 a11035a <=( (not A167)  and  (not A169) );
 a11038a <=( A202  and  (not A166) );
 a11039a <=( a11038a  and  a11035a );
 a11042a <=( A234  and  A233 );
 a11046a <=( A269  and  A266 );
 a11047a <=( (not A265)  and  a11046a );
 a11048a <=( a11047a  and  a11042a );
 a11051a <=( (not A167)  and  (not A169) );
 a11054a <=( A202  and  (not A166) );
 a11055a <=( a11054a  and  a11051a );
 a11058a <=( A234  and  A233 );
 a11062a <=( A269  and  (not A266) );
 a11063a <=( A265  and  a11062a );
 a11064a <=( a11063a  and  a11058a );
 a11067a <=( (not A167)  and  (not A169) );
 a11070a <=( A202  and  (not A166) );
 a11071a <=( a11070a  and  a11067a );
 a11074a <=( A233  and  (not A232) );
 a11078a <=( A267  and  A265 );
 a11079a <=( A236  and  a11078a );
 a11080a <=( a11079a  and  a11074a );
 a11083a <=( (not A167)  and  (not A169) );
 a11086a <=( A202  and  (not A166) );
 a11087a <=( a11086a  and  a11083a );
 a11090a <=( A233  and  (not A232) );
 a11094a <=( A267  and  A266 );
 a11095a <=( A236  and  a11094a );
 a11096a <=( a11095a  and  a11090a );
 a11099a <=( (not A167)  and  (not A169) );
 a11102a <=( A202  and  (not A166) );
 a11103a <=( a11102a  and  a11099a );
 a11106a <=( (not A233)  and  A232 );
 a11110a <=( A267  and  A265 );
 a11111a <=( A236  and  a11110a );
 a11112a <=( a11111a  and  a11106a );
 a11115a <=( (not A167)  and  (not A169) );
 a11118a <=( A202  and  (not A166) );
 a11119a <=( a11118a  and  a11115a );
 a11122a <=( (not A233)  and  A232 );
 a11126a <=( A267  and  A266 );
 a11127a <=( A236  and  a11126a );
 a11128a <=( a11127a  and  a11122a );
 a11131a <=( (not A167)  and  (not A169) );
 a11134a <=( A199  and  (not A166) );
 a11135a <=( a11134a  and  a11131a );
 a11138a <=( A235  and  A201 );
 a11142a <=( (not A302)  and  (not A301) );
 a11143a <=( (not A300)  and  a11142a );
 a11144a <=( a11143a  and  a11138a );
 a11147a <=( (not A167)  and  (not A169) );
 a11150a <=( A199  and  (not A166) );
 a11151a <=( a11150a  and  a11147a );
 a11154a <=( A235  and  A201 );
 a11158a <=( (not A301)  and  (not A299) );
 a11159a <=( (not A298)  and  a11158a );
 a11160a <=( a11159a  and  a11154a );
 a11163a <=( (not A167)  and  (not A169) );
 a11166a <=( A199  and  (not A166) );
 a11167a <=( a11166a  and  a11163a );
 a11170a <=( A235  and  A201 );
 a11174a <=( A269  and  A266 );
 a11175a <=( (not A265)  and  a11174a );
 a11176a <=( a11175a  and  a11170a );
 a11179a <=( (not A167)  and  (not A169) );
 a11182a <=( A199  and  (not A166) );
 a11183a <=( a11182a  and  a11179a );
 a11186a <=( A235  and  A201 );
 a11190a <=( A269  and  (not A266) );
 a11191a <=( A265  and  a11190a );
 a11192a <=( a11191a  and  a11186a );
 a11195a <=( (not A167)  and  (not A169) );
 a11198a <=( A199  and  (not A166) );
 a11199a <=( a11198a  and  a11195a );
 a11202a <=( A232  and  A201 );
 a11206a <=( A267  and  A265 );
 a11207a <=( A234  and  a11206a );
 a11208a <=( a11207a  and  a11202a );
 a11211a <=( (not A167)  and  (not A169) );
 a11214a <=( A199  and  (not A166) );
 a11215a <=( a11214a  and  a11211a );
 a11218a <=( A232  and  A201 );
 a11222a <=( A267  and  A266 );
 a11223a <=( A234  and  a11222a );
 a11224a <=( a11223a  and  a11218a );
 a11227a <=( (not A167)  and  (not A169) );
 a11230a <=( A199  and  (not A166) );
 a11231a <=( a11230a  and  a11227a );
 a11234a <=( A233  and  A201 );
 a11238a <=( A267  and  A265 );
 a11239a <=( A234  and  a11238a );
 a11240a <=( a11239a  and  a11234a );
 a11243a <=( (not A167)  and  (not A169) );
 a11246a <=( A199  and  (not A166) );
 a11247a <=( a11246a  and  a11243a );
 a11250a <=( A233  and  A201 );
 a11254a <=( A267  and  A266 );
 a11255a <=( A234  and  a11254a );
 a11256a <=( a11255a  and  a11250a );
 a11259a <=( (not A167)  and  (not A169) );
 a11262a <=( A199  and  (not A166) );
 a11263a <=( a11262a  and  a11259a );
 a11266a <=( (not A232)  and  A201 );
 a11270a <=( A268  and  A236 );
 a11271a <=( A233  and  a11270a );
 a11272a <=( a11271a  and  a11266a );
 a11275a <=( (not A167)  and  (not A169) );
 a11278a <=( A199  and  (not A166) );
 a11279a <=( a11278a  and  a11275a );
 a11282a <=( A232  and  A201 );
 a11286a <=( A268  and  A236 );
 a11287a <=( (not A233)  and  a11286a );
 a11288a <=( a11287a  and  a11282a );
 a11291a <=( (not A167)  and  (not A169) );
 a11294a <=( A200  and  (not A166) );
 a11295a <=( a11294a  and  a11291a );
 a11298a <=( A235  and  A201 );
 a11302a <=( (not A302)  and  (not A301) );
 a11303a <=( (not A300)  and  a11302a );
 a11304a <=( a11303a  and  a11298a );
 a11307a <=( (not A167)  and  (not A169) );
 a11310a <=( A200  and  (not A166) );
 a11311a <=( a11310a  and  a11307a );
 a11314a <=( A235  and  A201 );
 a11318a <=( (not A301)  and  (not A299) );
 a11319a <=( (not A298)  and  a11318a );
 a11320a <=( a11319a  and  a11314a );
 a11323a <=( (not A167)  and  (not A169) );
 a11326a <=( A200  and  (not A166) );
 a11327a <=( a11326a  and  a11323a );
 a11330a <=( A235  and  A201 );
 a11334a <=( A269  and  A266 );
 a11335a <=( (not A265)  and  a11334a );
 a11336a <=( a11335a  and  a11330a );
 a11339a <=( (not A167)  and  (not A169) );
 a11342a <=( A200  and  (not A166) );
 a11343a <=( a11342a  and  a11339a );
 a11346a <=( A235  and  A201 );
 a11350a <=( A269  and  (not A266) );
 a11351a <=( A265  and  a11350a );
 a11352a <=( a11351a  and  a11346a );
 a11355a <=( (not A167)  and  (not A169) );
 a11358a <=( A200  and  (not A166) );
 a11359a <=( a11358a  and  a11355a );
 a11362a <=( A232  and  A201 );
 a11366a <=( A267  and  A265 );
 a11367a <=( A234  and  a11366a );
 a11368a <=( a11367a  and  a11362a );
 a11371a <=( (not A167)  and  (not A169) );
 a11374a <=( A200  and  (not A166) );
 a11375a <=( a11374a  and  a11371a );
 a11378a <=( A232  and  A201 );
 a11382a <=( A267  and  A266 );
 a11383a <=( A234  and  a11382a );
 a11384a <=( a11383a  and  a11378a );
 a11387a <=( (not A167)  and  (not A169) );
 a11390a <=( A200  and  (not A166) );
 a11391a <=( a11390a  and  a11387a );
 a11394a <=( A233  and  A201 );
 a11398a <=( A267  and  A265 );
 a11399a <=( A234  and  a11398a );
 a11400a <=( a11399a  and  a11394a );
 a11403a <=( (not A167)  and  (not A169) );
 a11406a <=( A200  and  (not A166) );
 a11407a <=( a11406a  and  a11403a );
 a11410a <=( A233  and  A201 );
 a11414a <=( A267  and  A266 );
 a11415a <=( A234  and  a11414a );
 a11416a <=( a11415a  and  a11410a );
 a11419a <=( (not A167)  and  (not A169) );
 a11422a <=( A200  and  (not A166) );
 a11423a <=( a11422a  and  a11419a );
 a11426a <=( (not A232)  and  A201 );
 a11430a <=( A268  and  A236 );
 a11431a <=( A233  and  a11430a );
 a11432a <=( a11431a  and  a11426a );
 a11435a <=( (not A167)  and  (not A169) );
 a11438a <=( A200  and  (not A166) );
 a11439a <=( a11438a  and  a11435a );
 a11442a <=( A232  and  A201 );
 a11446a <=( A268  and  A236 );
 a11447a <=( (not A233)  and  a11446a );
 a11448a <=( a11447a  and  a11442a );
 a11451a <=( (not A167)  and  (not A169) );
 a11454a <=( (not A199)  and  (not A166) );
 a11455a <=( a11454a  and  a11451a );
 a11458a <=( A203  and  A200 );
 a11462a <=( A267  and  A265 );
 a11463a <=( A235  and  a11462a );
 a11464a <=( a11463a  and  a11458a );
 a11467a <=( (not A167)  and  (not A169) );
 a11470a <=( (not A199)  and  (not A166) );
 a11471a <=( a11470a  and  a11467a );
 a11474a <=( A203  and  A200 );
 a11478a <=( A267  and  A266 );
 a11479a <=( A235  and  a11478a );
 a11480a <=( a11479a  and  a11474a );
 a11483a <=( (not A167)  and  (not A169) );
 a11486a <=( (not A199)  and  (not A166) );
 a11487a <=( a11486a  and  a11483a );
 a11490a <=( A203  and  A200 );
 a11494a <=( A268  and  A234 );
 a11495a <=( A232  and  a11494a );
 a11496a <=( a11495a  and  a11490a );
 a11499a <=( (not A167)  and  (not A169) );
 a11502a <=( (not A199)  and  (not A166) );
 a11503a <=( a11502a  and  a11499a );
 a11506a <=( A203  and  A200 );
 a11510a <=( A268  and  A234 );
 a11511a <=( A233  and  a11510a );
 a11512a <=( a11511a  and  a11506a );
 a11515a <=( (not A167)  and  (not A169) );
 a11518a <=( A199  and  (not A166) );
 a11519a <=( a11518a  and  a11515a );
 a11522a <=( A203  and  (not A200) );
 a11526a <=( A267  and  A265 );
 a11527a <=( A235  and  a11526a );
 a11528a <=( a11527a  and  a11522a );
 a11531a <=( (not A167)  and  (not A169) );
 a11534a <=( A199  and  (not A166) );
 a11535a <=( a11534a  and  a11531a );
 a11538a <=( A203  and  (not A200) );
 a11542a <=( A267  and  A266 );
 a11543a <=( A235  and  a11542a );
 a11544a <=( a11543a  and  a11538a );
 a11547a <=( (not A167)  and  (not A169) );
 a11550a <=( A199  and  (not A166) );
 a11551a <=( a11550a  and  a11547a );
 a11554a <=( A203  and  (not A200) );
 a11558a <=( A268  and  A234 );
 a11559a <=( A232  and  a11558a );
 a11560a <=( a11559a  and  a11554a );
 a11563a <=( (not A167)  and  (not A169) );
 a11566a <=( A199  and  (not A166) );
 a11567a <=( a11566a  and  a11563a );
 a11570a <=( A203  and  (not A200) );
 a11574a <=( A268  and  A234 );
 a11575a <=( A233  and  a11574a );
 a11576a <=( a11575a  and  a11570a );
 a11579a <=( (not A168)  and  (not A169) );
 a11582a <=( A166  and  A167 );
 a11583a <=( a11582a  and  a11579a );
 a11586a <=( A235  and  A202 );
 a11590a <=( (not A302)  and  (not A301) );
 a11591a <=( (not A300)  and  a11590a );
 a11592a <=( a11591a  and  a11586a );
 a11595a <=( (not A168)  and  (not A169) );
 a11598a <=( A166  and  A167 );
 a11599a <=( a11598a  and  a11595a );
 a11602a <=( A235  and  A202 );
 a11606a <=( (not A301)  and  (not A299) );
 a11607a <=( (not A298)  and  a11606a );
 a11608a <=( a11607a  and  a11602a );
 a11611a <=( (not A168)  and  (not A169) );
 a11614a <=( A166  and  A167 );
 a11615a <=( a11614a  and  a11611a );
 a11618a <=( A235  and  A202 );
 a11622a <=( A269  and  A266 );
 a11623a <=( (not A265)  and  a11622a );
 a11624a <=( a11623a  and  a11618a );
 a11627a <=( (not A168)  and  (not A169) );
 a11630a <=( A166  and  A167 );
 a11631a <=( a11630a  and  a11627a );
 a11634a <=( A235  and  A202 );
 a11638a <=( A269  and  (not A266) );
 a11639a <=( A265  and  a11638a );
 a11640a <=( a11639a  and  a11634a );
 a11643a <=( (not A168)  and  (not A169) );
 a11646a <=( A166  and  A167 );
 a11647a <=( a11646a  and  a11643a );
 a11650a <=( A232  and  A202 );
 a11654a <=( A267  and  A265 );
 a11655a <=( A234  and  a11654a );
 a11656a <=( a11655a  and  a11650a );
 a11659a <=( (not A168)  and  (not A169) );
 a11662a <=( A166  and  A167 );
 a11663a <=( a11662a  and  a11659a );
 a11666a <=( A232  and  A202 );
 a11670a <=( A267  and  A266 );
 a11671a <=( A234  and  a11670a );
 a11672a <=( a11671a  and  a11666a );
 a11675a <=( (not A168)  and  (not A169) );
 a11678a <=( A166  and  A167 );
 a11679a <=( a11678a  and  a11675a );
 a11682a <=( A233  and  A202 );
 a11686a <=( A267  and  A265 );
 a11687a <=( A234  and  a11686a );
 a11688a <=( a11687a  and  a11682a );
 a11691a <=( (not A168)  and  (not A169) );
 a11694a <=( A166  and  A167 );
 a11695a <=( a11694a  and  a11691a );
 a11698a <=( A233  and  A202 );
 a11702a <=( A267  and  A266 );
 a11703a <=( A234  and  a11702a );
 a11704a <=( a11703a  and  a11698a );
 a11707a <=( (not A168)  and  (not A169) );
 a11710a <=( A166  and  A167 );
 a11711a <=( a11710a  and  a11707a );
 a11714a <=( (not A232)  and  A202 );
 a11718a <=( A268  and  A236 );
 a11719a <=( A233  and  a11718a );
 a11720a <=( a11719a  and  a11714a );
 a11723a <=( (not A168)  and  (not A169) );
 a11726a <=( A166  and  A167 );
 a11727a <=( a11726a  and  a11723a );
 a11730a <=( A232  and  A202 );
 a11734a <=( A268  and  A236 );
 a11735a <=( (not A233)  and  a11734a );
 a11736a <=( a11735a  and  a11730a );
 a11739a <=( (not A168)  and  (not A169) );
 a11742a <=( A166  and  A167 );
 a11743a <=( a11742a  and  a11739a );
 a11746a <=( A201  and  A199 );
 a11750a <=( A267  and  A265 );
 a11751a <=( A235  and  a11750a );
 a11752a <=( a11751a  and  a11746a );
 a11755a <=( (not A168)  and  (not A169) );
 a11758a <=( A166  and  A167 );
 a11759a <=( a11758a  and  a11755a );
 a11762a <=( A201  and  A199 );
 a11766a <=( A267  and  A266 );
 a11767a <=( A235  and  a11766a );
 a11768a <=( a11767a  and  a11762a );
 a11771a <=( (not A168)  and  (not A169) );
 a11774a <=( A166  and  A167 );
 a11775a <=( a11774a  and  a11771a );
 a11778a <=( A201  and  A199 );
 a11782a <=( A268  and  A234 );
 a11783a <=( A232  and  a11782a );
 a11784a <=( a11783a  and  a11778a );
 a11787a <=( (not A168)  and  (not A169) );
 a11790a <=( A166  and  A167 );
 a11791a <=( a11790a  and  a11787a );
 a11794a <=( A201  and  A199 );
 a11798a <=( A268  and  A234 );
 a11799a <=( A233  and  a11798a );
 a11800a <=( a11799a  and  a11794a );
 a11803a <=( (not A168)  and  (not A169) );
 a11806a <=( A166  and  A167 );
 a11807a <=( a11806a  and  a11803a );
 a11810a <=( A201  and  A200 );
 a11814a <=( A267  and  A265 );
 a11815a <=( A235  and  a11814a );
 a11816a <=( a11815a  and  a11810a );
 a11819a <=( (not A168)  and  (not A169) );
 a11822a <=( A166  and  A167 );
 a11823a <=( a11822a  and  a11819a );
 a11826a <=( A201  and  A200 );
 a11830a <=( A267  and  A266 );
 a11831a <=( A235  and  a11830a );
 a11832a <=( a11831a  and  a11826a );
 a11835a <=( (not A168)  and  (not A169) );
 a11838a <=( A166  and  A167 );
 a11839a <=( a11838a  and  a11835a );
 a11842a <=( A201  and  A200 );
 a11846a <=( A268  and  A234 );
 a11847a <=( A232  and  a11846a );
 a11848a <=( a11847a  and  a11842a );
 a11851a <=( (not A168)  and  (not A169) );
 a11854a <=( A166  and  A167 );
 a11855a <=( a11854a  and  a11851a );
 a11858a <=( A201  and  A200 );
 a11862a <=( A268  and  A234 );
 a11863a <=( A233  and  a11862a );
 a11864a <=( a11863a  and  a11858a );
 a11867a <=( (not A168)  and  (not A169) );
 a11870a <=( A166  and  A167 );
 a11871a <=( a11870a  and  a11867a );
 a11874a <=( A200  and  (not A199) );
 a11878a <=( A268  and  A235 );
 a11879a <=( A203  and  a11878a );
 a11880a <=( a11879a  and  a11874a );
 a11883a <=( (not A168)  and  (not A169) );
 a11886a <=( A166  and  A167 );
 a11887a <=( a11886a  and  a11883a );
 a11890a <=( (not A200)  and  A199 );
 a11894a <=( A268  and  A235 );
 a11895a <=( A203  and  a11894a );
 a11896a <=( a11895a  and  a11890a );
 a11899a <=( (not A169)  and  (not A170) );
 a11902a <=( A202  and  (not A168) );
 a11903a <=( a11902a  and  a11899a );
 a11906a <=( A298  and  A235 );
 a11910a <=( (not A301)  and  (not A300) );
 a11911a <=( A299  and  a11910a );
 a11912a <=( a11911a  and  a11906a );
 a11915a <=( (not A169)  and  (not A170) );
 a11918a <=( A202  and  (not A168) );
 a11919a <=( a11918a  and  a11915a );
 a11922a <=( A234  and  A232 );
 a11926a <=( (not A302)  and  (not A301) );
 a11927a <=( (not A300)  and  a11926a );
 a11928a <=( a11927a  and  a11922a );
 a11931a <=( (not A169)  and  (not A170) );
 a11934a <=( A202  and  (not A168) );
 a11935a <=( a11934a  and  a11931a );
 a11938a <=( A234  and  A232 );
 a11942a <=( (not A301)  and  (not A299) );
 a11943a <=( (not A298)  and  a11942a );
 a11944a <=( a11943a  and  a11938a );
 a11947a <=( (not A169)  and  (not A170) );
 a11950a <=( A202  and  (not A168) );
 a11951a <=( a11950a  and  a11947a );
 a11954a <=( A234  and  A232 );
 a11958a <=( A269  and  A266 );
 a11959a <=( (not A265)  and  a11958a );
 a11960a <=( a11959a  and  a11954a );
 a11963a <=( (not A169)  and  (not A170) );
 a11966a <=( A202  and  (not A168) );
 a11967a <=( a11966a  and  a11963a );
 a11970a <=( A234  and  A232 );
 a11974a <=( A269  and  (not A266) );
 a11975a <=( A265  and  a11974a );
 a11976a <=( a11975a  and  a11970a );
 a11979a <=( (not A169)  and  (not A170) );
 a11982a <=( A202  and  (not A168) );
 a11983a <=( a11982a  and  a11979a );
 a11986a <=( A234  and  A233 );
 a11990a <=( (not A302)  and  (not A301) );
 a11991a <=( (not A300)  and  a11990a );
 a11992a <=( a11991a  and  a11986a );
 a11995a <=( (not A169)  and  (not A170) );
 a11998a <=( A202  and  (not A168) );
 a11999a <=( a11998a  and  a11995a );
 a12002a <=( A234  and  A233 );
 a12006a <=( (not A301)  and  (not A299) );
 a12007a <=( (not A298)  and  a12006a );
 a12008a <=( a12007a  and  a12002a );
 a12011a <=( (not A169)  and  (not A170) );
 a12014a <=( A202  and  (not A168) );
 a12015a <=( a12014a  and  a12011a );
 a12018a <=( A234  and  A233 );
 a12022a <=( A269  and  A266 );
 a12023a <=( (not A265)  and  a12022a );
 a12024a <=( a12023a  and  a12018a );
 a12027a <=( (not A169)  and  (not A170) );
 a12030a <=( A202  and  (not A168) );
 a12031a <=( a12030a  and  a12027a );
 a12034a <=( A234  and  A233 );
 a12038a <=( A269  and  (not A266) );
 a12039a <=( A265  and  a12038a );
 a12040a <=( a12039a  and  a12034a );
 a12043a <=( (not A169)  and  (not A170) );
 a12046a <=( A202  and  (not A168) );
 a12047a <=( a12046a  and  a12043a );
 a12050a <=( A233  and  (not A232) );
 a12054a <=( A267  and  A265 );
 a12055a <=( A236  and  a12054a );
 a12056a <=( a12055a  and  a12050a );
 a12059a <=( (not A169)  and  (not A170) );
 a12062a <=( A202  and  (not A168) );
 a12063a <=( a12062a  and  a12059a );
 a12066a <=( A233  and  (not A232) );
 a12070a <=( A267  and  A266 );
 a12071a <=( A236  and  a12070a );
 a12072a <=( a12071a  and  a12066a );
 a12075a <=( (not A169)  and  (not A170) );
 a12078a <=( A202  and  (not A168) );
 a12079a <=( a12078a  and  a12075a );
 a12082a <=( (not A233)  and  A232 );
 a12086a <=( A267  and  A265 );
 a12087a <=( A236  and  a12086a );
 a12088a <=( a12087a  and  a12082a );
 a12091a <=( (not A169)  and  (not A170) );
 a12094a <=( A202  and  (not A168) );
 a12095a <=( a12094a  and  a12091a );
 a12098a <=( (not A233)  and  A232 );
 a12102a <=( A267  and  A266 );
 a12103a <=( A236  and  a12102a );
 a12104a <=( a12103a  and  a12098a );
 a12107a <=( (not A169)  and  (not A170) );
 a12110a <=( A199  and  (not A168) );
 a12111a <=( a12110a  and  a12107a );
 a12114a <=( A235  and  A201 );
 a12118a <=( (not A302)  and  (not A301) );
 a12119a <=( (not A300)  and  a12118a );
 a12120a <=( a12119a  and  a12114a );
 a12123a <=( (not A169)  and  (not A170) );
 a12126a <=( A199  and  (not A168) );
 a12127a <=( a12126a  and  a12123a );
 a12130a <=( A235  and  A201 );
 a12134a <=( (not A301)  and  (not A299) );
 a12135a <=( (not A298)  and  a12134a );
 a12136a <=( a12135a  and  a12130a );
 a12139a <=( (not A169)  and  (not A170) );
 a12142a <=( A199  and  (not A168) );
 a12143a <=( a12142a  and  a12139a );
 a12146a <=( A235  and  A201 );
 a12150a <=( A269  and  A266 );
 a12151a <=( (not A265)  and  a12150a );
 a12152a <=( a12151a  and  a12146a );
 a12155a <=( (not A169)  and  (not A170) );
 a12158a <=( A199  and  (not A168) );
 a12159a <=( a12158a  and  a12155a );
 a12162a <=( A235  and  A201 );
 a12166a <=( A269  and  (not A266) );
 a12167a <=( A265  and  a12166a );
 a12168a <=( a12167a  and  a12162a );
 a12171a <=( (not A169)  and  (not A170) );
 a12174a <=( A199  and  (not A168) );
 a12175a <=( a12174a  and  a12171a );
 a12178a <=( A232  and  A201 );
 a12182a <=( A267  and  A265 );
 a12183a <=( A234  and  a12182a );
 a12184a <=( a12183a  and  a12178a );
 a12187a <=( (not A169)  and  (not A170) );
 a12190a <=( A199  and  (not A168) );
 a12191a <=( a12190a  and  a12187a );
 a12194a <=( A232  and  A201 );
 a12198a <=( A267  and  A266 );
 a12199a <=( A234  and  a12198a );
 a12200a <=( a12199a  and  a12194a );
 a12203a <=( (not A169)  and  (not A170) );
 a12206a <=( A199  and  (not A168) );
 a12207a <=( a12206a  and  a12203a );
 a12210a <=( A233  and  A201 );
 a12214a <=( A267  and  A265 );
 a12215a <=( A234  and  a12214a );
 a12216a <=( a12215a  and  a12210a );
 a12219a <=( (not A169)  and  (not A170) );
 a12222a <=( A199  and  (not A168) );
 a12223a <=( a12222a  and  a12219a );
 a12226a <=( A233  and  A201 );
 a12230a <=( A267  and  A266 );
 a12231a <=( A234  and  a12230a );
 a12232a <=( a12231a  and  a12226a );
 a12235a <=( (not A169)  and  (not A170) );
 a12238a <=( A199  and  (not A168) );
 a12239a <=( a12238a  and  a12235a );
 a12242a <=( (not A232)  and  A201 );
 a12246a <=( A268  and  A236 );
 a12247a <=( A233  and  a12246a );
 a12248a <=( a12247a  and  a12242a );
 a12251a <=( (not A169)  and  (not A170) );
 a12254a <=( A199  and  (not A168) );
 a12255a <=( a12254a  and  a12251a );
 a12258a <=( A232  and  A201 );
 a12262a <=( A268  and  A236 );
 a12263a <=( (not A233)  and  a12262a );
 a12264a <=( a12263a  and  a12258a );
 a12267a <=( (not A169)  and  (not A170) );
 a12270a <=( A200  and  (not A168) );
 a12271a <=( a12270a  and  a12267a );
 a12274a <=( A235  and  A201 );
 a12278a <=( (not A302)  and  (not A301) );
 a12279a <=( (not A300)  and  a12278a );
 a12280a <=( a12279a  and  a12274a );
 a12283a <=( (not A169)  and  (not A170) );
 a12286a <=( A200  and  (not A168) );
 a12287a <=( a12286a  and  a12283a );
 a12290a <=( A235  and  A201 );
 a12294a <=( (not A301)  and  (not A299) );
 a12295a <=( (not A298)  and  a12294a );
 a12296a <=( a12295a  and  a12290a );
 a12299a <=( (not A169)  and  (not A170) );
 a12302a <=( A200  and  (not A168) );
 a12303a <=( a12302a  and  a12299a );
 a12306a <=( A235  and  A201 );
 a12310a <=( A269  and  A266 );
 a12311a <=( (not A265)  and  a12310a );
 a12312a <=( a12311a  and  a12306a );
 a12315a <=( (not A169)  and  (not A170) );
 a12318a <=( A200  and  (not A168) );
 a12319a <=( a12318a  and  a12315a );
 a12322a <=( A235  and  A201 );
 a12326a <=( A269  and  (not A266) );
 a12327a <=( A265  and  a12326a );
 a12328a <=( a12327a  and  a12322a );
 a12331a <=( (not A169)  and  (not A170) );
 a12334a <=( A200  and  (not A168) );
 a12335a <=( a12334a  and  a12331a );
 a12338a <=( A232  and  A201 );
 a12342a <=( A267  and  A265 );
 a12343a <=( A234  and  a12342a );
 a12344a <=( a12343a  and  a12338a );
 a12347a <=( (not A169)  and  (not A170) );
 a12350a <=( A200  and  (not A168) );
 a12351a <=( a12350a  and  a12347a );
 a12354a <=( A232  and  A201 );
 a12358a <=( A267  and  A266 );
 a12359a <=( A234  and  a12358a );
 a12360a <=( a12359a  and  a12354a );
 a12363a <=( (not A169)  and  (not A170) );
 a12366a <=( A200  and  (not A168) );
 a12367a <=( a12366a  and  a12363a );
 a12370a <=( A233  and  A201 );
 a12374a <=( A267  and  A265 );
 a12375a <=( A234  and  a12374a );
 a12376a <=( a12375a  and  a12370a );
 a12379a <=( (not A169)  and  (not A170) );
 a12382a <=( A200  and  (not A168) );
 a12383a <=( a12382a  and  a12379a );
 a12386a <=( A233  and  A201 );
 a12390a <=( A267  and  A266 );
 a12391a <=( A234  and  a12390a );
 a12392a <=( a12391a  and  a12386a );
 a12395a <=( (not A169)  and  (not A170) );
 a12398a <=( A200  and  (not A168) );
 a12399a <=( a12398a  and  a12395a );
 a12402a <=( (not A232)  and  A201 );
 a12406a <=( A268  and  A236 );
 a12407a <=( A233  and  a12406a );
 a12408a <=( a12407a  and  a12402a );
 a12411a <=( (not A169)  and  (not A170) );
 a12414a <=( A200  and  (not A168) );
 a12415a <=( a12414a  and  a12411a );
 a12418a <=( A232  and  A201 );
 a12422a <=( A268  and  A236 );
 a12423a <=( (not A233)  and  a12422a );
 a12424a <=( a12423a  and  a12418a );
 a12427a <=( (not A169)  and  (not A170) );
 a12430a <=( (not A199)  and  (not A168) );
 a12431a <=( a12430a  and  a12427a );
 a12434a <=( A203  and  A200 );
 a12438a <=( A267  and  A265 );
 a12439a <=( A235  and  a12438a );
 a12440a <=( a12439a  and  a12434a );
 a12443a <=( (not A169)  and  (not A170) );
 a12446a <=( (not A199)  and  (not A168) );
 a12447a <=( a12446a  and  a12443a );
 a12450a <=( A203  and  A200 );
 a12454a <=( A267  and  A266 );
 a12455a <=( A235  and  a12454a );
 a12456a <=( a12455a  and  a12450a );
 a12459a <=( (not A169)  and  (not A170) );
 a12462a <=( (not A199)  and  (not A168) );
 a12463a <=( a12462a  and  a12459a );
 a12466a <=( A203  and  A200 );
 a12470a <=( A268  and  A234 );
 a12471a <=( A232  and  a12470a );
 a12472a <=( a12471a  and  a12466a );
 a12475a <=( (not A169)  and  (not A170) );
 a12478a <=( (not A199)  and  (not A168) );
 a12479a <=( a12478a  and  a12475a );
 a12482a <=( A203  and  A200 );
 a12486a <=( A268  and  A234 );
 a12487a <=( A233  and  a12486a );
 a12488a <=( a12487a  and  a12482a );
 a12491a <=( (not A169)  and  (not A170) );
 a12494a <=( A199  and  (not A168) );
 a12495a <=( a12494a  and  a12491a );
 a12498a <=( A203  and  (not A200) );
 a12502a <=( A267  and  A265 );
 a12503a <=( A235  and  a12502a );
 a12504a <=( a12503a  and  a12498a );
 a12507a <=( (not A169)  and  (not A170) );
 a12510a <=( A199  and  (not A168) );
 a12511a <=( a12510a  and  a12507a );
 a12514a <=( A203  and  (not A200) );
 a12518a <=( A267  and  A266 );
 a12519a <=( A235  and  a12518a );
 a12520a <=( a12519a  and  a12514a );
 a12523a <=( (not A169)  and  (not A170) );
 a12526a <=( A199  and  (not A168) );
 a12527a <=( a12526a  and  a12523a );
 a12530a <=( A203  and  (not A200) );
 a12534a <=( A268  and  A234 );
 a12535a <=( A232  and  a12534a );
 a12536a <=( a12535a  and  a12530a );
 a12539a <=( (not A169)  and  (not A170) );
 a12542a <=( A199  and  (not A168) );
 a12543a <=( a12542a  and  a12539a );
 a12546a <=( A203  and  (not A200) );
 a12550a <=( A268  and  A234 );
 a12551a <=( A233  and  a12550a );
 a12552a <=( a12551a  and  a12546a );
 a12555a <=( A166  and  A168 );
 a12559a <=( (not A203)  and  (not A202) );
 a12560a <=( (not A201)  and  a12559a );
 a12561a <=( a12560a  and  a12555a );
 a12564a <=( A298  and  A235 );
 a12568a <=( (not A301)  and  (not A300) );
 a12569a <=( A299  and  a12568a );
 a12570a <=( a12569a  and  a12564a );
 a12573a <=( A166  and  A168 );
 a12577a <=( (not A203)  and  (not A202) );
 a12578a <=( (not A201)  and  a12577a );
 a12579a <=( a12578a  and  a12573a );
 a12582a <=( A234  and  A232 );
 a12586a <=( (not A302)  and  (not A301) );
 a12587a <=( (not A300)  and  a12586a );
 a12588a <=( a12587a  and  a12582a );
 a12591a <=( A166  and  A168 );
 a12595a <=( (not A203)  and  (not A202) );
 a12596a <=( (not A201)  and  a12595a );
 a12597a <=( a12596a  and  a12591a );
 a12600a <=( A234  and  A232 );
 a12604a <=( (not A301)  and  (not A299) );
 a12605a <=( (not A298)  and  a12604a );
 a12606a <=( a12605a  and  a12600a );
 a12609a <=( A166  and  A168 );
 a12613a <=( (not A203)  and  (not A202) );
 a12614a <=( (not A201)  and  a12613a );
 a12615a <=( a12614a  and  a12609a );
 a12618a <=( A234  and  A232 );
 a12622a <=( A269  and  A266 );
 a12623a <=( (not A265)  and  a12622a );
 a12624a <=( a12623a  and  a12618a );
 a12627a <=( A166  and  A168 );
 a12631a <=( (not A203)  and  (not A202) );
 a12632a <=( (not A201)  and  a12631a );
 a12633a <=( a12632a  and  a12627a );
 a12636a <=( A234  and  A232 );
 a12640a <=( A269  and  (not A266) );
 a12641a <=( A265  and  a12640a );
 a12642a <=( a12641a  and  a12636a );
 a12645a <=( A166  and  A168 );
 a12649a <=( (not A203)  and  (not A202) );
 a12650a <=( (not A201)  and  a12649a );
 a12651a <=( a12650a  and  a12645a );
 a12654a <=( A234  and  A233 );
 a12658a <=( (not A302)  and  (not A301) );
 a12659a <=( (not A300)  and  a12658a );
 a12660a <=( a12659a  and  a12654a );
 a12663a <=( A166  and  A168 );
 a12667a <=( (not A203)  and  (not A202) );
 a12668a <=( (not A201)  and  a12667a );
 a12669a <=( a12668a  and  a12663a );
 a12672a <=( A234  and  A233 );
 a12676a <=( (not A301)  and  (not A299) );
 a12677a <=( (not A298)  and  a12676a );
 a12678a <=( a12677a  and  a12672a );
 a12681a <=( A166  and  A168 );
 a12685a <=( (not A203)  and  (not A202) );
 a12686a <=( (not A201)  and  a12685a );
 a12687a <=( a12686a  and  a12681a );
 a12690a <=( A234  and  A233 );
 a12694a <=( A269  and  A266 );
 a12695a <=( (not A265)  and  a12694a );
 a12696a <=( a12695a  and  a12690a );
 a12699a <=( A166  and  A168 );
 a12703a <=( (not A203)  and  (not A202) );
 a12704a <=( (not A201)  and  a12703a );
 a12705a <=( a12704a  and  a12699a );
 a12708a <=( A234  and  A233 );
 a12712a <=( A269  and  (not A266) );
 a12713a <=( A265  and  a12712a );
 a12714a <=( a12713a  and  a12708a );
 a12717a <=( A166  and  A168 );
 a12721a <=( (not A203)  and  (not A202) );
 a12722a <=( (not A201)  and  a12721a );
 a12723a <=( a12722a  and  a12717a );
 a12726a <=( A233  and  (not A232) );
 a12730a <=( A267  and  A265 );
 a12731a <=( A236  and  a12730a );
 a12732a <=( a12731a  and  a12726a );
 a12735a <=( A166  and  A168 );
 a12739a <=( (not A203)  and  (not A202) );
 a12740a <=( (not A201)  and  a12739a );
 a12741a <=( a12740a  and  a12735a );
 a12744a <=( A233  and  (not A232) );
 a12748a <=( A267  and  A266 );
 a12749a <=( A236  and  a12748a );
 a12750a <=( a12749a  and  a12744a );
 a12753a <=( A166  and  A168 );
 a12757a <=( (not A203)  and  (not A202) );
 a12758a <=( (not A201)  and  a12757a );
 a12759a <=( a12758a  and  a12753a );
 a12762a <=( (not A233)  and  A232 );
 a12766a <=( A267  and  A265 );
 a12767a <=( A236  and  a12766a );
 a12768a <=( a12767a  and  a12762a );
 a12771a <=( A166  and  A168 );
 a12775a <=( (not A203)  and  (not A202) );
 a12776a <=( (not A201)  and  a12775a );
 a12777a <=( a12776a  and  a12771a );
 a12780a <=( (not A233)  and  A232 );
 a12784a <=( A267  and  A266 );
 a12785a <=( A236  and  a12784a );
 a12786a <=( a12785a  and  a12780a );
 a12789a <=( A166  and  A168 );
 a12793a <=( (not A201)  and  A200 );
 a12794a <=( A199  and  a12793a );
 a12795a <=( a12794a  and  a12789a );
 a12798a <=( A235  and  (not A202) );
 a12802a <=( (not A302)  and  (not A301) );
 a12803a <=( (not A300)  and  a12802a );
 a12804a <=( a12803a  and  a12798a );
 a12807a <=( A166  and  A168 );
 a12811a <=( (not A201)  and  A200 );
 a12812a <=( A199  and  a12811a );
 a12813a <=( a12812a  and  a12807a );
 a12816a <=( A235  and  (not A202) );
 a12820a <=( (not A301)  and  (not A299) );
 a12821a <=( (not A298)  and  a12820a );
 a12822a <=( a12821a  and  a12816a );
 a12825a <=( A166  and  A168 );
 a12829a <=( (not A201)  and  A200 );
 a12830a <=( A199  and  a12829a );
 a12831a <=( a12830a  and  a12825a );
 a12834a <=( A235  and  (not A202) );
 a12838a <=( A269  and  A266 );
 a12839a <=( (not A265)  and  a12838a );
 a12840a <=( a12839a  and  a12834a );
 a12843a <=( A166  and  A168 );
 a12847a <=( (not A201)  and  A200 );
 a12848a <=( A199  and  a12847a );
 a12849a <=( a12848a  and  a12843a );
 a12852a <=( A235  and  (not A202) );
 a12856a <=( A269  and  (not A266) );
 a12857a <=( A265  and  a12856a );
 a12858a <=( a12857a  and  a12852a );
 a12861a <=( A166  and  A168 );
 a12865a <=( (not A201)  and  A200 );
 a12866a <=( A199  and  a12865a );
 a12867a <=( a12866a  and  a12861a );
 a12870a <=( A232  and  (not A202) );
 a12874a <=( A267  and  A265 );
 a12875a <=( A234  and  a12874a );
 a12876a <=( a12875a  and  a12870a );
 a12879a <=( A166  and  A168 );
 a12883a <=( (not A201)  and  A200 );
 a12884a <=( A199  and  a12883a );
 a12885a <=( a12884a  and  a12879a );
 a12888a <=( A232  and  (not A202) );
 a12892a <=( A267  and  A266 );
 a12893a <=( A234  and  a12892a );
 a12894a <=( a12893a  and  a12888a );
 a12897a <=( A166  and  A168 );
 a12901a <=( (not A201)  and  A200 );
 a12902a <=( A199  and  a12901a );
 a12903a <=( a12902a  and  a12897a );
 a12906a <=( A233  and  (not A202) );
 a12910a <=( A267  and  A265 );
 a12911a <=( A234  and  a12910a );
 a12912a <=( a12911a  and  a12906a );
 a12915a <=( A166  and  A168 );
 a12919a <=( (not A201)  and  A200 );
 a12920a <=( A199  and  a12919a );
 a12921a <=( a12920a  and  a12915a );
 a12924a <=( A233  and  (not A202) );
 a12928a <=( A267  and  A266 );
 a12929a <=( A234  and  a12928a );
 a12930a <=( a12929a  and  a12924a );
 a12933a <=( A166  and  A168 );
 a12937a <=( (not A201)  and  A200 );
 a12938a <=( A199  and  a12937a );
 a12939a <=( a12938a  and  a12933a );
 a12942a <=( (not A232)  and  (not A202) );
 a12946a <=( A268  and  A236 );
 a12947a <=( A233  and  a12946a );
 a12948a <=( a12947a  and  a12942a );
 a12951a <=( A166  and  A168 );
 a12955a <=( (not A201)  and  A200 );
 a12956a <=( A199  and  a12955a );
 a12957a <=( a12956a  and  a12951a );
 a12960a <=( A232  and  (not A202) );
 a12964a <=( A268  and  A236 );
 a12965a <=( (not A233)  and  a12964a );
 a12966a <=( a12965a  and  a12960a );
 a12969a <=( A166  and  A168 );
 a12973a <=( (not A202)  and  (not A200) );
 a12974a <=( (not A199)  and  a12973a );
 a12975a <=( a12974a  and  a12969a );
 a12978a <=( A298  and  A235 );
 a12982a <=( (not A301)  and  (not A300) );
 a12983a <=( A299  and  a12982a );
 a12984a <=( a12983a  and  a12978a );
 a12987a <=( A166  and  A168 );
 a12991a <=( (not A202)  and  (not A200) );
 a12992a <=( (not A199)  and  a12991a );
 a12993a <=( a12992a  and  a12987a );
 a12996a <=( A234  and  A232 );
 a13000a <=( (not A302)  and  (not A301) );
 a13001a <=( (not A300)  and  a13000a );
 a13002a <=( a13001a  and  a12996a );
 a13005a <=( A166  and  A168 );
 a13009a <=( (not A202)  and  (not A200) );
 a13010a <=( (not A199)  and  a13009a );
 a13011a <=( a13010a  and  a13005a );
 a13014a <=( A234  and  A232 );
 a13018a <=( (not A301)  and  (not A299) );
 a13019a <=( (not A298)  and  a13018a );
 a13020a <=( a13019a  and  a13014a );
 a13023a <=( A166  and  A168 );
 a13027a <=( (not A202)  and  (not A200) );
 a13028a <=( (not A199)  and  a13027a );
 a13029a <=( a13028a  and  a13023a );
 a13032a <=( A234  and  A232 );
 a13036a <=( A269  and  A266 );
 a13037a <=( (not A265)  and  a13036a );
 a13038a <=( a13037a  and  a13032a );
 a13041a <=( A166  and  A168 );
 a13045a <=( (not A202)  and  (not A200) );
 a13046a <=( (not A199)  and  a13045a );
 a13047a <=( a13046a  and  a13041a );
 a13050a <=( A234  and  A232 );
 a13054a <=( A269  and  (not A266) );
 a13055a <=( A265  and  a13054a );
 a13056a <=( a13055a  and  a13050a );
 a13059a <=( A166  and  A168 );
 a13063a <=( (not A202)  and  (not A200) );
 a13064a <=( (not A199)  and  a13063a );
 a13065a <=( a13064a  and  a13059a );
 a13068a <=( A234  and  A233 );
 a13072a <=( (not A302)  and  (not A301) );
 a13073a <=( (not A300)  and  a13072a );
 a13074a <=( a13073a  and  a13068a );
 a13077a <=( A166  and  A168 );
 a13081a <=( (not A202)  and  (not A200) );
 a13082a <=( (not A199)  and  a13081a );
 a13083a <=( a13082a  and  a13077a );
 a13086a <=( A234  and  A233 );
 a13090a <=( (not A301)  and  (not A299) );
 a13091a <=( (not A298)  and  a13090a );
 a13092a <=( a13091a  and  a13086a );
 a13095a <=( A166  and  A168 );
 a13099a <=( (not A202)  and  (not A200) );
 a13100a <=( (not A199)  and  a13099a );
 a13101a <=( a13100a  and  a13095a );
 a13104a <=( A234  and  A233 );
 a13108a <=( A269  and  A266 );
 a13109a <=( (not A265)  and  a13108a );
 a13110a <=( a13109a  and  a13104a );
 a13113a <=( A166  and  A168 );
 a13117a <=( (not A202)  and  (not A200) );
 a13118a <=( (not A199)  and  a13117a );
 a13119a <=( a13118a  and  a13113a );
 a13122a <=( A234  and  A233 );
 a13126a <=( A269  and  (not A266) );
 a13127a <=( A265  and  a13126a );
 a13128a <=( a13127a  and  a13122a );
 a13131a <=( A166  and  A168 );
 a13135a <=( (not A202)  and  (not A200) );
 a13136a <=( (not A199)  and  a13135a );
 a13137a <=( a13136a  and  a13131a );
 a13140a <=( A233  and  (not A232) );
 a13144a <=( A267  and  A265 );
 a13145a <=( A236  and  a13144a );
 a13146a <=( a13145a  and  a13140a );
 a13149a <=( A166  and  A168 );
 a13153a <=( (not A202)  and  (not A200) );
 a13154a <=( (not A199)  and  a13153a );
 a13155a <=( a13154a  and  a13149a );
 a13158a <=( A233  and  (not A232) );
 a13162a <=( A267  and  A266 );
 a13163a <=( A236  and  a13162a );
 a13164a <=( a13163a  and  a13158a );
 a13167a <=( A166  and  A168 );
 a13171a <=( (not A202)  and  (not A200) );
 a13172a <=( (not A199)  and  a13171a );
 a13173a <=( a13172a  and  a13167a );
 a13176a <=( (not A233)  and  A232 );
 a13180a <=( A267  and  A265 );
 a13181a <=( A236  and  a13180a );
 a13182a <=( a13181a  and  a13176a );
 a13185a <=( A166  and  A168 );
 a13189a <=( (not A202)  and  (not A200) );
 a13190a <=( (not A199)  and  a13189a );
 a13191a <=( a13190a  and  a13185a );
 a13194a <=( (not A233)  and  A232 );
 a13198a <=( A267  and  A266 );
 a13199a <=( A236  and  a13198a );
 a13200a <=( a13199a  and  a13194a );
 a13203a <=( A167  and  A168 );
 a13207a <=( (not A203)  and  (not A202) );
 a13208a <=( (not A201)  and  a13207a );
 a13209a <=( a13208a  and  a13203a );
 a13212a <=( A298  and  A235 );
 a13216a <=( (not A301)  and  (not A300) );
 a13217a <=( A299  and  a13216a );
 a13218a <=( a13217a  and  a13212a );
 a13221a <=( A167  and  A168 );
 a13225a <=( (not A203)  and  (not A202) );
 a13226a <=( (not A201)  and  a13225a );
 a13227a <=( a13226a  and  a13221a );
 a13230a <=( A234  and  A232 );
 a13234a <=( (not A302)  and  (not A301) );
 a13235a <=( (not A300)  and  a13234a );
 a13236a <=( a13235a  and  a13230a );
 a13239a <=( A167  and  A168 );
 a13243a <=( (not A203)  and  (not A202) );
 a13244a <=( (not A201)  and  a13243a );
 a13245a <=( a13244a  and  a13239a );
 a13248a <=( A234  and  A232 );
 a13252a <=( (not A301)  and  (not A299) );
 a13253a <=( (not A298)  and  a13252a );
 a13254a <=( a13253a  and  a13248a );
 a13257a <=( A167  and  A168 );
 a13261a <=( (not A203)  and  (not A202) );
 a13262a <=( (not A201)  and  a13261a );
 a13263a <=( a13262a  and  a13257a );
 a13266a <=( A234  and  A232 );
 a13270a <=( A269  and  A266 );
 a13271a <=( (not A265)  and  a13270a );
 a13272a <=( a13271a  and  a13266a );
 a13275a <=( A167  and  A168 );
 a13279a <=( (not A203)  and  (not A202) );
 a13280a <=( (not A201)  and  a13279a );
 a13281a <=( a13280a  and  a13275a );
 a13284a <=( A234  and  A232 );
 a13288a <=( A269  and  (not A266) );
 a13289a <=( A265  and  a13288a );
 a13290a <=( a13289a  and  a13284a );
 a13293a <=( A167  and  A168 );
 a13297a <=( (not A203)  and  (not A202) );
 a13298a <=( (not A201)  and  a13297a );
 a13299a <=( a13298a  and  a13293a );
 a13302a <=( A234  and  A233 );
 a13306a <=( (not A302)  and  (not A301) );
 a13307a <=( (not A300)  and  a13306a );
 a13308a <=( a13307a  and  a13302a );
 a13311a <=( A167  and  A168 );
 a13315a <=( (not A203)  and  (not A202) );
 a13316a <=( (not A201)  and  a13315a );
 a13317a <=( a13316a  and  a13311a );
 a13320a <=( A234  and  A233 );
 a13324a <=( (not A301)  and  (not A299) );
 a13325a <=( (not A298)  and  a13324a );
 a13326a <=( a13325a  and  a13320a );
 a13329a <=( A167  and  A168 );
 a13333a <=( (not A203)  and  (not A202) );
 a13334a <=( (not A201)  and  a13333a );
 a13335a <=( a13334a  and  a13329a );
 a13338a <=( A234  and  A233 );
 a13342a <=( A269  and  A266 );
 a13343a <=( (not A265)  and  a13342a );
 a13344a <=( a13343a  and  a13338a );
 a13347a <=( A167  and  A168 );
 a13351a <=( (not A203)  and  (not A202) );
 a13352a <=( (not A201)  and  a13351a );
 a13353a <=( a13352a  and  a13347a );
 a13356a <=( A234  and  A233 );
 a13360a <=( A269  and  (not A266) );
 a13361a <=( A265  and  a13360a );
 a13362a <=( a13361a  and  a13356a );
 a13365a <=( A167  and  A168 );
 a13369a <=( (not A203)  and  (not A202) );
 a13370a <=( (not A201)  and  a13369a );
 a13371a <=( a13370a  and  a13365a );
 a13374a <=( A233  and  (not A232) );
 a13378a <=( A267  and  A265 );
 a13379a <=( A236  and  a13378a );
 a13380a <=( a13379a  and  a13374a );
 a13383a <=( A167  and  A168 );
 a13387a <=( (not A203)  and  (not A202) );
 a13388a <=( (not A201)  and  a13387a );
 a13389a <=( a13388a  and  a13383a );
 a13392a <=( A233  and  (not A232) );
 a13396a <=( A267  and  A266 );
 a13397a <=( A236  and  a13396a );
 a13398a <=( a13397a  and  a13392a );
 a13401a <=( A167  and  A168 );
 a13405a <=( (not A203)  and  (not A202) );
 a13406a <=( (not A201)  and  a13405a );
 a13407a <=( a13406a  and  a13401a );
 a13410a <=( (not A233)  and  A232 );
 a13414a <=( A267  and  A265 );
 a13415a <=( A236  and  a13414a );
 a13416a <=( a13415a  and  a13410a );
 a13419a <=( A167  and  A168 );
 a13423a <=( (not A203)  and  (not A202) );
 a13424a <=( (not A201)  and  a13423a );
 a13425a <=( a13424a  and  a13419a );
 a13428a <=( (not A233)  and  A232 );
 a13432a <=( A267  and  A266 );
 a13433a <=( A236  and  a13432a );
 a13434a <=( a13433a  and  a13428a );
 a13437a <=( A167  and  A168 );
 a13441a <=( (not A201)  and  A200 );
 a13442a <=( A199  and  a13441a );
 a13443a <=( a13442a  and  a13437a );
 a13446a <=( A235  and  (not A202) );
 a13450a <=( (not A302)  and  (not A301) );
 a13451a <=( (not A300)  and  a13450a );
 a13452a <=( a13451a  and  a13446a );
 a13455a <=( A167  and  A168 );
 a13459a <=( (not A201)  and  A200 );
 a13460a <=( A199  and  a13459a );
 a13461a <=( a13460a  and  a13455a );
 a13464a <=( A235  and  (not A202) );
 a13468a <=( (not A301)  and  (not A299) );
 a13469a <=( (not A298)  and  a13468a );
 a13470a <=( a13469a  and  a13464a );
 a13473a <=( A167  and  A168 );
 a13477a <=( (not A201)  and  A200 );
 a13478a <=( A199  and  a13477a );
 a13479a <=( a13478a  and  a13473a );
 a13482a <=( A235  and  (not A202) );
 a13486a <=( A269  and  A266 );
 a13487a <=( (not A265)  and  a13486a );
 a13488a <=( a13487a  and  a13482a );
 a13491a <=( A167  and  A168 );
 a13495a <=( (not A201)  and  A200 );
 a13496a <=( A199  and  a13495a );
 a13497a <=( a13496a  and  a13491a );
 a13500a <=( A235  and  (not A202) );
 a13504a <=( A269  and  (not A266) );
 a13505a <=( A265  and  a13504a );
 a13506a <=( a13505a  and  a13500a );
 a13509a <=( A167  and  A168 );
 a13513a <=( (not A201)  and  A200 );
 a13514a <=( A199  and  a13513a );
 a13515a <=( a13514a  and  a13509a );
 a13518a <=( A232  and  (not A202) );
 a13522a <=( A267  and  A265 );
 a13523a <=( A234  and  a13522a );
 a13524a <=( a13523a  and  a13518a );
 a13527a <=( A167  and  A168 );
 a13531a <=( (not A201)  and  A200 );
 a13532a <=( A199  and  a13531a );
 a13533a <=( a13532a  and  a13527a );
 a13536a <=( A232  and  (not A202) );
 a13540a <=( A267  and  A266 );
 a13541a <=( A234  and  a13540a );
 a13542a <=( a13541a  and  a13536a );
 a13545a <=( A167  and  A168 );
 a13549a <=( (not A201)  and  A200 );
 a13550a <=( A199  and  a13549a );
 a13551a <=( a13550a  and  a13545a );
 a13554a <=( A233  and  (not A202) );
 a13558a <=( A267  and  A265 );
 a13559a <=( A234  and  a13558a );
 a13560a <=( a13559a  and  a13554a );
 a13563a <=( A167  and  A168 );
 a13567a <=( (not A201)  and  A200 );
 a13568a <=( A199  and  a13567a );
 a13569a <=( a13568a  and  a13563a );
 a13572a <=( A233  and  (not A202) );
 a13576a <=( A267  and  A266 );
 a13577a <=( A234  and  a13576a );
 a13578a <=( a13577a  and  a13572a );
 a13581a <=( A167  and  A168 );
 a13585a <=( (not A201)  and  A200 );
 a13586a <=( A199  and  a13585a );
 a13587a <=( a13586a  and  a13581a );
 a13590a <=( (not A232)  and  (not A202) );
 a13594a <=( A268  and  A236 );
 a13595a <=( A233  and  a13594a );
 a13596a <=( a13595a  and  a13590a );
 a13599a <=( A167  and  A168 );
 a13603a <=( (not A201)  and  A200 );
 a13604a <=( A199  and  a13603a );
 a13605a <=( a13604a  and  a13599a );
 a13608a <=( A232  and  (not A202) );
 a13612a <=( A268  and  A236 );
 a13613a <=( (not A233)  and  a13612a );
 a13614a <=( a13613a  and  a13608a );
 a13617a <=( A167  and  A168 );
 a13621a <=( (not A202)  and  (not A200) );
 a13622a <=( (not A199)  and  a13621a );
 a13623a <=( a13622a  and  a13617a );
 a13626a <=( A298  and  A235 );
 a13630a <=( (not A301)  and  (not A300) );
 a13631a <=( A299  and  a13630a );
 a13632a <=( a13631a  and  a13626a );
 a13635a <=( A167  and  A168 );
 a13639a <=( (not A202)  and  (not A200) );
 a13640a <=( (not A199)  and  a13639a );
 a13641a <=( a13640a  and  a13635a );
 a13644a <=( A234  and  A232 );
 a13648a <=( (not A302)  and  (not A301) );
 a13649a <=( (not A300)  and  a13648a );
 a13650a <=( a13649a  and  a13644a );
 a13653a <=( A167  and  A168 );
 a13657a <=( (not A202)  and  (not A200) );
 a13658a <=( (not A199)  and  a13657a );
 a13659a <=( a13658a  and  a13653a );
 a13662a <=( A234  and  A232 );
 a13666a <=( (not A301)  and  (not A299) );
 a13667a <=( (not A298)  and  a13666a );
 a13668a <=( a13667a  and  a13662a );
 a13671a <=( A167  and  A168 );
 a13675a <=( (not A202)  and  (not A200) );
 a13676a <=( (not A199)  and  a13675a );
 a13677a <=( a13676a  and  a13671a );
 a13680a <=( A234  and  A232 );
 a13684a <=( A269  and  A266 );
 a13685a <=( (not A265)  and  a13684a );
 a13686a <=( a13685a  and  a13680a );
 a13689a <=( A167  and  A168 );
 a13693a <=( (not A202)  and  (not A200) );
 a13694a <=( (not A199)  and  a13693a );
 a13695a <=( a13694a  and  a13689a );
 a13698a <=( A234  and  A232 );
 a13702a <=( A269  and  (not A266) );
 a13703a <=( A265  and  a13702a );
 a13704a <=( a13703a  and  a13698a );
 a13707a <=( A167  and  A168 );
 a13711a <=( (not A202)  and  (not A200) );
 a13712a <=( (not A199)  and  a13711a );
 a13713a <=( a13712a  and  a13707a );
 a13716a <=( A234  and  A233 );
 a13720a <=( (not A302)  and  (not A301) );
 a13721a <=( (not A300)  and  a13720a );
 a13722a <=( a13721a  and  a13716a );
 a13725a <=( A167  and  A168 );
 a13729a <=( (not A202)  and  (not A200) );
 a13730a <=( (not A199)  and  a13729a );
 a13731a <=( a13730a  and  a13725a );
 a13734a <=( A234  and  A233 );
 a13738a <=( (not A301)  and  (not A299) );
 a13739a <=( (not A298)  and  a13738a );
 a13740a <=( a13739a  and  a13734a );
 a13743a <=( A167  and  A168 );
 a13747a <=( (not A202)  and  (not A200) );
 a13748a <=( (not A199)  and  a13747a );
 a13749a <=( a13748a  and  a13743a );
 a13752a <=( A234  and  A233 );
 a13756a <=( A269  and  A266 );
 a13757a <=( (not A265)  and  a13756a );
 a13758a <=( a13757a  and  a13752a );
 a13761a <=( A167  and  A168 );
 a13765a <=( (not A202)  and  (not A200) );
 a13766a <=( (not A199)  and  a13765a );
 a13767a <=( a13766a  and  a13761a );
 a13770a <=( A234  and  A233 );
 a13774a <=( A269  and  (not A266) );
 a13775a <=( A265  and  a13774a );
 a13776a <=( a13775a  and  a13770a );
 a13779a <=( A167  and  A168 );
 a13783a <=( (not A202)  and  (not A200) );
 a13784a <=( (not A199)  and  a13783a );
 a13785a <=( a13784a  and  a13779a );
 a13788a <=( A233  and  (not A232) );
 a13792a <=( A267  and  A265 );
 a13793a <=( A236  and  a13792a );
 a13794a <=( a13793a  and  a13788a );
 a13797a <=( A167  and  A168 );
 a13801a <=( (not A202)  and  (not A200) );
 a13802a <=( (not A199)  and  a13801a );
 a13803a <=( a13802a  and  a13797a );
 a13806a <=( A233  and  (not A232) );
 a13810a <=( A267  and  A266 );
 a13811a <=( A236  and  a13810a );
 a13812a <=( a13811a  and  a13806a );
 a13815a <=( A167  and  A168 );
 a13819a <=( (not A202)  and  (not A200) );
 a13820a <=( (not A199)  and  a13819a );
 a13821a <=( a13820a  and  a13815a );
 a13824a <=( (not A233)  and  A232 );
 a13828a <=( A267  and  A265 );
 a13829a <=( A236  and  a13828a );
 a13830a <=( a13829a  and  a13824a );
 a13833a <=( A167  and  A168 );
 a13837a <=( (not A202)  and  (not A200) );
 a13838a <=( (not A199)  and  a13837a );
 a13839a <=( a13838a  and  a13833a );
 a13842a <=( (not A233)  and  A232 );
 a13846a <=( A267  and  A266 );
 a13847a <=( A236  and  a13846a );
 a13848a <=( a13847a  and  a13842a );
 a13851a <=( A167  and  A170 );
 a13855a <=( (not A202)  and  (not A201) );
 a13856a <=( (not A166)  and  a13855a );
 a13857a <=( a13856a  and  a13851a );
 a13860a <=( A235  and  (not A203) );
 a13864a <=( (not A302)  and  (not A301) );
 a13865a <=( (not A300)  and  a13864a );
 a13866a <=( a13865a  and  a13860a );
 a13869a <=( A167  and  A170 );
 a13873a <=( (not A202)  and  (not A201) );
 a13874a <=( (not A166)  and  a13873a );
 a13875a <=( a13874a  and  a13869a );
 a13878a <=( A235  and  (not A203) );
 a13882a <=( (not A301)  and  (not A299) );
 a13883a <=( (not A298)  and  a13882a );
 a13884a <=( a13883a  and  a13878a );
 a13887a <=( A167  and  A170 );
 a13891a <=( (not A202)  and  (not A201) );
 a13892a <=( (not A166)  and  a13891a );
 a13893a <=( a13892a  and  a13887a );
 a13896a <=( A235  and  (not A203) );
 a13900a <=( A269  and  A266 );
 a13901a <=( (not A265)  and  a13900a );
 a13902a <=( a13901a  and  a13896a );
 a13905a <=( A167  and  A170 );
 a13909a <=( (not A202)  and  (not A201) );
 a13910a <=( (not A166)  and  a13909a );
 a13911a <=( a13910a  and  a13905a );
 a13914a <=( A235  and  (not A203) );
 a13918a <=( A269  and  (not A266) );
 a13919a <=( A265  and  a13918a );
 a13920a <=( a13919a  and  a13914a );
 a13923a <=( A167  and  A170 );
 a13927a <=( (not A202)  and  (not A201) );
 a13928a <=( (not A166)  and  a13927a );
 a13929a <=( a13928a  and  a13923a );
 a13932a <=( A232  and  (not A203) );
 a13936a <=( A267  and  A265 );
 a13937a <=( A234  and  a13936a );
 a13938a <=( a13937a  and  a13932a );
 a13941a <=( A167  and  A170 );
 a13945a <=( (not A202)  and  (not A201) );
 a13946a <=( (not A166)  and  a13945a );
 a13947a <=( a13946a  and  a13941a );
 a13950a <=( A232  and  (not A203) );
 a13954a <=( A267  and  A266 );
 a13955a <=( A234  and  a13954a );
 a13956a <=( a13955a  and  a13950a );
 a13959a <=( A167  and  A170 );
 a13963a <=( (not A202)  and  (not A201) );
 a13964a <=( (not A166)  and  a13963a );
 a13965a <=( a13964a  and  a13959a );
 a13968a <=( A233  and  (not A203) );
 a13972a <=( A267  and  A265 );
 a13973a <=( A234  and  a13972a );
 a13974a <=( a13973a  and  a13968a );
 a13977a <=( A167  and  A170 );
 a13981a <=( (not A202)  and  (not A201) );
 a13982a <=( (not A166)  and  a13981a );
 a13983a <=( a13982a  and  a13977a );
 a13986a <=( A233  and  (not A203) );
 a13990a <=( A267  and  A266 );
 a13991a <=( A234  and  a13990a );
 a13992a <=( a13991a  and  a13986a );
 a13995a <=( A167  and  A170 );
 a13999a <=( (not A202)  and  (not A201) );
 a14000a <=( (not A166)  and  a13999a );
 a14001a <=( a14000a  and  a13995a );
 a14004a <=( (not A232)  and  (not A203) );
 a14008a <=( A268  and  A236 );
 a14009a <=( A233  and  a14008a );
 a14010a <=( a14009a  and  a14004a );
 a14013a <=( A167  and  A170 );
 a14017a <=( (not A202)  and  (not A201) );
 a14018a <=( (not A166)  and  a14017a );
 a14019a <=( a14018a  and  a14013a );
 a14022a <=( A232  and  (not A203) );
 a14026a <=( A268  and  A236 );
 a14027a <=( (not A233)  and  a14026a );
 a14028a <=( a14027a  and  a14022a );
 a14031a <=( A167  and  A170 );
 a14035a <=( A200  and  A199 );
 a14036a <=( (not A166)  and  a14035a );
 a14037a <=( a14036a  and  a14031a );
 a14040a <=( (not A202)  and  (not A201) );
 a14044a <=( A267  and  A265 );
 a14045a <=( A235  and  a14044a );
 a14046a <=( a14045a  and  a14040a );
 a14049a <=( A167  and  A170 );
 a14053a <=( A200  and  A199 );
 a14054a <=( (not A166)  and  a14053a );
 a14055a <=( a14054a  and  a14049a );
 a14058a <=( (not A202)  and  (not A201) );
 a14062a <=( A267  and  A266 );
 a14063a <=( A235  and  a14062a );
 a14064a <=( a14063a  and  a14058a );
 a14067a <=( A167  and  A170 );
 a14071a <=( A200  and  A199 );
 a14072a <=( (not A166)  and  a14071a );
 a14073a <=( a14072a  and  a14067a );
 a14076a <=( (not A202)  and  (not A201) );
 a14080a <=( A268  and  A234 );
 a14081a <=( A232  and  a14080a );
 a14082a <=( a14081a  and  a14076a );
 a14085a <=( A167  and  A170 );
 a14089a <=( A200  and  A199 );
 a14090a <=( (not A166)  and  a14089a );
 a14091a <=( a14090a  and  a14085a );
 a14094a <=( (not A202)  and  (not A201) );
 a14098a <=( A268  and  A234 );
 a14099a <=( A233  and  a14098a );
 a14100a <=( a14099a  and  a14094a );
 a14103a <=( A167  and  A170 );
 a14107a <=( (not A200)  and  (not A199) );
 a14108a <=( (not A166)  and  a14107a );
 a14109a <=( a14108a  and  a14103a );
 a14112a <=( A235  and  (not A202) );
 a14116a <=( (not A302)  and  (not A301) );
 a14117a <=( (not A300)  and  a14116a );
 a14118a <=( a14117a  and  a14112a );
 a14121a <=( A167  and  A170 );
 a14125a <=( (not A200)  and  (not A199) );
 a14126a <=( (not A166)  and  a14125a );
 a14127a <=( a14126a  and  a14121a );
 a14130a <=( A235  and  (not A202) );
 a14134a <=( (not A301)  and  (not A299) );
 a14135a <=( (not A298)  and  a14134a );
 a14136a <=( a14135a  and  a14130a );
 a14139a <=( A167  and  A170 );
 a14143a <=( (not A200)  and  (not A199) );
 a14144a <=( (not A166)  and  a14143a );
 a14145a <=( a14144a  and  a14139a );
 a14148a <=( A235  and  (not A202) );
 a14152a <=( A269  and  A266 );
 a14153a <=( (not A265)  and  a14152a );
 a14154a <=( a14153a  and  a14148a );
 a14157a <=( A167  and  A170 );
 a14161a <=( (not A200)  and  (not A199) );
 a14162a <=( (not A166)  and  a14161a );
 a14163a <=( a14162a  and  a14157a );
 a14166a <=( A235  and  (not A202) );
 a14170a <=( A269  and  (not A266) );
 a14171a <=( A265  and  a14170a );
 a14172a <=( a14171a  and  a14166a );
 a14175a <=( A167  and  A170 );
 a14179a <=( (not A200)  and  (not A199) );
 a14180a <=( (not A166)  and  a14179a );
 a14181a <=( a14180a  and  a14175a );
 a14184a <=( A232  and  (not A202) );
 a14188a <=( A267  and  A265 );
 a14189a <=( A234  and  a14188a );
 a14190a <=( a14189a  and  a14184a );
 a14193a <=( A167  and  A170 );
 a14197a <=( (not A200)  and  (not A199) );
 a14198a <=( (not A166)  and  a14197a );
 a14199a <=( a14198a  and  a14193a );
 a14202a <=( A232  and  (not A202) );
 a14206a <=( A267  and  A266 );
 a14207a <=( A234  and  a14206a );
 a14208a <=( a14207a  and  a14202a );
 a14211a <=( A167  and  A170 );
 a14215a <=( (not A200)  and  (not A199) );
 a14216a <=( (not A166)  and  a14215a );
 a14217a <=( a14216a  and  a14211a );
 a14220a <=( A233  and  (not A202) );
 a14224a <=( A267  and  A265 );
 a14225a <=( A234  and  a14224a );
 a14226a <=( a14225a  and  a14220a );
 a14229a <=( A167  and  A170 );
 a14233a <=( (not A200)  and  (not A199) );
 a14234a <=( (not A166)  and  a14233a );
 a14235a <=( a14234a  and  a14229a );
 a14238a <=( A233  and  (not A202) );
 a14242a <=( A267  and  A266 );
 a14243a <=( A234  and  a14242a );
 a14244a <=( a14243a  and  a14238a );
 a14247a <=( A167  and  A170 );
 a14251a <=( (not A200)  and  (not A199) );
 a14252a <=( (not A166)  and  a14251a );
 a14253a <=( a14252a  and  a14247a );
 a14256a <=( (not A232)  and  (not A202) );
 a14260a <=( A268  and  A236 );
 a14261a <=( A233  and  a14260a );
 a14262a <=( a14261a  and  a14256a );
 a14265a <=( A167  and  A170 );
 a14269a <=( (not A200)  and  (not A199) );
 a14270a <=( (not A166)  and  a14269a );
 a14271a <=( a14270a  and  a14265a );
 a14274a <=( A232  and  (not A202) );
 a14278a <=( A268  and  A236 );
 a14279a <=( (not A233)  and  a14278a );
 a14280a <=( a14279a  and  a14274a );
 a14283a <=( (not A167)  and  A170 );
 a14287a <=( (not A202)  and  (not A201) );
 a14288a <=( A166  and  a14287a );
 a14289a <=( a14288a  and  a14283a );
 a14292a <=( A235  and  (not A203) );
 a14296a <=( (not A302)  and  (not A301) );
 a14297a <=( (not A300)  and  a14296a );
 a14298a <=( a14297a  and  a14292a );
 a14301a <=( (not A167)  and  A170 );
 a14305a <=( (not A202)  and  (not A201) );
 a14306a <=( A166  and  a14305a );
 a14307a <=( a14306a  and  a14301a );
 a14310a <=( A235  and  (not A203) );
 a14314a <=( (not A301)  and  (not A299) );
 a14315a <=( (not A298)  and  a14314a );
 a14316a <=( a14315a  and  a14310a );
 a14319a <=( (not A167)  and  A170 );
 a14323a <=( (not A202)  and  (not A201) );
 a14324a <=( A166  and  a14323a );
 a14325a <=( a14324a  and  a14319a );
 a14328a <=( A235  and  (not A203) );
 a14332a <=( A269  and  A266 );
 a14333a <=( (not A265)  and  a14332a );
 a14334a <=( a14333a  and  a14328a );
 a14337a <=( (not A167)  and  A170 );
 a14341a <=( (not A202)  and  (not A201) );
 a14342a <=( A166  and  a14341a );
 a14343a <=( a14342a  and  a14337a );
 a14346a <=( A235  and  (not A203) );
 a14350a <=( A269  and  (not A266) );
 a14351a <=( A265  and  a14350a );
 a14352a <=( a14351a  and  a14346a );
 a14355a <=( (not A167)  and  A170 );
 a14359a <=( (not A202)  and  (not A201) );
 a14360a <=( A166  and  a14359a );
 a14361a <=( a14360a  and  a14355a );
 a14364a <=( A232  and  (not A203) );
 a14368a <=( A267  and  A265 );
 a14369a <=( A234  and  a14368a );
 a14370a <=( a14369a  and  a14364a );
 a14373a <=( (not A167)  and  A170 );
 a14377a <=( (not A202)  and  (not A201) );
 a14378a <=( A166  and  a14377a );
 a14379a <=( a14378a  and  a14373a );
 a14382a <=( A232  and  (not A203) );
 a14386a <=( A267  and  A266 );
 a14387a <=( A234  and  a14386a );
 a14388a <=( a14387a  and  a14382a );
 a14391a <=( (not A167)  and  A170 );
 a14395a <=( (not A202)  and  (not A201) );
 a14396a <=( A166  and  a14395a );
 a14397a <=( a14396a  and  a14391a );
 a14400a <=( A233  and  (not A203) );
 a14404a <=( A267  and  A265 );
 a14405a <=( A234  and  a14404a );
 a14406a <=( a14405a  and  a14400a );
 a14409a <=( (not A167)  and  A170 );
 a14413a <=( (not A202)  and  (not A201) );
 a14414a <=( A166  and  a14413a );
 a14415a <=( a14414a  and  a14409a );
 a14418a <=( A233  and  (not A203) );
 a14422a <=( A267  and  A266 );
 a14423a <=( A234  and  a14422a );
 a14424a <=( a14423a  and  a14418a );
 a14427a <=( (not A167)  and  A170 );
 a14431a <=( (not A202)  and  (not A201) );
 a14432a <=( A166  and  a14431a );
 a14433a <=( a14432a  and  a14427a );
 a14436a <=( (not A232)  and  (not A203) );
 a14440a <=( A268  and  A236 );
 a14441a <=( A233  and  a14440a );
 a14442a <=( a14441a  and  a14436a );
 a14445a <=( (not A167)  and  A170 );
 a14449a <=( (not A202)  and  (not A201) );
 a14450a <=( A166  and  a14449a );
 a14451a <=( a14450a  and  a14445a );
 a14454a <=( A232  and  (not A203) );
 a14458a <=( A268  and  A236 );
 a14459a <=( (not A233)  and  a14458a );
 a14460a <=( a14459a  and  a14454a );
 a14463a <=( (not A167)  and  A170 );
 a14467a <=( A200  and  A199 );
 a14468a <=( A166  and  a14467a );
 a14469a <=( a14468a  and  a14463a );
 a14472a <=( (not A202)  and  (not A201) );
 a14476a <=( A267  and  A265 );
 a14477a <=( A235  and  a14476a );
 a14478a <=( a14477a  and  a14472a );
 a14481a <=( (not A167)  and  A170 );
 a14485a <=( A200  and  A199 );
 a14486a <=( A166  and  a14485a );
 a14487a <=( a14486a  and  a14481a );
 a14490a <=( (not A202)  and  (not A201) );
 a14494a <=( A267  and  A266 );
 a14495a <=( A235  and  a14494a );
 a14496a <=( a14495a  and  a14490a );
 a14499a <=( (not A167)  and  A170 );
 a14503a <=( A200  and  A199 );
 a14504a <=( A166  and  a14503a );
 a14505a <=( a14504a  and  a14499a );
 a14508a <=( (not A202)  and  (not A201) );
 a14512a <=( A268  and  A234 );
 a14513a <=( A232  and  a14512a );
 a14514a <=( a14513a  and  a14508a );
 a14517a <=( (not A167)  and  A170 );
 a14521a <=( A200  and  A199 );
 a14522a <=( A166  and  a14521a );
 a14523a <=( a14522a  and  a14517a );
 a14526a <=( (not A202)  and  (not A201) );
 a14530a <=( A268  and  A234 );
 a14531a <=( A233  and  a14530a );
 a14532a <=( a14531a  and  a14526a );
 a14535a <=( (not A167)  and  A170 );
 a14539a <=( (not A200)  and  (not A199) );
 a14540a <=( A166  and  a14539a );
 a14541a <=( a14540a  and  a14535a );
 a14544a <=( A235  and  (not A202) );
 a14548a <=( (not A302)  and  (not A301) );
 a14549a <=( (not A300)  and  a14548a );
 a14550a <=( a14549a  and  a14544a );
 a14553a <=( (not A167)  and  A170 );
 a14557a <=( (not A200)  and  (not A199) );
 a14558a <=( A166  and  a14557a );
 a14559a <=( a14558a  and  a14553a );
 a14562a <=( A235  and  (not A202) );
 a14566a <=( (not A301)  and  (not A299) );
 a14567a <=( (not A298)  and  a14566a );
 a14568a <=( a14567a  and  a14562a );
 a14571a <=( (not A167)  and  A170 );
 a14575a <=( (not A200)  and  (not A199) );
 a14576a <=( A166  and  a14575a );
 a14577a <=( a14576a  and  a14571a );
 a14580a <=( A235  and  (not A202) );
 a14584a <=( A269  and  A266 );
 a14585a <=( (not A265)  and  a14584a );
 a14586a <=( a14585a  and  a14580a );
 a14589a <=( (not A167)  and  A170 );
 a14593a <=( (not A200)  and  (not A199) );
 a14594a <=( A166  and  a14593a );
 a14595a <=( a14594a  and  a14589a );
 a14598a <=( A235  and  (not A202) );
 a14602a <=( A269  and  (not A266) );
 a14603a <=( A265  and  a14602a );
 a14604a <=( a14603a  and  a14598a );
 a14607a <=( (not A167)  and  A170 );
 a14611a <=( (not A200)  and  (not A199) );
 a14612a <=( A166  and  a14611a );
 a14613a <=( a14612a  and  a14607a );
 a14616a <=( A232  and  (not A202) );
 a14620a <=( A267  and  A265 );
 a14621a <=( A234  and  a14620a );
 a14622a <=( a14621a  and  a14616a );
 a14625a <=( (not A167)  and  A170 );
 a14629a <=( (not A200)  and  (not A199) );
 a14630a <=( A166  and  a14629a );
 a14631a <=( a14630a  and  a14625a );
 a14634a <=( A232  and  (not A202) );
 a14638a <=( A267  and  A266 );
 a14639a <=( A234  and  a14638a );
 a14640a <=( a14639a  and  a14634a );
 a14643a <=( (not A167)  and  A170 );
 a14647a <=( (not A200)  and  (not A199) );
 a14648a <=( A166  and  a14647a );
 a14649a <=( a14648a  and  a14643a );
 a14652a <=( A233  and  (not A202) );
 a14656a <=( A267  and  A265 );
 a14657a <=( A234  and  a14656a );
 a14658a <=( a14657a  and  a14652a );
 a14661a <=( (not A167)  and  A170 );
 a14665a <=( (not A200)  and  (not A199) );
 a14666a <=( A166  and  a14665a );
 a14667a <=( a14666a  and  a14661a );
 a14670a <=( A233  and  (not A202) );
 a14674a <=( A267  and  A266 );
 a14675a <=( A234  and  a14674a );
 a14676a <=( a14675a  and  a14670a );
 a14679a <=( (not A167)  and  A170 );
 a14683a <=( (not A200)  and  (not A199) );
 a14684a <=( A166  and  a14683a );
 a14685a <=( a14684a  and  a14679a );
 a14688a <=( (not A232)  and  (not A202) );
 a14692a <=( A268  and  A236 );
 a14693a <=( A233  and  a14692a );
 a14694a <=( a14693a  and  a14688a );
 a14697a <=( (not A167)  and  A170 );
 a14701a <=( (not A200)  and  (not A199) );
 a14702a <=( A166  and  a14701a );
 a14703a <=( a14702a  and  a14697a );
 a14706a <=( A232  and  (not A202) );
 a14710a <=( A268  and  A236 );
 a14711a <=( (not A233)  and  a14710a );
 a14712a <=( a14711a  and  a14706a );
 a14715a <=( (not A201)  and  A169 );
 a14719a <=( A232  and  (not A203) );
 a14720a <=( (not A202)  and  a14719a );
 a14721a <=( a14720a  and  a14715a );
 a14724a <=( A298  and  A234 );
 a14728a <=( (not A301)  and  (not A300) );
 a14729a <=( A299  and  a14728a );
 a14730a <=( a14729a  and  a14724a );
 a14733a <=( (not A201)  and  A169 );
 a14737a <=( A233  and  (not A203) );
 a14738a <=( (not A202)  and  a14737a );
 a14739a <=( a14738a  and  a14733a );
 a14742a <=( A298  and  A234 );
 a14746a <=( (not A301)  and  (not A300) );
 a14747a <=( A299  and  a14746a );
 a14748a <=( a14747a  and  a14742a );
 a14751a <=( (not A201)  and  A169 );
 a14755a <=( (not A232)  and  (not A203) );
 a14756a <=( (not A202)  and  a14755a );
 a14757a <=( a14756a  and  a14751a );
 a14760a <=( A236  and  A233 );
 a14764a <=( (not A302)  and  (not A301) );
 a14765a <=( (not A300)  and  a14764a );
 a14766a <=( a14765a  and  a14760a );
 a14769a <=( (not A201)  and  A169 );
 a14773a <=( (not A232)  and  (not A203) );
 a14774a <=( (not A202)  and  a14773a );
 a14775a <=( a14774a  and  a14769a );
 a14778a <=( A236  and  A233 );
 a14782a <=( (not A301)  and  (not A299) );
 a14783a <=( (not A298)  and  a14782a );
 a14784a <=( a14783a  and  a14778a );
 a14787a <=( (not A201)  and  A169 );
 a14791a <=( (not A232)  and  (not A203) );
 a14792a <=( (not A202)  and  a14791a );
 a14793a <=( a14792a  and  a14787a );
 a14796a <=( A236  and  A233 );
 a14800a <=( A269  and  A266 );
 a14801a <=( (not A265)  and  a14800a );
 a14802a <=( a14801a  and  a14796a );
 a14805a <=( (not A201)  and  A169 );
 a14809a <=( (not A232)  and  (not A203) );
 a14810a <=( (not A202)  and  a14809a );
 a14811a <=( a14810a  and  a14805a );
 a14814a <=( A236  and  A233 );
 a14818a <=( A269  and  (not A266) );
 a14819a <=( A265  and  a14818a );
 a14820a <=( a14819a  and  a14814a );
 a14823a <=( (not A201)  and  A169 );
 a14827a <=( A232  and  (not A203) );
 a14828a <=( (not A202)  and  a14827a );
 a14829a <=( a14828a  and  a14823a );
 a14832a <=( A236  and  (not A233) );
 a14836a <=( (not A302)  and  (not A301) );
 a14837a <=( (not A300)  and  a14836a );
 a14838a <=( a14837a  and  a14832a );
 a14841a <=( (not A201)  and  A169 );
 a14845a <=( A232  and  (not A203) );
 a14846a <=( (not A202)  and  a14845a );
 a14847a <=( a14846a  and  a14841a );
 a14850a <=( A236  and  (not A233) );
 a14854a <=( (not A301)  and  (not A299) );
 a14855a <=( (not A298)  and  a14854a );
 a14856a <=( a14855a  and  a14850a );
 a14859a <=( (not A201)  and  A169 );
 a14863a <=( A232  and  (not A203) );
 a14864a <=( (not A202)  and  a14863a );
 a14865a <=( a14864a  and  a14859a );
 a14868a <=( A236  and  (not A233) );
 a14872a <=( A269  and  A266 );
 a14873a <=( (not A265)  and  a14872a );
 a14874a <=( a14873a  and  a14868a );
 a14877a <=( (not A201)  and  A169 );
 a14881a <=( A232  and  (not A203) );
 a14882a <=( (not A202)  and  a14881a );
 a14883a <=( a14882a  and  a14877a );
 a14886a <=( A236  and  (not A233) );
 a14890a <=( A269  and  (not A266) );
 a14891a <=( A265  and  a14890a );
 a14892a <=( a14891a  and  a14886a );
 a14895a <=( A199  and  A169 );
 a14899a <=( (not A202)  and  (not A201) );
 a14900a <=( A200  and  a14899a );
 a14901a <=( a14900a  and  a14895a );
 a14904a <=( A298  and  A235 );
 a14908a <=( (not A301)  and  (not A300) );
 a14909a <=( A299  and  a14908a );
 a14910a <=( a14909a  and  a14904a );
 a14913a <=( A199  and  A169 );
 a14917a <=( (not A202)  and  (not A201) );
 a14918a <=( A200  and  a14917a );
 a14919a <=( a14918a  and  a14913a );
 a14922a <=( A234  and  A232 );
 a14926a <=( (not A302)  and  (not A301) );
 a14927a <=( (not A300)  and  a14926a );
 a14928a <=( a14927a  and  a14922a );
 a14931a <=( A199  and  A169 );
 a14935a <=( (not A202)  and  (not A201) );
 a14936a <=( A200  and  a14935a );
 a14937a <=( a14936a  and  a14931a );
 a14940a <=( A234  and  A232 );
 a14944a <=( (not A301)  and  (not A299) );
 a14945a <=( (not A298)  and  a14944a );
 a14946a <=( a14945a  and  a14940a );
 a14949a <=( A199  and  A169 );
 a14953a <=( (not A202)  and  (not A201) );
 a14954a <=( A200  and  a14953a );
 a14955a <=( a14954a  and  a14949a );
 a14958a <=( A234  and  A232 );
 a14962a <=( A269  and  A266 );
 a14963a <=( (not A265)  and  a14962a );
 a14964a <=( a14963a  and  a14958a );
 a14967a <=( A199  and  A169 );
 a14971a <=( (not A202)  and  (not A201) );
 a14972a <=( A200  and  a14971a );
 a14973a <=( a14972a  and  a14967a );
 a14976a <=( A234  and  A232 );
 a14980a <=( A269  and  (not A266) );
 a14981a <=( A265  and  a14980a );
 a14982a <=( a14981a  and  a14976a );
 a14985a <=( A199  and  A169 );
 a14989a <=( (not A202)  and  (not A201) );
 a14990a <=( A200  and  a14989a );
 a14991a <=( a14990a  and  a14985a );
 a14994a <=( A234  and  A233 );
 a14998a <=( (not A302)  and  (not A301) );
 a14999a <=( (not A300)  and  a14998a );
 a15000a <=( a14999a  and  a14994a );
 a15003a <=( A199  and  A169 );
 a15007a <=( (not A202)  and  (not A201) );
 a15008a <=( A200  and  a15007a );
 a15009a <=( a15008a  and  a15003a );
 a15012a <=( A234  and  A233 );
 a15016a <=( (not A301)  and  (not A299) );
 a15017a <=( (not A298)  and  a15016a );
 a15018a <=( a15017a  and  a15012a );
 a15021a <=( A199  and  A169 );
 a15025a <=( (not A202)  and  (not A201) );
 a15026a <=( A200  and  a15025a );
 a15027a <=( a15026a  and  a15021a );
 a15030a <=( A234  and  A233 );
 a15034a <=( A269  and  A266 );
 a15035a <=( (not A265)  and  a15034a );
 a15036a <=( a15035a  and  a15030a );
 a15039a <=( A199  and  A169 );
 a15043a <=( (not A202)  and  (not A201) );
 a15044a <=( A200  and  a15043a );
 a15045a <=( a15044a  and  a15039a );
 a15048a <=( A234  and  A233 );
 a15052a <=( A269  and  (not A266) );
 a15053a <=( A265  and  a15052a );
 a15054a <=( a15053a  and  a15048a );
 a15057a <=( A199  and  A169 );
 a15061a <=( (not A202)  and  (not A201) );
 a15062a <=( A200  and  a15061a );
 a15063a <=( a15062a  and  a15057a );
 a15066a <=( A233  and  (not A232) );
 a15070a <=( A267  and  A265 );
 a15071a <=( A236  and  a15070a );
 a15072a <=( a15071a  and  a15066a );
 a15075a <=( A199  and  A169 );
 a15079a <=( (not A202)  and  (not A201) );
 a15080a <=( A200  and  a15079a );
 a15081a <=( a15080a  and  a15075a );
 a15084a <=( A233  and  (not A232) );
 a15088a <=( A267  and  A266 );
 a15089a <=( A236  and  a15088a );
 a15090a <=( a15089a  and  a15084a );
 a15093a <=( A199  and  A169 );
 a15097a <=( (not A202)  and  (not A201) );
 a15098a <=( A200  and  a15097a );
 a15099a <=( a15098a  and  a15093a );
 a15102a <=( (not A233)  and  A232 );
 a15106a <=( A267  and  A265 );
 a15107a <=( A236  and  a15106a );
 a15108a <=( a15107a  and  a15102a );
 a15111a <=( A199  and  A169 );
 a15115a <=( (not A202)  and  (not A201) );
 a15116a <=( A200  and  a15115a );
 a15117a <=( a15116a  and  a15111a );
 a15120a <=( (not A233)  and  A232 );
 a15124a <=( A267  and  A266 );
 a15125a <=( A236  and  a15124a );
 a15126a <=( a15125a  and  a15120a );
 a15129a <=( (not A199)  and  A169 );
 a15133a <=( A232  and  (not A202) );
 a15134a <=( (not A200)  and  a15133a );
 a15135a <=( a15134a  and  a15129a );
 a15138a <=( A298  and  A234 );
 a15142a <=( (not A301)  and  (not A300) );
 a15143a <=( A299  and  a15142a );
 a15144a <=( a15143a  and  a15138a );
 a15147a <=( (not A199)  and  A169 );
 a15151a <=( A233  and  (not A202) );
 a15152a <=( (not A200)  and  a15151a );
 a15153a <=( a15152a  and  a15147a );
 a15156a <=( A298  and  A234 );
 a15160a <=( (not A301)  and  (not A300) );
 a15161a <=( A299  and  a15160a );
 a15162a <=( a15161a  and  a15156a );
 a15165a <=( (not A199)  and  A169 );
 a15169a <=( (not A232)  and  (not A202) );
 a15170a <=( (not A200)  and  a15169a );
 a15171a <=( a15170a  and  a15165a );
 a15174a <=( A236  and  A233 );
 a15178a <=( (not A302)  and  (not A301) );
 a15179a <=( (not A300)  and  a15178a );
 a15180a <=( a15179a  and  a15174a );
 a15183a <=( (not A199)  and  A169 );
 a15187a <=( (not A232)  and  (not A202) );
 a15188a <=( (not A200)  and  a15187a );
 a15189a <=( a15188a  and  a15183a );
 a15192a <=( A236  and  A233 );
 a15196a <=( (not A301)  and  (not A299) );
 a15197a <=( (not A298)  and  a15196a );
 a15198a <=( a15197a  and  a15192a );
 a15201a <=( (not A199)  and  A169 );
 a15205a <=( (not A232)  and  (not A202) );
 a15206a <=( (not A200)  and  a15205a );
 a15207a <=( a15206a  and  a15201a );
 a15210a <=( A236  and  A233 );
 a15214a <=( A269  and  A266 );
 a15215a <=( (not A265)  and  a15214a );
 a15216a <=( a15215a  and  a15210a );
 a15219a <=( (not A199)  and  A169 );
 a15223a <=( (not A232)  and  (not A202) );
 a15224a <=( (not A200)  and  a15223a );
 a15225a <=( a15224a  and  a15219a );
 a15228a <=( A236  and  A233 );
 a15232a <=( A269  and  (not A266) );
 a15233a <=( A265  and  a15232a );
 a15234a <=( a15233a  and  a15228a );
 a15237a <=( (not A199)  and  A169 );
 a15241a <=( A232  and  (not A202) );
 a15242a <=( (not A200)  and  a15241a );
 a15243a <=( a15242a  and  a15237a );
 a15246a <=( A236  and  (not A233) );
 a15250a <=( (not A302)  and  (not A301) );
 a15251a <=( (not A300)  and  a15250a );
 a15252a <=( a15251a  and  a15246a );
 a15255a <=( (not A199)  and  A169 );
 a15259a <=( A232  and  (not A202) );
 a15260a <=( (not A200)  and  a15259a );
 a15261a <=( a15260a  and  a15255a );
 a15264a <=( A236  and  (not A233) );
 a15268a <=( (not A301)  and  (not A299) );
 a15269a <=( (not A298)  and  a15268a );
 a15270a <=( a15269a  and  a15264a );
 a15273a <=( (not A199)  and  A169 );
 a15277a <=( A232  and  (not A202) );
 a15278a <=( (not A200)  and  a15277a );
 a15279a <=( a15278a  and  a15273a );
 a15282a <=( A236  and  (not A233) );
 a15286a <=( A269  and  A266 );
 a15287a <=( (not A265)  and  a15286a );
 a15288a <=( a15287a  and  a15282a );
 a15291a <=( (not A199)  and  A169 );
 a15295a <=( A232  and  (not A202) );
 a15296a <=( (not A200)  and  a15295a );
 a15297a <=( a15296a  and  a15291a );
 a15300a <=( A236  and  (not A233) );
 a15304a <=( A269  and  (not A266) );
 a15305a <=( A265  and  a15304a );
 a15306a <=( a15305a  and  a15300a );
 a15309a <=( (not A167)  and  (not A169) );
 a15313a <=( A232  and  A202 );
 a15314a <=( (not A166)  and  a15313a );
 a15315a <=( a15314a  and  a15309a );
 a15318a <=( A298  and  A234 );
 a15322a <=( (not A301)  and  (not A300) );
 a15323a <=( A299  and  a15322a );
 a15324a <=( a15323a  and  a15318a );
 a15327a <=( (not A167)  and  (not A169) );
 a15331a <=( A233  and  A202 );
 a15332a <=( (not A166)  and  a15331a );
 a15333a <=( a15332a  and  a15327a );
 a15336a <=( A298  and  A234 );
 a15340a <=( (not A301)  and  (not A300) );
 a15341a <=( A299  and  a15340a );
 a15342a <=( a15341a  and  a15336a );
 a15345a <=( (not A167)  and  (not A169) );
 a15349a <=( (not A232)  and  A202 );
 a15350a <=( (not A166)  and  a15349a );
 a15351a <=( a15350a  and  a15345a );
 a15354a <=( A236  and  A233 );
 a15358a <=( (not A302)  and  (not A301) );
 a15359a <=( (not A300)  and  a15358a );
 a15360a <=( a15359a  and  a15354a );
 a15363a <=( (not A167)  and  (not A169) );
 a15367a <=( (not A232)  and  A202 );
 a15368a <=( (not A166)  and  a15367a );
 a15369a <=( a15368a  and  a15363a );
 a15372a <=( A236  and  A233 );
 a15376a <=( (not A301)  and  (not A299) );
 a15377a <=( (not A298)  and  a15376a );
 a15378a <=( a15377a  and  a15372a );
 a15381a <=( (not A167)  and  (not A169) );
 a15385a <=( (not A232)  and  A202 );
 a15386a <=( (not A166)  and  a15385a );
 a15387a <=( a15386a  and  a15381a );
 a15390a <=( A236  and  A233 );
 a15394a <=( A269  and  A266 );
 a15395a <=( (not A265)  and  a15394a );
 a15396a <=( a15395a  and  a15390a );
 a15399a <=( (not A167)  and  (not A169) );
 a15403a <=( (not A232)  and  A202 );
 a15404a <=( (not A166)  and  a15403a );
 a15405a <=( a15404a  and  a15399a );
 a15408a <=( A236  and  A233 );
 a15412a <=( A269  and  (not A266) );
 a15413a <=( A265  and  a15412a );
 a15414a <=( a15413a  and  a15408a );
 a15417a <=( (not A167)  and  (not A169) );
 a15421a <=( A232  and  A202 );
 a15422a <=( (not A166)  and  a15421a );
 a15423a <=( a15422a  and  a15417a );
 a15426a <=( A236  and  (not A233) );
 a15430a <=( (not A302)  and  (not A301) );
 a15431a <=( (not A300)  and  a15430a );
 a15432a <=( a15431a  and  a15426a );
 a15435a <=( (not A167)  and  (not A169) );
 a15439a <=( A232  and  A202 );
 a15440a <=( (not A166)  and  a15439a );
 a15441a <=( a15440a  and  a15435a );
 a15444a <=( A236  and  (not A233) );
 a15448a <=( (not A301)  and  (not A299) );
 a15449a <=( (not A298)  and  a15448a );
 a15450a <=( a15449a  and  a15444a );
 a15453a <=( (not A167)  and  (not A169) );
 a15457a <=( A232  and  A202 );
 a15458a <=( (not A166)  and  a15457a );
 a15459a <=( a15458a  and  a15453a );
 a15462a <=( A236  and  (not A233) );
 a15466a <=( A269  and  A266 );
 a15467a <=( (not A265)  and  a15466a );
 a15468a <=( a15467a  and  a15462a );
 a15471a <=( (not A167)  and  (not A169) );
 a15475a <=( A232  and  A202 );
 a15476a <=( (not A166)  and  a15475a );
 a15477a <=( a15476a  and  a15471a );
 a15480a <=( A236  and  (not A233) );
 a15484a <=( A269  and  (not A266) );
 a15485a <=( A265  and  a15484a );
 a15486a <=( a15485a  and  a15480a );
 a15489a <=( (not A167)  and  (not A169) );
 a15493a <=( A201  and  A199 );
 a15494a <=( (not A166)  and  a15493a );
 a15495a <=( a15494a  and  a15489a );
 a15498a <=( A298  and  A235 );
 a15502a <=( (not A301)  and  (not A300) );
 a15503a <=( A299  and  a15502a );
 a15504a <=( a15503a  and  a15498a );
 a15507a <=( (not A167)  and  (not A169) );
 a15511a <=( A201  and  A199 );
 a15512a <=( (not A166)  and  a15511a );
 a15513a <=( a15512a  and  a15507a );
 a15516a <=( A234  and  A232 );
 a15520a <=( (not A302)  and  (not A301) );
 a15521a <=( (not A300)  and  a15520a );
 a15522a <=( a15521a  and  a15516a );
 a15525a <=( (not A167)  and  (not A169) );
 a15529a <=( A201  and  A199 );
 a15530a <=( (not A166)  and  a15529a );
 a15531a <=( a15530a  and  a15525a );
 a15534a <=( A234  and  A232 );
 a15538a <=( (not A301)  and  (not A299) );
 a15539a <=( (not A298)  and  a15538a );
 a15540a <=( a15539a  and  a15534a );
 a15543a <=( (not A167)  and  (not A169) );
 a15547a <=( A201  and  A199 );
 a15548a <=( (not A166)  and  a15547a );
 a15549a <=( a15548a  and  a15543a );
 a15552a <=( A234  and  A232 );
 a15556a <=( A269  and  A266 );
 a15557a <=( (not A265)  and  a15556a );
 a15558a <=( a15557a  and  a15552a );
 a15561a <=( (not A167)  and  (not A169) );
 a15565a <=( A201  and  A199 );
 a15566a <=( (not A166)  and  a15565a );
 a15567a <=( a15566a  and  a15561a );
 a15570a <=( A234  and  A232 );
 a15574a <=( A269  and  (not A266) );
 a15575a <=( A265  and  a15574a );
 a15576a <=( a15575a  and  a15570a );
 a15579a <=( (not A167)  and  (not A169) );
 a15583a <=( A201  and  A199 );
 a15584a <=( (not A166)  and  a15583a );
 a15585a <=( a15584a  and  a15579a );
 a15588a <=( A234  and  A233 );
 a15592a <=( (not A302)  and  (not A301) );
 a15593a <=( (not A300)  and  a15592a );
 a15594a <=( a15593a  and  a15588a );
 a15597a <=( (not A167)  and  (not A169) );
 a15601a <=( A201  and  A199 );
 a15602a <=( (not A166)  and  a15601a );
 a15603a <=( a15602a  and  a15597a );
 a15606a <=( A234  and  A233 );
 a15610a <=( (not A301)  and  (not A299) );
 a15611a <=( (not A298)  and  a15610a );
 a15612a <=( a15611a  and  a15606a );
 a15615a <=( (not A167)  and  (not A169) );
 a15619a <=( A201  and  A199 );
 a15620a <=( (not A166)  and  a15619a );
 a15621a <=( a15620a  and  a15615a );
 a15624a <=( A234  and  A233 );
 a15628a <=( A269  and  A266 );
 a15629a <=( (not A265)  and  a15628a );
 a15630a <=( a15629a  and  a15624a );
 a15633a <=( (not A167)  and  (not A169) );
 a15637a <=( A201  and  A199 );
 a15638a <=( (not A166)  and  a15637a );
 a15639a <=( a15638a  and  a15633a );
 a15642a <=( A234  and  A233 );
 a15646a <=( A269  and  (not A266) );
 a15647a <=( A265  and  a15646a );
 a15648a <=( a15647a  and  a15642a );
 a15651a <=( (not A167)  and  (not A169) );
 a15655a <=( A201  and  A199 );
 a15656a <=( (not A166)  and  a15655a );
 a15657a <=( a15656a  and  a15651a );
 a15660a <=( A233  and  (not A232) );
 a15664a <=( A267  and  A265 );
 a15665a <=( A236  and  a15664a );
 a15666a <=( a15665a  and  a15660a );
 a15669a <=( (not A167)  and  (not A169) );
 a15673a <=( A201  and  A199 );
 a15674a <=( (not A166)  and  a15673a );
 a15675a <=( a15674a  and  a15669a );
 a15678a <=( A233  and  (not A232) );
 a15682a <=( A267  and  A266 );
 a15683a <=( A236  and  a15682a );
 a15684a <=( a15683a  and  a15678a );
 a15687a <=( (not A167)  and  (not A169) );
 a15691a <=( A201  and  A199 );
 a15692a <=( (not A166)  and  a15691a );
 a15693a <=( a15692a  and  a15687a );
 a15696a <=( (not A233)  and  A232 );
 a15700a <=( A267  and  A265 );
 a15701a <=( A236  and  a15700a );
 a15702a <=( a15701a  and  a15696a );
 a15705a <=( (not A167)  and  (not A169) );
 a15709a <=( A201  and  A199 );
 a15710a <=( (not A166)  and  a15709a );
 a15711a <=( a15710a  and  a15705a );
 a15714a <=( (not A233)  and  A232 );
 a15718a <=( A267  and  A266 );
 a15719a <=( A236  and  a15718a );
 a15720a <=( a15719a  and  a15714a );
 a15723a <=( (not A167)  and  (not A169) );
 a15727a <=( A201  and  A200 );
 a15728a <=( (not A166)  and  a15727a );
 a15729a <=( a15728a  and  a15723a );
 a15732a <=( A298  and  A235 );
 a15736a <=( (not A301)  and  (not A300) );
 a15737a <=( A299  and  a15736a );
 a15738a <=( a15737a  and  a15732a );
 a15741a <=( (not A167)  and  (not A169) );
 a15745a <=( A201  and  A200 );
 a15746a <=( (not A166)  and  a15745a );
 a15747a <=( a15746a  and  a15741a );
 a15750a <=( A234  and  A232 );
 a15754a <=( (not A302)  and  (not A301) );
 a15755a <=( (not A300)  and  a15754a );
 a15756a <=( a15755a  and  a15750a );
 a15759a <=( (not A167)  and  (not A169) );
 a15763a <=( A201  and  A200 );
 a15764a <=( (not A166)  and  a15763a );
 a15765a <=( a15764a  and  a15759a );
 a15768a <=( A234  and  A232 );
 a15772a <=( (not A301)  and  (not A299) );
 a15773a <=( (not A298)  and  a15772a );
 a15774a <=( a15773a  and  a15768a );
 a15777a <=( (not A167)  and  (not A169) );
 a15781a <=( A201  and  A200 );
 a15782a <=( (not A166)  and  a15781a );
 a15783a <=( a15782a  and  a15777a );
 a15786a <=( A234  and  A232 );
 a15790a <=( A269  and  A266 );
 a15791a <=( (not A265)  and  a15790a );
 a15792a <=( a15791a  and  a15786a );
 a15795a <=( (not A167)  and  (not A169) );
 a15799a <=( A201  and  A200 );
 a15800a <=( (not A166)  and  a15799a );
 a15801a <=( a15800a  and  a15795a );
 a15804a <=( A234  and  A232 );
 a15808a <=( A269  and  (not A266) );
 a15809a <=( A265  and  a15808a );
 a15810a <=( a15809a  and  a15804a );
 a15813a <=( (not A167)  and  (not A169) );
 a15817a <=( A201  and  A200 );
 a15818a <=( (not A166)  and  a15817a );
 a15819a <=( a15818a  and  a15813a );
 a15822a <=( A234  and  A233 );
 a15826a <=( (not A302)  and  (not A301) );
 a15827a <=( (not A300)  and  a15826a );
 a15828a <=( a15827a  and  a15822a );
 a15831a <=( (not A167)  and  (not A169) );
 a15835a <=( A201  and  A200 );
 a15836a <=( (not A166)  and  a15835a );
 a15837a <=( a15836a  and  a15831a );
 a15840a <=( A234  and  A233 );
 a15844a <=( (not A301)  and  (not A299) );
 a15845a <=( (not A298)  and  a15844a );
 a15846a <=( a15845a  and  a15840a );
 a15849a <=( (not A167)  and  (not A169) );
 a15853a <=( A201  and  A200 );
 a15854a <=( (not A166)  and  a15853a );
 a15855a <=( a15854a  and  a15849a );
 a15858a <=( A234  and  A233 );
 a15862a <=( A269  and  A266 );
 a15863a <=( (not A265)  and  a15862a );
 a15864a <=( a15863a  and  a15858a );
 a15867a <=( (not A167)  and  (not A169) );
 a15871a <=( A201  and  A200 );
 a15872a <=( (not A166)  and  a15871a );
 a15873a <=( a15872a  and  a15867a );
 a15876a <=( A234  and  A233 );
 a15880a <=( A269  and  (not A266) );
 a15881a <=( A265  and  a15880a );
 a15882a <=( a15881a  and  a15876a );
 a15885a <=( (not A167)  and  (not A169) );
 a15889a <=( A201  and  A200 );
 a15890a <=( (not A166)  and  a15889a );
 a15891a <=( a15890a  and  a15885a );
 a15894a <=( A233  and  (not A232) );
 a15898a <=( A267  and  A265 );
 a15899a <=( A236  and  a15898a );
 a15900a <=( a15899a  and  a15894a );
 a15903a <=( (not A167)  and  (not A169) );
 a15907a <=( A201  and  A200 );
 a15908a <=( (not A166)  and  a15907a );
 a15909a <=( a15908a  and  a15903a );
 a15912a <=( A233  and  (not A232) );
 a15916a <=( A267  and  A266 );
 a15917a <=( A236  and  a15916a );
 a15918a <=( a15917a  and  a15912a );
 a15921a <=( (not A167)  and  (not A169) );
 a15925a <=( A201  and  A200 );
 a15926a <=( (not A166)  and  a15925a );
 a15927a <=( a15926a  and  a15921a );
 a15930a <=( (not A233)  and  A232 );
 a15934a <=( A267  and  A265 );
 a15935a <=( A236  and  a15934a );
 a15936a <=( a15935a  and  a15930a );
 a15939a <=( (not A167)  and  (not A169) );
 a15943a <=( A201  and  A200 );
 a15944a <=( (not A166)  and  a15943a );
 a15945a <=( a15944a  and  a15939a );
 a15948a <=( (not A233)  and  A232 );
 a15952a <=( A267  and  A266 );
 a15953a <=( A236  and  a15952a );
 a15954a <=( a15953a  and  a15948a );
 a15957a <=( (not A167)  and  (not A169) );
 a15961a <=( A200  and  (not A199) );
 a15962a <=( (not A166)  and  a15961a );
 a15963a <=( a15962a  and  a15957a );
 a15966a <=( A235  and  A203 );
 a15970a <=( (not A302)  and  (not A301) );
 a15971a <=( (not A300)  and  a15970a );
 a15972a <=( a15971a  and  a15966a );
 a15975a <=( (not A167)  and  (not A169) );
 a15979a <=( A200  and  (not A199) );
 a15980a <=( (not A166)  and  a15979a );
 a15981a <=( a15980a  and  a15975a );
 a15984a <=( A235  and  A203 );
 a15988a <=( (not A301)  and  (not A299) );
 a15989a <=( (not A298)  and  a15988a );
 a15990a <=( a15989a  and  a15984a );
 a15993a <=( (not A167)  and  (not A169) );
 a15997a <=( A200  and  (not A199) );
 a15998a <=( (not A166)  and  a15997a );
 a15999a <=( a15998a  and  a15993a );
 a16002a <=( A235  and  A203 );
 a16006a <=( A269  and  A266 );
 a16007a <=( (not A265)  and  a16006a );
 a16008a <=( a16007a  and  a16002a );
 a16011a <=( (not A167)  and  (not A169) );
 a16015a <=( A200  and  (not A199) );
 a16016a <=( (not A166)  and  a16015a );
 a16017a <=( a16016a  and  a16011a );
 a16020a <=( A235  and  A203 );
 a16024a <=( A269  and  (not A266) );
 a16025a <=( A265  and  a16024a );
 a16026a <=( a16025a  and  a16020a );
 a16029a <=( (not A167)  and  (not A169) );
 a16033a <=( A200  and  (not A199) );
 a16034a <=( (not A166)  and  a16033a );
 a16035a <=( a16034a  and  a16029a );
 a16038a <=( A232  and  A203 );
 a16042a <=( A267  and  A265 );
 a16043a <=( A234  and  a16042a );
 a16044a <=( a16043a  and  a16038a );
 a16047a <=( (not A167)  and  (not A169) );
 a16051a <=( A200  and  (not A199) );
 a16052a <=( (not A166)  and  a16051a );
 a16053a <=( a16052a  and  a16047a );
 a16056a <=( A232  and  A203 );
 a16060a <=( A267  and  A266 );
 a16061a <=( A234  and  a16060a );
 a16062a <=( a16061a  and  a16056a );
 a16065a <=( (not A167)  and  (not A169) );
 a16069a <=( A200  and  (not A199) );
 a16070a <=( (not A166)  and  a16069a );
 a16071a <=( a16070a  and  a16065a );
 a16074a <=( A233  and  A203 );
 a16078a <=( A267  and  A265 );
 a16079a <=( A234  and  a16078a );
 a16080a <=( a16079a  and  a16074a );
 a16083a <=( (not A167)  and  (not A169) );
 a16087a <=( A200  and  (not A199) );
 a16088a <=( (not A166)  and  a16087a );
 a16089a <=( a16088a  and  a16083a );
 a16092a <=( A233  and  A203 );
 a16096a <=( A267  and  A266 );
 a16097a <=( A234  and  a16096a );
 a16098a <=( a16097a  and  a16092a );
 a16101a <=( (not A167)  and  (not A169) );
 a16105a <=( A200  and  (not A199) );
 a16106a <=( (not A166)  and  a16105a );
 a16107a <=( a16106a  and  a16101a );
 a16110a <=( (not A232)  and  A203 );
 a16114a <=( A268  and  A236 );
 a16115a <=( A233  and  a16114a );
 a16116a <=( a16115a  and  a16110a );
 a16119a <=( (not A167)  and  (not A169) );
 a16123a <=( A200  and  (not A199) );
 a16124a <=( (not A166)  and  a16123a );
 a16125a <=( a16124a  and  a16119a );
 a16128a <=( A232  and  A203 );
 a16132a <=( A268  and  A236 );
 a16133a <=( (not A233)  and  a16132a );
 a16134a <=( a16133a  and  a16128a );
 a16137a <=( (not A167)  and  (not A169) );
 a16141a <=( (not A200)  and  A199 );
 a16142a <=( (not A166)  and  a16141a );
 a16143a <=( a16142a  and  a16137a );
 a16146a <=( A235  and  A203 );
 a16150a <=( (not A302)  and  (not A301) );
 a16151a <=( (not A300)  and  a16150a );
 a16152a <=( a16151a  and  a16146a );
 a16155a <=( (not A167)  and  (not A169) );
 a16159a <=( (not A200)  and  A199 );
 a16160a <=( (not A166)  and  a16159a );
 a16161a <=( a16160a  and  a16155a );
 a16164a <=( A235  and  A203 );
 a16168a <=( (not A301)  and  (not A299) );
 a16169a <=( (not A298)  and  a16168a );
 a16170a <=( a16169a  and  a16164a );
 a16173a <=( (not A167)  and  (not A169) );
 a16177a <=( (not A200)  and  A199 );
 a16178a <=( (not A166)  and  a16177a );
 a16179a <=( a16178a  and  a16173a );
 a16182a <=( A235  and  A203 );
 a16186a <=( A269  and  A266 );
 a16187a <=( (not A265)  and  a16186a );
 a16188a <=( a16187a  and  a16182a );
 a16191a <=( (not A167)  and  (not A169) );
 a16195a <=( (not A200)  and  A199 );
 a16196a <=( (not A166)  and  a16195a );
 a16197a <=( a16196a  and  a16191a );
 a16200a <=( A235  and  A203 );
 a16204a <=( A269  and  (not A266) );
 a16205a <=( A265  and  a16204a );
 a16206a <=( a16205a  and  a16200a );
 a16209a <=( (not A167)  and  (not A169) );
 a16213a <=( (not A200)  and  A199 );
 a16214a <=( (not A166)  and  a16213a );
 a16215a <=( a16214a  and  a16209a );
 a16218a <=( A232  and  A203 );
 a16222a <=( A267  and  A265 );
 a16223a <=( A234  and  a16222a );
 a16224a <=( a16223a  and  a16218a );
 a16227a <=( (not A167)  and  (not A169) );
 a16231a <=( (not A200)  and  A199 );
 a16232a <=( (not A166)  and  a16231a );
 a16233a <=( a16232a  and  a16227a );
 a16236a <=( A232  and  A203 );
 a16240a <=( A267  and  A266 );
 a16241a <=( A234  and  a16240a );
 a16242a <=( a16241a  and  a16236a );
 a16245a <=( (not A167)  and  (not A169) );
 a16249a <=( (not A200)  and  A199 );
 a16250a <=( (not A166)  and  a16249a );
 a16251a <=( a16250a  and  a16245a );
 a16254a <=( A233  and  A203 );
 a16258a <=( A267  and  A265 );
 a16259a <=( A234  and  a16258a );
 a16260a <=( a16259a  and  a16254a );
 a16263a <=( (not A167)  and  (not A169) );
 a16267a <=( (not A200)  and  A199 );
 a16268a <=( (not A166)  and  a16267a );
 a16269a <=( a16268a  and  a16263a );
 a16272a <=( A233  and  A203 );
 a16276a <=( A267  and  A266 );
 a16277a <=( A234  and  a16276a );
 a16278a <=( a16277a  and  a16272a );
 a16281a <=( (not A167)  and  (not A169) );
 a16285a <=( (not A200)  and  A199 );
 a16286a <=( (not A166)  and  a16285a );
 a16287a <=( a16286a  and  a16281a );
 a16290a <=( (not A232)  and  A203 );
 a16294a <=( A268  and  A236 );
 a16295a <=( A233  and  a16294a );
 a16296a <=( a16295a  and  a16290a );
 a16299a <=( (not A167)  and  (not A169) );
 a16303a <=( (not A200)  and  A199 );
 a16304a <=( (not A166)  and  a16303a );
 a16305a <=( a16304a  and  a16299a );
 a16308a <=( A232  and  A203 );
 a16312a <=( A268  and  A236 );
 a16313a <=( (not A233)  and  a16312a );
 a16314a <=( a16313a  and  a16308a );
 a16317a <=( (not A168)  and  (not A169) );
 a16321a <=( A202  and  A166 );
 a16322a <=( A167  and  a16321a );
 a16323a <=( a16322a  and  a16317a );
 a16326a <=( A298  and  A235 );
 a16330a <=( (not A301)  and  (not A300) );
 a16331a <=( A299  and  a16330a );
 a16332a <=( a16331a  and  a16326a );
 a16335a <=( (not A168)  and  (not A169) );
 a16339a <=( A202  and  A166 );
 a16340a <=( A167  and  a16339a );
 a16341a <=( a16340a  and  a16335a );
 a16344a <=( A234  and  A232 );
 a16348a <=( (not A302)  and  (not A301) );
 a16349a <=( (not A300)  and  a16348a );
 a16350a <=( a16349a  and  a16344a );
 a16353a <=( (not A168)  and  (not A169) );
 a16357a <=( A202  and  A166 );
 a16358a <=( A167  and  a16357a );
 a16359a <=( a16358a  and  a16353a );
 a16362a <=( A234  and  A232 );
 a16366a <=( (not A301)  and  (not A299) );
 a16367a <=( (not A298)  and  a16366a );
 a16368a <=( a16367a  and  a16362a );
 a16371a <=( (not A168)  and  (not A169) );
 a16375a <=( A202  and  A166 );
 a16376a <=( A167  and  a16375a );
 a16377a <=( a16376a  and  a16371a );
 a16380a <=( A234  and  A232 );
 a16384a <=( A269  and  A266 );
 a16385a <=( (not A265)  and  a16384a );
 a16386a <=( a16385a  and  a16380a );
 a16389a <=( (not A168)  and  (not A169) );
 a16393a <=( A202  and  A166 );
 a16394a <=( A167  and  a16393a );
 a16395a <=( a16394a  and  a16389a );
 a16398a <=( A234  and  A232 );
 a16402a <=( A269  and  (not A266) );
 a16403a <=( A265  and  a16402a );
 a16404a <=( a16403a  and  a16398a );
 a16407a <=( (not A168)  and  (not A169) );
 a16411a <=( A202  and  A166 );
 a16412a <=( A167  and  a16411a );
 a16413a <=( a16412a  and  a16407a );
 a16416a <=( A234  and  A233 );
 a16420a <=( (not A302)  and  (not A301) );
 a16421a <=( (not A300)  and  a16420a );
 a16422a <=( a16421a  and  a16416a );
 a16425a <=( (not A168)  and  (not A169) );
 a16429a <=( A202  and  A166 );
 a16430a <=( A167  and  a16429a );
 a16431a <=( a16430a  and  a16425a );
 a16434a <=( A234  and  A233 );
 a16438a <=( (not A301)  and  (not A299) );
 a16439a <=( (not A298)  and  a16438a );
 a16440a <=( a16439a  and  a16434a );
 a16443a <=( (not A168)  and  (not A169) );
 a16447a <=( A202  and  A166 );
 a16448a <=( A167  and  a16447a );
 a16449a <=( a16448a  and  a16443a );
 a16452a <=( A234  and  A233 );
 a16456a <=( A269  and  A266 );
 a16457a <=( (not A265)  and  a16456a );
 a16458a <=( a16457a  and  a16452a );
 a16461a <=( (not A168)  and  (not A169) );
 a16465a <=( A202  and  A166 );
 a16466a <=( A167  and  a16465a );
 a16467a <=( a16466a  and  a16461a );
 a16470a <=( A234  and  A233 );
 a16474a <=( A269  and  (not A266) );
 a16475a <=( A265  and  a16474a );
 a16476a <=( a16475a  and  a16470a );
 a16479a <=( (not A168)  and  (not A169) );
 a16483a <=( A202  and  A166 );
 a16484a <=( A167  and  a16483a );
 a16485a <=( a16484a  and  a16479a );
 a16488a <=( A233  and  (not A232) );
 a16492a <=( A267  and  A265 );
 a16493a <=( A236  and  a16492a );
 a16494a <=( a16493a  and  a16488a );
 a16497a <=( (not A168)  and  (not A169) );
 a16501a <=( A202  and  A166 );
 a16502a <=( A167  and  a16501a );
 a16503a <=( a16502a  and  a16497a );
 a16506a <=( A233  and  (not A232) );
 a16510a <=( A267  and  A266 );
 a16511a <=( A236  and  a16510a );
 a16512a <=( a16511a  and  a16506a );
 a16515a <=( (not A168)  and  (not A169) );
 a16519a <=( A202  and  A166 );
 a16520a <=( A167  and  a16519a );
 a16521a <=( a16520a  and  a16515a );
 a16524a <=( (not A233)  and  A232 );
 a16528a <=( A267  and  A265 );
 a16529a <=( A236  and  a16528a );
 a16530a <=( a16529a  and  a16524a );
 a16533a <=( (not A168)  and  (not A169) );
 a16537a <=( A202  and  A166 );
 a16538a <=( A167  and  a16537a );
 a16539a <=( a16538a  and  a16533a );
 a16542a <=( (not A233)  and  A232 );
 a16546a <=( A267  and  A266 );
 a16547a <=( A236  and  a16546a );
 a16548a <=( a16547a  and  a16542a );
 a16551a <=( (not A168)  and  (not A169) );
 a16555a <=( A199  and  A166 );
 a16556a <=( A167  and  a16555a );
 a16557a <=( a16556a  and  a16551a );
 a16560a <=( A235  and  A201 );
 a16564a <=( (not A302)  and  (not A301) );
 a16565a <=( (not A300)  and  a16564a );
 a16566a <=( a16565a  and  a16560a );
 a16569a <=( (not A168)  and  (not A169) );
 a16573a <=( A199  and  A166 );
 a16574a <=( A167  and  a16573a );
 a16575a <=( a16574a  and  a16569a );
 a16578a <=( A235  and  A201 );
 a16582a <=( (not A301)  and  (not A299) );
 a16583a <=( (not A298)  and  a16582a );
 a16584a <=( a16583a  and  a16578a );
 a16587a <=( (not A168)  and  (not A169) );
 a16591a <=( A199  and  A166 );
 a16592a <=( A167  and  a16591a );
 a16593a <=( a16592a  and  a16587a );
 a16596a <=( A235  and  A201 );
 a16600a <=( A269  and  A266 );
 a16601a <=( (not A265)  and  a16600a );
 a16602a <=( a16601a  and  a16596a );
 a16605a <=( (not A168)  and  (not A169) );
 a16609a <=( A199  and  A166 );
 a16610a <=( A167  and  a16609a );
 a16611a <=( a16610a  and  a16605a );
 a16614a <=( A235  and  A201 );
 a16618a <=( A269  and  (not A266) );
 a16619a <=( A265  and  a16618a );
 a16620a <=( a16619a  and  a16614a );
 a16623a <=( (not A168)  and  (not A169) );
 a16627a <=( A199  and  A166 );
 a16628a <=( A167  and  a16627a );
 a16629a <=( a16628a  and  a16623a );
 a16632a <=( A232  and  A201 );
 a16636a <=( A267  and  A265 );
 a16637a <=( A234  and  a16636a );
 a16638a <=( a16637a  and  a16632a );
 a16641a <=( (not A168)  and  (not A169) );
 a16645a <=( A199  and  A166 );
 a16646a <=( A167  and  a16645a );
 a16647a <=( a16646a  and  a16641a );
 a16650a <=( A232  and  A201 );
 a16654a <=( A267  and  A266 );
 a16655a <=( A234  and  a16654a );
 a16656a <=( a16655a  and  a16650a );
 a16659a <=( (not A168)  and  (not A169) );
 a16663a <=( A199  and  A166 );
 a16664a <=( A167  and  a16663a );
 a16665a <=( a16664a  and  a16659a );
 a16668a <=( A233  and  A201 );
 a16672a <=( A267  and  A265 );
 a16673a <=( A234  and  a16672a );
 a16674a <=( a16673a  and  a16668a );
 a16677a <=( (not A168)  and  (not A169) );
 a16681a <=( A199  and  A166 );
 a16682a <=( A167  and  a16681a );
 a16683a <=( a16682a  and  a16677a );
 a16686a <=( A233  and  A201 );
 a16690a <=( A267  and  A266 );
 a16691a <=( A234  and  a16690a );
 a16692a <=( a16691a  and  a16686a );
 a16695a <=( (not A168)  and  (not A169) );
 a16699a <=( A199  and  A166 );
 a16700a <=( A167  and  a16699a );
 a16701a <=( a16700a  and  a16695a );
 a16704a <=( (not A232)  and  A201 );
 a16708a <=( A268  and  A236 );
 a16709a <=( A233  and  a16708a );
 a16710a <=( a16709a  and  a16704a );
 a16713a <=( (not A168)  and  (not A169) );
 a16717a <=( A199  and  A166 );
 a16718a <=( A167  and  a16717a );
 a16719a <=( a16718a  and  a16713a );
 a16722a <=( A232  and  A201 );
 a16726a <=( A268  and  A236 );
 a16727a <=( (not A233)  and  a16726a );
 a16728a <=( a16727a  and  a16722a );
 a16731a <=( (not A168)  and  (not A169) );
 a16735a <=( A200  and  A166 );
 a16736a <=( A167  and  a16735a );
 a16737a <=( a16736a  and  a16731a );
 a16740a <=( A235  and  A201 );
 a16744a <=( (not A302)  and  (not A301) );
 a16745a <=( (not A300)  and  a16744a );
 a16746a <=( a16745a  and  a16740a );
 a16749a <=( (not A168)  and  (not A169) );
 a16753a <=( A200  and  A166 );
 a16754a <=( A167  and  a16753a );
 a16755a <=( a16754a  and  a16749a );
 a16758a <=( A235  and  A201 );
 a16762a <=( (not A301)  and  (not A299) );
 a16763a <=( (not A298)  and  a16762a );
 a16764a <=( a16763a  and  a16758a );
 a16767a <=( (not A168)  and  (not A169) );
 a16771a <=( A200  and  A166 );
 a16772a <=( A167  and  a16771a );
 a16773a <=( a16772a  and  a16767a );
 a16776a <=( A235  and  A201 );
 a16780a <=( A269  and  A266 );
 a16781a <=( (not A265)  and  a16780a );
 a16782a <=( a16781a  and  a16776a );
 a16785a <=( (not A168)  and  (not A169) );
 a16789a <=( A200  and  A166 );
 a16790a <=( A167  and  a16789a );
 a16791a <=( a16790a  and  a16785a );
 a16794a <=( A235  and  A201 );
 a16798a <=( A269  and  (not A266) );
 a16799a <=( A265  and  a16798a );
 a16800a <=( a16799a  and  a16794a );
 a16803a <=( (not A168)  and  (not A169) );
 a16807a <=( A200  and  A166 );
 a16808a <=( A167  and  a16807a );
 a16809a <=( a16808a  and  a16803a );
 a16812a <=( A232  and  A201 );
 a16816a <=( A267  and  A265 );
 a16817a <=( A234  and  a16816a );
 a16818a <=( a16817a  and  a16812a );
 a16821a <=( (not A168)  and  (not A169) );
 a16825a <=( A200  and  A166 );
 a16826a <=( A167  and  a16825a );
 a16827a <=( a16826a  and  a16821a );
 a16830a <=( A232  and  A201 );
 a16834a <=( A267  and  A266 );
 a16835a <=( A234  and  a16834a );
 a16836a <=( a16835a  and  a16830a );
 a16839a <=( (not A168)  and  (not A169) );
 a16843a <=( A200  and  A166 );
 a16844a <=( A167  and  a16843a );
 a16845a <=( a16844a  and  a16839a );
 a16848a <=( A233  and  A201 );
 a16852a <=( A267  and  A265 );
 a16853a <=( A234  and  a16852a );
 a16854a <=( a16853a  and  a16848a );
 a16857a <=( (not A168)  and  (not A169) );
 a16861a <=( A200  and  A166 );
 a16862a <=( A167  and  a16861a );
 a16863a <=( a16862a  and  a16857a );
 a16866a <=( A233  and  A201 );
 a16870a <=( A267  and  A266 );
 a16871a <=( A234  and  a16870a );
 a16872a <=( a16871a  and  a16866a );
 a16875a <=( (not A168)  and  (not A169) );
 a16879a <=( A200  and  A166 );
 a16880a <=( A167  and  a16879a );
 a16881a <=( a16880a  and  a16875a );
 a16884a <=( (not A232)  and  A201 );
 a16888a <=( A268  and  A236 );
 a16889a <=( A233  and  a16888a );
 a16890a <=( a16889a  and  a16884a );
 a16893a <=( (not A168)  and  (not A169) );
 a16897a <=( A200  and  A166 );
 a16898a <=( A167  and  a16897a );
 a16899a <=( a16898a  and  a16893a );
 a16902a <=( A232  and  A201 );
 a16906a <=( A268  and  A236 );
 a16907a <=( (not A233)  and  a16906a );
 a16908a <=( a16907a  and  a16902a );
 a16911a <=( (not A168)  and  (not A169) );
 a16915a <=( (not A199)  and  A166 );
 a16916a <=( A167  and  a16915a );
 a16917a <=( a16916a  and  a16911a );
 a16920a <=( A203  and  A200 );
 a16924a <=( A267  and  A265 );
 a16925a <=( A235  and  a16924a );
 a16926a <=( a16925a  and  a16920a );
 a16929a <=( (not A168)  and  (not A169) );
 a16933a <=( (not A199)  and  A166 );
 a16934a <=( A167  and  a16933a );
 a16935a <=( a16934a  and  a16929a );
 a16938a <=( A203  and  A200 );
 a16942a <=( A267  and  A266 );
 a16943a <=( A235  and  a16942a );
 a16944a <=( a16943a  and  a16938a );
 a16947a <=( (not A168)  and  (not A169) );
 a16951a <=( (not A199)  and  A166 );
 a16952a <=( A167  and  a16951a );
 a16953a <=( a16952a  and  a16947a );
 a16956a <=( A203  and  A200 );
 a16960a <=( A268  and  A234 );
 a16961a <=( A232  and  a16960a );
 a16962a <=( a16961a  and  a16956a );
 a16965a <=( (not A168)  and  (not A169) );
 a16969a <=( (not A199)  and  A166 );
 a16970a <=( A167  and  a16969a );
 a16971a <=( a16970a  and  a16965a );
 a16974a <=( A203  and  A200 );
 a16978a <=( A268  and  A234 );
 a16979a <=( A233  and  a16978a );
 a16980a <=( a16979a  and  a16974a );
 a16983a <=( (not A168)  and  (not A169) );
 a16987a <=( A199  and  A166 );
 a16988a <=( A167  and  a16987a );
 a16989a <=( a16988a  and  a16983a );
 a16992a <=( A203  and  (not A200) );
 a16996a <=( A267  and  A265 );
 a16997a <=( A235  and  a16996a );
 a16998a <=( a16997a  and  a16992a );
 a17001a <=( (not A168)  and  (not A169) );
 a17005a <=( A199  and  A166 );
 a17006a <=( A167  and  a17005a );
 a17007a <=( a17006a  and  a17001a );
 a17010a <=( A203  and  (not A200) );
 a17014a <=( A267  and  A266 );
 a17015a <=( A235  and  a17014a );
 a17016a <=( a17015a  and  a17010a );
 a17019a <=( (not A168)  and  (not A169) );
 a17023a <=( A199  and  A166 );
 a17024a <=( A167  and  a17023a );
 a17025a <=( a17024a  and  a17019a );
 a17028a <=( A203  and  (not A200) );
 a17032a <=( A268  and  A234 );
 a17033a <=( A232  and  a17032a );
 a17034a <=( a17033a  and  a17028a );
 a17037a <=( (not A168)  and  (not A169) );
 a17041a <=( A199  and  A166 );
 a17042a <=( A167  and  a17041a );
 a17043a <=( a17042a  and  a17037a );
 a17046a <=( A203  and  (not A200) );
 a17050a <=( A268  and  A234 );
 a17051a <=( A233  and  a17050a );
 a17052a <=( a17051a  and  a17046a );
 a17055a <=( (not A169)  and  (not A170) );
 a17059a <=( A232  and  A202 );
 a17060a <=( (not A168)  and  a17059a );
 a17061a <=( a17060a  and  a17055a );
 a17064a <=( A298  and  A234 );
 a17068a <=( (not A301)  and  (not A300) );
 a17069a <=( A299  and  a17068a );
 a17070a <=( a17069a  and  a17064a );
 a17073a <=( (not A169)  and  (not A170) );
 a17077a <=( A233  and  A202 );
 a17078a <=( (not A168)  and  a17077a );
 a17079a <=( a17078a  and  a17073a );
 a17082a <=( A298  and  A234 );
 a17086a <=( (not A301)  and  (not A300) );
 a17087a <=( A299  and  a17086a );
 a17088a <=( a17087a  and  a17082a );
 a17091a <=( (not A169)  and  (not A170) );
 a17095a <=( (not A232)  and  A202 );
 a17096a <=( (not A168)  and  a17095a );
 a17097a <=( a17096a  and  a17091a );
 a17100a <=( A236  and  A233 );
 a17104a <=( (not A302)  and  (not A301) );
 a17105a <=( (not A300)  and  a17104a );
 a17106a <=( a17105a  and  a17100a );
 a17109a <=( (not A169)  and  (not A170) );
 a17113a <=( (not A232)  and  A202 );
 a17114a <=( (not A168)  and  a17113a );
 a17115a <=( a17114a  and  a17109a );
 a17118a <=( A236  and  A233 );
 a17122a <=( (not A301)  and  (not A299) );
 a17123a <=( (not A298)  and  a17122a );
 a17124a <=( a17123a  and  a17118a );
 a17127a <=( (not A169)  and  (not A170) );
 a17131a <=( (not A232)  and  A202 );
 a17132a <=( (not A168)  and  a17131a );
 a17133a <=( a17132a  and  a17127a );
 a17136a <=( A236  and  A233 );
 a17140a <=( A269  and  A266 );
 a17141a <=( (not A265)  and  a17140a );
 a17142a <=( a17141a  and  a17136a );
 a17145a <=( (not A169)  and  (not A170) );
 a17149a <=( (not A232)  and  A202 );
 a17150a <=( (not A168)  and  a17149a );
 a17151a <=( a17150a  and  a17145a );
 a17154a <=( A236  and  A233 );
 a17158a <=( A269  and  (not A266) );
 a17159a <=( A265  and  a17158a );
 a17160a <=( a17159a  and  a17154a );
 a17163a <=( (not A169)  and  (not A170) );
 a17167a <=( A232  and  A202 );
 a17168a <=( (not A168)  and  a17167a );
 a17169a <=( a17168a  and  a17163a );
 a17172a <=( A236  and  (not A233) );
 a17176a <=( (not A302)  and  (not A301) );
 a17177a <=( (not A300)  and  a17176a );
 a17178a <=( a17177a  and  a17172a );
 a17181a <=( (not A169)  and  (not A170) );
 a17185a <=( A232  and  A202 );
 a17186a <=( (not A168)  and  a17185a );
 a17187a <=( a17186a  and  a17181a );
 a17190a <=( A236  and  (not A233) );
 a17194a <=( (not A301)  and  (not A299) );
 a17195a <=( (not A298)  and  a17194a );
 a17196a <=( a17195a  and  a17190a );
 a17199a <=( (not A169)  and  (not A170) );
 a17203a <=( A232  and  A202 );
 a17204a <=( (not A168)  and  a17203a );
 a17205a <=( a17204a  and  a17199a );
 a17208a <=( A236  and  (not A233) );
 a17212a <=( A269  and  A266 );
 a17213a <=( (not A265)  and  a17212a );
 a17214a <=( a17213a  and  a17208a );
 a17217a <=( (not A169)  and  (not A170) );
 a17221a <=( A232  and  A202 );
 a17222a <=( (not A168)  and  a17221a );
 a17223a <=( a17222a  and  a17217a );
 a17226a <=( A236  and  (not A233) );
 a17230a <=( A269  and  (not A266) );
 a17231a <=( A265  and  a17230a );
 a17232a <=( a17231a  and  a17226a );
 a17235a <=( (not A169)  and  (not A170) );
 a17239a <=( A201  and  A199 );
 a17240a <=( (not A168)  and  a17239a );
 a17241a <=( a17240a  and  a17235a );
 a17244a <=( A298  and  A235 );
 a17248a <=( (not A301)  and  (not A300) );
 a17249a <=( A299  and  a17248a );
 a17250a <=( a17249a  and  a17244a );
 a17253a <=( (not A169)  and  (not A170) );
 a17257a <=( A201  and  A199 );
 a17258a <=( (not A168)  and  a17257a );
 a17259a <=( a17258a  and  a17253a );
 a17262a <=( A234  and  A232 );
 a17266a <=( (not A302)  and  (not A301) );
 a17267a <=( (not A300)  and  a17266a );
 a17268a <=( a17267a  and  a17262a );
 a17271a <=( (not A169)  and  (not A170) );
 a17275a <=( A201  and  A199 );
 a17276a <=( (not A168)  and  a17275a );
 a17277a <=( a17276a  and  a17271a );
 a17280a <=( A234  and  A232 );
 a17284a <=( (not A301)  and  (not A299) );
 a17285a <=( (not A298)  and  a17284a );
 a17286a <=( a17285a  and  a17280a );
 a17289a <=( (not A169)  and  (not A170) );
 a17293a <=( A201  and  A199 );
 a17294a <=( (not A168)  and  a17293a );
 a17295a <=( a17294a  and  a17289a );
 a17298a <=( A234  and  A232 );
 a17302a <=( A269  and  A266 );
 a17303a <=( (not A265)  and  a17302a );
 a17304a <=( a17303a  and  a17298a );
 a17307a <=( (not A169)  and  (not A170) );
 a17311a <=( A201  and  A199 );
 a17312a <=( (not A168)  and  a17311a );
 a17313a <=( a17312a  and  a17307a );
 a17316a <=( A234  and  A232 );
 a17320a <=( A269  and  (not A266) );
 a17321a <=( A265  and  a17320a );
 a17322a <=( a17321a  and  a17316a );
 a17325a <=( (not A169)  and  (not A170) );
 a17329a <=( A201  and  A199 );
 a17330a <=( (not A168)  and  a17329a );
 a17331a <=( a17330a  and  a17325a );
 a17334a <=( A234  and  A233 );
 a17338a <=( (not A302)  and  (not A301) );
 a17339a <=( (not A300)  and  a17338a );
 a17340a <=( a17339a  and  a17334a );
 a17343a <=( (not A169)  and  (not A170) );
 a17347a <=( A201  and  A199 );
 a17348a <=( (not A168)  and  a17347a );
 a17349a <=( a17348a  and  a17343a );
 a17352a <=( A234  and  A233 );
 a17356a <=( (not A301)  and  (not A299) );
 a17357a <=( (not A298)  and  a17356a );
 a17358a <=( a17357a  and  a17352a );
 a17361a <=( (not A169)  and  (not A170) );
 a17365a <=( A201  and  A199 );
 a17366a <=( (not A168)  and  a17365a );
 a17367a <=( a17366a  and  a17361a );
 a17370a <=( A234  and  A233 );
 a17374a <=( A269  and  A266 );
 a17375a <=( (not A265)  and  a17374a );
 a17376a <=( a17375a  and  a17370a );
 a17379a <=( (not A169)  and  (not A170) );
 a17383a <=( A201  and  A199 );
 a17384a <=( (not A168)  and  a17383a );
 a17385a <=( a17384a  and  a17379a );
 a17388a <=( A234  and  A233 );
 a17392a <=( A269  and  (not A266) );
 a17393a <=( A265  and  a17392a );
 a17394a <=( a17393a  and  a17388a );
 a17397a <=( (not A169)  and  (not A170) );
 a17401a <=( A201  and  A199 );
 a17402a <=( (not A168)  and  a17401a );
 a17403a <=( a17402a  and  a17397a );
 a17406a <=( A233  and  (not A232) );
 a17410a <=( A267  and  A265 );
 a17411a <=( A236  and  a17410a );
 a17412a <=( a17411a  and  a17406a );
 a17415a <=( (not A169)  and  (not A170) );
 a17419a <=( A201  and  A199 );
 a17420a <=( (not A168)  and  a17419a );
 a17421a <=( a17420a  and  a17415a );
 a17424a <=( A233  and  (not A232) );
 a17428a <=( A267  and  A266 );
 a17429a <=( A236  and  a17428a );
 a17430a <=( a17429a  and  a17424a );
 a17433a <=( (not A169)  and  (not A170) );
 a17437a <=( A201  and  A199 );
 a17438a <=( (not A168)  and  a17437a );
 a17439a <=( a17438a  and  a17433a );
 a17442a <=( (not A233)  and  A232 );
 a17446a <=( A267  and  A265 );
 a17447a <=( A236  and  a17446a );
 a17448a <=( a17447a  and  a17442a );
 a17451a <=( (not A169)  and  (not A170) );
 a17455a <=( A201  and  A199 );
 a17456a <=( (not A168)  and  a17455a );
 a17457a <=( a17456a  and  a17451a );
 a17460a <=( (not A233)  and  A232 );
 a17464a <=( A267  and  A266 );
 a17465a <=( A236  and  a17464a );
 a17466a <=( a17465a  and  a17460a );
 a17469a <=( (not A169)  and  (not A170) );
 a17473a <=( A201  and  A200 );
 a17474a <=( (not A168)  and  a17473a );
 a17475a <=( a17474a  and  a17469a );
 a17478a <=( A298  and  A235 );
 a17482a <=( (not A301)  and  (not A300) );
 a17483a <=( A299  and  a17482a );
 a17484a <=( a17483a  and  a17478a );
 a17487a <=( (not A169)  and  (not A170) );
 a17491a <=( A201  and  A200 );
 a17492a <=( (not A168)  and  a17491a );
 a17493a <=( a17492a  and  a17487a );
 a17496a <=( A234  and  A232 );
 a17500a <=( (not A302)  and  (not A301) );
 a17501a <=( (not A300)  and  a17500a );
 a17502a <=( a17501a  and  a17496a );
 a17505a <=( (not A169)  and  (not A170) );
 a17509a <=( A201  and  A200 );
 a17510a <=( (not A168)  and  a17509a );
 a17511a <=( a17510a  and  a17505a );
 a17514a <=( A234  and  A232 );
 a17518a <=( (not A301)  and  (not A299) );
 a17519a <=( (not A298)  and  a17518a );
 a17520a <=( a17519a  and  a17514a );
 a17523a <=( (not A169)  and  (not A170) );
 a17527a <=( A201  and  A200 );
 a17528a <=( (not A168)  and  a17527a );
 a17529a <=( a17528a  and  a17523a );
 a17532a <=( A234  and  A232 );
 a17536a <=( A269  and  A266 );
 a17537a <=( (not A265)  and  a17536a );
 a17538a <=( a17537a  and  a17532a );
 a17541a <=( (not A169)  and  (not A170) );
 a17545a <=( A201  and  A200 );
 a17546a <=( (not A168)  and  a17545a );
 a17547a <=( a17546a  and  a17541a );
 a17550a <=( A234  and  A232 );
 a17554a <=( A269  and  (not A266) );
 a17555a <=( A265  and  a17554a );
 a17556a <=( a17555a  and  a17550a );
 a17559a <=( (not A169)  and  (not A170) );
 a17563a <=( A201  and  A200 );
 a17564a <=( (not A168)  and  a17563a );
 a17565a <=( a17564a  and  a17559a );
 a17568a <=( A234  and  A233 );
 a17572a <=( (not A302)  and  (not A301) );
 a17573a <=( (not A300)  and  a17572a );
 a17574a <=( a17573a  and  a17568a );
 a17577a <=( (not A169)  and  (not A170) );
 a17581a <=( A201  and  A200 );
 a17582a <=( (not A168)  and  a17581a );
 a17583a <=( a17582a  and  a17577a );
 a17586a <=( A234  and  A233 );
 a17590a <=( (not A301)  and  (not A299) );
 a17591a <=( (not A298)  and  a17590a );
 a17592a <=( a17591a  and  a17586a );
 a17595a <=( (not A169)  and  (not A170) );
 a17599a <=( A201  and  A200 );
 a17600a <=( (not A168)  and  a17599a );
 a17601a <=( a17600a  and  a17595a );
 a17604a <=( A234  and  A233 );
 a17608a <=( A269  and  A266 );
 a17609a <=( (not A265)  and  a17608a );
 a17610a <=( a17609a  and  a17604a );
 a17613a <=( (not A169)  and  (not A170) );
 a17617a <=( A201  and  A200 );
 a17618a <=( (not A168)  and  a17617a );
 a17619a <=( a17618a  and  a17613a );
 a17622a <=( A234  and  A233 );
 a17626a <=( A269  and  (not A266) );
 a17627a <=( A265  and  a17626a );
 a17628a <=( a17627a  and  a17622a );
 a17631a <=( (not A169)  and  (not A170) );
 a17635a <=( A201  and  A200 );
 a17636a <=( (not A168)  and  a17635a );
 a17637a <=( a17636a  and  a17631a );
 a17640a <=( A233  and  (not A232) );
 a17644a <=( A267  and  A265 );
 a17645a <=( A236  and  a17644a );
 a17646a <=( a17645a  and  a17640a );
 a17649a <=( (not A169)  and  (not A170) );
 a17653a <=( A201  and  A200 );
 a17654a <=( (not A168)  and  a17653a );
 a17655a <=( a17654a  and  a17649a );
 a17658a <=( A233  and  (not A232) );
 a17662a <=( A267  and  A266 );
 a17663a <=( A236  and  a17662a );
 a17664a <=( a17663a  and  a17658a );
 a17667a <=( (not A169)  and  (not A170) );
 a17671a <=( A201  and  A200 );
 a17672a <=( (not A168)  and  a17671a );
 a17673a <=( a17672a  and  a17667a );
 a17676a <=( (not A233)  and  A232 );
 a17680a <=( A267  and  A265 );
 a17681a <=( A236  and  a17680a );
 a17682a <=( a17681a  and  a17676a );
 a17685a <=( (not A169)  and  (not A170) );
 a17689a <=( A201  and  A200 );
 a17690a <=( (not A168)  and  a17689a );
 a17691a <=( a17690a  and  a17685a );
 a17694a <=( (not A233)  and  A232 );
 a17698a <=( A267  and  A266 );
 a17699a <=( A236  and  a17698a );
 a17700a <=( a17699a  and  a17694a );
 a17703a <=( (not A169)  and  (not A170) );
 a17707a <=( A200  and  (not A199) );
 a17708a <=( (not A168)  and  a17707a );
 a17709a <=( a17708a  and  a17703a );
 a17712a <=( A235  and  A203 );
 a17716a <=( (not A302)  and  (not A301) );
 a17717a <=( (not A300)  and  a17716a );
 a17718a <=( a17717a  and  a17712a );
 a17721a <=( (not A169)  and  (not A170) );
 a17725a <=( A200  and  (not A199) );
 a17726a <=( (not A168)  and  a17725a );
 a17727a <=( a17726a  and  a17721a );
 a17730a <=( A235  and  A203 );
 a17734a <=( (not A301)  and  (not A299) );
 a17735a <=( (not A298)  and  a17734a );
 a17736a <=( a17735a  and  a17730a );
 a17739a <=( (not A169)  and  (not A170) );
 a17743a <=( A200  and  (not A199) );
 a17744a <=( (not A168)  and  a17743a );
 a17745a <=( a17744a  and  a17739a );
 a17748a <=( A235  and  A203 );
 a17752a <=( A269  and  A266 );
 a17753a <=( (not A265)  and  a17752a );
 a17754a <=( a17753a  and  a17748a );
 a17757a <=( (not A169)  and  (not A170) );
 a17761a <=( A200  and  (not A199) );
 a17762a <=( (not A168)  and  a17761a );
 a17763a <=( a17762a  and  a17757a );
 a17766a <=( A235  and  A203 );
 a17770a <=( A269  and  (not A266) );
 a17771a <=( A265  and  a17770a );
 a17772a <=( a17771a  and  a17766a );
 a17775a <=( (not A169)  and  (not A170) );
 a17779a <=( A200  and  (not A199) );
 a17780a <=( (not A168)  and  a17779a );
 a17781a <=( a17780a  and  a17775a );
 a17784a <=( A232  and  A203 );
 a17788a <=( A267  and  A265 );
 a17789a <=( A234  and  a17788a );
 a17790a <=( a17789a  and  a17784a );
 a17793a <=( (not A169)  and  (not A170) );
 a17797a <=( A200  and  (not A199) );
 a17798a <=( (not A168)  and  a17797a );
 a17799a <=( a17798a  and  a17793a );
 a17802a <=( A232  and  A203 );
 a17806a <=( A267  and  A266 );
 a17807a <=( A234  and  a17806a );
 a17808a <=( a17807a  and  a17802a );
 a17811a <=( (not A169)  and  (not A170) );
 a17815a <=( A200  and  (not A199) );
 a17816a <=( (not A168)  and  a17815a );
 a17817a <=( a17816a  and  a17811a );
 a17820a <=( A233  and  A203 );
 a17824a <=( A267  and  A265 );
 a17825a <=( A234  and  a17824a );
 a17826a <=( a17825a  and  a17820a );
 a17829a <=( (not A169)  and  (not A170) );
 a17833a <=( A200  and  (not A199) );
 a17834a <=( (not A168)  and  a17833a );
 a17835a <=( a17834a  and  a17829a );
 a17838a <=( A233  and  A203 );
 a17842a <=( A267  and  A266 );
 a17843a <=( A234  and  a17842a );
 a17844a <=( a17843a  and  a17838a );
 a17847a <=( (not A169)  and  (not A170) );
 a17851a <=( A200  and  (not A199) );
 a17852a <=( (not A168)  and  a17851a );
 a17853a <=( a17852a  and  a17847a );
 a17856a <=( (not A232)  and  A203 );
 a17860a <=( A268  and  A236 );
 a17861a <=( A233  and  a17860a );
 a17862a <=( a17861a  and  a17856a );
 a17865a <=( (not A169)  and  (not A170) );
 a17869a <=( A200  and  (not A199) );
 a17870a <=( (not A168)  and  a17869a );
 a17871a <=( a17870a  and  a17865a );
 a17874a <=( A232  and  A203 );
 a17878a <=( A268  and  A236 );
 a17879a <=( (not A233)  and  a17878a );
 a17880a <=( a17879a  and  a17874a );
 a17883a <=( (not A169)  and  (not A170) );
 a17887a <=( (not A200)  and  A199 );
 a17888a <=( (not A168)  and  a17887a );
 a17889a <=( a17888a  and  a17883a );
 a17892a <=( A235  and  A203 );
 a17896a <=( (not A302)  and  (not A301) );
 a17897a <=( (not A300)  and  a17896a );
 a17898a <=( a17897a  and  a17892a );
 a17901a <=( (not A169)  and  (not A170) );
 a17905a <=( (not A200)  and  A199 );
 a17906a <=( (not A168)  and  a17905a );
 a17907a <=( a17906a  and  a17901a );
 a17910a <=( A235  and  A203 );
 a17914a <=( (not A301)  and  (not A299) );
 a17915a <=( (not A298)  and  a17914a );
 a17916a <=( a17915a  and  a17910a );
 a17919a <=( (not A169)  and  (not A170) );
 a17923a <=( (not A200)  and  A199 );
 a17924a <=( (not A168)  and  a17923a );
 a17925a <=( a17924a  and  a17919a );
 a17928a <=( A235  and  A203 );
 a17932a <=( A269  and  A266 );
 a17933a <=( (not A265)  and  a17932a );
 a17934a <=( a17933a  and  a17928a );
 a17937a <=( (not A169)  and  (not A170) );
 a17941a <=( (not A200)  and  A199 );
 a17942a <=( (not A168)  and  a17941a );
 a17943a <=( a17942a  and  a17937a );
 a17946a <=( A235  and  A203 );
 a17950a <=( A269  and  (not A266) );
 a17951a <=( A265  and  a17950a );
 a17952a <=( a17951a  and  a17946a );
 a17955a <=( (not A169)  and  (not A170) );
 a17959a <=( (not A200)  and  A199 );
 a17960a <=( (not A168)  and  a17959a );
 a17961a <=( a17960a  and  a17955a );
 a17964a <=( A232  and  A203 );
 a17968a <=( A267  and  A265 );
 a17969a <=( A234  and  a17968a );
 a17970a <=( a17969a  and  a17964a );
 a17973a <=( (not A169)  and  (not A170) );
 a17977a <=( (not A200)  and  A199 );
 a17978a <=( (not A168)  and  a17977a );
 a17979a <=( a17978a  and  a17973a );
 a17982a <=( A232  and  A203 );
 a17986a <=( A267  and  A266 );
 a17987a <=( A234  and  a17986a );
 a17988a <=( a17987a  and  a17982a );
 a17991a <=( (not A169)  and  (not A170) );
 a17995a <=( (not A200)  and  A199 );
 a17996a <=( (not A168)  and  a17995a );
 a17997a <=( a17996a  and  a17991a );
 a18000a <=( A233  and  A203 );
 a18004a <=( A267  and  A265 );
 a18005a <=( A234  and  a18004a );
 a18006a <=( a18005a  and  a18000a );
 a18009a <=( (not A169)  and  (not A170) );
 a18013a <=( (not A200)  and  A199 );
 a18014a <=( (not A168)  and  a18013a );
 a18015a <=( a18014a  and  a18009a );
 a18018a <=( A233  and  A203 );
 a18022a <=( A267  and  A266 );
 a18023a <=( A234  and  a18022a );
 a18024a <=( a18023a  and  a18018a );
 a18027a <=( (not A169)  and  (not A170) );
 a18031a <=( (not A200)  and  A199 );
 a18032a <=( (not A168)  and  a18031a );
 a18033a <=( a18032a  and  a18027a );
 a18036a <=( (not A232)  and  A203 );
 a18040a <=( A268  and  A236 );
 a18041a <=( A233  and  a18040a );
 a18042a <=( a18041a  and  a18036a );
 a18045a <=( (not A169)  and  (not A170) );
 a18049a <=( (not A200)  and  A199 );
 a18050a <=( (not A168)  and  a18049a );
 a18051a <=( a18050a  and  a18045a );
 a18054a <=( A232  and  A203 );
 a18058a <=( A268  and  A236 );
 a18059a <=( (not A233)  and  a18058a );
 a18060a <=( a18059a  and  a18054a );
 a18063a <=( A166  and  A168 );
 a18067a <=( (not A203)  and  (not A202) );
 a18068a <=( (not A201)  and  a18067a );
 a18069a <=( a18068a  and  a18063a );
 a18073a <=( A298  and  A234 );
 a18074a <=( A232  and  a18073a );
 a18078a <=( (not A301)  and  (not A300) );
 a18079a <=( A299  and  a18078a );
 a18080a <=( a18079a  and  a18074a );
 a18083a <=( A166  and  A168 );
 a18087a <=( (not A203)  and  (not A202) );
 a18088a <=( (not A201)  and  a18087a );
 a18089a <=( a18088a  and  a18083a );
 a18093a <=( A298  and  A234 );
 a18094a <=( A233  and  a18093a );
 a18098a <=( (not A301)  and  (not A300) );
 a18099a <=( A299  and  a18098a );
 a18100a <=( a18099a  and  a18094a );
 a18103a <=( A166  and  A168 );
 a18107a <=( (not A203)  and  (not A202) );
 a18108a <=( (not A201)  and  a18107a );
 a18109a <=( a18108a  and  a18103a );
 a18113a <=( A236  and  A233 );
 a18114a <=( (not A232)  and  a18113a );
 a18118a <=( (not A302)  and  (not A301) );
 a18119a <=( (not A300)  and  a18118a );
 a18120a <=( a18119a  and  a18114a );
 a18123a <=( A166  and  A168 );
 a18127a <=( (not A203)  and  (not A202) );
 a18128a <=( (not A201)  and  a18127a );
 a18129a <=( a18128a  and  a18123a );
 a18133a <=( A236  and  A233 );
 a18134a <=( (not A232)  and  a18133a );
 a18138a <=( (not A301)  and  (not A299) );
 a18139a <=( (not A298)  and  a18138a );
 a18140a <=( a18139a  and  a18134a );
 a18143a <=( A166  and  A168 );
 a18147a <=( (not A203)  and  (not A202) );
 a18148a <=( (not A201)  and  a18147a );
 a18149a <=( a18148a  and  a18143a );
 a18153a <=( A236  and  A233 );
 a18154a <=( (not A232)  and  a18153a );
 a18158a <=( A269  and  A266 );
 a18159a <=( (not A265)  and  a18158a );
 a18160a <=( a18159a  and  a18154a );
 a18163a <=( A166  and  A168 );
 a18167a <=( (not A203)  and  (not A202) );
 a18168a <=( (not A201)  and  a18167a );
 a18169a <=( a18168a  and  a18163a );
 a18173a <=( A236  and  A233 );
 a18174a <=( (not A232)  and  a18173a );
 a18178a <=( A269  and  (not A266) );
 a18179a <=( A265  and  a18178a );
 a18180a <=( a18179a  and  a18174a );
 a18183a <=( A166  and  A168 );
 a18187a <=( (not A203)  and  (not A202) );
 a18188a <=( (not A201)  and  a18187a );
 a18189a <=( a18188a  and  a18183a );
 a18193a <=( A236  and  (not A233) );
 a18194a <=( A232  and  a18193a );
 a18198a <=( (not A302)  and  (not A301) );
 a18199a <=( (not A300)  and  a18198a );
 a18200a <=( a18199a  and  a18194a );
 a18203a <=( A166  and  A168 );
 a18207a <=( (not A203)  and  (not A202) );
 a18208a <=( (not A201)  and  a18207a );
 a18209a <=( a18208a  and  a18203a );
 a18213a <=( A236  and  (not A233) );
 a18214a <=( A232  and  a18213a );
 a18218a <=( (not A301)  and  (not A299) );
 a18219a <=( (not A298)  and  a18218a );
 a18220a <=( a18219a  and  a18214a );
 a18223a <=( A166  and  A168 );
 a18227a <=( (not A203)  and  (not A202) );
 a18228a <=( (not A201)  and  a18227a );
 a18229a <=( a18228a  and  a18223a );
 a18233a <=( A236  and  (not A233) );
 a18234a <=( A232  and  a18233a );
 a18238a <=( A269  and  A266 );
 a18239a <=( (not A265)  and  a18238a );
 a18240a <=( a18239a  and  a18234a );
 a18243a <=( A166  and  A168 );
 a18247a <=( (not A203)  and  (not A202) );
 a18248a <=( (not A201)  and  a18247a );
 a18249a <=( a18248a  and  a18243a );
 a18253a <=( A236  and  (not A233) );
 a18254a <=( A232  and  a18253a );
 a18258a <=( A269  and  (not A266) );
 a18259a <=( A265  and  a18258a );
 a18260a <=( a18259a  and  a18254a );
 a18263a <=( A166  and  A168 );
 a18267a <=( (not A201)  and  A200 );
 a18268a <=( A199  and  a18267a );
 a18269a <=( a18268a  and  a18263a );
 a18273a <=( A298  and  A235 );
 a18274a <=( (not A202)  and  a18273a );
 a18278a <=( (not A301)  and  (not A300) );
 a18279a <=( A299  and  a18278a );
 a18280a <=( a18279a  and  a18274a );
 a18283a <=( A166  and  A168 );
 a18287a <=( (not A201)  and  A200 );
 a18288a <=( A199  and  a18287a );
 a18289a <=( a18288a  and  a18283a );
 a18293a <=( A234  and  A232 );
 a18294a <=( (not A202)  and  a18293a );
 a18298a <=( (not A302)  and  (not A301) );
 a18299a <=( (not A300)  and  a18298a );
 a18300a <=( a18299a  and  a18294a );
 a18303a <=( A166  and  A168 );
 a18307a <=( (not A201)  and  A200 );
 a18308a <=( A199  and  a18307a );
 a18309a <=( a18308a  and  a18303a );
 a18313a <=( A234  and  A232 );
 a18314a <=( (not A202)  and  a18313a );
 a18318a <=( (not A301)  and  (not A299) );
 a18319a <=( (not A298)  and  a18318a );
 a18320a <=( a18319a  and  a18314a );
 a18323a <=( A166  and  A168 );
 a18327a <=( (not A201)  and  A200 );
 a18328a <=( A199  and  a18327a );
 a18329a <=( a18328a  and  a18323a );
 a18333a <=( A234  and  A232 );
 a18334a <=( (not A202)  and  a18333a );
 a18338a <=( A269  and  A266 );
 a18339a <=( (not A265)  and  a18338a );
 a18340a <=( a18339a  and  a18334a );
 a18343a <=( A166  and  A168 );
 a18347a <=( (not A201)  and  A200 );
 a18348a <=( A199  and  a18347a );
 a18349a <=( a18348a  and  a18343a );
 a18353a <=( A234  and  A232 );
 a18354a <=( (not A202)  and  a18353a );
 a18358a <=( A269  and  (not A266) );
 a18359a <=( A265  and  a18358a );
 a18360a <=( a18359a  and  a18354a );
 a18363a <=( A166  and  A168 );
 a18367a <=( (not A201)  and  A200 );
 a18368a <=( A199  and  a18367a );
 a18369a <=( a18368a  and  a18363a );
 a18373a <=( A234  and  A233 );
 a18374a <=( (not A202)  and  a18373a );
 a18378a <=( (not A302)  and  (not A301) );
 a18379a <=( (not A300)  and  a18378a );
 a18380a <=( a18379a  and  a18374a );
 a18383a <=( A166  and  A168 );
 a18387a <=( (not A201)  and  A200 );
 a18388a <=( A199  and  a18387a );
 a18389a <=( a18388a  and  a18383a );
 a18393a <=( A234  and  A233 );
 a18394a <=( (not A202)  and  a18393a );
 a18398a <=( (not A301)  and  (not A299) );
 a18399a <=( (not A298)  and  a18398a );
 a18400a <=( a18399a  and  a18394a );
 a18403a <=( A166  and  A168 );
 a18407a <=( (not A201)  and  A200 );
 a18408a <=( A199  and  a18407a );
 a18409a <=( a18408a  and  a18403a );
 a18413a <=( A234  and  A233 );
 a18414a <=( (not A202)  and  a18413a );
 a18418a <=( A269  and  A266 );
 a18419a <=( (not A265)  and  a18418a );
 a18420a <=( a18419a  and  a18414a );
 a18423a <=( A166  and  A168 );
 a18427a <=( (not A201)  and  A200 );
 a18428a <=( A199  and  a18427a );
 a18429a <=( a18428a  and  a18423a );
 a18433a <=( A234  and  A233 );
 a18434a <=( (not A202)  and  a18433a );
 a18438a <=( A269  and  (not A266) );
 a18439a <=( A265  and  a18438a );
 a18440a <=( a18439a  and  a18434a );
 a18443a <=( A166  and  A168 );
 a18447a <=( (not A201)  and  A200 );
 a18448a <=( A199  and  a18447a );
 a18449a <=( a18448a  and  a18443a );
 a18453a <=( A233  and  (not A232) );
 a18454a <=( (not A202)  and  a18453a );
 a18458a <=( A267  and  A265 );
 a18459a <=( A236  and  a18458a );
 a18460a <=( a18459a  and  a18454a );
 a18463a <=( A166  and  A168 );
 a18467a <=( (not A201)  and  A200 );
 a18468a <=( A199  and  a18467a );
 a18469a <=( a18468a  and  a18463a );
 a18473a <=( A233  and  (not A232) );
 a18474a <=( (not A202)  and  a18473a );
 a18478a <=( A267  and  A266 );
 a18479a <=( A236  and  a18478a );
 a18480a <=( a18479a  and  a18474a );
 a18483a <=( A166  and  A168 );
 a18487a <=( (not A201)  and  A200 );
 a18488a <=( A199  and  a18487a );
 a18489a <=( a18488a  and  a18483a );
 a18493a <=( (not A233)  and  A232 );
 a18494a <=( (not A202)  and  a18493a );
 a18498a <=( A267  and  A265 );
 a18499a <=( A236  and  a18498a );
 a18500a <=( a18499a  and  a18494a );
 a18503a <=( A166  and  A168 );
 a18507a <=( (not A201)  and  A200 );
 a18508a <=( A199  and  a18507a );
 a18509a <=( a18508a  and  a18503a );
 a18513a <=( (not A233)  and  A232 );
 a18514a <=( (not A202)  and  a18513a );
 a18518a <=( A267  and  A266 );
 a18519a <=( A236  and  a18518a );
 a18520a <=( a18519a  and  a18514a );
 a18523a <=( A166  and  A168 );
 a18527a <=( (not A202)  and  (not A200) );
 a18528a <=( (not A199)  and  a18527a );
 a18529a <=( a18528a  and  a18523a );
 a18533a <=( A298  and  A234 );
 a18534a <=( A232  and  a18533a );
 a18538a <=( (not A301)  and  (not A300) );
 a18539a <=( A299  and  a18538a );
 a18540a <=( a18539a  and  a18534a );
 a18543a <=( A166  and  A168 );
 a18547a <=( (not A202)  and  (not A200) );
 a18548a <=( (not A199)  and  a18547a );
 a18549a <=( a18548a  and  a18543a );
 a18553a <=( A298  and  A234 );
 a18554a <=( A233  and  a18553a );
 a18558a <=( (not A301)  and  (not A300) );
 a18559a <=( A299  and  a18558a );
 a18560a <=( a18559a  and  a18554a );
 a18563a <=( A166  and  A168 );
 a18567a <=( (not A202)  and  (not A200) );
 a18568a <=( (not A199)  and  a18567a );
 a18569a <=( a18568a  and  a18563a );
 a18573a <=( A236  and  A233 );
 a18574a <=( (not A232)  and  a18573a );
 a18578a <=( (not A302)  and  (not A301) );
 a18579a <=( (not A300)  and  a18578a );
 a18580a <=( a18579a  and  a18574a );
 a18583a <=( A166  and  A168 );
 a18587a <=( (not A202)  and  (not A200) );
 a18588a <=( (not A199)  and  a18587a );
 a18589a <=( a18588a  and  a18583a );
 a18593a <=( A236  and  A233 );
 a18594a <=( (not A232)  and  a18593a );
 a18598a <=( (not A301)  and  (not A299) );
 a18599a <=( (not A298)  and  a18598a );
 a18600a <=( a18599a  and  a18594a );
 a18603a <=( A166  and  A168 );
 a18607a <=( (not A202)  and  (not A200) );
 a18608a <=( (not A199)  and  a18607a );
 a18609a <=( a18608a  and  a18603a );
 a18613a <=( A236  and  A233 );
 a18614a <=( (not A232)  and  a18613a );
 a18618a <=( A269  and  A266 );
 a18619a <=( (not A265)  and  a18618a );
 a18620a <=( a18619a  and  a18614a );
 a18623a <=( A166  and  A168 );
 a18627a <=( (not A202)  and  (not A200) );
 a18628a <=( (not A199)  and  a18627a );
 a18629a <=( a18628a  and  a18623a );
 a18633a <=( A236  and  A233 );
 a18634a <=( (not A232)  and  a18633a );
 a18638a <=( A269  and  (not A266) );
 a18639a <=( A265  and  a18638a );
 a18640a <=( a18639a  and  a18634a );
 a18643a <=( A166  and  A168 );
 a18647a <=( (not A202)  and  (not A200) );
 a18648a <=( (not A199)  and  a18647a );
 a18649a <=( a18648a  and  a18643a );
 a18653a <=( A236  and  (not A233) );
 a18654a <=( A232  and  a18653a );
 a18658a <=( (not A302)  and  (not A301) );
 a18659a <=( (not A300)  and  a18658a );
 a18660a <=( a18659a  and  a18654a );
 a18663a <=( A166  and  A168 );
 a18667a <=( (not A202)  and  (not A200) );
 a18668a <=( (not A199)  and  a18667a );
 a18669a <=( a18668a  and  a18663a );
 a18673a <=( A236  and  (not A233) );
 a18674a <=( A232  and  a18673a );
 a18678a <=( (not A301)  and  (not A299) );
 a18679a <=( (not A298)  and  a18678a );
 a18680a <=( a18679a  and  a18674a );
 a18683a <=( A166  and  A168 );
 a18687a <=( (not A202)  and  (not A200) );
 a18688a <=( (not A199)  and  a18687a );
 a18689a <=( a18688a  and  a18683a );
 a18693a <=( A236  and  (not A233) );
 a18694a <=( A232  and  a18693a );
 a18698a <=( A269  and  A266 );
 a18699a <=( (not A265)  and  a18698a );
 a18700a <=( a18699a  and  a18694a );
 a18703a <=( A166  and  A168 );
 a18707a <=( (not A202)  and  (not A200) );
 a18708a <=( (not A199)  and  a18707a );
 a18709a <=( a18708a  and  a18703a );
 a18713a <=( A236  and  (not A233) );
 a18714a <=( A232  and  a18713a );
 a18718a <=( A269  and  (not A266) );
 a18719a <=( A265  and  a18718a );
 a18720a <=( a18719a  and  a18714a );
 a18723a <=( A167  and  A168 );
 a18727a <=( (not A203)  and  (not A202) );
 a18728a <=( (not A201)  and  a18727a );
 a18729a <=( a18728a  and  a18723a );
 a18733a <=( A298  and  A234 );
 a18734a <=( A232  and  a18733a );
 a18738a <=( (not A301)  and  (not A300) );
 a18739a <=( A299  and  a18738a );
 a18740a <=( a18739a  and  a18734a );
 a18743a <=( A167  and  A168 );
 a18747a <=( (not A203)  and  (not A202) );
 a18748a <=( (not A201)  and  a18747a );
 a18749a <=( a18748a  and  a18743a );
 a18753a <=( A298  and  A234 );
 a18754a <=( A233  and  a18753a );
 a18758a <=( (not A301)  and  (not A300) );
 a18759a <=( A299  and  a18758a );
 a18760a <=( a18759a  and  a18754a );
 a18763a <=( A167  and  A168 );
 a18767a <=( (not A203)  and  (not A202) );
 a18768a <=( (not A201)  and  a18767a );
 a18769a <=( a18768a  and  a18763a );
 a18773a <=( A236  and  A233 );
 a18774a <=( (not A232)  and  a18773a );
 a18778a <=( (not A302)  and  (not A301) );
 a18779a <=( (not A300)  and  a18778a );
 a18780a <=( a18779a  and  a18774a );
 a18783a <=( A167  and  A168 );
 a18787a <=( (not A203)  and  (not A202) );
 a18788a <=( (not A201)  and  a18787a );
 a18789a <=( a18788a  and  a18783a );
 a18793a <=( A236  and  A233 );
 a18794a <=( (not A232)  and  a18793a );
 a18798a <=( (not A301)  and  (not A299) );
 a18799a <=( (not A298)  and  a18798a );
 a18800a <=( a18799a  and  a18794a );
 a18803a <=( A167  and  A168 );
 a18807a <=( (not A203)  and  (not A202) );
 a18808a <=( (not A201)  and  a18807a );
 a18809a <=( a18808a  and  a18803a );
 a18813a <=( A236  and  A233 );
 a18814a <=( (not A232)  and  a18813a );
 a18818a <=( A269  and  A266 );
 a18819a <=( (not A265)  and  a18818a );
 a18820a <=( a18819a  and  a18814a );
 a18823a <=( A167  and  A168 );
 a18827a <=( (not A203)  and  (not A202) );
 a18828a <=( (not A201)  and  a18827a );
 a18829a <=( a18828a  and  a18823a );
 a18833a <=( A236  and  A233 );
 a18834a <=( (not A232)  and  a18833a );
 a18838a <=( A269  and  (not A266) );
 a18839a <=( A265  and  a18838a );
 a18840a <=( a18839a  and  a18834a );
 a18843a <=( A167  and  A168 );
 a18847a <=( (not A203)  and  (not A202) );
 a18848a <=( (not A201)  and  a18847a );
 a18849a <=( a18848a  and  a18843a );
 a18853a <=( A236  and  (not A233) );
 a18854a <=( A232  and  a18853a );
 a18858a <=( (not A302)  and  (not A301) );
 a18859a <=( (not A300)  and  a18858a );
 a18860a <=( a18859a  and  a18854a );
 a18863a <=( A167  and  A168 );
 a18867a <=( (not A203)  and  (not A202) );
 a18868a <=( (not A201)  and  a18867a );
 a18869a <=( a18868a  and  a18863a );
 a18873a <=( A236  and  (not A233) );
 a18874a <=( A232  and  a18873a );
 a18878a <=( (not A301)  and  (not A299) );
 a18879a <=( (not A298)  and  a18878a );
 a18880a <=( a18879a  and  a18874a );
 a18883a <=( A167  and  A168 );
 a18887a <=( (not A203)  and  (not A202) );
 a18888a <=( (not A201)  and  a18887a );
 a18889a <=( a18888a  and  a18883a );
 a18893a <=( A236  and  (not A233) );
 a18894a <=( A232  and  a18893a );
 a18898a <=( A269  and  A266 );
 a18899a <=( (not A265)  and  a18898a );
 a18900a <=( a18899a  and  a18894a );
 a18903a <=( A167  and  A168 );
 a18907a <=( (not A203)  and  (not A202) );
 a18908a <=( (not A201)  and  a18907a );
 a18909a <=( a18908a  and  a18903a );
 a18913a <=( A236  and  (not A233) );
 a18914a <=( A232  and  a18913a );
 a18918a <=( A269  and  (not A266) );
 a18919a <=( A265  and  a18918a );
 a18920a <=( a18919a  and  a18914a );
 a18923a <=( A167  and  A168 );
 a18927a <=( (not A201)  and  A200 );
 a18928a <=( A199  and  a18927a );
 a18929a <=( a18928a  and  a18923a );
 a18933a <=( A298  and  A235 );
 a18934a <=( (not A202)  and  a18933a );
 a18938a <=( (not A301)  and  (not A300) );
 a18939a <=( A299  and  a18938a );
 a18940a <=( a18939a  and  a18934a );
 a18943a <=( A167  and  A168 );
 a18947a <=( (not A201)  and  A200 );
 a18948a <=( A199  and  a18947a );
 a18949a <=( a18948a  and  a18943a );
 a18953a <=( A234  and  A232 );
 a18954a <=( (not A202)  and  a18953a );
 a18958a <=( (not A302)  and  (not A301) );
 a18959a <=( (not A300)  and  a18958a );
 a18960a <=( a18959a  and  a18954a );
 a18963a <=( A167  and  A168 );
 a18967a <=( (not A201)  and  A200 );
 a18968a <=( A199  and  a18967a );
 a18969a <=( a18968a  and  a18963a );
 a18973a <=( A234  and  A232 );
 a18974a <=( (not A202)  and  a18973a );
 a18978a <=( (not A301)  and  (not A299) );
 a18979a <=( (not A298)  and  a18978a );
 a18980a <=( a18979a  and  a18974a );
 a18983a <=( A167  and  A168 );
 a18987a <=( (not A201)  and  A200 );
 a18988a <=( A199  and  a18987a );
 a18989a <=( a18988a  and  a18983a );
 a18993a <=( A234  and  A232 );
 a18994a <=( (not A202)  and  a18993a );
 a18998a <=( A269  and  A266 );
 a18999a <=( (not A265)  and  a18998a );
 a19000a <=( a18999a  and  a18994a );
 a19003a <=( A167  and  A168 );
 a19007a <=( (not A201)  and  A200 );
 a19008a <=( A199  and  a19007a );
 a19009a <=( a19008a  and  a19003a );
 a19013a <=( A234  and  A232 );
 a19014a <=( (not A202)  and  a19013a );
 a19018a <=( A269  and  (not A266) );
 a19019a <=( A265  and  a19018a );
 a19020a <=( a19019a  and  a19014a );
 a19023a <=( A167  and  A168 );
 a19027a <=( (not A201)  and  A200 );
 a19028a <=( A199  and  a19027a );
 a19029a <=( a19028a  and  a19023a );
 a19033a <=( A234  and  A233 );
 a19034a <=( (not A202)  and  a19033a );
 a19038a <=( (not A302)  and  (not A301) );
 a19039a <=( (not A300)  and  a19038a );
 a19040a <=( a19039a  and  a19034a );
 a19043a <=( A167  and  A168 );
 a19047a <=( (not A201)  and  A200 );
 a19048a <=( A199  and  a19047a );
 a19049a <=( a19048a  and  a19043a );
 a19053a <=( A234  and  A233 );
 a19054a <=( (not A202)  and  a19053a );
 a19058a <=( (not A301)  and  (not A299) );
 a19059a <=( (not A298)  and  a19058a );
 a19060a <=( a19059a  and  a19054a );
 a19063a <=( A167  and  A168 );
 a19067a <=( (not A201)  and  A200 );
 a19068a <=( A199  and  a19067a );
 a19069a <=( a19068a  and  a19063a );
 a19073a <=( A234  and  A233 );
 a19074a <=( (not A202)  and  a19073a );
 a19078a <=( A269  and  A266 );
 a19079a <=( (not A265)  and  a19078a );
 a19080a <=( a19079a  and  a19074a );
 a19083a <=( A167  and  A168 );
 a19087a <=( (not A201)  and  A200 );
 a19088a <=( A199  and  a19087a );
 a19089a <=( a19088a  and  a19083a );
 a19093a <=( A234  and  A233 );
 a19094a <=( (not A202)  and  a19093a );
 a19098a <=( A269  and  (not A266) );
 a19099a <=( A265  and  a19098a );
 a19100a <=( a19099a  and  a19094a );
 a19103a <=( A167  and  A168 );
 a19107a <=( (not A201)  and  A200 );
 a19108a <=( A199  and  a19107a );
 a19109a <=( a19108a  and  a19103a );
 a19113a <=( A233  and  (not A232) );
 a19114a <=( (not A202)  and  a19113a );
 a19118a <=( A267  and  A265 );
 a19119a <=( A236  and  a19118a );
 a19120a <=( a19119a  and  a19114a );
 a19123a <=( A167  and  A168 );
 a19127a <=( (not A201)  and  A200 );
 a19128a <=( A199  and  a19127a );
 a19129a <=( a19128a  and  a19123a );
 a19133a <=( A233  and  (not A232) );
 a19134a <=( (not A202)  and  a19133a );
 a19138a <=( A267  and  A266 );
 a19139a <=( A236  and  a19138a );
 a19140a <=( a19139a  and  a19134a );
 a19143a <=( A167  and  A168 );
 a19147a <=( (not A201)  and  A200 );
 a19148a <=( A199  and  a19147a );
 a19149a <=( a19148a  and  a19143a );
 a19153a <=( (not A233)  and  A232 );
 a19154a <=( (not A202)  and  a19153a );
 a19158a <=( A267  and  A265 );
 a19159a <=( A236  and  a19158a );
 a19160a <=( a19159a  and  a19154a );
 a19163a <=( A167  and  A168 );
 a19167a <=( (not A201)  and  A200 );
 a19168a <=( A199  and  a19167a );
 a19169a <=( a19168a  and  a19163a );
 a19173a <=( (not A233)  and  A232 );
 a19174a <=( (not A202)  and  a19173a );
 a19178a <=( A267  and  A266 );
 a19179a <=( A236  and  a19178a );
 a19180a <=( a19179a  and  a19174a );
 a19183a <=( A167  and  A168 );
 a19187a <=( (not A202)  and  (not A200) );
 a19188a <=( (not A199)  and  a19187a );
 a19189a <=( a19188a  and  a19183a );
 a19193a <=( A298  and  A234 );
 a19194a <=( A232  and  a19193a );
 a19198a <=( (not A301)  and  (not A300) );
 a19199a <=( A299  and  a19198a );
 a19200a <=( a19199a  and  a19194a );
 a19203a <=( A167  and  A168 );
 a19207a <=( (not A202)  and  (not A200) );
 a19208a <=( (not A199)  and  a19207a );
 a19209a <=( a19208a  and  a19203a );
 a19213a <=( A298  and  A234 );
 a19214a <=( A233  and  a19213a );
 a19218a <=( (not A301)  and  (not A300) );
 a19219a <=( A299  and  a19218a );
 a19220a <=( a19219a  and  a19214a );
 a19223a <=( A167  and  A168 );
 a19227a <=( (not A202)  and  (not A200) );
 a19228a <=( (not A199)  and  a19227a );
 a19229a <=( a19228a  and  a19223a );
 a19233a <=( A236  and  A233 );
 a19234a <=( (not A232)  and  a19233a );
 a19238a <=( (not A302)  and  (not A301) );
 a19239a <=( (not A300)  and  a19238a );
 a19240a <=( a19239a  and  a19234a );
 a19243a <=( A167  and  A168 );
 a19247a <=( (not A202)  and  (not A200) );
 a19248a <=( (not A199)  and  a19247a );
 a19249a <=( a19248a  and  a19243a );
 a19253a <=( A236  and  A233 );
 a19254a <=( (not A232)  and  a19253a );
 a19258a <=( (not A301)  and  (not A299) );
 a19259a <=( (not A298)  and  a19258a );
 a19260a <=( a19259a  and  a19254a );
 a19263a <=( A167  and  A168 );
 a19267a <=( (not A202)  and  (not A200) );
 a19268a <=( (not A199)  and  a19267a );
 a19269a <=( a19268a  and  a19263a );
 a19273a <=( A236  and  A233 );
 a19274a <=( (not A232)  and  a19273a );
 a19278a <=( A269  and  A266 );
 a19279a <=( (not A265)  and  a19278a );
 a19280a <=( a19279a  and  a19274a );
 a19283a <=( A167  and  A168 );
 a19287a <=( (not A202)  and  (not A200) );
 a19288a <=( (not A199)  and  a19287a );
 a19289a <=( a19288a  and  a19283a );
 a19293a <=( A236  and  A233 );
 a19294a <=( (not A232)  and  a19293a );
 a19298a <=( A269  and  (not A266) );
 a19299a <=( A265  and  a19298a );
 a19300a <=( a19299a  and  a19294a );
 a19303a <=( A167  and  A168 );
 a19307a <=( (not A202)  and  (not A200) );
 a19308a <=( (not A199)  and  a19307a );
 a19309a <=( a19308a  and  a19303a );
 a19313a <=( A236  and  (not A233) );
 a19314a <=( A232  and  a19313a );
 a19318a <=( (not A302)  and  (not A301) );
 a19319a <=( (not A300)  and  a19318a );
 a19320a <=( a19319a  and  a19314a );
 a19323a <=( A167  and  A168 );
 a19327a <=( (not A202)  and  (not A200) );
 a19328a <=( (not A199)  and  a19327a );
 a19329a <=( a19328a  and  a19323a );
 a19333a <=( A236  and  (not A233) );
 a19334a <=( A232  and  a19333a );
 a19338a <=( (not A301)  and  (not A299) );
 a19339a <=( (not A298)  and  a19338a );
 a19340a <=( a19339a  and  a19334a );
 a19343a <=( A167  and  A168 );
 a19347a <=( (not A202)  and  (not A200) );
 a19348a <=( (not A199)  and  a19347a );
 a19349a <=( a19348a  and  a19343a );
 a19353a <=( A236  and  (not A233) );
 a19354a <=( A232  and  a19353a );
 a19358a <=( A269  and  A266 );
 a19359a <=( (not A265)  and  a19358a );
 a19360a <=( a19359a  and  a19354a );
 a19363a <=( A167  and  A168 );
 a19367a <=( (not A202)  and  (not A200) );
 a19368a <=( (not A199)  and  a19367a );
 a19369a <=( a19368a  and  a19363a );
 a19373a <=( A236  and  (not A233) );
 a19374a <=( A232  and  a19373a );
 a19378a <=( A269  and  (not A266) );
 a19379a <=( A265  and  a19378a );
 a19380a <=( a19379a  and  a19374a );
 a19383a <=( A167  and  A170 );
 a19387a <=( (not A202)  and  (not A201) );
 a19388a <=( (not A166)  and  a19387a );
 a19389a <=( a19388a  and  a19383a );
 a19393a <=( A298  and  A235 );
 a19394a <=( (not A203)  and  a19393a );
 a19398a <=( (not A301)  and  (not A300) );
 a19399a <=( A299  and  a19398a );
 a19400a <=( a19399a  and  a19394a );
 a19403a <=( A167  and  A170 );
 a19407a <=( (not A202)  and  (not A201) );
 a19408a <=( (not A166)  and  a19407a );
 a19409a <=( a19408a  and  a19403a );
 a19413a <=( A234  and  A232 );
 a19414a <=( (not A203)  and  a19413a );
 a19418a <=( (not A302)  and  (not A301) );
 a19419a <=( (not A300)  and  a19418a );
 a19420a <=( a19419a  and  a19414a );
 a19423a <=( A167  and  A170 );
 a19427a <=( (not A202)  and  (not A201) );
 a19428a <=( (not A166)  and  a19427a );
 a19429a <=( a19428a  and  a19423a );
 a19433a <=( A234  and  A232 );
 a19434a <=( (not A203)  and  a19433a );
 a19438a <=( (not A301)  and  (not A299) );
 a19439a <=( (not A298)  and  a19438a );
 a19440a <=( a19439a  and  a19434a );
 a19443a <=( A167  and  A170 );
 a19447a <=( (not A202)  and  (not A201) );
 a19448a <=( (not A166)  and  a19447a );
 a19449a <=( a19448a  and  a19443a );
 a19453a <=( A234  and  A232 );
 a19454a <=( (not A203)  and  a19453a );
 a19458a <=( A269  and  A266 );
 a19459a <=( (not A265)  and  a19458a );
 a19460a <=( a19459a  and  a19454a );
 a19463a <=( A167  and  A170 );
 a19467a <=( (not A202)  and  (not A201) );
 a19468a <=( (not A166)  and  a19467a );
 a19469a <=( a19468a  and  a19463a );
 a19473a <=( A234  and  A232 );
 a19474a <=( (not A203)  and  a19473a );
 a19478a <=( A269  and  (not A266) );
 a19479a <=( A265  and  a19478a );
 a19480a <=( a19479a  and  a19474a );
 a19483a <=( A167  and  A170 );
 a19487a <=( (not A202)  and  (not A201) );
 a19488a <=( (not A166)  and  a19487a );
 a19489a <=( a19488a  and  a19483a );
 a19493a <=( A234  and  A233 );
 a19494a <=( (not A203)  and  a19493a );
 a19498a <=( (not A302)  and  (not A301) );
 a19499a <=( (not A300)  and  a19498a );
 a19500a <=( a19499a  and  a19494a );
 a19503a <=( A167  and  A170 );
 a19507a <=( (not A202)  and  (not A201) );
 a19508a <=( (not A166)  and  a19507a );
 a19509a <=( a19508a  and  a19503a );
 a19513a <=( A234  and  A233 );
 a19514a <=( (not A203)  and  a19513a );
 a19518a <=( (not A301)  and  (not A299) );
 a19519a <=( (not A298)  and  a19518a );
 a19520a <=( a19519a  and  a19514a );
 a19523a <=( A167  and  A170 );
 a19527a <=( (not A202)  and  (not A201) );
 a19528a <=( (not A166)  and  a19527a );
 a19529a <=( a19528a  and  a19523a );
 a19533a <=( A234  and  A233 );
 a19534a <=( (not A203)  and  a19533a );
 a19538a <=( A269  and  A266 );
 a19539a <=( (not A265)  and  a19538a );
 a19540a <=( a19539a  and  a19534a );
 a19543a <=( A167  and  A170 );
 a19547a <=( (not A202)  and  (not A201) );
 a19548a <=( (not A166)  and  a19547a );
 a19549a <=( a19548a  and  a19543a );
 a19553a <=( A234  and  A233 );
 a19554a <=( (not A203)  and  a19553a );
 a19558a <=( A269  and  (not A266) );
 a19559a <=( A265  and  a19558a );
 a19560a <=( a19559a  and  a19554a );
 a19563a <=( A167  and  A170 );
 a19567a <=( (not A202)  and  (not A201) );
 a19568a <=( (not A166)  and  a19567a );
 a19569a <=( a19568a  and  a19563a );
 a19573a <=( A233  and  (not A232) );
 a19574a <=( (not A203)  and  a19573a );
 a19578a <=( A267  and  A265 );
 a19579a <=( A236  and  a19578a );
 a19580a <=( a19579a  and  a19574a );
 a19583a <=( A167  and  A170 );
 a19587a <=( (not A202)  and  (not A201) );
 a19588a <=( (not A166)  and  a19587a );
 a19589a <=( a19588a  and  a19583a );
 a19593a <=( A233  and  (not A232) );
 a19594a <=( (not A203)  and  a19593a );
 a19598a <=( A267  and  A266 );
 a19599a <=( A236  and  a19598a );
 a19600a <=( a19599a  and  a19594a );
 a19603a <=( A167  and  A170 );
 a19607a <=( (not A202)  and  (not A201) );
 a19608a <=( (not A166)  and  a19607a );
 a19609a <=( a19608a  and  a19603a );
 a19613a <=( (not A233)  and  A232 );
 a19614a <=( (not A203)  and  a19613a );
 a19618a <=( A267  and  A265 );
 a19619a <=( A236  and  a19618a );
 a19620a <=( a19619a  and  a19614a );
 a19623a <=( A167  and  A170 );
 a19627a <=( (not A202)  and  (not A201) );
 a19628a <=( (not A166)  and  a19627a );
 a19629a <=( a19628a  and  a19623a );
 a19633a <=( (not A233)  and  A232 );
 a19634a <=( (not A203)  and  a19633a );
 a19638a <=( A267  and  A266 );
 a19639a <=( A236  and  a19638a );
 a19640a <=( a19639a  and  a19634a );
 a19643a <=( A167  and  A170 );
 a19647a <=( A200  and  A199 );
 a19648a <=( (not A166)  and  a19647a );
 a19649a <=( a19648a  and  a19643a );
 a19653a <=( A235  and  (not A202) );
 a19654a <=( (not A201)  and  a19653a );
 a19658a <=( (not A302)  and  (not A301) );
 a19659a <=( (not A300)  and  a19658a );
 a19660a <=( a19659a  and  a19654a );
 a19663a <=( A167  and  A170 );
 a19667a <=( A200  and  A199 );
 a19668a <=( (not A166)  and  a19667a );
 a19669a <=( a19668a  and  a19663a );
 a19673a <=( A235  and  (not A202) );
 a19674a <=( (not A201)  and  a19673a );
 a19678a <=( (not A301)  and  (not A299) );
 a19679a <=( (not A298)  and  a19678a );
 a19680a <=( a19679a  and  a19674a );
 a19683a <=( A167  and  A170 );
 a19687a <=( A200  and  A199 );
 a19688a <=( (not A166)  and  a19687a );
 a19689a <=( a19688a  and  a19683a );
 a19693a <=( A235  and  (not A202) );
 a19694a <=( (not A201)  and  a19693a );
 a19698a <=( A269  and  A266 );
 a19699a <=( (not A265)  and  a19698a );
 a19700a <=( a19699a  and  a19694a );
 a19703a <=( A167  and  A170 );
 a19707a <=( A200  and  A199 );
 a19708a <=( (not A166)  and  a19707a );
 a19709a <=( a19708a  and  a19703a );
 a19713a <=( A235  and  (not A202) );
 a19714a <=( (not A201)  and  a19713a );
 a19718a <=( A269  and  (not A266) );
 a19719a <=( A265  and  a19718a );
 a19720a <=( a19719a  and  a19714a );
 a19723a <=( A167  and  A170 );
 a19727a <=( A200  and  A199 );
 a19728a <=( (not A166)  and  a19727a );
 a19729a <=( a19728a  and  a19723a );
 a19733a <=( A232  and  (not A202) );
 a19734a <=( (not A201)  and  a19733a );
 a19738a <=( A267  and  A265 );
 a19739a <=( A234  and  a19738a );
 a19740a <=( a19739a  and  a19734a );
 a19743a <=( A167  and  A170 );
 a19747a <=( A200  and  A199 );
 a19748a <=( (not A166)  and  a19747a );
 a19749a <=( a19748a  and  a19743a );
 a19753a <=( A232  and  (not A202) );
 a19754a <=( (not A201)  and  a19753a );
 a19758a <=( A267  and  A266 );
 a19759a <=( A234  and  a19758a );
 a19760a <=( a19759a  and  a19754a );
 a19763a <=( A167  and  A170 );
 a19767a <=( A200  and  A199 );
 a19768a <=( (not A166)  and  a19767a );
 a19769a <=( a19768a  and  a19763a );
 a19773a <=( A233  and  (not A202) );
 a19774a <=( (not A201)  and  a19773a );
 a19778a <=( A267  and  A265 );
 a19779a <=( A234  and  a19778a );
 a19780a <=( a19779a  and  a19774a );
 a19783a <=( A167  and  A170 );
 a19787a <=( A200  and  A199 );
 a19788a <=( (not A166)  and  a19787a );
 a19789a <=( a19788a  and  a19783a );
 a19793a <=( A233  and  (not A202) );
 a19794a <=( (not A201)  and  a19793a );
 a19798a <=( A267  and  A266 );
 a19799a <=( A234  and  a19798a );
 a19800a <=( a19799a  and  a19794a );
 a19803a <=( A167  and  A170 );
 a19807a <=( A200  and  A199 );
 a19808a <=( (not A166)  and  a19807a );
 a19809a <=( a19808a  and  a19803a );
 a19813a <=( (not A232)  and  (not A202) );
 a19814a <=( (not A201)  and  a19813a );
 a19818a <=( A268  and  A236 );
 a19819a <=( A233  and  a19818a );
 a19820a <=( a19819a  and  a19814a );
 a19823a <=( A167  and  A170 );
 a19827a <=( A200  and  A199 );
 a19828a <=( (not A166)  and  a19827a );
 a19829a <=( a19828a  and  a19823a );
 a19833a <=( A232  and  (not A202) );
 a19834a <=( (not A201)  and  a19833a );
 a19838a <=( A268  and  A236 );
 a19839a <=( (not A233)  and  a19838a );
 a19840a <=( a19839a  and  a19834a );
 a19843a <=( A167  and  A170 );
 a19847a <=( (not A200)  and  (not A199) );
 a19848a <=( (not A166)  and  a19847a );
 a19849a <=( a19848a  and  a19843a );
 a19853a <=( A298  and  A235 );
 a19854a <=( (not A202)  and  a19853a );
 a19858a <=( (not A301)  and  (not A300) );
 a19859a <=( A299  and  a19858a );
 a19860a <=( a19859a  and  a19854a );
 a19863a <=( A167  and  A170 );
 a19867a <=( (not A200)  and  (not A199) );
 a19868a <=( (not A166)  and  a19867a );
 a19869a <=( a19868a  and  a19863a );
 a19873a <=( A234  and  A232 );
 a19874a <=( (not A202)  and  a19873a );
 a19878a <=( (not A302)  and  (not A301) );
 a19879a <=( (not A300)  and  a19878a );
 a19880a <=( a19879a  and  a19874a );
 a19883a <=( A167  and  A170 );
 a19887a <=( (not A200)  and  (not A199) );
 a19888a <=( (not A166)  and  a19887a );
 a19889a <=( a19888a  and  a19883a );
 a19893a <=( A234  and  A232 );
 a19894a <=( (not A202)  and  a19893a );
 a19898a <=( (not A301)  and  (not A299) );
 a19899a <=( (not A298)  and  a19898a );
 a19900a <=( a19899a  and  a19894a );
 a19903a <=( A167  and  A170 );
 a19907a <=( (not A200)  and  (not A199) );
 a19908a <=( (not A166)  and  a19907a );
 a19909a <=( a19908a  and  a19903a );
 a19913a <=( A234  and  A232 );
 a19914a <=( (not A202)  and  a19913a );
 a19918a <=( A269  and  A266 );
 a19919a <=( (not A265)  and  a19918a );
 a19920a <=( a19919a  and  a19914a );
 a19923a <=( A167  and  A170 );
 a19927a <=( (not A200)  and  (not A199) );
 a19928a <=( (not A166)  and  a19927a );
 a19929a <=( a19928a  and  a19923a );
 a19933a <=( A234  and  A232 );
 a19934a <=( (not A202)  and  a19933a );
 a19938a <=( A269  and  (not A266) );
 a19939a <=( A265  and  a19938a );
 a19940a <=( a19939a  and  a19934a );
 a19943a <=( A167  and  A170 );
 a19947a <=( (not A200)  and  (not A199) );
 a19948a <=( (not A166)  and  a19947a );
 a19949a <=( a19948a  and  a19943a );
 a19953a <=( A234  and  A233 );
 a19954a <=( (not A202)  and  a19953a );
 a19958a <=( (not A302)  and  (not A301) );
 a19959a <=( (not A300)  and  a19958a );
 a19960a <=( a19959a  and  a19954a );
 a19963a <=( A167  and  A170 );
 a19967a <=( (not A200)  and  (not A199) );
 a19968a <=( (not A166)  and  a19967a );
 a19969a <=( a19968a  and  a19963a );
 a19973a <=( A234  and  A233 );
 a19974a <=( (not A202)  and  a19973a );
 a19978a <=( (not A301)  and  (not A299) );
 a19979a <=( (not A298)  and  a19978a );
 a19980a <=( a19979a  and  a19974a );
 a19983a <=( A167  and  A170 );
 a19987a <=( (not A200)  and  (not A199) );
 a19988a <=( (not A166)  and  a19987a );
 a19989a <=( a19988a  and  a19983a );
 a19993a <=( A234  and  A233 );
 a19994a <=( (not A202)  and  a19993a );
 a19998a <=( A269  and  A266 );
 a19999a <=( (not A265)  and  a19998a );
 a20000a <=( a19999a  and  a19994a );
 a20003a <=( A167  and  A170 );
 a20007a <=( (not A200)  and  (not A199) );
 a20008a <=( (not A166)  and  a20007a );
 a20009a <=( a20008a  and  a20003a );
 a20013a <=( A234  and  A233 );
 a20014a <=( (not A202)  and  a20013a );
 a20018a <=( A269  and  (not A266) );
 a20019a <=( A265  and  a20018a );
 a20020a <=( a20019a  and  a20014a );
 a20023a <=( A167  and  A170 );
 a20027a <=( (not A200)  and  (not A199) );
 a20028a <=( (not A166)  and  a20027a );
 a20029a <=( a20028a  and  a20023a );
 a20033a <=( A233  and  (not A232) );
 a20034a <=( (not A202)  and  a20033a );
 a20038a <=( A267  and  A265 );
 a20039a <=( A236  and  a20038a );
 a20040a <=( a20039a  and  a20034a );
 a20043a <=( A167  and  A170 );
 a20047a <=( (not A200)  and  (not A199) );
 a20048a <=( (not A166)  and  a20047a );
 a20049a <=( a20048a  and  a20043a );
 a20053a <=( A233  and  (not A232) );
 a20054a <=( (not A202)  and  a20053a );
 a20058a <=( A267  and  A266 );
 a20059a <=( A236  and  a20058a );
 a20060a <=( a20059a  and  a20054a );
 a20063a <=( A167  and  A170 );
 a20067a <=( (not A200)  and  (not A199) );
 a20068a <=( (not A166)  and  a20067a );
 a20069a <=( a20068a  and  a20063a );
 a20073a <=( (not A233)  and  A232 );
 a20074a <=( (not A202)  and  a20073a );
 a20078a <=( A267  and  A265 );
 a20079a <=( A236  and  a20078a );
 a20080a <=( a20079a  and  a20074a );
 a20083a <=( A167  and  A170 );
 a20087a <=( (not A200)  and  (not A199) );
 a20088a <=( (not A166)  and  a20087a );
 a20089a <=( a20088a  and  a20083a );
 a20093a <=( (not A233)  and  A232 );
 a20094a <=( (not A202)  and  a20093a );
 a20098a <=( A267  and  A266 );
 a20099a <=( A236  and  a20098a );
 a20100a <=( a20099a  and  a20094a );
 a20103a <=( (not A167)  and  A170 );
 a20107a <=( (not A202)  and  (not A201) );
 a20108a <=( A166  and  a20107a );
 a20109a <=( a20108a  and  a20103a );
 a20113a <=( A298  and  A235 );
 a20114a <=( (not A203)  and  a20113a );
 a20118a <=( (not A301)  and  (not A300) );
 a20119a <=( A299  and  a20118a );
 a20120a <=( a20119a  and  a20114a );
 a20123a <=( (not A167)  and  A170 );
 a20127a <=( (not A202)  and  (not A201) );
 a20128a <=( A166  and  a20127a );
 a20129a <=( a20128a  and  a20123a );
 a20133a <=( A234  and  A232 );
 a20134a <=( (not A203)  and  a20133a );
 a20138a <=( (not A302)  and  (not A301) );
 a20139a <=( (not A300)  and  a20138a );
 a20140a <=( a20139a  and  a20134a );
 a20143a <=( (not A167)  and  A170 );
 a20147a <=( (not A202)  and  (not A201) );
 a20148a <=( A166  and  a20147a );
 a20149a <=( a20148a  and  a20143a );
 a20153a <=( A234  and  A232 );
 a20154a <=( (not A203)  and  a20153a );
 a20158a <=( (not A301)  and  (not A299) );
 a20159a <=( (not A298)  and  a20158a );
 a20160a <=( a20159a  and  a20154a );
 a20163a <=( (not A167)  and  A170 );
 a20167a <=( (not A202)  and  (not A201) );
 a20168a <=( A166  and  a20167a );
 a20169a <=( a20168a  and  a20163a );
 a20173a <=( A234  and  A232 );
 a20174a <=( (not A203)  and  a20173a );
 a20178a <=( A269  and  A266 );
 a20179a <=( (not A265)  and  a20178a );
 a20180a <=( a20179a  and  a20174a );
 a20183a <=( (not A167)  and  A170 );
 a20187a <=( (not A202)  and  (not A201) );
 a20188a <=( A166  and  a20187a );
 a20189a <=( a20188a  and  a20183a );
 a20193a <=( A234  and  A232 );
 a20194a <=( (not A203)  and  a20193a );
 a20198a <=( A269  and  (not A266) );
 a20199a <=( A265  and  a20198a );
 a20200a <=( a20199a  and  a20194a );
 a20203a <=( (not A167)  and  A170 );
 a20207a <=( (not A202)  and  (not A201) );
 a20208a <=( A166  and  a20207a );
 a20209a <=( a20208a  and  a20203a );
 a20213a <=( A234  and  A233 );
 a20214a <=( (not A203)  and  a20213a );
 a20218a <=( (not A302)  and  (not A301) );
 a20219a <=( (not A300)  and  a20218a );
 a20220a <=( a20219a  and  a20214a );
 a20223a <=( (not A167)  and  A170 );
 a20227a <=( (not A202)  and  (not A201) );
 a20228a <=( A166  and  a20227a );
 a20229a <=( a20228a  and  a20223a );
 a20233a <=( A234  and  A233 );
 a20234a <=( (not A203)  and  a20233a );
 a20238a <=( (not A301)  and  (not A299) );
 a20239a <=( (not A298)  and  a20238a );
 a20240a <=( a20239a  and  a20234a );
 a20243a <=( (not A167)  and  A170 );
 a20247a <=( (not A202)  and  (not A201) );
 a20248a <=( A166  and  a20247a );
 a20249a <=( a20248a  and  a20243a );
 a20253a <=( A234  and  A233 );
 a20254a <=( (not A203)  and  a20253a );
 a20258a <=( A269  and  A266 );
 a20259a <=( (not A265)  and  a20258a );
 a20260a <=( a20259a  and  a20254a );
 a20263a <=( (not A167)  and  A170 );
 a20267a <=( (not A202)  and  (not A201) );
 a20268a <=( A166  and  a20267a );
 a20269a <=( a20268a  and  a20263a );
 a20273a <=( A234  and  A233 );
 a20274a <=( (not A203)  and  a20273a );
 a20278a <=( A269  and  (not A266) );
 a20279a <=( A265  and  a20278a );
 a20280a <=( a20279a  and  a20274a );
 a20283a <=( (not A167)  and  A170 );
 a20287a <=( (not A202)  and  (not A201) );
 a20288a <=( A166  and  a20287a );
 a20289a <=( a20288a  and  a20283a );
 a20293a <=( A233  and  (not A232) );
 a20294a <=( (not A203)  and  a20293a );
 a20298a <=( A267  and  A265 );
 a20299a <=( A236  and  a20298a );
 a20300a <=( a20299a  and  a20294a );
 a20303a <=( (not A167)  and  A170 );
 a20307a <=( (not A202)  and  (not A201) );
 a20308a <=( A166  and  a20307a );
 a20309a <=( a20308a  and  a20303a );
 a20313a <=( A233  and  (not A232) );
 a20314a <=( (not A203)  and  a20313a );
 a20318a <=( A267  and  A266 );
 a20319a <=( A236  and  a20318a );
 a20320a <=( a20319a  and  a20314a );
 a20323a <=( (not A167)  and  A170 );
 a20327a <=( (not A202)  and  (not A201) );
 a20328a <=( A166  and  a20327a );
 a20329a <=( a20328a  and  a20323a );
 a20333a <=( (not A233)  and  A232 );
 a20334a <=( (not A203)  and  a20333a );
 a20338a <=( A267  and  A265 );
 a20339a <=( A236  and  a20338a );
 a20340a <=( a20339a  and  a20334a );
 a20343a <=( (not A167)  and  A170 );
 a20347a <=( (not A202)  and  (not A201) );
 a20348a <=( A166  and  a20347a );
 a20349a <=( a20348a  and  a20343a );
 a20353a <=( (not A233)  and  A232 );
 a20354a <=( (not A203)  and  a20353a );
 a20358a <=( A267  and  A266 );
 a20359a <=( A236  and  a20358a );
 a20360a <=( a20359a  and  a20354a );
 a20363a <=( (not A167)  and  A170 );
 a20367a <=( A200  and  A199 );
 a20368a <=( A166  and  a20367a );
 a20369a <=( a20368a  and  a20363a );
 a20373a <=( A235  and  (not A202) );
 a20374a <=( (not A201)  and  a20373a );
 a20378a <=( (not A302)  and  (not A301) );
 a20379a <=( (not A300)  and  a20378a );
 a20380a <=( a20379a  and  a20374a );
 a20383a <=( (not A167)  and  A170 );
 a20387a <=( A200  and  A199 );
 a20388a <=( A166  and  a20387a );
 a20389a <=( a20388a  and  a20383a );
 a20393a <=( A235  and  (not A202) );
 a20394a <=( (not A201)  and  a20393a );
 a20398a <=( (not A301)  and  (not A299) );
 a20399a <=( (not A298)  and  a20398a );
 a20400a <=( a20399a  and  a20394a );
 a20403a <=( (not A167)  and  A170 );
 a20407a <=( A200  and  A199 );
 a20408a <=( A166  and  a20407a );
 a20409a <=( a20408a  and  a20403a );
 a20413a <=( A235  and  (not A202) );
 a20414a <=( (not A201)  and  a20413a );
 a20418a <=( A269  and  A266 );
 a20419a <=( (not A265)  and  a20418a );
 a20420a <=( a20419a  and  a20414a );
 a20423a <=( (not A167)  and  A170 );
 a20427a <=( A200  and  A199 );
 a20428a <=( A166  and  a20427a );
 a20429a <=( a20428a  and  a20423a );
 a20433a <=( A235  and  (not A202) );
 a20434a <=( (not A201)  and  a20433a );
 a20438a <=( A269  and  (not A266) );
 a20439a <=( A265  and  a20438a );
 a20440a <=( a20439a  and  a20434a );
 a20443a <=( (not A167)  and  A170 );
 a20447a <=( A200  and  A199 );
 a20448a <=( A166  and  a20447a );
 a20449a <=( a20448a  and  a20443a );
 a20453a <=( A232  and  (not A202) );
 a20454a <=( (not A201)  and  a20453a );
 a20458a <=( A267  and  A265 );
 a20459a <=( A234  and  a20458a );
 a20460a <=( a20459a  and  a20454a );
 a20463a <=( (not A167)  and  A170 );
 a20467a <=( A200  and  A199 );
 a20468a <=( A166  and  a20467a );
 a20469a <=( a20468a  and  a20463a );
 a20473a <=( A232  and  (not A202) );
 a20474a <=( (not A201)  and  a20473a );
 a20478a <=( A267  and  A266 );
 a20479a <=( A234  and  a20478a );
 a20480a <=( a20479a  and  a20474a );
 a20483a <=( (not A167)  and  A170 );
 a20487a <=( A200  and  A199 );
 a20488a <=( A166  and  a20487a );
 a20489a <=( a20488a  and  a20483a );
 a20493a <=( A233  and  (not A202) );
 a20494a <=( (not A201)  and  a20493a );
 a20498a <=( A267  and  A265 );
 a20499a <=( A234  and  a20498a );
 a20500a <=( a20499a  and  a20494a );
 a20503a <=( (not A167)  and  A170 );
 a20507a <=( A200  and  A199 );
 a20508a <=( A166  and  a20507a );
 a20509a <=( a20508a  and  a20503a );
 a20513a <=( A233  and  (not A202) );
 a20514a <=( (not A201)  and  a20513a );
 a20518a <=( A267  and  A266 );
 a20519a <=( A234  and  a20518a );
 a20520a <=( a20519a  and  a20514a );
 a20523a <=( (not A167)  and  A170 );
 a20527a <=( A200  and  A199 );
 a20528a <=( A166  and  a20527a );
 a20529a <=( a20528a  and  a20523a );
 a20533a <=( (not A232)  and  (not A202) );
 a20534a <=( (not A201)  and  a20533a );
 a20538a <=( A268  and  A236 );
 a20539a <=( A233  and  a20538a );
 a20540a <=( a20539a  and  a20534a );
 a20543a <=( (not A167)  and  A170 );
 a20547a <=( A200  and  A199 );
 a20548a <=( A166  and  a20547a );
 a20549a <=( a20548a  and  a20543a );
 a20553a <=( A232  and  (not A202) );
 a20554a <=( (not A201)  and  a20553a );
 a20558a <=( A268  and  A236 );
 a20559a <=( (not A233)  and  a20558a );
 a20560a <=( a20559a  and  a20554a );
 a20563a <=( (not A167)  and  A170 );
 a20567a <=( (not A200)  and  (not A199) );
 a20568a <=( A166  and  a20567a );
 a20569a <=( a20568a  and  a20563a );
 a20573a <=( A298  and  A235 );
 a20574a <=( (not A202)  and  a20573a );
 a20578a <=( (not A301)  and  (not A300) );
 a20579a <=( A299  and  a20578a );
 a20580a <=( a20579a  and  a20574a );
 a20583a <=( (not A167)  and  A170 );
 a20587a <=( (not A200)  and  (not A199) );
 a20588a <=( A166  and  a20587a );
 a20589a <=( a20588a  and  a20583a );
 a20593a <=( A234  and  A232 );
 a20594a <=( (not A202)  and  a20593a );
 a20598a <=( (not A302)  and  (not A301) );
 a20599a <=( (not A300)  and  a20598a );
 a20600a <=( a20599a  and  a20594a );
 a20603a <=( (not A167)  and  A170 );
 a20607a <=( (not A200)  and  (not A199) );
 a20608a <=( A166  and  a20607a );
 a20609a <=( a20608a  and  a20603a );
 a20613a <=( A234  and  A232 );
 a20614a <=( (not A202)  and  a20613a );
 a20618a <=( (not A301)  and  (not A299) );
 a20619a <=( (not A298)  and  a20618a );
 a20620a <=( a20619a  and  a20614a );
 a20623a <=( (not A167)  and  A170 );
 a20627a <=( (not A200)  and  (not A199) );
 a20628a <=( A166  and  a20627a );
 a20629a <=( a20628a  and  a20623a );
 a20633a <=( A234  and  A232 );
 a20634a <=( (not A202)  and  a20633a );
 a20638a <=( A269  and  A266 );
 a20639a <=( (not A265)  and  a20638a );
 a20640a <=( a20639a  and  a20634a );
 a20643a <=( (not A167)  and  A170 );
 a20647a <=( (not A200)  and  (not A199) );
 a20648a <=( A166  and  a20647a );
 a20649a <=( a20648a  and  a20643a );
 a20653a <=( A234  and  A232 );
 a20654a <=( (not A202)  and  a20653a );
 a20658a <=( A269  and  (not A266) );
 a20659a <=( A265  and  a20658a );
 a20660a <=( a20659a  and  a20654a );
 a20663a <=( (not A167)  and  A170 );
 a20667a <=( (not A200)  and  (not A199) );
 a20668a <=( A166  and  a20667a );
 a20669a <=( a20668a  and  a20663a );
 a20673a <=( A234  and  A233 );
 a20674a <=( (not A202)  and  a20673a );
 a20678a <=( (not A302)  and  (not A301) );
 a20679a <=( (not A300)  and  a20678a );
 a20680a <=( a20679a  and  a20674a );
 a20683a <=( (not A167)  and  A170 );
 a20687a <=( (not A200)  and  (not A199) );
 a20688a <=( A166  and  a20687a );
 a20689a <=( a20688a  and  a20683a );
 a20693a <=( A234  and  A233 );
 a20694a <=( (not A202)  and  a20693a );
 a20698a <=( (not A301)  and  (not A299) );
 a20699a <=( (not A298)  and  a20698a );
 a20700a <=( a20699a  and  a20694a );
 a20703a <=( (not A167)  and  A170 );
 a20707a <=( (not A200)  and  (not A199) );
 a20708a <=( A166  and  a20707a );
 a20709a <=( a20708a  and  a20703a );
 a20713a <=( A234  and  A233 );
 a20714a <=( (not A202)  and  a20713a );
 a20718a <=( A269  and  A266 );
 a20719a <=( (not A265)  and  a20718a );
 a20720a <=( a20719a  and  a20714a );
 a20723a <=( (not A167)  and  A170 );
 a20727a <=( (not A200)  and  (not A199) );
 a20728a <=( A166  and  a20727a );
 a20729a <=( a20728a  and  a20723a );
 a20733a <=( A234  and  A233 );
 a20734a <=( (not A202)  and  a20733a );
 a20738a <=( A269  and  (not A266) );
 a20739a <=( A265  and  a20738a );
 a20740a <=( a20739a  and  a20734a );
 a20743a <=( (not A167)  and  A170 );
 a20747a <=( (not A200)  and  (not A199) );
 a20748a <=( A166  and  a20747a );
 a20749a <=( a20748a  and  a20743a );
 a20753a <=( A233  and  (not A232) );
 a20754a <=( (not A202)  and  a20753a );
 a20758a <=( A267  and  A265 );
 a20759a <=( A236  and  a20758a );
 a20760a <=( a20759a  and  a20754a );
 a20763a <=( (not A167)  and  A170 );
 a20767a <=( (not A200)  and  (not A199) );
 a20768a <=( A166  and  a20767a );
 a20769a <=( a20768a  and  a20763a );
 a20773a <=( A233  and  (not A232) );
 a20774a <=( (not A202)  and  a20773a );
 a20778a <=( A267  and  A266 );
 a20779a <=( A236  and  a20778a );
 a20780a <=( a20779a  and  a20774a );
 a20783a <=( (not A167)  and  A170 );
 a20787a <=( (not A200)  and  (not A199) );
 a20788a <=( A166  and  a20787a );
 a20789a <=( a20788a  and  a20783a );
 a20793a <=( (not A233)  and  A232 );
 a20794a <=( (not A202)  and  a20793a );
 a20798a <=( A267  and  A265 );
 a20799a <=( A236  and  a20798a );
 a20800a <=( a20799a  and  a20794a );
 a20803a <=( (not A167)  and  A170 );
 a20807a <=( (not A200)  and  (not A199) );
 a20808a <=( A166  and  a20807a );
 a20809a <=( a20808a  and  a20803a );
 a20813a <=( (not A233)  and  A232 );
 a20814a <=( (not A202)  and  a20813a );
 a20818a <=( A267  and  A266 );
 a20819a <=( A236  and  a20818a );
 a20820a <=( a20819a  and  a20814a );
 a20823a <=( (not A201)  and  A169 );
 a20827a <=( (not A234)  and  (not A203) );
 a20828a <=( (not A202)  and  a20827a );
 a20829a <=( a20828a  and  a20823a );
 a20833a <=( (not A267)  and  (not A236) );
 a20834a <=( (not A235)  and  a20833a );
 a20838a <=( A301  and  (not A269) );
 a20839a <=( (not A268)  and  a20838a );
 a20840a <=( a20839a  and  a20834a );
 a20843a <=( (not A201)  and  A169 );
 a20847a <=( (not A234)  and  (not A203) );
 a20848a <=( (not A202)  and  a20847a );
 a20849a <=( a20848a  and  a20843a );
 a20853a <=( (not A265)  and  (not A236) );
 a20854a <=( (not A235)  and  a20853a );
 a20858a <=( A301  and  (not A268) );
 a20859a <=( (not A266)  and  a20858a );
 a20860a <=( a20859a  and  a20854a );
 a20863a <=( (not A201)  and  A169 );
 a20867a <=( (not A232)  and  (not A203) );
 a20868a <=( (not A202)  and  a20867a );
 a20869a <=( a20868a  and  a20863a );
 a20873a <=( A298  and  A236 );
 a20874a <=( A233  and  a20873a );
 a20878a <=( (not A301)  and  (not A300) );
 a20879a <=( A299  and  a20878a );
 a20880a <=( a20879a  and  a20874a );
 a20883a <=( (not A201)  and  A169 );
 a20887a <=( A232  and  (not A203) );
 a20888a <=( (not A202)  and  a20887a );
 a20889a <=( a20888a  and  a20883a );
 a20893a <=( A298  and  A236 );
 a20894a <=( (not A233)  and  a20893a );
 a20898a <=( (not A301)  and  (not A300) );
 a20899a <=( A299  and  a20898a );
 a20900a <=( a20899a  and  a20894a );
 a20903a <=( (not A201)  and  A169 );
 a20907a <=( (not A232)  and  (not A203) );
 a20908a <=( (not A202)  and  a20907a );
 a20909a <=( a20908a  and  a20903a );
 a20913a <=( (not A267)  and  (not A235) );
 a20914a <=( (not A233)  and  a20913a );
 a20918a <=( A301  and  (not A269) );
 a20919a <=( (not A268)  and  a20918a );
 a20920a <=( a20919a  and  a20914a );
 a20923a <=( (not A201)  and  A169 );
 a20927a <=( (not A232)  and  (not A203) );
 a20928a <=( (not A202)  and  a20927a );
 a20929a <=( a20928a  and  a20923a );
 a20933a <=( (not A265)  and  (not A235) );
 a20934a <=( (not A233)  and  a20933a );
 a20938a <=( A301  and  (not A268) );
 a20939a <=( (not A266)  and  a20938a );
 a20940a <=( a20939a  and  a20934a );
 a20943a <=( A199  and  A169 );
 a20947a <=( (not A202)  and  (not A201) );
 a20948a <=( A200  and  a20947a );
 a20949a <=( a20948a  and  a20943a );
 a20953a <=( A298  and  A234 );
 a20954a <=( A232  and  a20953a );
 a20958a <=( (not A301)  and  (not A300) );
 a20959a <=( A299  and  a20958a );
 a20960a <=( a20959a  and  a20954a );
 a20963a <=( A199  and  A169 );
 a20967a <=( (not A202)  and  (not A201) );
 a20968a <=( A200  and  a20967a );
 a20969a <=( a20968a  and  a20963a );
 a20973a <=( A298  and  A234 );
 a20974a <=( A233  and  a20973a );
 a20978a <=( (not A301)  and  (not A300) );
 a20979a <=( A299  and  a20978a );
 a20980a <=( a20979a  and  a20974a );
 a20983a <=( A199  and  A169 );
 a20987a <=( (not A202)  and  (not A201) );
 a20988a <=( A200  and  a20987a );
 a20989a <=( a20988a  and  a20983a );
 a20993a <=( A236  and  A233 );
 a20994a <=( (not A232)  and  a20993a );
 a20998a <=( (not A302)  and  (not A301) );
 a20999a <=( (not A300)  and  a20998a );
 a21000a <=( a20999a  and  a20994a );
 a21003a <=( A199  and  A169 );
 a21007a <=( (not A202)  and  (not A201) );
 a21008a <=( A200  and  a21007a );
 a21009a <=( a21008a  and  a21003a );
 a21013a <=( A236  and  A233 );
 a21014a <=( (not A232)  and  a21013a );
 a21018a <=( (not A301)  and  (not A299) );
 a21019a <=( (not A298)  and  a21018a );
 a21020a <=( a21019a  and  a21014a );
 a21023a <=( A199  and  A169 );
 a21027a <=( (not A202)  and  (not A201) );
 a21028a <=( A200  and  a21027a );
 a21029a <=( a21028a  and  a21023a );
 a21033a <=( A236  and  A233 );
 a21034a <=( (not A232)  and  a21033a );
 a21038a <=( A269  and  A266 );
 a21039a <=( (not A265)  and  a21038a );
 a21040a <=( a21039a  and  a21034a );
 a21043a <=( A199  and  A169 );
 a21047a <=( (not A202)  and  (not A201) );
 a21048a <=( A200  and  a21047a );
 a21049a <=( a21048a  and  a21043a );
 a21053a <=( A236  and  A233 );
 a21054a <=( (not A232)  and  a21053a );
 a21058a <=( A269  and  (not A266) );
 a21059a <=( A265  and  a21058a );
 a21060a <=( a21059a  and  a21054a );
 a21063a <=( A199  and  A169 );
 a21067a <=( (not A202)  and  (not A201) );
 a21068a <=( A200  and  a21067a );
 a21069a <=( a21068a  and  a21063a );
 a21073a <=( A236  and  (not A233) );
 a21074a <=( A232  and  a21073a );
 a21078a <=( (not A302)  and  (not A301) );
 a21079a <=( (not A300)  and  a21078a );
 a21080a <=( a21079a  and  a21074a );
 a21083a <=( A199  and  A169 );
 a21087a <=( (not A202)  and  (not A201) );
 a21088a <=( A200  and  a21087a );
 a21089a <=( a21088a  and  a21083a );
 a21093a <=( A236  and  (not A233) );
 a21094a <=( A232  and  a21093a );
 a21098a <=( (not A301)  and  (not A299) );
 a21099a <=( (not A298)  and  a21098a );
 a21100a <=( a21099a  and  a21094a );
 a21103a <=( A199  and  A169 );
 a21107a <=( (not A202)  and  (not A201) );
 a21108a <=( A200  and  a21107a );
 a21109a <=( a21108a  and  a21103a );
 a21113a <=( A236  and  (not A233) );
 a21114a <=( A232  and  a21113a );
 a21118a <=( A269  and  A266 );
 a21119a <=( (not A265)  and  a21118a );
 a21120a <=( a21119a  and  a21114a );
 a21123a <=( A199  and  A169 );
 a21127a <=( (not A202)  and  (not A201) );
 a21128a <=( A200  and  a21127a );
 a21129a <=( a21128a  and  a21123a );
 a21133a <=( A236  and  (not A233) );
 a21134a <=( A232  and  a21133a );
 a21138a <=( A269  and  (not A266) );
 a21139a <=( A265  and  a21138a );
 a21140a <=( a21139a  and  a21134a );
 a21143a <=( (not A199)  and  A169 );
 a21147a <=( (not A234)  and  (not A202) );
 a21148a <=( (not A200)  and  a21147a );
 a21149a <=( a21148a  and  a21143a );
 a21153a <=( (not A267)  and  (not A236) );
 a21154a <=( (not A235)  and  a21153a );
 a21158a <=( A301  and  (not A269) );
 a21159a <=( (not A268)  and  a21158a );
 a21160a <=( a21159a  and  a21154a );
 a21163a <=( (not A199)  and  A169 );
 a21167a <=( (not A234)  and  (not A202) );
 a21168a <=( (not A200)  and  a21167a );
 a21169a <=( a21168a  and  a21163a );
 a21173a <=( (not A265)  and  (not A236) );
 a21174a <=( (not A235)  and  a21173a );
 a21178a <=( A301  and  (not A268) );
 a21179a <=( (not A266)  and  a21178a );
 a21180a <=( a21179a  and  a21174a );
 a21183a <=( (not A199)  and  A169 );
 a21187a <=( (not A232)  and  (not A202) );
 a21188a <=( (not A200)  and  a21187a );
 a21189a <=( a21188a  and  a21183a );
 a21193a <=( A298  and  A236 );
 a21194a <=( A233  and  a21193a );
 a21198a <=( (not A301)  and  (not A300) );
 a21199a <=( A299  and  a21198a );
 a21200a <=( a21199a  and  a21194a );
 a21203a <=( (not A199)  and  A169 );
 a21207a <=( A232  and  (not A202) );
 a21208a <=( (not A200)  and  a21207a );
 a21209a <=( a21208a  and  a21203a );
 a21213a <=( A298  and  A236 );
 a21214a <=( (not A233)  and  a21213a );
 a21218a <=( (not A301)  and  (not A300) );
 a21219a <=( A299  and  a21218a );
 a21220a <=( a21219a  and  a21214a );
 a21223a <=( (not A199)  and  A169 );
 a21227a <=( (not A232)  and  (not A202) );
 a21228a <=( (not A200)  and  a21227a );
 a21229a <=( a21228a  and  a21223a );
 a21233a <=( (not A267)  and  (not A235) );
 a21234a <=( (not A233)  and  a21233a );
 a21238a <=( A301  and  (not A269) );
 a21239a <=( (not A268)  and  a21238a );
 a21240a <=( a21239a  and  a21234a );
 a21243a <=( (not A199)  and  A169 );
 a21247a <=( (not A232)  and  (not A202) );
 a21248a <=( (not A200)  and  a21247a );
 a21249a <=( a21248a  and  a21243a );
 a21253a <=( (not A265)  and  (not A235) );
 a21254a <=( (not A233)  and  a21253a );
 a21258a <=( A301  and  (not A268) );
 a21259a <=( (not A266)  and  a21258a );
 a21260a <=( a21259a  and  a21254a );
 a21263a <=( (not A167)  and  (not A169) );
 a21267a <=( (not A234)  and  A202 );
 a21268a <=( (not A166)  and  a21267a );
 a21269a <=( a21268a  and  a21263a );
 a21273a <=( (not A267)  and  (not A236) );
 a21274a <=( (not A235)  and  a21273a );
 a21278a <=( A301  and  (not A269) );
 a21279a <=( (not A268)  and  a21278a );
 a21280a <=( a21279a  and  a21274a );
 a21283a <=( (not A167)  and  (not A169) );
 a21287a <=( (not A234)  and  A202 );
 a21288a <=( (not A166)  and  a21287a );
 a21289a <=( a21288a  and  a21283a );
 a21293a <=( (not A265)  and  (not A236) );
 a21294a <=( (not A235)  and  a21293a );
 a21298a <=( A301  and  (not A268) );
 a21299a <=( (not A266)  and  a21298a );
 a21300a <=( a21299a  and  a21294a );
 a21303a <=( (not A167)  and  (not A169) );
 a21307a <=( (not A232)  and  A202 );
 a21308a <=( (not A166)  and  a21307a );
 a21309a <=( a21308a  and  a21303a );
 a21313a <=( A298  and  A236 );
 a21314a <=( A233  and  a21313a );
 a21318a <=( (not A301)  and  (not A300) );
 a21319a <=( A299  and  a21318a );
 a21320a <=( a21319a  and  a21314a );
 a21323a <=( (not A167)  and  (not A169) );
 a21327a <=( A232  and  A202 );
 a21328a <=( (not A166)  and  a21327a );
 a21329a <=( a21328a  and  a21323a );
 a21333a <=( A298  and  A236 );
 a21334a <=( (not A233)  and  a21333a );
 a21338a <=( (not A301)  and  (not A300) );
 a21339a <=( A299  and  a21338a );
 a21340a <=( a21339a  and  a21334a );
 a21343a <=( (not A167)  and  (not A169) );
 a21347a <=( (not A232)  and  A202 );
 a21348a <=( (not A166)  and  a21347a );
 a21349a <=( a21348a  and  a21343a );
 a21353a <=( (not A267)  and  (not A235) );
 a21354a <=( (not A233)  and  a21353a );
 a21358a <=( A301  and  (not A269) );
 a21359a <=( (not A268)  and  a21358a );
 a21360a <=( a21359a  and  a21354a );
 a21363a <=( (not A167)  and  (not A169) );
 a21367a <=( (not A232)  and  A202 );
 a21368a <=( (not A166)  and  a21367a );
 a21369a <=( a21368a  and  a21363a );
 a21373a <=( (not A265)  and  (not A235) );
 a21374a <=( (not A233)  and  a21373a );
 a21378a <=( A301  and  (not A268) );
 a21379a <=( (not A266)  and  a21378a );
 a21380a <=( a21379a  and  a21374a );
 a21383a <=( (not A167)  and  (not A169) );
 a21387a <=( A201  and  A199 );
 a21388a <=( (not A166)  and  a21387a );
 a21389a <=( a21388a  and  a21383a );
 a21393a <=( A298  and  A234 );
 a21394a <=( A232  and  a21393a );
 a21398a <=( (not A301)  and  (not A300) );
 a21399a <=( A299  and  a21398a );
 a21400a <=( a21399a  and  a21394a );
 a21403a <=( (not A167)  and  (not A169) );
 a21407a <=( A201  and  A199 );
 a21408a <=( (not A166)  and  a21407a );
 a21409a <=( a21408a  and  a21403a );
 a21413a <=( A298  and  A234 );
 a21414a <=( A233  and  a21413a );
 a21418a <=( (not A301)  and  (not A300) );
 a21419a <=( A299  and  a21418a );
 a21420a <=( a21419a  and  a21414a );
 a21423a <=( (not A167)  and  (not A169) );
 a21427a <=( A201  and  A199 );
 a21428a <=( (not A166)  and  a21427a );
 a21429a <=( a21428a  and  a21423a );
 a21433a <=( A236  and  A233 );
 a21434a <=( (not A232)  and  a21433a );
 a21438a <=( (not A302)  and  (not A301) );
 a21439a <=( (not A300)  and  a21438a );
 a21440a <=( a21439a  and  a21434a );
 a21443a <=( (not A167)  and  (not A169) );
 a21447a <=( A201  and  A199 );
 a21448a <=( (not A166)  and  a21447a );
 a21449a <=( a21448a  and  a21443a );
 a21453a <=( A236  and  A233 );
 a21454a <=( (not A232)  and  a21453a );
 a21458a <=( (not A301)  and  (not A299) );
 a21459a <=( (not A298)  and  a21458a );
 a21460a <=( a21459a  and  a21454a );
 a21463a <=( (not A167)  and  (not A169) );
 a21467a <=( A201  and  A199 );
 a21468a <=( (not A166)  and  a21467a );
 a21469a <=( a21468a  and  a21463a );
 a21473a <=( A236  and  A233 );
 a21474a <=( (not A232)  and  a21473a );
 a21478a <=( A269  and  A266 );
 a21479a <=( (not A265)  and  a21478a );
 a21480a <=( a21479a  and  a21474a );
 a21483a <=( (not A167)  and  (not A169) );
 a21487a <=( A201  and  A199 );
 a21488a <=( (not A166)  and  a21487a );
 a21489a <=( a21488a  and  a21483a );
 a21493a <=( A236  and  A233 );
 a21494a <=( (not A232)  and  a21493a );
 a21498a <=( A269  and  (not A266) );
 a21499a <=( A265  and  a21498a );
 a21500a <=( a21499a  and  a21494a );
 a21503a <=( (not A167)  and  (not A169) );
 a21507a <=( A201  and  A199 );
 a21508a <=( (not A166)  and  a21507a );
 a21509a <=( a21508a  and  a21503a );
 a21513a <=( A236  and  (not A233) );
 a21514a <=( A232  and  a21513a );
 a21518a <=( (not A302)  and  (not A301) );
 a21519a <=( (not A300)  and  a21518a );
 a21520a <=( a21519a  and  a21514a );
 a21523a <=( (not A167)  and  (not A169) );
 a21527a <=( A201  and  A199 );
 a21528a <=( (not A166)  and  a21527a );
 a21529a <=( a21528a  and  a21523a );
 a21533a <=( A236  and  (not A233) );
 a21534a <=( A232  and  a21533a );
 a21538a <=( (not A301)  and  (not A299) );
 a21539a <=( (not A298)  and  a21538a );
 a21540a <=( a21539a  and  a21534a );
 a21543a <=( (not A167)  and  (not A169) );
 a21547a <=( A201  and  A199 );
 a21548a <=( (not A166)  and  a21547a );
 a21549a <=( a21548a  and  a21543a );
 a21553a <=( A236  and  (not A233) );
 a21554a <=( A232  and  a21553a );
 a21558a <=( A269  and  A266 );
 a21559a <=( (not A265)  and  a21558a );
 a21560a <=( a21559a  and  a21554a );
 a21563a <=( (not A167)  and  (not A169) );
 a21567a <=( A201  and  A199 );
 a21568a <=( (not A166)  and  a21567a );
 a21569a <=( a21568a  and  a21563a );
 a21573a <=( A236  and  (not A233) );
 a21574a <=( A232  and  a21573a );
 a21578a <=( A269  and  (not A266) );
 a21579a <=( A265  and  a21578a );
 a21580a <=( a21579a  and  a21574a );
 a21583a <=( (not A167)  and  (not A169) );
 a21587a <=( A201  and  A200 );
 a21588a <=( (not A166)  and  a21587a );
 a21589a <=( a21588a  and  a21583a );
 a21593a <=( A298  and  A234 );
 a21594a <=( A232  and  a21593a );
 a21598a <=( (not A301)  and  (not A300) );
 a21599a <=( A299  and  a21598a );
 a21600a <=( a21599a  and  a21594a );
 a21603a <=( (not A167)  and  (not A169) );
 a21607a <=( A201  and  A200 );
 a21608a <=( (not A166)  and  a21607a );
 a21609a <=( a21608a  and  a21603a );
 a21613a <=( A298  and  A234 );
 a21614a <=( A233  and  a21613a );
 a21618a <=( (not A301)  and  (not A300) );
 a21619a <=( A299  and  a21618a );
 a21620a <=( a21619a  and  a21614a );
 a21623a <=( (not A167)  and  (not A169) );
 a21627a <=( A201  and  A200 );
 a21628a <=( (not A166)  and  a21627a );
 a21629a <=( a21628a  and  a21623a );
 a21633a <=( A236  and  A233 );
 a21634a <=( (not A232)  and  a21633a );
 a21638a <=( (not A302)  and  (not A301) );
 a21639a <=( (not A300)  and  a21638a );
 a21640a <=( a21639a  and  a21634a );
 a21643a <=( (not A167)  and  (not A169) );
 a21647a <=( A201  and  A200 );
 a21648a <=( (not A166)  and  a21647a );
 a21649a <=( a21648a  and  a21643a );
 a21653a <=( A236  and  A233 );
 a21654a <=( (not A232)  and  a21653a );
 a21658a <=( (not A301)  and  (not A299) );
 a21659a <=( (not A298)  and  a21658a );
 a21660a <=( a21659a  and  a21654a );
 a21663a <=( (not A167)  and  (not A169) );
 a21667a <=( A201  and  A200 );
 a21668a <=( (not A166)  and  a21667a );
 a21669a <=( a21668a  and  a21663a );
 a21673a <=( A236  and  A233 );
 a21674a <=( (not A232)  and  a21673a );
 a21678a <=( A269  and  A266 );
 a21679a <=( (not A265)  and  a21678a );
 a21680a <=( a21679a  and  a21674a );
 a21683a <=( (not A167)  and  (not A169) );
 a21687a <=( A201  and  A200 );
 a21688a <=( (not A166)  and  a21687a );
 a21689a <=( a21688a  and  a21683a );
 a21693a <=( A236  and  A233 );
 a21694a <=( (not A232)  and  a21693a );
 a21698a <=( A269  and  (not A266) );
 a21699a <=( A265  and  a21698a );
 a21700a <=( a21699a  and  a21694a );
 a21703a <=( (not A167)  and  (not A169) );
 a21707a <=( A201  and  A200 );
 a21708a <=( (not A166)  and  a21707a );
 a21709a <=( a21708a  and  a21703a );
 a21713a <=( A236  and  (not A233) );
 a21714a <=( A232  and  a21713a );
 a21718a <=( (not A302)  and  (not A301) );
 a21719a <=( (not A300)  and  a21718a );
 a21720a <=( a21719a  and  a21714a );
 a21723a <=( (not A167)  and  (not A169) );
 a21727a <=( A201  and  A200 );
 a21728a <=( (not A166)  and  a21727a );
 a21729a <=( a21728a  and  a21723a );
 a21733a <=( A236  and  (not A233) );
 a21734a <=( A232  and  a21733a );
 a21738a <=( (not A301)  and  (not A299) );
 a21739a <=( (not A298)  and  a21738a );
 a21740a <=( a21739a  and  a21734a );
 a21743a <=( (not A167)  and  (not A169) );
 a21747a <=( A201  and  A200 );
 a21748a <=( (not A166)  and  a21747a );
 a21749a <=( a21748a  and  a21743a );
 a21753a <=( A236  and  (not A233) );
 a21754a <=( A232  and  a21753a );
 a21758a <=( A269  and  A266 );
 a21759a <=( (not A265)  and  a21758a );
 a21760a <=( a21759a  and  a21754a );
 a21763a <=( (not A167)  and  (not A169) );
 a21767a <=( A201  and  A200 );
 a21768a <=( (not A166)  and  a21767a );
 a21769a <=( a21768a  and  a21763a );
 a21773a <=( A236  and  (not A233) );
 a21774a <=( A232  and  a21773a );
 a21778a <=( A269  and  (not A266) );
 a21779a <=( A265  and  a21778a );
 a21780a <=( a21779a  and  a21774a );
 a21783a <=( (not A167)  and  (not A169) );
 a21787a <=( A200  and  (not A199) );
 a21788a <=( (not A166)  and  a21787a );
 a21789a <=( a21788a  and  a21783a );
 a21793a <=( A298  and  A235 );
 a21794a <=( A203  and  a21793a );
 a21798a <=( (not A301)  and  (not A300) );
 a21799a <=( A299  and  a21798a );
 a21800a <=( a21799a  and  a21794a );
 a21803a <=( (not A167)  and  (not A169) );
 a21807a <=( A200  and  (not A199) );
 a21808a <=( (not A166)  and  a21807a );
 a21809a <=( a21808a  and  a21803a );
 a21813a <=( A234  and  A232 );
 a21814a <=( A203  and  a21813a );
 a21818a <=( (not A302)  and  (not A301) );
 a21819a <=( (not A300)  and  a21818a );
 a21820a <=( a21819a  and  a21814a );
 a21823a <=( (not A167)  and  (not A169) );
 a21827a <=( A200  and  (not A199) );
 a21828a <=( (not A166)  and  a21827a );
 a21829a <=( a21828a  and  a21823a );
 a21833a <=( A234  and  A232 );
 a21834a <=( A203  and  a21833a );
 a21838a <=( (not A301)  and  (not A299) );
 a21839a <=( (not A298)  and  a21838a );
 a21840a <=( a21839a  and  a21834a );
 a21843a <=( (not A167)  and  (not A169) );
 a21847a <=( A200  and  (not A199) );
 a21848a <=( (not A166)  and  a21847a );
 a21849a <=( a21848a  and  a21843a );
 a21853a <=( A234  and  A232 );
 a21854a <=( A203  and  a21853a );
 a21858a <=( A269  and  A266 );
 a21859a <=( (not A265)  and  a21858a );
 a21860a <=( a21859a  and  a21854a );
 a21863a <=( (not A167)  and  (not A169) );
 a21867a <=( A200  and  (not A199) );
 a21868a <=( (not A166)  and  a21867a );
 a21869a <=( a21868a  and  a21863a );
 a21873a <=( A234  and  A232 );
 a21874a <=( A203  and  a21873a );
 a21878a <=( A269  and  (not A266) );
 a21879a <=( A265  and  a21878a );
 a21880a <=( a21879a  and  a21874a );
 a21883a <=( (not A167)  and  (not A169) );
 a21887a <=( A200  and  (not A199) );
 a21888a <=( (not A166)  and  a21887a );
 a21889a <=( a21888a  and  a21883a );
 a21893a <=( A234  and  A233 );
 a21894a <=( A203  and  a21893a );
 a21898a <=( (not A302)  and  (not A301) );
 a21899a <=( (not A300)  and  a21898a );
 a21900a <=( a21899a  and  a21894a );
 a21903a <=( (not A167)  and  (not A169) );
 a21907a <=( A200  and  (not A199) );
 a21908a <=( (not A166)  and  a21907a );
 a21909a <=( a21908a  and  a21903a );
 a21913a <=( A234  and  A233 );
 a21914a <=( A203  and  a21913a );
 a21918a <=( (not A301)  and  (not A299) );
 a21919a <=( (not A298)  and  a21918a );
 a21920a <=( a21919a  and  a21914a );
 a21923a <=( (not A167)  and  (not A169) );
 a21927a <=( A200  and  (not A199) );
 a21928a <=( (not A166)  and  a21927a );
 a21929a <=( a21928a  and  a21923a );
 a21933a <=( A234  and  A233 );
 a21934a <=( A203  and  a21933a );
 a21938a <=( A269  and  A266 );
 a21939a <=( (not A265)  and  a21938a );
 a21940a <=( a21939a  and  a21934a );
 a21943a <=( (not A167)  and  (not A169) );
 a21947a <=( A200  and  (not A199) );
 a21948a <=( (not A166)  and  a21947a );
 a21949a <=( a21948a  and  a21943a );
 a21953a <=( A234  and  A233 );
 a21954a <=( A203  and  a21953a );
 a21958a <=( A269  and  (not A266) );
 a21959a <=( A265  and  a21958a );
 a21960a <=( a21959a  and  a21954a );
 a21963a <=( (not A167)  and  (not A169) );
 a21967a <=( A200  and  (not A199) );
 a21968a <=( (not A166)  and  a21967a );
 a21969a <=( a21968a  and  a21963a );
 a21973a <=( A233  and  (not A232) );
 a21974a <=( A203  and  a21973a );
 a21978a <=( A267  and  A265 );
 a21979a <=( A236  and  a21978a );
 a21980a <=( a21979a  and  a21974a );
 a21983a <=( (not A167)  and  (not A169) );
 a21987a <=( A200  and  (not A199) );
 a21988a <=( (not A166)  and  a21987a );
 a21989a <=( a21988a  and  a21983a );
 a21993a <=( A233  and  (not A232) );
 a21994a <=( A203  and  a21993a );
 a21998a <=( A267  and  A266 );
 a21999a <=( A236  and  a21998a );
 a22000a <=( a21999a  and  a21994a );
 a22003a <=( (not A167)  and  (not A169) );
 a22007a <=( A200  and  (not A199) );
 a22008a <=( (not A166)  and  a22007a );
 a22009a <=( a22008a  and  a22003a );
 a22013a <=( (not A233)  and  A232 );
 a22014a <=( A203  and  a22013a );
 a22018a <=( A267  and  A265 );
 a22019a <=( A236  and  a22018a );
 a22020a <=( a22019a  and  a22014a );
 a22023a <=( (not A167)  and  (not A169) );
 a22027a <=( A200  and  (not A199) );
 a22028a <=( (not A166)  and  a22027a );
 a22029a <=( a22028a  and  a22023a );
 a22033a <=( (not A233)  and  A232 );
 a22034a <=( A203  and  a22033a );
 a22038a <=( A267  and  A266 );
 a22039a <=( A236  and  a22038a );
 a22040a <=( a22039a  and  a22034a );
 a22043a <=( (not A167)  and  (not A169) );
 a22047a <=( (not A200)  and  A199 );
 a22048a <=( (not A166)  and  a22047a );
 a22049a <=( a22048a  and  a22043a );
 a22053a <=( A298  and  A235 );
 a22054a <=( A203  and  a22053a );
 a22058a <=( (not A301)  and  (not A300) );
 a22059a <=( A299  and  a22058a );
 a22060a <=( a22059a  and  a22054a );
 a22063a <=( (not A167)  and  (not A169) );
 a22067a <=( (not A200)  and  A199 );
 a22068a <=( (not A166)  and  a22067a );
 a22069a <=( a22068a  and  a22063a );
 a22073a <=( A234  and  A232 );
 a22074a <=( A203  and  a22073a );
 a22078a <=( (not A302)  and  (not A301) );
 a22079a <=( (not A300)  and  a22078a );
 a22080a <=( a22079a  and  a22074a );
 a22083a <=( (not A167)  and  (not A169) );
 a22087a <=( (not A200)  and  A199 );
 a22088a <=( (not A166)  and  a22087a );
 a22089a <=( a22088a  and  a22083a );
 a22093a <=( A234  and  A232 );
 a22094a <=( A203  and  a22093a );
 a22098a <=( (not A301)  and  (not A299) );
 a22099a <=( (not A298)  and  a22098a );
 a22100a <=( a22099a  and  a22094a );
 a22103a <=( (not A167)  and  (not A169) );
 a22107a <=( (not A200)  and  A199 );
 a22108a <=( (not A166)  and  a22107a );
 a22109a <=( a22108a  and  a22103a );
 a22113a <=( A234  and  A232 );
 a22114a <=( A203  and  a22113a );
 a22118a <=( A269  and  A266 );
 a22119a <=( (not A265)  and  a22118a );
 a22120a <=( a22119a  and  a22114a );
 a22123a <=( (not A167)  and  (not A169) );
 a22127a <=( (not A200)  and  A199 );
 a22128a <=( (not A166)  and  a22127a );
 a22129a <=( a22128a  and  a22123a );
 a22133a <=( A234  and  A232 );
 a22134a <=( A203  and  a22133a );
 a22138a <=( A269  and  (not A266) );
 a22139a <=( A265  and  a22138a );
 a22140a <=( a22139a  and  a22134a );
 a22143a <=( (not A167)  and  (not A169) );
 a22147a <=( (not A200)  and  A199 );
 a22148a <=( (not A166)  and  a22147a );
 a22149a <=( a22148a  and  a22143a );
 a22153a <=( A234  and  A233 );
 a22154a <=( A203  and  a22153a );
 a22158a <=( (not A302)  and  (not A301) );
 a22159a <=( (not A300)  and  a22158a );
 a22160a <=( a22159a  and  a22154a );
 a22163a <=( (not A167)  and  (not A169) );
 a22167a <=( (not A200)  and  A199 );
 a22168a <=( (not A166)  and  a22167a );
 a22169a <=( a22168a  and  a22163a );
 a22173a <=( A234  and  A233 );
 a22174a <=( A203  and  a22173a );
 a22178a <=( (not A301)  and  (not A299) );
 a22179a <=( (not A298)  and  a22178a );
 a22180a <=( a22179a  and  a22174a );
 a22183a <=( (not A167)  and  (not A169) );
 a22187a <=( (not A200)  and  A199 );
 a22188a <=( (not A166)  and  a22187a );
 a22189a <=( a22188a  and  a22183a );
 a22193a <=( A234  and  A233 );
 a22194a <=( A203  and  a22193a );
 a22198a <=( A269  and  A266 );
 a22199a <=( (not A265)  and  a22198a );
 a22200a <=( a22199a  and  a22194a );
 a22203a <=( (not A167)  and  (not A169) );
 a22207a <=( (not A200)  and  A199 );
 a22208a <=( (not A166)  and  a22207a );
 a22209a <=( a22208a  and  a22203a );
 a22213a <=( A234  and  A233 );
 a22214a <=( A203  and  a22213a );
 a22218a <=( A269  and  (not A266) );
 a22219a <=( A265  and  a22218a );
 a22220a <=( a22219a  and  a22214a );
 a22223a <=( (not A167)  and  (not A169) );
 a22227a <=( (not A200)  and  A199 );
 a22228a <=( (not A166)  and  a22227a );
 a22229a <=( a22228a  and  a22223a );
 a22233a <=( A233  and  (not A232) );
 a22234a <=( A203  and  a22233a );
 a22238a <=( A267  and  A265 );
 a22239a <=( A236  and  a22238a );
 a22240a <=( a22239a  and  a22234a );
 a22243a <=( (not A167)  and  (not A169) );
 a22247a <=( (not A200)  and  A199 );
 a22248a <=( (not A166)  and  a22247a );
 a22249a <=( a22248a  and  a22243a );
 a22253a <=( A233  and  (not A232) );
 a22254a <=( A203  and  a22253a );
 a22258a <=( A267  and  A266 );
 a22259a <=( A236  and  a22258a );
 a22260a <=( a22259a  and  a22254a );
 a22263a <=( (not A167)  and  (not A169) );
 a22267a <=( (not A200)  and  A199 );
 a22268a <=( (not A166)  and  a22267a );
 a22269a <=( a22268a  and  a22263a );
 a22273a <=( (not A233)  and  A232 );
 a22274a <=( A203  and  a22273a );
 a22278a <=( A267  and  A265 );
 a22279a <=( A236  and  a22278a );
 a22280a <=( a22279a  and  a22274a );
 a22283a <=( (not A167)  and  (not A169) );
 a22287a <=( (not A200)  and  A199 );
 a22288a <=( (not A166)  and  a22287a );
 a22289a <=( a22288a  and  a22283a );
 a22293a <=( (not A233)  and  A232 );
 a22294a <=( A203  and  a22293a );
 a22298a <=( A267  and  A266 );
 a22299a <=( A236  and  a22298a );
 a22300a <=( a22299a  and  a22294a );
 a22303a <=( (not A168)  and  (not A169) );
 a22307a <=( A202  and  A166 );
 a22308a <=( A167  and  a22307a );
 a22309a <=( a22308a  and  a22303a );
 a22313a <=( A298  and  A234 );
 a22314a <=( A232  and  a22313a );
 a22318a <=( (not A301)  and  (not A300) );
 a22319a <=( A299  and  a22318a );
 a22320a <=( a22319a  and  a22314a );
 a22323a <=( (not A168)  and  (not A169) );
 a22327a <=( A202  and  A166 );
 a22328a <=( A167  and  a22327a );
 a22329a <=( a22328a  and  a22323a );
 a22333a <=( A298  and  A234 );
 a22334a <=( A233  and  a22333a );
 a22338a <=( (not A301)  and  (not A300) );
 a22339a <=( A299  and  a22338a );
 a22340a <=( a22339a  and  a22334a );
 a22343a <=( (not A168)  and  (not A169) );
 a22347a <=( A202  and  A166 );
 a22348a <=( A167  and  a22347a );
 a22349a <=( a22348a  and  a22343a );
 a22353a <=( A236  and  A233 );
 a22354a <=( (not A232)  and  a22353a );
 a22358a <=( (not A302)  and  (not A301) );
 a22359a <=( (not A300)  and  a22358a );
 a22360a <=( a22359a  and  a22354a );
 a22363a <=( (not A168)  and  (not A169) );
 a22367a <=( A202  and  A166 );
 a22368a <=( A167  and  a22367a );
 a22369a <=( a22368a  and  a22363a );
 a22373a <=( A236  and  A233 );
 a22374a <=( (not A232)  and  a22373a );
 a22378a <=( (not A301)  and  (not A299) );
 a22379a <=( (not A298)  and  a22378a );
 a22380a <=( a22379a  and  a22374a );
 a22383a <=( (not A168)  and  (not A169) );
 a22387a <=( A202  and  A166 );
 a22388a <=( A167  and  a22387a );
 a22389a <=( a22388a  and  a22383a );
 a22393a <=( A236  and  A233 );
 a22394a <=( (not A232)  and  a22393a );
 a22398a <=( A269  and  A266 );
 a22399a <=( (not A265)  and  a22398a );
 a22400a <=( a22399a  and  a22394a );
 a22403a <=( (not A168)  and  (not A169) );
 a22407a <=( A202  and  A166 );
 a22408a <=( A167  and  a22407a );
 a22409a <=( a22408a  and  a22403a );
 a22413a <=( A236  and  A233 );
 a22414a <=( (not A232)  and  a22413a );
 a22418a <=( A269  and  (not A266) );
 a22419a <=( A265  and  a22418a );
 a22420a <=( a22419a  and  a22414a );
 a22423a <=( (not A168)  and  (not A169) );
 a22427a <=( A202  and  A166 );
 a22428a <=( A167  and  a22427a );
 a22429a <=( a22428a  and  a22423a );
 a22433a <=( A236  and  (not A233) );
 a22434a <=( A232  and  a22433a );
 a22438a <=( (not A302)  and  (not A301) );
 a22439a <=( (not A300)  and  a22438a );
 a22440a <=( a22439a  and  a22434a );
 a22443a <=( (not A168)  and  (not A169) );
 a22447a <=( A202  and  A166 );
 a22448a <=( A167  and  a22447a );
 a22449a <=( a22448a  and  a22443a );
 a22453a <=( A236  and  (not A233) );
 a22454a <=( A232  and  a22453a );
 a22458a <=( (not A301)  and  (not A299) );
 a22459a <=( (not A298)  and  a22458a );
 a22460a <=( a22459a  and  a22454a );
 a22463a <=( (not A168)  and  (not A169) );
 a22467a <=( A202  and  A166 );
 a22468a <=( A167  and  a22467a );
 a22469a <=( a22468a  and  a22463a );
 a22473a <=( A236  and  (not A233) );
 a22474a <=( A232  and  a22473a );
 a22478a <=( A269  and  A266 );
 a22479a <=( (not A265)  and  a22478a );
 a22480a <=( a22479a  and  a22474a );
 a22483a <=( (not A168)  and  (not A169) );
 a22487a <=( A202  and  A166 );
 a22488a <=( A167  and  a22487a );
 a22489a <=( a22488a  and  a22483a );
 a22493a <=( A236  and  (not A233) );
 a22494a <=( A232  and  a22493a );
 a22498a <=( A269  and  (not A266) );
 a22499a <=( A265  and  a22498a );
 a22500a <=( a22499a  and  a22494a );
 a22503a <=( (not A168)  and  (not A169) );
 a22507a <=( A199  and  A166 );
 a22508a <=( A167  and  a22507a );
 a22509a <=( a22508a  and  a22503a );
 a22513a <=( A298  and  A235 );
 a22514a <=( A201  and  a22513a );
 a22518a <=( (not A301)  and  (not A300) );
 a22519a <=( A299  and  a22518a );
 a22520a <=( a22519a  and  a22514a );
 a22523a <=( (not A168)  and  (not A169) );
 a22527a <=( A199  and  A166 );
 a22528a <=( A167  and  a22527a );
 a22529a <=( a22528a  and  a22523a );
 a22533a <=( A234  and  A232 );
 a22534a <=( A201  and  a22533a );
 a22538a <=( (not A302)  and  (not A301) );
 a22539a <=( (not A300)  and  a22538a );
 a22540a <=( a22539a  and  a22534a );
 a22543a <=( (not A168)  and  (not A169) );
 a22547a <=( A199  and  A166 );
 a22548a <=( A167  and  a22547a );
 a22549a <=( a22548a  and  a22543a );
 a22553a <=( A234  and  A232 );
 a22554a <=( A201  and  a22553a );
 a22558a <=( (not A301)  and  (not A299) );
 a22559a <=( (not A298)  and  a22558a );
 a22560a <=( a22559a  and  a22554a );
 a22563a <=( (not A168)  and  (not A169) );
 a22567a <=( A199  and  A166 );
 a22568a <=( A167  and  a22567a );
 a22569a <=( a22568a  and  a22563a );
 a22573a <=( A234  and  A232 );
 a22574a <=( A201  and  a22573a );
 a22578a <=( A269  and  A266 );
 a22579a <=( (not A265)  and  a22578a );
 a22580a <=( a22579a  and  a22574a );
 a22583a <=( (not A168)  and  (not A169) );
 a22587a <=( A199  and  A166 );
 a22588a <=( A167  and  a22587a );
 a22589a <=( a22588a  and  a22583a );
 a22593a <=( A234  and  A232 );
 a22594a <=( A201  and  a22593a );
 a22598a <=( A269  and  (not A266) );
 a22599a <=( A265  and  a22598a );
 a22600a <=( a22599a  and  a22594a );
 a22603a <=( (not A168)  and  (not A169) );
 a22607a <=( A199  and  A166 );
 a22608a <=( A167  and  a22607a );
 a22609a <=( a22608a  and  a22603a );
 a22613a <=( A234  and  A233 );
 a22614a <=( A201  and  a22613a );
 a22618a <=( (not A302)  and  (not A301) );
 a22619a <=( (not A300)  and  a22618a );
 a22620a <=( a22619a  and  a22614a );
 a22623a <=( (not A168)  and  (not A169) );
 a22627a <=( A199  and  A166 );
 a22628a <=( A167  and  a22627a );
 a22629a <=( a22628a  and  a22623a );
 a22633a <=( A234  and  A233 );
 a22634a <=( A201  and  a22633a );
 a22638a <=( (not A301)  and  (not A299) );
 a22639a <=( (not A298)  and  a22638a );
 a22640a <=( a22639a  and  a22634a );
 a22643a <=( (not A168)  and  (not A169) );
 a22647a <=( A199  and  A166 );
 a22648a <=( A167  and  a22647a );
 a22649a <=( a22648a  and  a22643a );
 a22653a <=( A234  and  A233 );
 a22654a <=( A201  and  a22653a );
 a22658a <=( A269  and  A266 );
 a22659a <=( (not A265)  and  a22658a );
 a22660a <=( a22659a  and  a22654a );
 a22663a <=( (not A168)  and  (not A169) );
 a22667a <=( A199  and  A166 );
 a22668a <=( A167  and  a22667a );
 a22669a <=( a22668a  and  a22663a );
 a22673a <=( A234  and  A233 );
 a22674a <=( A201  and  a22673a );
 a22678a <=( A269  and  (not A266) );
 a22679a <=( A265  and  a22678a );
 a22680a <=( a22679a  and  a22674a );
 a22683a <=( (not A168)  and  (not A169) );
 a22687a <=( A199  and  A166 );
 a22688a <=( A167  and  a22687a );
 a22689a <=( a22688a  and  a22683a );
 a22693a <=( A233  and  (not A232) );
 a22694a <=( A201  and  a22693a );
 a22698a <=( A267  and  A265 );
 a22699a <=( A236  and  a22698a );
 a22700a <=( a22699a  and  a22694a );
 a22703a <=( (not A168)  and  (not A169) );
 a22707a <=( A199  and  A166 );
 a22708a <=( A167  and  a22707a );
 a22709a <=( a22708a  and  a22703a );
 a22713a <=( A233  and  (not A232) );
 a22714a <=( A201  and  a22713a );
 a22718a <=( A267  and  A266 );
 a22719a <=( A236  and  a22718a );
 a22720a <=( a22719a  and  a22714a );
 a22723a <=( (not A168)  and  (not A169) );
 a22727a <=( A199  and  A166 );
 a22728a <=( A167  and  a22727a );
 a22729a <=( a22728a  and  a22723a );
 a22733a <=( (not A233)  and  A232 );
 a22734a <=( A201  and  a22733a );
 a22738a <=( A267  and  A265 );
 a22739a <=( A236  and  a22738a );
 a22740a <=( a22739a  and  a22734a );
 a22743a <=( (not A168)  and  (not A169) );
 a22747a <=( A199  and  A166 );
 a22748a <=( A167  and  a22747a );
 a22749a <=( a22748a  and  a22743a );
 a22753a <=( (not A233)  and  A232 );
 a22754a <=( A201  and  a22753a );
 a22758a <=( A267  and  A266 );
 a22759a <=( A236  and  a22758a );
 a22760a <=( a22759a  and  a22754a );
 a22763a <=( (not A168)  and  (not A169) );
 a22767a <=( A200  and  A166 );
 a22768a <=( A167  and  a22767a );
 a22769a <=( a22768a  and  a22763a );
 a22773a <=( A298  and  A235 );
 a22774a <=( A201  and  a22773a );
 a22778a <=( (not A301)  and  (not A300) );
 a22779a <=( A299  and  a22778a );
 a22780a <=( a22779a  and  a22774a );
 a22783a <=( (not A168)  and  (not A169) );
 a22787a <=( A200  and  A166 );
 a22788a <=( A167  and  a22787a );
 a22789a <=( a22788a  and  a22783a );
 a22793a <=( A234  and  A232 );
 a22794a <=( A201  and  a22793a );
 a22798a <=( (not A302)  and  (not A301) );
 a22799a <=( (not A300)  and  a22798a );
 a22800a <=( a22799a  and  a22794a );
 a22803a <=( (not A168)  and  (not A169) );
 a22807a <=( A200  and  A166 );
 a22808a <=( A167  and  a22807a );
 a22809a <=( a22808a  and  a22803a );
 a22813a <=( A234  and  A232 );
 a22814a <=( A201  and  a22813a );
 a22818a <=( (not A301)  and  (not A299) );
 a22819a <=( (not A298)  and  a22818a );
 a22820a <=( a22819a  and  a22814a );
 a22823a <=( (not A168)  and  (not A169) );
 a22827a <=( A200  and  A166 );
 a22828a <=( A167  and  a22827a );
 a22829a <=( a22828a  and  a22823a );
 a22833a <=( A234  and  A232 );
 a22834a <=( A201  and  a22833a );
 a22838a <=( A269  and  A266 );
 a22839a <=( (not A265)  and  a22838a );
 a22840a <=( a22839a  and  a22834a );
 a22843a <=( (not A168)  and  (not A169) );
 a22847a <=( A200  and  A166 );
 a22848a <=( A167  and  a22847a );
 a22849a <=( a22848a  and  a22843a );
 a22853a <=( A234  and  A232 );
 a22854a <=( A201  and  a22853a );
 a22858a <=( A269  and  (not A266) );
 a22859a <=( A265  and  a22858a );
 a22860a <=( a22859a  and  a22854a );
 a22863a <=( (not A168)  and  (not A169) );
 a22867a <=( A200  and  A166 );
 a22868a <=( A167  and  a22867a );
 a22869a <=( a22868a  and  a22863a );
 a22873a <=( A234  and  A233 );
 a22874a <=( A201  and  a22873a );
 a22878a <=( (not A302)  and  (not A301) );
 a22879a <=( (not A300)  and  a22878a );
 a22880a <=( a22879a  and  a22874a );
 a22883a <=( (not A168)  and  (not A169) );
 a22887a <=( A200  and  A166 );
 a22888a <=( A167  and  a22887a );
 a22889a <=( a22888a  and  a22883a );
 a22893a <=( A234  and  A233 );
 a22894a <=( A201  and  a22893a );
 a22898a <=( (not A301)  and  (not A299) );
 a22899a <=( (not A298)  and  a22898a );
 a22900a <=( a22899a  and  a22894a );
 a22903a <=( (not A168)  and  (not A169) );
 a22907a <=( A200  and  A166 );
 a22908a <=( A167  and  a22907a );
 a22909a <=( a22908a  and  a22903a );
 a22913a <=( A234  and  A233 );
 a22914a <=( A201  and  a22913a );
 a22918a <=( A269  and  A266 );
 a22919a <=( (not A265)  and  a22918a );
 a22920a <=( a22919a  and  a22914a );
 a22923a <=( (not A168)  and  (not A169) );
 a22927a <=( A200  and  A166 );
 a22928a <=( A167  and  a22927a );
 a22929a <=( a22928a  and  a22923a );
 a22933a <=( A234  and  A233 );
 a22934a <=( A201  and  a22933a );
 a22938a <=( A269  and  (not A266) );
 a22939a <=( A265  and  a22938a );
 a22940a <=( a22939a  and  a22934a );
 a22943a <=( (not A168)  and  (not A169) );
 a22947a <=( A200  and  A166 );
 a22948a <=( A167  and  a22947a );
 a22949a <=( a22948a  and  a22943a );
 a22953a <=( A233  and  (not A232) );
 a22954a <=( A201  and  a22953a );
 a22958a <=( A267  and  A265 );
 a22959a <=( A236  and  a22958a );
 a22960a <=( a22959a  and  a22954a );
 a22963a <=( (not A168)  and  (not A169) );
 a22967a <=( A200  and  A166 );
 a22968a <=( A167  and  a22967a );
 a22969a <=( a22968a  and  a22963a );
 a22973a <=( A233  and  (not A232) );
 a22974a <=( A201  and  a22973a );
 a22978a <=( A267  and  A266 );
 a22979a <=( A236  and  a22978a );
 a22980a <=( a22979a  and  a22974a );
 a22983a <=( (not A168)  and  (not A169) );
 a22987a <=( A200  and  A166 );
 a22988a <=( A167  and  a22987a );
 a22989a <=( a22988a  and  a22983a );
 a22993a <=( (not A233)  and  A232 );
 a22994a <=( A201  and  a22993a );
 a22998a <=( A267  and  A265 );
 a22999a <=( A236  and  a22998a );
 a23000a <=( a22999a  and  a22994a );
 a23003a <=( (not A168)  and  (not A169) );
 a23007a <=( A200  and  A166 );
 a23008a <=( A167  and  a23007a );
 a23009a <=( a23008a  and  a23003a );
 a23013a <=( (not A233)  and  A232 );
 a23014a <=( A201  and  a23013a );
 a23018a <=( A267  and  A266 );
 a23019a <=( A236  and  a23018a );
 a23020a <=( a23019a  and  a23014a );
 a23023a <=( (not A168)  and  (not A169) );
 a23027a <=( (not A199)  and  A166 );
 a23028a <=( A167  and  a23027a );
 a23029a <=( a23028a  and  a23023a );
 a23033a <=( A235  and  A203 );
 a23034a <=( A200  and  a23033a );
 a23038a <=( (not A302)  and  (not A301) );
 a23039a <=( (not A300)  and  a23038a );
 a23040a <=( a23039a  and  a23034a );
 a23043a <=( (not A168)  and  (not A169) );
 a23047a <=( (not A199)  and  A166 );
 a23048a <=( A167  and  a23047a );
 a23049a <=( a23048a  and  a23043a );
 a23053a <=( A235  and  A203 );
 a23054a <=( A200  and  a23053a );
 a23058a <=( (not A301)  and  (not A299) );
 a23059a <=( (not A298)  and  a23058a );
 a23060a <=( a23059a  and  a23054a );
 a23063a <=( (not A168)  and  (not A169) );
 a23067a <=( (not A199)  and  A166 );
 a23068a <=( A167  and  a23067a );
 a23069a <=( a23068a  and  a23063a );
 a23073a <=( A235  and  A203 );
 a23074a <=( A200  and  a23073a );
 a23078a <=( A269  and  A266 );
 a23079a <=( (not A265)  and  a23078a );
 a23080a <=( a23079a  and  a23074a );
 a23083a <=( (not A168)  and  (not A169) );
 a23087a <=( (not A199)  and  A166 );
 a23088a <=( A167  and  a23087a );
 a23089a <=( a23088a  and  a23083a );
 a23093a <=( A235  and  A203 );
 a23094a <=( A200  and  a23093a );
 a23098a <=( A269  and  (not A266) );
 a23099a <=( A265  and  a23098a );
 a23100a <=( a23099a  and  a23094a );
 a23103a <=( (not A168)  and  (not A169) );
 a23107a <=( (not A199)  and  A166 );
 a23108a <=( A167  and  a23107a );
 a23109a <=( a23108a  and  a23103a );
 a23113a <=( A232  and  A203 );
 a23114a <=( A200  and  a23113a );
 a23118a <=( A267  and  A265 );
 a23119a <=( A234  and  a23118a );
 a23120a <=( a23119a  and  a23114a );
 a23123a <=( (not A168)  and  (not A169) );
 a23127a <=( (not A199)  and  A166 );
 a23128a <=( A167  and  a23127a );
 a23129a <=( a23128a  and  a23123a );
 a23133a <=( A232  and  A203 );
 a23134a <=( A200  and  a23133a );
 a23138a <=( A267  and  A266 );
 a23139a <=( A234  and  a23138a );
 a23140a <=( a23139a  and  a23134a );
 a23143a <=( (not A168)  and  (not A169) );
 a23147a <=( (not A199)  and  A166 );
 a23148a <=( A167  and  a23147a );
 a23149a <=( a23148a  and  a23143a );
 a23153a <=( A233  and  A203 );
 a23154a <=( A200  and  a23153a );
 a23158a <=( A267  and  A265 );
 a23159a <=( A234  and  a23158a );
 a23160a <=( a23159a  and  a23154a );
 a23163a <=( (not A168)  and  (not A169) );
 a23167a <=( (not A199)  and  A166 );
 a23168a <=( A167  and  a23167a );
 a23169a <=( a23168a  and  a23163a );
 a23173a <=( A233  and  A203 );
 a23174a <=( A200  and  a23173a );
 a23178a <=( A267  and  A266 );
 a23179a <=( A234  and  a23178a );
 a23180a <=( a23179a  and  a23174a );
 a23183a <=( (not A168)  and  (not A169) );
 a23187a <=( (not A199)  and  A166 );
 a23188a <=( A167  and  a23187a );
 a23189a <=( a23188a  and  a23183a );
 a23193a <=( (not A232)  and  A203 );
 a23194a <=( A200  and  a23193a );
 a23198a <=( A268  and  A236 );
 a23199a <=( A233  and  a23198a );
 a23200a <=( a23199a  and  a23194a );
 a23203a <=( (not A168)  and  (not A169) );
 a23207a <=( (not A199)  and  A166 );
 a23208a <=( A167  and  a23207a );
 a23209a <=( a23208a  and  a23203a );
 a23213a <=( A232  and  A203 );
 a23214a <=( A200  and  a23213a );
 a23218a <=( A268  and  A236 );
 a23219a <=( (not A233)  and  a23218a );
 a23220a <=( a23219a  and  a23214a );
 a23223a <=( (not A168)  and  (not A169) );
 a23227a <=( A199  and  A166 );
 a23228a <=( A167  and  a23227a );
 a23229a <=( a23228a  and  a23223a );
 a23233a <=( A235  and  A203 );
 a23234a <=( (not A200)  and  a23233a );
 a23238a <=( (not A302)  and  (not A301) );
 a23239a <=( (not A300)  and  a23238a );
 a23240a <=( a23239a  and  a23234a );
 a23243a <=( (not A168)  and  (not A169) );
 a23247a <=( A199  and  A166 );
 a23248a <=( A167  and  a23247a );
 a23249a <=( a23248a  and  a23243a );
 a23253a <=( A235  and  A203 );
 a23254a <=( (not A200)  and  a23253a );
 a23258a <=( (not A301)  and  (not A299) );
 a23259a <=( (not A298)  and  a23258a );
 a23260a <=( a23259a  and  a23254a );
 a23263a <=( (not A168)  and  (not A169) );
 a23267a <=( A199  and  A166 );
 a23268a <=( A167  and  a23267a );
 a23269a <=( a23268a  and  a23263a );
 a23273a <=( A235  and  A203 );
 a23274a <=( (not A200)  and  a23273a );
 a23278a <=( A269  and  A266 );
 a23279a <=( (not A265)  and  a23278a );
 a23280a <=( a23279a  and  a23274a );
 a23283a <=( (not A168)  and  (not A169) );
 a23287a <=( A199  and  A166 );
 a23288a <=( A167  and  a23287a );
 a23289a <=( a23288a  and  a23283a );
 a23293a <=( A235  and  A203 );
 a23294a <=( (not A200)  and  a23293a );
 a23298a <=( A269  and  (not A266) );
 a23299a <=( A265  and  a23298a );
 a23300a <=( a23299a  and  a23294a );
 a23303a <=( (not A168)  and  (not A169) );
 a23307a <=( A199  and  A166 );
 a23308a <=( A167  and  a23307a );
 a23309a <=( a23308a  and  a23303a );
 a23313a <=( A232  and  A203 );
 a23314a <=( (not A200)  and  a23313a );
 a23318a <=( A267  and  A265 );
 a23319a <=( A234  and  a23318a );
 a23320a <=( a23319a  and  a23314a );
 a23323a <=( (not A168)  and  (not A169) );
 a23327a <=( A199  and  A166 );
 a23328a <=( A167  and  a23327a );
 a23329a <=( a23328a  and  a23323a );
 a23333a <=( A232  and  A203 );
 a23334a <=( (not A200)  and  a23333a );
 a23338a <=( A267  and  A266 );
 a23339a <=( A234  and  a23338a );
 a23340a <=( a23339a  and  a23334a );
 a23343a <=( (not A168)  and  (not A169) );
 a23347a <=( A199  and  A166 );
 a23348a <=( A167  and  a23347a );
 a23349a <=( a23348a  and  a23343a );
 a23353a <=( A233  and  A203 );
 a23354a <=( (not A200)  and  a23353a );
 a23358a <=( A267  and  A265 );
 a23359a <=( A234  and  a23358a );
 a23360a <=( a23359a  and  a23354a );
 a23363a <=( (not A168)  and  (not A169) );
 a23367a <=( A199  and  A166 );
 a23368a <=( A167  and  a23367a );
 a23369a <=( a23368a  and  a23363a );
 a23373a <=( A233  and  A203 );
 a23374a <=( (not A200)  and  a23373a );
 a23378a <=( A267  and  A266 );
 a23379a <=( A234  and  a23378a );
 a23380a <=( a23379a  and  a23374a );
 a23383a <=( (not A168)  and  (not A169) );
 a23387a <=( A199  and  A166 );
 a23388a <=( A167  and  a23387a );
 a23389a <=( a23388a  and  a23383a );
 a23393a <=( (not A232)  and  A203 );
 a23394a <=( (not A200)  and  a23393a );
 a23398a <=( A268  and  A236 );
 a23399a <=( A233  and  a23398a );
 a23400a <=( a23399a  and  a23394a );
 a23403a <=( (not A168)  and  (not A169) );
 a23407a <=( A199  and  A166 );
 a23408a <=( A167  and  a23407a );
 a23409a <=( a23408a  and  a23403a );
 a23413a <=( A232  and  A203 );
 a23414a <=( (not A200)  and  a23413a );
 a23418a <=( A268  and  A236 );
 a23419a <=( (not A233)  and  a23418a );
 a23420a <=( a23419a  and  a23414a );
 a23423a <=( (not A169)  and  (not A170) );
 a23427a <=( (not A234)  and  A202 );
 a23428a <=( (not A168)  and  a23427a );
 a23429a <=( a23428a  and  a23423a );
 a23433a <=( (not A267)  and  (not A236) );
 a23434a <=( (not A235)  and  a23433a );
 a23438a <=( A301  and  (not A269) );
 a23439a <=( (not A268)  and  a23438a );
 a23440a <=( a23439a  and  a23434a );
 a23443a <=( (not A169)  and  (not A170) );
 a23447a <=( (not A234)  and  A202 );
 a23448a <=( (not A168)  and  a23447a );
 a23449a <=( a23448a  and  a23443a );
 a23453a <=( (not A265)  and  (not A236) );
 a23454a <=( (not A235)  and  a23453a );
 a23458a <=( A301  and  (not A268) );
 a23459a <=( (not A266)  and  a23458a );
 a23460a <=( a23459a  and  a23454a );
 a23463a <=( (not A169)  and  (not A170) );
 a23467a <=( (not A232)  and  A202 );
 a23468a <=( (not A168)  and  a23467a );
 a23469a <=( a23468a  and  a23463a );
 a23473a <=( A298  and  A236 );
 a23474a <=( A233  and  a23473a );
 a23478a <=( (not A301)  and  (not A300) );
 a23479a <=( A299  and  a23478a );
 a23480a <=( a23479a  and  a23474a );
 a23483a <=( (not A169)  and  (not A170) );
 a23487a <=( A232  and  A202 );
 a23488a <=( (not A168)  and  a23487a );
 a23489a <=( a23488a  and  a23483a );
 a23493a <=( A298  and  A236 );
 a23494a <=( (not A233)  and  a23493a );
 a23498a <=( (not A301)  and  (not A300) );
 a23499a <=( A299  and  a23498a );
 a23500a <=( a23499a  and  a23494a );
 a23503a <=( (not A169)  and  (not A170) );
 a23507a <=( (not A232)  and  A202 );
 a23508a <=( (not A168)  and  a23507a );
 a23509a <=( a23508a  and  a23503a );
 a23513a <=( (not A267)  and  (not A235) );
 a23514a <=( (not A233)  and  a23513a );
 a23518a <=( A301  and  (not A269) );
 a23519a <=( (not A268)  and  a23518a );
 a23520a <=( a23519a  and  a23514a );
 a23523a <=( (not A169)  and  (not A170) );
 a23527a <=( (not A232)  and  A202 );
 a23528a <=( (not A168)  and  a23527a );
 a23529a <=( a23528a  and  a23523a );
 a23533a <=( (not A265)  and  (not A235) );
 a23534a <=( (not A233)  and  a23533a );
 a23538a <=( A301  and  (not A268) );
 a23539a <=( (not A266)  and  a23538a );
 a23540a <=( a23539a  and  a23534a );
 a23543a <=( (not A169)  and  (not A170) );
 a23547a <=( A201  and  A199 );
 a23548a <=( (not A168)  and  a23547a );
 a23549a <=( a23548a  and  a23543a );
 a23553a <=( A298  and  A234 );
 a23554a <=( A232  and  a23553a );
 a23558a <=( (not A301)  and  (not A300) );
 a23559a <=( A299  and  a23558a );
 a23560a <=( a23559a  and  a23554a );
 a23563a <=( (not A169)  and  (not A170) );
 a23567a <=( A201  and  A199 );
 a23568a <=( (not A168)  and  a23567a );
 a23569a <=( a23568a  and  a23563a );
 a23573a <=( A298  and  A234 );
 a23574a <=( A233  and  a23573a );
 a23578a <=( (not A301)  and  (not A300) );
 a23579a <=( A299  and  a23578a );
 a23580a <=( a23579a  and  a23574a );
 a23583a <=( (not A169)  and  (not A170) );
 a23587a <=( A201  and  A199 );
 a23588a <=( (not A168)  and  a23587a );
 a23589a <=( a23588a  and  a23583a );
 a23593a <=( A236  and  A233 );
 a23594a <=( (not A232)  and  a23593a );
 a23598a <=( (not A302)  and  (not A301) );
 a23599a <=( (not A300)  and  a23598a );
 a23600a <=( a23599a  and  a23594a );
 a23603a <=( (not A169)  and  (not A170) );
 a23607a <=( A201  and  A199 );
 a23608a <=( (not A168)  and  a23607a );
 a23609a <=( a23608a  and  a23603a );
 a23613a <=( A236  and  A233 );
 a23614a <=( (not A232)  and  a23613a );
 a23618a <=( (not A301)  and  (not A299) );
 a23619a <=( (not A298)  and  a23618a );
 a23620a <=( a23619a  and  a23614a );
 a23623a <=( (not A169)  and  (not A170) );
 a23627a <=( A201  and  A199 );
 a23628a <=( (not A168)  and  a23627a );
 a23629a <=( a23628a  and  a23623a );
 a23633a <=( A236  and  A233 );
 a23634a <=( (not A232)  and  a23633a );
 a23638a <=( A269  and  A266 );
 a23639a <=( (not A265)  and  a23638a );
 a23640a <=( a23639a  and  a23634a );
 a23643a <=( (not A169)  and  (not A170) );
 a23647a <=( A201  and  A199 );
 a23648a <=( (not A168)  and  a23647a );
 a23649a <=( a23648a  and  a23643a );
 a23653a <=( A236  and  A233 );
 a23654a <=( (not A232)  and  a23653a );
 a23658a <=( A269  and  (not A266) );
 a23659a <=( A265  and  a23658a );
 a23660a <=( a23659a  and  a23654a );
 a23663a <=( (not A169)  and  (not A170) );
 a23667a <=( A201  and  A199 );
 a23668a <=( (not A168)  and  a23667a );
 a23669a <=( a23668a  and  a23663a );
 a23673a <=( A236  and  (not A233) );
 a23674a <=( A232  and  a23673a );
 a23678a <=( (not A302)  and  (not A301) );
 a23679a <=( (not A300)  and  a23678a );
 a23680a <=( a23679a  and  a23674a );
 a23683a <=( (not A169)  and  (not A170) );
 a23687a <=( A201  and  A199 );
 a23688a <=( (not A168)  and  a23687a );
 a23689a <=( a23688a  and  a23683a );
 a23693a <=( A236  and  (not A233) );
 a23694a <=( A232  and  a23693a );
 a23698a <=( (not A301)  and  (not A299) );
 a23699a <=( (not A298)  and  a23698a );
 a23700a <=( a23699a  and  a23694a );
 a23703a <=( (not A169)  and  (not A170) );
 a23707a <=( A201  and  A199 );
 a23708a <=( (not A168)  and  a23707a );
 a23709a <=( a23708a  and  a23703a );
 a23713a <=( A236  and  (not A233) );
 a23714a <=( A232  and  a23713a );
 a23718a <=( A269  and  A266 );
 a23719a <=( (not A265)  and  a23718a );
 a23720a <=( a23719a  and  a23714a );
 a23723a <=( (not A169)  and  (not A170) );
 a23727a <=( A201  and  A199 );
 a23728a <=( (not A168)  and  a23727a );
 a23729a <=( a23728a  and  a23723a );
 a23733a <=( A236  and  (not A233) );
 a23734a <=( A232  and  a23733a );
 a23738a <=( A269  and  (not A266) );
 a23739a <=( A265  and  a23738a );
 a23740a <=( a23739a  and  a23734a );
 a23743a <=( (not A169)  and  (not A170) );
 a23747a <=( A201  and  A200 );
 a23748a <=( (not A168)  and  a23747a );
 a23749a <=( a23748a  and  a23743a );
 a23753a <=( A298  and  A234 );
 a23754a <=( A232  and  a23753a );
 a23758a <=( (not A301)  and  (not A300) );
 a23759a <=( A299  and  a23758a );
 a23760a <=( a23759a  and  a23754a );
 a23763a <=( (not A169)  and  (not A170) );
 a23767a <=( A201  and  A200 );
 a23768a <=( (not A168)  and  a23767a );
 a23769a <=( a23768a  and  a23763a );
 a23773a <=( A298  and  A234 );
 a23774a <=( A233  and  a23773a );
 a23778a <=( (not A301)  and  (not A300) );
 a23779a <=( A299  and  a23778a );
 a23780a <=( a23779a  and  a23774a );
 a23783a <=( (not A169)  and  (not A170) );
 a23787a <=( A201  and  A200 );
 a23788a <=( (not A168)  and  a23787a );
 a23789a <=( a23788a  and  a23783a );
 a23793a <=( A236  and  A233 );
 a23794a <=( (not A232)  and  a23793a );
 a23798a <=( (not A302)  and  (not A301) );
 a23799a <=( (not A300)  and  a23798a );
 a23800a <=( a23799a  and  a23794a );
 a23803a <=( (not A169)  and  (not A170) );
 a23807a <=( A201  and  A200 );
 a23808a <=( (not A168)  and  a23807a );
 a23809a <=( a23808a  and  a23803a );
 a23813a <=( A236  and  A233 );
 a23814a <=( (not A232)  and  a23813a );
 a23818a <=( (not A301)  and  (not A299) );
 a23819a <=( (not A298)  and  a23818a );
 a23820a <=( a23819a  and  a23814a );
 a23823a <=( (not A169)  and  (not A170) );
 a23827a <=( A201  and  A200 );
 a23828a <=( (not A168)  and  a23827a );
 a23829a <=( a23828a  and  a23823a );
 a23833a <=( A236  and  A233 );
 a23834a <=( (not A232)  and  a23833a );
 a23838a <=( A269  and  A266 );
 a23839a <=( (not A265)  and  a23838a );
 a23840a <=( a23839a  and  a23834a );
 a23843a <=( (not A169)  and  (not A170) );
 a23847a <=( A201  and  A200 );
 a23848a <=( (not A168)  and  a23847a );
 a23849a <=( a23848a  and  a23843a );
 a23853a <=( A236  and  A233 );
 a23854a <=( (not A232)  and  a23853a );
 a23858a <=( A269  and  (not A266) );
 a23859a <=( A265  and  a23858a );
 a23860a <=( a23859a  and  a23854a );
 a23863a <=( (not A169)  and  (not A170) );
 a23867a <=( A201  and  A200 );
 a23868a <=( (not A168)  and  a23867a );
 a23869a <=( a23868a  and  a23863a );
 a23873a <=( A236  and  (not A233) );
 a23874a <=( A232  and  a23873a );
 a23878a <=( (not A302)  and  (not A301) );
 a23879a <=( (not A300)  and  a23878a );
 a23880a <=( a23879a  and  a23874a );
 a23883a <=( (not A169)  and  (not A170) );
 a23887a <=( A201  and  A200 );
 a23888a <=( (not A168)  and  a23887a );
 a23889a <=( a23888a  and  a23883a );
 a23893a <=( A236  and  (not A233) );
 a23894a <=( A232  and  a23893a );
 a23898a <=( (not A301)  and  (not A299) );
 a23899a <=( (not A298)  and  a23898a );
 a23900a <=( a23899a  and  a23894a );
 a23903a <=( (not A169)  and  (not A170) );
 a23907a <=( A201  and  A200 );
 a23908a <=( (not A168)  and  a23907a );
 a23909a <=( a23908a  and  a23903a );
 a23913a <=( A236  and  (not A233) );
 a23914a <=( A232  and  a23913a );
 a23918a <=( A269  and  A266 );
 a23919a <=( (not A265)  and  a23918a );
 a23920a <=( a23919a  and  a23914a );
 a23923a <=( (not A169)  and  (not A170) );
 a23927a <=( A201  and  A200 );
 a23928a <=( (not A168)  and  a23927a );
 a23929a <=( a23928a  and  a23923a );
 a23933a <=( A236  and  (not A233) );
 a23934a <=( A232  and  a23933a );
 a23938a <=( A269  and  (not A266) );
 a23939a <=( A265  and  a23938a );
 a23940a <=( a23939a  and  a23934a );
 a23943a <=( (not A169)  and  (not A170) );
 a23947a <=( A200  and  (not A199) );
 a23948a <=( (not A168)  and  a23947a );
 a23949a <=( a23948a  and  a23943a );
 a23953a <=( A298  and  A235 );
 a23954a <=( A203  and  a23953a );
 a23958a <=( (not A301)  and  (not A300) );
 a23959a <=( A299  and  a23958a );
 a23960a <=( a23959a  and  a23954a );
 a23963a <=( (not A169)  and  (not A170) );
 a23967a <=( A200  and  (not A199) );
 a23968a <=( (not A168)  and  a23967a );
 a23969a <=( a23968a  and  a23963a );
 a23973a <=( A234  and  A232 );
 a23974a <=( A203  and  a23973a );
 a23978a <=( (not A302)  and  (not A301) );
 a23979a <=( (not A300)  and  a23978a );
 a23980a <=( a23979a  and  a23974a );
 a23983a <=( (not A169)  and  (not A170) );
 a23987a <=( A200  and  (not A199) );
 a23988a <=( (not A168)  and  a23987a );
 a23989a <=( a23988a  and  a23983a );
 a23993a <=( A234  and  A232 );
 a23994a <=( A203  and  a23993a );
 a23998a <=( (not A301)  and  (not A299) );
 a23999a <=( (not A298)  and  a23998a );
 a24000a <=( a23999a  and  a23994a );
 a24003a <=( (not A169)  and  (not A170) );
 a24007a <=( A200  and  (not A199) );
 a24008a <=( (not A168)  and  a24007a );
 a24009a <=( a24008a  and  a24003a );
 a24013a <=( A234  and  A232 );
 a24014a <=( A203  and  a24013a );
 a24018a <=( A269  and  A266 );
 a24019a <=( (not A265)  and  a24018a );
 a24020a <=( a24019a  and  a24014a );
 a24023a <=( (not A169)  and  (not A170) );
 a24027a <=( A200  and  (not A199) );
 a24028a <=( (not A168)  and  a24027a );
 a24029a <=( a24028a  and  a24023a );
 a24033a <=( A234  and  A232 );
 a24034a <=( A203  and  a24033a );
 a24038a <=( A269  and  (not A266) );
 a24039a <=( A265  and  a24038a );
 a24040a <=( a24039a  and  a24034a );
 a24043a <=( (not A169)  and  (not A170) );
 a24047a <=( A200  and  (not A199) );
 a24048a <=( (not A168)  and  a24047a );
 a24049a <=( a24048a  and  a24043a );
 a24053a <=( A234  and  A233 );
 a24054a <=( A203  and  a24053a );
 a24058a <=( (not A302)  and  (not A301) );
 a24059a <=( (not A300)  and  a24058a );
 a24060a <=( a24059a  and  a24054a );
 a24063a <=( (not A169)  and  (not A170) );
 a24067a <=( A200  and  (not A199) );
 a24068a <=( (not A168)  and  a24067a );
 a24069a <=( a24068a  and  a24063a );
 a24073a <=( A234  and  A233 );
 a24074a <=( A203  and  a24073a );
 a24078a <=( (not A301)  and  (not A299) );
 a24079a <=( (not A298)  and  a24078a );
 a24080a <=( a24079a  and  a24074a );
 a24083a <=( (not A169)  and  (not A170) );
 a24087a <=( A200  and  (not A199) );
 a24088a <=( (not A168)  and  a24087a );
 a24089a <=( a24088a  and  a24083a );
 a24093a <=( A234  and  A233 );
 a24094a <=( A203  and  a24093a );
 a24098a <=( A269  and  A266 );
 a24099a <=( (not A265)  and  a24098a );
 a24100a <=( a24099a  and  a24094a );
 a24103a <=( (not A169)  and  (not A170) );
 a24107a <=( A200  and  (not A199) );
 a24108a <=( (not A168)  and  a24107a );
 a24109a <=( a24108a  and  a24103a );
 a24113a <=( A234  and  A233 );
 a24114a <=( A203  and  a24113a );
 a24118a <=( A269  and  (not A266) );
 a24119a <=( A265  and  a24118a );
 a24120a <=( a24119a  and  a24114a );
 a24123a <=( (not A169)  and  (not A170) );
 a24127a <=( A200  and  (not A199) );
 a24128a <=( (not A168)  and  a24127a );
 a24129a <=( a24128a  and  a24123a );
 a24133a <=( A233  and  (not A232) );
 a24134a <=( A203  and  a24133a );
 a24138a <=( A267  and  A265 );
 a24139a <=( A236  and  a24138a );
 a24140a <=( a24139a  and  a24134a );
 a24143a <=( (not A169)  and  (not A170) );
 a24147a <=( A200  and  (not A199) );
 a24148a <=( (not A168)  and  a24147a );
 a24149a <=( a24148a  and  a24143a );
 a24153a <=( A233  and  (not A232) );
 a24154a <=( A203  and  a24153a );
 a24158a <=( A267  and  A266 );
 a24159a <=( A236  and  a24158a );
 a24160a <=( a24159a  and  a24154a );
 a24163a <=( (not A169)  and  (not A170) );
 a24167a <=( A200  and  (not A199) );
 a24168a <=( (not A168)  and  a24167a );
 a24169a <=( a24168a  and  a24163a );
 a24173a <=( (not A233)  and  A232 );
 a24174a <=( A203  and  a24173a );
 a24178a <=( A267  and  A265 );
 a24179a <=( A236  and  a24178a );
 a24180a <=( a24179a  and  a24174a );
 a24183a <=( (not A169)  and  (not A170) );
 a24187a <=( A200  and  (not A199) );
 a24188a <=( (not A168)  and  a24187a );
 a24189a <=( a24188a  and  a24183a );
 a24193a <=( (not A233)  and  A232 );
 a24194a <=( A203  and  a24193a );
 a24198a <=( A267  and  A266 );
 a24199a <=( A236  and  a24198a );
 a24200a <=( a24199a  and  a24194a );
 a24203a <=( (not A169)  and  (not A170) );
 a24207a <=( (not A200)  and  A199 );
 a24208a <=( (not A168)  and  a24207a );
 a24209a <=( a24208a  and  a24203a );
 a24213a <=( A298  and  A235 );
 a24214a <=( A203  and  a24213a );
 a24218a <=( (not A301)  and  (not A300) );
 a24219a <=( A299  and  a24218a );
 a24220a <=( a24219a  and  a24214a );
 a24223a <=( (not A169)  and  (not A170) );
 a24227a <=( (not A200)  and  A199 );
 a24228a <=( (not A168)  and  a24227a );
 a24229a <=( a24228a  and  a24223a );
 a24233a <=( A234  and  A232 );
 a24234a <=( A203  and  a24233a );
 a24238a <=( (not A302)  and  (not A301) );
 a24239a <=( (not A300)  and  a24238a );
 a24240a <=( a24239a  and  a24234a );
 a24243a <=( (not A169)  and  (not A170) );
 a24247a <=( (not A200)  and  A199 );
 a24248a <=( (not A168)  and  a24247a );
 a24249a <=( a24248a  and  a24243a );
 a24253a <=( A234  and  A232 );
 a24254a <=( A203  and  a24253a );
 a24258a <=( (not A301)  and  (not A299) );
 a24259a <=( (not A298)  and  a24258a );
 a24260a <=( a24259a  and  a24254a );
 a24263a <=( (not A169)  and  (not A170) );
 a24267a <=( (not A200)  and  A199 );
 a24268a <=( (not A168)  and  a24267a );
 a24269a <=( a24268a  and  a24263a );
 a24273a <=( A234  and  A232 );
 a24274a <=( A203  and  a24273a );
 a24278a <=( A269  and  A266 );
 a24279a <=( (not A265)  and  a24278a );
 a24280a <=( a24279a  and  a24274a );
 a24283a <=( (not A169)  and  (not A170) );
 a24287a <=( (not A200)  and  A199 );
 a24288a <=( (not A168)  and  a24287a );
 a24289a <=( a24288a  and  a24283a );
 a24293a <=( A234  and  A232 );
 a24294a <=( A203  and  a24293a );
 a24298a <=( A269  and  (not A266) );
 a24299a <=( A265  and  a24298a );
 a24300a <=( a24299a  and  a24294a );
 a24303a <=( (not A169)  and  (not A170) );
 a24307a <=( (not A200)  and  A199 );
 a24308a <=( (not A168)  and  a24307a );
 a24309a <=( a24308a  and  a24303a );
 a24313a <=( A234  and  A233 );
 a24314a <=( A203  and  a24313a );
 a24318a <=( (not A302)  and  (not A301) );
 a24319a <=( (not A300)  and  a24318a );
 a24320a <=( a24319a  and  a24314a );
 a24323a <=( (not A169)  and  (not A170) );
 a24327a <=( (not A200)  and  A199 );
 a24328a <=( (not A168)  and  a24327a );
 a24329a <=( a24328a  and  a24323a );
 a24333a <=( A234  and  A233 );
 a24334a <=( A203  and  a24333a );
 a24338a <=( (not A301)  and  (not A299) );
 a24339a <=( (not A298)  and  a24338a );
 a24340a <=( a24339a  and  a24334a );
 a24343a <=( (not A169)  and  (not A170) );
 a24347a <=( (not A200)  and  A199 );
 a24348a <=( (not A168)  and  a24347a );
 a24349a <=( a24348a  and  a24343a );
 a24353a <=( A234  and  A233 );
 a24354a <=( A203  and  a24353a );
 a24358a <=( A269  and  A266 );
 a24359a <=( (not A265)  and  a24358a );
 a24360a <=( a24359a  and  a24354a );
 a24363a <=( (not A169)  and  (not A170) );
 a24367a <=( (not A200)  and  A199 );
 a24368a <=( (not A168)  and  a24367a );
 a24369a <=( a24368a  and  a24363a );
 a24373a <=( A234  and  A233 );
 a24374a <=( A203  and  a24373a );
 a24378a <=( A269  and  (not A266) );
 a24379a <=( A265  and  a24378a );
 a24380a <=( a24379a  and  a24374a );
 a24383a <=( (not A169)  and  (not A170) );
 a24387a <=( (not A200)  and  A199 );
 a24388a <=( (not A168)  and  a24387a );
 a24389a <=( a24388a  and  a24383a );
 a24393a <=( A233  and  (not A232) );
 a24394a <=( A203  and  a24393a );
 a24398a <=( A267  and  A265 );
 a24399a <=( A236  and  a24398a );
 a24400a <=( a24399a  and  a24394a );
 a24403a <=( (not A169)  and  (not A170) );
 a24407a <=( (not A200)  and  A199 );
 a24408a <=( (not A168)  and  a24407a );
 a24409a <=( a24408a  and  a24403a );
 a24413a <=( A233  and  (not A232) );
 a24414a <=( A203  and  a24413a );
 a24418a <=( A267  and  A266 );
 a24419a <=( A236  and  a24418a );
 a24420a <=( a24419a  and  a24414a );
 a24423a <=( (not A169)  and  (not A170) );
 a24427a <=( (not A200)  and  A199 );
 a24428a <=( (not A168)  and  a24427a );
 a24429a <=( a24428a  and  a24423a );
 a24433a <=( (not A233)  and  A232 );
 a24434a <=( A203  and  a24433a );
 a24438a <=( A267  and  A265 );
 a24439a <=( A236  and  a24438a );
 a24440a <=( a24439a  and  a24434a );
 a24443a <=( (not A169)  and  (not A170) );
 a24447a <=( (not A200)  and  A199 );
 a24448a <=( (not A168)  and  a24447a );
 a24449a <=( a24448a  and  a24443a );
 a24453a <=( (not A233)  and  A232 );
 a24454a <=( A203  and  a24453a );
 a24458a <=( A267  and  A266 );
 a24459a <=( A236  and  a24458a );
 a24460a <=( a24459a  and  a24454a );
 a24464a <=( (not A201)  and  A166 );
 a24465a <=( A168  and  a24464a );
 a24469a <=( (not A234)  and  (not A203) );
 a24470a <=( (not A202)  and  a24469a );
 a24471a <=( a24470a  and  a24465a );
 a24475a <=( (not A267)  and  (not A236) );
 a24476a <=( (not A235)  and  a24475a );
 a24480a <=( A301  and  (not A269) );
 a24481a <=( (not A268)  and  a24480a );
 a24482a <=( a24481a  and  a24476a );
 a24486a <=( (not A201)  and  A166 );
 a24487a <=( A168  and  a24486a );
 a24491a <=( (not A234)  and  (not A203) );
 a24492a <=( (not A202)  and  a24491a );
 a24493a <=( a24492a  and  a24487a );
 a24497a <=( (not A265)  and  (not A236) );
 a24498a <=( (not A235)  and  a24497a );
 a24502a <=( A301  and  (not A268) );
 a24503a <=( (not A266)  and  a24502a );
 a24504a <=( a24503a  and  a24498a );
 a24508a <=( (not A201)  and  A166 );
 a24509a <=( A168  and  a24508a );
 a24513a <=( (not A232)  and  (not A203) );
 a24514a <=( (not A202)  and  a24513a );
 a24515a <=( a24514a  and  a24509a );
 a24519a <=( A298  and  A236 );
 a24520a <=( A233  and  a24519a );
 a24524a <=( (not A301)  and  (not A300) );
 a24525a <=( A299  and  a24524a );
 a24526a <=( a24525a  and  a24520a );
 a24530a <=( (not A201)  and  A166 );
 a24531a <=( A168  and  a24530a );
 a24535a <=( A232  and  (not A203) );
 a24536a <=( (not A202)  and  a24535a );
 a24537a <=( a24536a  and  a24531a );
 a24541a <=( A298  and  A236 );
 a24542a <=( (not A233)  and  a24541a );
 a24546a <=( (not A301)  and  (not A300) );
 a24547a <=( A299  and  a24546a );
 a24548a <=( a24547a  and  a24542a );
 a24552a <=( (not A201)  and  A166 );
 a24553a <=( A168  and  a24552a );
 a24557a <=( (not A232)  and  (not A203) );
 a24558a <=( (not A202)  and  a24557a );
 a24559a <=( a24558a  and  a24553a );
 a24563a <=( (not A267)  and  (not A235) );
 a24564a <=( (not A233)  and  a24563a );
 a24568a <=( A301  and  (not A269) );
 a24569a <=( (not A268)  and  a24568a );
 a24570a <=( a24569a  and  a24564a );
 a24574a <=( (not A201)  and  A166 );
 a24575a <=( A168  and  a24574a );
 a24579a <=( (not A232)  and  (not A203) );
 a24580a <=( (not A202)  and  a24579a );
 a24581a <=( a24580a  and  a24575a );
 a24585a <=( (not A265)  and  (not A235) );
 a24586a <=( (not A233)  and  a24585a );
 a24590a <=( A301  and  (not A268) );
 a24591a <=( (not A266)  and  a24590a );
 a24592a <=( a24591a  and  a24586a );
 a24596a <=( A199  and  A166 );
 a24597a <=( A168  and  a24596a );
 a24601a <=( (not A202)  and  (not A201) );
 a24602a <=( A200  and  a24601a );
 a24603a <=( a24602a  and  a24597a );
 a24607a <=( A298  and  A234 );
 a24608a <=( A232  and  a24607a );
 a24612a <=( (not A301)  and  (not A300) );
 a24613a <=( A299  and  a24612a );
 a24614a <=( a24613a  and  a24608a );
 a24618a <=( A199  and  A166 );
 a24619a <=( A168  and  a24618a );
 a24623a <=( (not A202)  and  (not A201) );
 a24624a <=( A200  and  a24623a );
 a24625a <=( a24624a  and  a24619a );
 a24629a <=( A298  and  A234 );
 a24630a <=( A233  and  a24629a );
 a24634a <=( (not A301)  and  (not A300) );
 a24635a <=( A299  and  a24634a );
 a24636a <=( a24635a  and  a24630a );
 a24640a <=( A199  and  A166 );
 a24641a <=( A168  and  a24640a );
 a24645a <=( (not A202)  and  (not A201) );
 a24646a <=( A200  and  a24645a );
 a24647a <=( a24646a  and  a24641a );
 a24651a <=( A236  and  A233 );
 a24652a <=( (not A232)  and  a24651a );
 a24656a <=( (not A302)  and  (not A301) );
 a24657a <=( (not A300)  and  a24656a );
 a24658a <=( a24657a  and  a24652a );
 a24662a <=( A199  and  A166 );
 a24663a <=( A168  and  a24662a );
 a24667a <=( (not A202)  and  (not A201) );
 a24668a <=( A200  and  a24667a );
 a24669a <=( a24668a  and  a24663a );
 a24673a <=( A236  and  A233 );
 a24674a <=( (not A232)  and  a24673a );
 a24678a <=( (not A301)  and  (not A299) );
 a24679a <=( (not A298)  and  a24678a );
 a24680a <=( a24679a  and  a24674a );
 a24684a <=( A199  and  A166 );
 a24685a <=( A168  and  a24684a );
 a24689a <=( (not A202)  and  (not A201) );
 a24690a <=( A200  and  a24689a );
 a24691a <=( a24690a  and  a24685a );
 a24695a <=( A236  and  A233 );
 a24696a <=( (not A232)  and  a24695a );
 a24700a <=( A269  and  A266 );
 a24701a <=( (not A265)  and  a24700a );
 a24702a <=( a24701a  and  a24696a );
 a24706a <=( A199  and  A166 );
 a24707a <=( A168  and  a24706a );
 a24711a <=( (not A202)  and  (not A201) );
 a24712a <=( A200  and  a24711a );
 a24713a <=( a24712a  and  a24707a );
 a24717a <=( A236  and  A233 );
 a24718a <=( (not A232)  and  a24717a );
 a24722a <=( A269  and  (not A266) );
 a24723a <=( A265  and  a24722a );
 a24724a <=( a24723a  and  a24718a );
 a24728a <=( A199  and  A166 );
 a24729a <=( A168  and  a24728a );
 a24733a <=( (not A202)  and  (not A201) );
 a24734a <=( A200  and  a24733a );
 a24735a <=( a24734a  and  a24729a );
 a24739a <=( A236  and  (not A233) );
 a24740a <=( A232  and  a24739a );
 a24744a <=( (not A302)  and  (not A301) );
 a24745a <=( (not A300)  and  a24744a );
 a24746a <=( a24745a  and  a24740a );
 a24750a <=( A199  and  A166 );
 a24751a <=( A168  and  a24750a );
 a24755a <=( (not A202)  and  (not A201) );
 a24756a <=( A200  and  a24755a );
 a24757a <=( a24756a  and  a24751a );
 a24761a <=( A236  and  (not A233) );
 a24762a <=( A232  and  a24761a );
 a24766a <=( (not A301)  and  (not A299) );
 a24767a <=( (not A298)  and  a24766a );
 a24768a <=( a24767a  and  a24762a );
 a24772a <=( A199  and  A166 );
 a24773a <=( A168  and  a24772a );
 a24777a <=( (not A202)  and  (not A201) );
 a24778a <=( A200  and  a24777a );
 a24779a <=( a24778a  and  a24773a );
 a24783a <=( A236  and  (not A233) );
 a24784a <=( A232  and  a24783a );
 a24788a <=( A269  and  A266 );
 a24789a <=( (not A265)  and  a24788a );
 a24790a <=( a24789a  and  a24784a );
 a24794a <=( A199  and  A166 );
 a24795a <=( A168  and  a24794a );
 a24799a <=( (not A202)  and  (not A201) );
 a24800a <=( A200  and  a24799a );
 a24801a <=( a24800a  and  a24795a );
 a24805a <=( A236  and  (not A233) );
 a24806a <=( A232  and  a24805a );
 a24810a <=( A269  and  (not A266) );
 a24811a <=( A265  and  a24810a );
 a24812a <=( a24811a  and  a24806a );
 a24816a <=( (not A199)  and  A166 );
 a24817a <=( A168  and  a24816a );
 a24821a <=( (not A234)  and  (not A202) );
 a24822a <=( (not A200)  and  a24821a );
 a24823a <=( a24822a  and  a24817a );
 a24827a <=( (not A267)  and  (not A236) );
 a24828a <=( (not A235)  and  a24827a );
 a24832a <=( A301  and  (not A269) );
 a24833a <=( (not A268)  and  a24832a );
 a24834a <=( a24833a  and  a24828a );
 a24838a <=( (not A199)  and  A166 );
 a24839a <=( A168  and  a24838a );
 a24843a <=( (not A234)  and  (not A202) );
 a24844a <=( (not A200)  and  a24843a );
 a24845a <=( a24844a  and  a24839a );
 a24849a <=( (not A265)  and  (not A236) );
 a24850a <=( (not A235)  and  a24849a );
 a24854a <=( A301  and  (not A268) );
 a24855a <=( (not A266)  and  a24854a );
 a24856a <=( a24855a  and  a24850a );
 a24860a <=( (not A199)  and  A166 );
 a24861a <=( A168  and  a24860a );
 a24865a <=( (not A232)  and  (not A202) );
 a24866a <=( (not A200)  and  a24865a );
 a24867a <=( a24866a  and  a24861a );
 a24871a <=( A298  and  A236 );
 a24872a <=( A233  and  a24871a );
 a24876a <=( (not A301)  and  (not A300) );
 a24877a <=( A299  and  a24876a );
 a24878a <=( a24877a  and  a24872a );
 a24882a <=( (not A199)  and  A166 );
 a24883a <=( A168  and  a24882a );
 a24887a <=( A232  and  (not A202) );
 a24888a <=( (not A200)  and  a24887a );
 a24889a <=( a24888a  and  a24883a );
 a24893a <=( A298  and  A236 );
 a24894a <=( (not A233)  and  a24893a );
 a24898a <=( (not A301)  and  (not A300) );
 a24899a <=( A299  and  a24898a );
 a24900a <=( a24899a  and  a24894a );
 a24904a <=( (not A199)  and  A166 );
 a24905a <=( A168  and  a24904a );
 a24909a <=( (not A232)  and  (not A202) );
 a24910a <=( (not A200)  and  a24909a );
 a24911a <=( a24910a  and  a24905a );
 a24915a <=( (not A267)  and  (not A235) );
 a24916a <=( (not A233)  and  a24915a );
 a24920a <=( A301  and  (not A269) );
 a24921a <=( (not A268)  and  a24920a );
 a24922a <=( a24921a  and  a24916a );
 a24926a <=( (not A199)  and  A166 );
 a24927a <=( A168  and  a24926a );
 a24931a <=( (not A232)  and  (not A202) );
 a24932a <=( (not A200)  and  a24931a );
 a24933a <=( a24932a  and  a24927a );
 a24937a <=( (not A265)  and  (not A235) );
 a24938a <=( (not A233)  and  a24937a );
 a24942a <=( A301  and  (not A268) );
 a24943a <=( (not A266)  and  a24942a );
 a24944a <=( a24943a  and  a24938a );
 a24948a <=( (not A201)  and  A167 );
 a24949a <=( A168  and  a24948a );
 a24953a <=( (not A234)  and  (not A203) );
 a24954a <=( (not A202)  and  a24953a );
 a24955a <=( a24954a  and  a24949a );
 a24959a <=( (not A267)  and  (not A236) );
 a24960a <=( (not A235)  and  a24959a );
 a24964a <=( A301  and  (not A269) );
 a24965a <=( (not A268)  and  a24964a );
 a24966a <=( a24965a  and  a24960a );
 a24970a <=( (not A201)  and  A167 );
 a24971a <=( A168  and  a24970a );
 a24975a <=( (not A234)  and  (not A203) );
 a24976a <=( (not A202)  and  a24975a );
 a24977a <=( a24976a  and  a24971a );
 a24981a <=( (not A265)  and  (not A236) );
 a24982a <=( (not A235)  and  a24981a );
 a24986a <=( A301  and  (not A268) );
 a24987a <=( (not A266)  and  a24986a );
 a24988a <=( a24987a  and  a24982a );
 a24992a <=( (not A201)  and  A167 );
 a24993a <=( A168  and  a24992a );
 a24997a <=( (not A232)  and  (not A203) );
 a24998a <=( (not A202)  and  a24997a );
 a24999a <=( a24998a  and  a24993a );
 a25003a <=( A298  and  A236 );
 a25004a <=( A233  and  a25003a );
 a25008a <=( (not A301)  and  (not A300) );
 a25009a <=( A299  and  a25008a );
 a25010a <=( a25009a  and  a25004a );
 a25014a <=( (not A201)  and  A167 );
 a25015a <=( A168  and  a25014a );
 a25019a <=( A232  and  (not A203) );
 a25020a <=( (not A202)  and  a25019a );
 a25021a <=( a25020a  and  a25015a );
 a25025a <=( A298  and  A236 );
 a25026a <=( (not A233)  and  a25025a );
 a25030a <=( (not A301)  and  (not A300) );
 a25031a <=( A299  and  a25030a );
 a25032a <=( a25031a  and  a25026a );
 a25036a <=( (not A201)  and  A167 );
 a25037a <=( A168  and  a25036a );
 a25041a <=( (not A232)  and  (not A203) );
 a25042a <=( (not A202)  and  a25041a );
 a25043a <=( a25042a  and  a25037a );
 a25047a <=( (not A267)  and  (not A235) );
 a25048a <=( (not A233)  and  a25047a );
 a25052a <=( A301  and  (not A269) );
 a25053a <=( (not A268)  and  a25052a );
 a25054a <=( a25053a  and  a25048a );
 a25058a <=( (not A201)  and  A167 );
 a25059a <=( A168  and  a25058a );
 a25063a <=( (not A232)  and  (not A203) );
 a25064a <=( (not A202)  and  a25063a );
 a25065a <=( a25064a  and  a25059a );
 a25069a <=( (not A265)  and  (not A235) );
 a25070a <=( (not A233)  and  a25069a );
 a25074a <=( A301  and  (not A268) );
 a25075a <=( (not A266)  and  a25074a );
 a25076a <=( a25075a  and  a25070a );
 a25080a <=( A199  and  A167 );
 a25081a <=( A168  and  a25080a );
 a25085a <=( (not A202)  and  (not A201) );
 a25086a <=( A200  and  a25085a );
 a25087a <=( a25086a  and  a25081a );
 a25091a <=( A298  and  A234 );
 a25092a <=( A232  and  a25091a );
 a25096a <=( (not A301)  and  (not A300) );
 a25097a <=( A299  and  a25096a );
 a25098a <=( a25097a  and  a25092a );
 a25102a <=( A199  and  A167 );
 a25103a <=( A168  and  a25102a );
 a25107a <=( (not A202)  and  (not A201) );
 a25108a <=( A200  and  a25107a );
 a25109a <=( a25108a  and  a25103a );
 a25113a <=( A298  and  A234 );
 a25114a <=( A233  and  a25113a );
 a25118a <=( (not A301)  and  (not A300) );
 a25119a <=( A299  and  a25118a );
 a25120a <=( a25119a  and  a25114a );
 a25124a <=( A199  and  A167 );
 a25125a <=( A168  and  a25124a );
 a25129a <=( (not A202)  and  (not A201) );
 a25130a <=( A200  and  a25129a );
 a25131a <=( a25130a  and  a25125a );
 a25135a <=( A236  and  A233 );
 a25136a <=( (not A232)  and  a25135a );
 a25140a <=( (not A302)  and  (not A301) );
 a25141a <=( (not A300)  and  a25140a );
 a25142a <=( a25141a  and  a25136a );
 a25146a <=( A199  and  A167 );
 a25147a <=( A168  and  a25146a );
 a25151a <=( (not A202)  and  (not A201) );
 a25152a <=( A200  and  a25151a );
 a25153a <=( a25152a  and  a25147a );
 a25157a <=( A236  and  A233 );
 a25158a <=( (not A232)  and  a25157a );
 a25162a <=( (not A301)  and  (not A299) );
 a25163a <=( (not A298)  and  a25162a );
 a25164a <=( a25163a  and  a25158a );
 a25168a <=( A199  and  A167 );
 a25169a <=( A168  and  a25168a );
 a25173a <=( (not A202)  and  (not A201) );
 a25174a <=( A200  and  a25173a );
 a25175a <=( a25174a  and  a25169a );
 a25179a <=( A236  and  A233 );
 a25180a <=( (not A232)  and  a25179a );
 a25184a <=( A269  and  A266 );
 a25185a <=( (not A265)  and  a25184a );
 a25186a <=( a25185a  and  a25180a );
 a25190a <=( A199  and  A167 );
 a25191a <=( A168  and  a25190a );
 a25195a <=( (not A202)  and  (not A201) );
 a25196a <=( A200  and  a25195a );
 a25197a <=( a25196a  and  a25191a );
 a25201a <=( A236  and  A233 );
 a25202a <=( (not A232)  and  a25201a );
 a25206a <=( A269  and  (not A266) );
 a25207a <=( A265  and  a25206a );
 a25208a <=( a25207a  and  a25202a );
 a25212a <=( A199  and  A167 );
 a25213a <=( A168  and  a25212a );
 a25217a <=( (not A202)  and  (not A201) );
 a25218a <=( A200  and  a25217a );
 a25219a <=( a25218a  and  a25213a );
 a25223a <=( A236  and  (not A233) );
 a25224a <=( A232  and  a25223a );
 a25228a <=( (not A302)  and  (not A301) );
 a25229a <=( (not A300)  and  a25228a );
 a25230a <=( a25229a  and  a25224a );
 a25234a <=( A199  and  A167 );
 a25235a <=( A168  and  a25234a );
 a25239a <=( (not A202)  and  (not A201) );
 a25240a <=( A200  and  a25239a );
 a25241a <=( a25240a  and  a25235a );
 a25245a <=( A236  and  (not A233) );
 a25246a <=( A232  and  a25245a );
 a25250a <=( (not A301)  and  (not A299) );
 a25251a <=( (not A298)  and  a25250a );
 a25252a <=( a25251a  and  a25246a );
 a25256a <=( A199  and  A167 );
 a25257a <=( A168  and  a25256a );
 a25261a <=( (not A202)  and  (not A201) );
 a25262a <=( A200  and  a25261a );
 a25263a <=( a25262a  and  a25257a );
 a25267a <=( A236  and  (not A233) );
 a25268a <=( A232  and  a25267a );
 a25272a <=( A269  and  A266 );
 a25273a <=( (not A265)  and  a25272a );
 a25274a <=( a25273a  and  a25268a );
 a25278a <=( A199  and  A167 );
 a25279a <=( A168  and  a25278a );
 a25283a <=( (not A202)  and  (not A201) );
 a25284a <=( A200  and  a25283a );
 a25285a <=( a25284a  and  a25279a );
 a25289a <=( A236  and  (not A233) );
 a25290a <=( A232  and  a25289a );
 a25294a <=( A269  and  (not A266) );
 a25295a <=( A265  and  a25294a );
 a25296a <=( a25295a  and  a25290a );
 a25300a <=( (not A199)  and  A167 );
 a25301a <=( A168  and  a25300a );
 a25305a <=( (not A234)  and  (not A202) );
 a25306a <=( (not A200)  and  a25305a );
 a25307a <=( a25306a  and  a25301a );
 a25311a <=( (not A267)  and  (not A236) );
 a25312a <=( (not A235)  and  a25311a );
 a25316a <=( A301  and  (not A269) );
 a25317a <=( (not A268)  and  a25316a );
 a25318a <=( a25317a  and  a25312a );
 a25322a <=( (not A199)  and  A167 );
 a25323a <=( A168  and  a25322a );
 a25327a <=( (not A234)  and  (not A202) );
 a25328a <=( (not A200)  and  a25327a );
 a25329a <=( a25328a  and  a25323a );
 a25333a <=( (not A265)  and  (not A236) );
 a25334a <=( (not A235)  and  a25333a );
 a25338a <=( A301  and  (not A268) );
 a25339a <=( (not A266)  and  a25338a );
 a25340a <=( a25339a  and  a25334a );
 a25344a <=( (not A199)  and  A167 );
 a25345a <=( A168  and  a25344a );
 a25349a <=( (not A232)  and  (not A202) );
 a25350a <=( (not A200)  and  a25349a );
 a25351a <=( a25350a  and  a25345a );
 a25355a <=( A298  and  A236 );
 a25356a <=( A233  and  a25355a );
 a25360a <=( (not A301)  and  (not A300) );
 a25361a <=( A299  and  a25360a );
 a25362a <=( a25361a  and  a25356a );
 a25366a <=( (not A199)  and  A167 );
 a25367a <=( A168  and  a25366a );
 a25371a <=( A232  and  (not A202) );
 a25372a <=( (not A200)  and  a25371a );
 a25373a <=( a25372a  and  a25367a );
 a25377a <=( A298  and  A236 );
 a25378a <=( (not A233)  and  a25377a );
 a25382a <=( (not A301)  and  (not A300) );
 a25383a <=( A299  and  a25382a );
 a25384a <=( a25383a  and  a25378a );
 a25388a <=( (not A199)  and  A167 );
 a25389a <=( A168  and  a25388a );
 a25393a <=( (not A232)  and  (not A202) );
 a25394a <=( (not A200)  and  a25393a );
 a25395a <=( a25394a  and  a25389a );
 a25399a <=( (not A267)  and  (not A235) );
 a25400a <=( (not A233)  and  a25399a );
 a25404a <=( A301  and  (not A269) );
 a25405a <=( (not A268)  and  a25404a );
 a25406a <=( a25405a  and  a25400a );
 a25410a <=( (not A199)  and  A167 );
 a25411a <=( A168  and  a25410a );
 a25415a <=( (not A232)  and  (not A202) );
 a25416a <=( (not A200)  and  a25415a );
 a25417a <=( a25416a  and  a25411a );
 a25421a <=( (not A265)  and  (not A235) );
 a25422a <=( (not A233)  and  a25421a );
 a25426a <=( A301  and  (not A268) );
 a25427a <=( (not A266)  and  a25426a );
 a25428a <=( a25427a  and  a25422a );
 a25432a <=( (not A166)  and  A167 );
 a25433a <=( A170  and  a25432a );
 a25437a <=( (not A203)  and  (not A202) );
 a25438a <=( (not A201)  and  a25437a );
 a25439a <=( a25438a  and  a25433a );
 a25443a <=( A298  and  A234 );
 a25444a <=( A232  and  a25443a );
 a25448a <=( (not A301)  and  (not A300) );
 a25449a <=( A299  and  a25448a );
 a25450a <=( a25449a  and  a25444a );
 a25454a <=( (not A166)  and  A167 );
 a25455a <=( A170  and  a25454a );
 a25459a <=( (not A203)  and  (not A202) );
 a25460a <=( (not A201)  and  a25459a );
 a25461a <=( a25460a  and  a25455a );
 a25465a <=( A298  and  A234 );
 a25466a <=( A233  and  a25465a );
 a25470a <=( (not A301)  and  (not A300) );
 a25471a <=( A299  and  a25470a );
 a25472a <=( a25471a  and  a25466a );
 a25476a <=( (not A166)  and  A167 );
 a25477a <=( A170  and  a25476a );
 a25481a <=( (not A203)  and  (not A202) );
 a25482a <=( (not A201)  and  a25481a );
 a25483a <=( a25482a  and  a25477a );
 a25487a <=( A236  and  A233 );
 a25488a <=( (not A232)  and  a25487a );
 a25492a <=( (not A302)  and  (not A301) );
 a25493a <=( (not A300)  and  a25492a );
 a25494a <=( a25493a  and  a25488a );
 a25498a <=( (not A166)  and  A167 );
 a25499a <=( A170  and  a25498a );
 a25503a <=( (not A203)  and  (not A202) );
 a25504a <=( (not A201)  and  a25503a );
 a25505a <=( a25504a  and  a25499a );
 a25509a <=( A236  and  A233 );
 a25510a <=( (not A232)  and  a25509a );
 a25514a <=( (not A301)  and  (not A299) );
 a25515a <=( (not A298)  and  a25514a );
 a25516a <=( a25515a  and  a25510a );
 a25520a <=( (not A166)  and  A167 );
 a25521a <=( A170  and  a25520a );
 a25525a <=( (not A203)  and  (not A202) );
 a25526a <=( (not A201)  and  a25525a );
 a25527a <=( a25526a  and  a25521a );
 a25531a <=( A236  and  A233 );
 a25532a <=( (not A232)  and  a25531a );
 a25536a <=( A269  and  A266 );
 a25537a <=( (not A265)  and  a25536a );
 a25538a <=( a25537a  and  a25532a );
 a25542a <=( (not A166)  and  A167 );
 a25543a <=( A170  and  a25542a );
 a25547a <=( (not A203)  and  (not A202) );
 a25548a <=( (not A201)  and  a25547a );
 a25549a <=( a25548a  and  a25543a );
 a25553a <=( A236  and  A233 );
 a25554a <=( (not A232)  and  a25553a );
 a25558a <=( A269  and  (not A266) );
 a25559a <=( A265  and  a25558a );
 a25560a <=( a25559a  and  a25554a );
 a25564a <=( (not A166)  and  A167 );
 a25565a <=( A170  and  a25564a );
 a25569a <=( (not A203)  and  (not A202) );
 a25570a <=( (not A201)  and  a25569a );
 a25571a <=( a25570a  and  a25565a );
 a25575a <=( A236  and  (not A233) );
 a25576a <=( A232  and  a25575a );
 a25580a <=( (not A302)  and  (not A301) );
 a25581a <=( (not A300)  and  a25580a );
 a25582a <=( a25581a  and  a25576a );
 a25586a <=( (not A166)  and  A167 );
 a25587a <=( A170  and  a25586a );
 a25591a <=( (not A203)  and  (not A202) );
 a25592a <=( (not A201)  and  a25591a );
 a25593a <=( a25592a  and  a25587a );
 a25597a <=( A236  and  (not A233) );
 a25598a <=( A232  and  a25597a );
 a25602a <=( (not A301)  and  (not A299) );
 a25603a <=( (not A298)  and  a25602a );
 a25604a <=( a25603a  and  a25598a );
 a25608a <=( (not A166)  and  A167 );
 a25609a <=( A170  and  a25608a );
 a25613a <=( (not A203)  and  (not A202) );
 a25614a <=( (not A201)  and  a25613a );
 a25615a <=( a25614a  and  a25609a );
 a25619a <=( A236  and  (not A233) );
 a25620a <=( A232  and  a25619a );
 a25624a <=( A269  and  A266 );
 a25625a <=( (not A265)  and  a25624a );
 a25626a <=( a25625a  and  a25620a );
 a25630a <=( (not A166)  and  A167 );
 a25631a <=( A170  and  a25630a );
 a25635a <=( (not A203)  and  (not A202) );
 a25636a <=( (not A201)  and  a25635a );
 a25637a <=( a25636a  and  a25631a );
 a25641a <=( A236  and  (not A233) );
 a25642a <=( A232  and  a25641a );
 a25646a <=( A269  and  (not A266) );
 a25647a <=( A265  and  a25646a );
 a25648a <=( a25647a  and  a25642a );
 a25652a <=( (not A166)  and  A167 );
 a25653a <=( A170  and  a25652a );
 a25657a <=( (not A201)  and  A200 );
 a25658a <=( A199  and  a25657a );
 a25659a <=( a25658a  and  a25653a );
 a25663a <=( A298  and  A235 );
 a25664a <=( (not A202)  and  a25663a );
 a25668a <=( (not A301)  and  (not A300) );
 a25669a <=( A299  and  a25668a );
 a25670a <=( a25669a  and  a25664a );
 a25674a <=( (not A166)  and  A167 );
 a25675a <=( A170  and  a25674a );
 a25679a <=( (not A201)  and  A200 );
 a25680a <=( A199  and  a25679a );
 a25681a <=( a25680a  and  a25675a );
 a25685a <=( A234  and  A232 );
 a25686a <=( (not A202)  and  a25685a );
 a25690a <=( (not A302)  and  (not A301) );
 a25691a <=( (not A300)  and  a25690a );
 a25692a <=( a25691a  and  a25686a );
 a25696a <=( (not A166)  and  A167 );
 a25697a <=( A170  and  a25696a );
 a25701a <=( (not A201)  and  A200 );
 a25702a <=( A199  and  a25701a );
 a25703a <=( a25702a  and  a25697a );
 a25707a <=( A234  and  A232 );
 a25708a <=( (not A202)  and  a25707a );
 a25712a <=( (not A301)  and  (not A299) );
 a25713a <=( (not A298)  and  a25712a );
 a25714a <=( a25713a  and  a25708a );
 a25718a <=( (not A166)  and  A167 );
 a25719a <=( A170  and  a25718a );
 a25723a <=( (not A201)  and  A200 );
 a25724a <=( A199  and  a25723a );
 a25725a <=( a25724a  and  a25719a );
 a25729a <=( A234  and  A232 );
 a25730a <=( (not A202)  and  a25729a );
 a25734a <=( A269  and  A266 );
 a25735a <=( (not A265)  and  a25734a );
 a25736a <=( a25735a  and  a25730a );
 a25740a <=( (not A166)  and  A167 );
 a25741a <=( A170  and  a25740a );
 a25745a <=( (not A201)  and  A200 );
 a25746a <=( A199  and  a25745a );
 a25747a <=( a25746a  and  a25741a );
 a25751a <=( A234  and  A232 );
 a25752a <=( (not A202)  and  a25751a );
 a25756a <=( A269  and  (not A266) );
 a25757a <=( A265  and  a25756a );
 a25758a <=( a25757a  and  a25752a );
 a25762a <=( (not A166)  and  A167 );
 a25763a <=( A170  and  a25762a );
 a25767a <=( (not A201)  and  A200 );
 a25768a <=( A199  and  a25767a );
 a25769a <=( a25768a  and  a25763a );
 a25773a <=( A234  and  A233 );
 a25774a <=( (not A202)  and  a25773a );
 a25778a <=( (not A302)  and  (not A301) );
 a25779a <=( (not A300)  and  a25778a );
 a25780a <=( a25779a  and  a25774a );
 a25784a <=( (not A166)  and  A167 );
 a25785a <=( A170  and  a25784a );
 a25789a <=( (not A201)  and  A200 );
 a25790a <=( A199  and  a25789a );
 a25791a <=( a25790a  and  a25785a );
 a25795a <=( A234  and  A233 );
 a25796a <=( (not A202)  and  a25795a );
 a25800a <=( (not A301)  and  (not A299) );
 a25801a <=( (not A298)  and  a25800a );
 a25802a <=( a25801a  and  a25796a );
 a25806a <=( (not A166)  and  A167 );
 a25807a <=( A170  and  a25806a );
 a25811a <=( (not A201)  and  A200 );
 a25812a <=( A199  and  a25811a );
 a25813a <=( a25812a  and  a25807a );
 a25817a <=( A234  and  A233 );
 a25818a <=( (not A202)  and  a25817a );
 a25822a <=( A269  and  A266 );
 a25823a <=( (not A265)  and  a25822a );
 a25824a <=( a25823a  and  a25818a );
 a25828a <=( (not A166)  and  A167 );
 a25829a <=( A170  and  a25828a );
 a25833a <=( (not A201)  and  A200 );
 a25834a <=( A199  and  a25833a );
 a25835a <=( a25834a  and  a25829a );
 a25839a <=( A234  and  A233 );
 a25840a <=( (not A202)  and  a25839a );
 a25844a <=( A269  and  (not A266) );
 a25845a <=( A265  and  a25844a );
 a25846a <=( a25845a  and  a25840a );
 a25850a <=( (not A166)  and  A167 );
 a25851a <=( A170  and  a25850a );
 a25855a <=( (not A201)  and  A200 );
 a25856a <=( A199  and  a25855a );
 a25857a <=( a25856a  and  a25851a );
 a25861a <=( A233  and  (not A232) );
 a25862a <=( (not A202)  and  a25861a );
 a25866a <=( A267  and  A265 );
 a25867a <=( A236  and  a25866a );
 a25868a <=( a25867a  and  a25862a );
 a25872a <=( (not A166)  and  A167 );
 a25873a <=( A170  and  a25872a );
 a25877a <=( (not A201)  and  A200 );
 a25878a <=( A199  and  a25877a );
 a25879a <=( a25878a  and  a25873a );
 a25883a <=( A233  and  (not A232) );
 a25884a <=( (not A202)  and  a25883a );
 a25888a <=( A267  and  A266 );
 a25889a <=( A236  and  a25888a );
 a25890a <=( a25889a  and  a25884a );
 a25894a <=( (not A166)  and  A167 );
 a25895a <=( A170  and  a25894a );
 a25899a <=( (not A201)  and  A200 );
 a25900a <=( A199  and  a25899a );
 a25901a <=( a25900a  and  a25895a );
 a25905a <=( (not A233)  and  A232 );
 a25906a <=( (not A202)  and  a25905a );
 a25910a <=( A267  and  A265 );
 a25911a <=( A236  and  a25910a );
 a25912a <=( a25911a  and  a25906a );
 a25916a <=( (not A166)  and  A167 );
 a25917a <=( A170  and  a25916a );
 a25921a <=( (not A201)  and  A200 );
 a25922a <=( A199  and  a25921a );
 a25923a <=( a25922a  and  a25917a );
 a25927a <=( (not A233)  and  A232 );
 a25928a <=( (not A202)  and  a25927a );
 a25932a <=( A267  and  A266 );
 a25933a <=( A236  and  a25932a );
 a25934a <=( a25933a  and  a25928a );
 a25938a <=( (not A166)  and  A167 );
 a25939a <=( A170  and  a25938a );
 a25943a <=( (not A202)  and  (not A200) );
 a25944a <=( (not A199)  and  a25943a );
 a25945a <=( a25944a  and  a25939a );
 a25949a <=( A298  and  A234 );
 a25950a <=( A232  and  a25949a );
 a25954a <=( (not A301)  and  (not A300) );
 a25955a <=( A299  and  a25954a );
 a25956a <=( a25955a  and  a25950a );
 a25960a <=( (not A166)  and  A167 );
 a25961a <=( A170  and  a25960a );
 a25965a <=( (not A202)  and  (not A200) );
 a25966a <=( (not A199)  and  a25965a );
 a25967a <=( a25966a  and  a25961a );
 a25971a <=( A298  and  A234 );
 a25972a <=( A233  and  a25971a );
 a25976a <=( (not A301)  and  (not A300) );
 a25977a <=( A299  and  a25976a );
 a25978a <=( a25977a  and  a25972a );
 a25982a <=( (not A166)  and  A167 );
 a25983a <=( A170  and  a25982a );
 a25987a <=( (not A202)  and  (not A200) );
 a25988a <=( (not A199)  and  a25987a );
 a25989a <=( a25988a  and  a25983a );
 a25993a <=( A236  and  A233 );
 a25994a <=( (not A232)  and  a25993a );
 a25998a <=( (not A302)  and  (not A301) );
 a25999a <=( (not A300)  and  a25998a );
 a26000a <=( a25999a  and  a25994a );
 a26004a <=( (not A166)  and  A167 );
 a26005a <=( A170  and  a26004a );
 a26009a <=( (not A202)  and  (not A200) );
 a26010a <=( (not A199)  and  a26009a );
 a26011a <=( a26010a  and  a26005a );
 a26015a <=( A236  and  A233 );
 a26016a <=( (not A232)  and  a26015a );
 a26020a <=( (not A301)  and  (not A299) );
 a26021a <=( (not A298)  and  a26020a );
 a26022a <=( a26021a  and  a26016a );
 a26026a <=( (not A166)  and  A167 );
 a26027a <=( A170  and  a26026a );
 a26031a <=( (not A202)  and  (not A200) );
 a26032a <=( (not A199)  and  a26031a );
 a26033a <=( a26032a  and  a26027a );
 a26037a <=( A236  and  A233 );
 a26038a <=( (not A232)  and  a26037a );
 a26042a <=( A269  and  A266 );
 a26043a <=( (not A265)  and  a26042a );
 a26044a <=( a26043a  and  a26038a );
 a26048a <=( (not A166)  and  A167 );
 a26049a <=( A170  and  a26048a );
 a26053a <=( (not A202)  and  (not A200) );
 a26054a <=( (not A199)  and  a26053a );
 a26055a <=( a26054a  and  a26049a );
 a26059a <=( A236  and  A233 );
 a26060a <=( (not A232)  and  a26059a );
 a26064a <=( A269  and  (not A266) );
 a26065a <=( A265  and  a26064a );
 a26066a <=( a26065a  and  a26060a );
 a26070a <=( (not A166)  and  A167 );
 a26071a <=( A170  and  a26070a );
 a26075a <=( (not A202)  and  (not A200) );
 a26076a <=( (not A199)  and  a26075a );
 a26077a <=( a26076a  and  a26071a );
 a26081a <=( A236  and  (not A233) );
 a26082a <=( A232  and  a26081a );
 a26086a <=( (not A302)  and  (not A301) );
 a26087a <=( (not A300)  and  a26086a );
 a26088a <=( a26087a  and  a26082a );
 a26092a <=( (not A166)  and  A167 );
 a26093a <=( A170  and  a26092a );
 a26097a <=( (not A202)  and  (not A200) );
 a26098a <=( (not A199)  and  a26097a );
 a26099a <=( a26098a  and  a26093a );
 a26103a <=( A236  and  (not A233) );
 a26104a <=( A232  and  a26103a );
 a26108a <=( (not A301)  and  (not A299) );
 a26109a <=( (not A298)  and  a26108a );
 a26110a <=( a26109a  and  a26104a );
 a26114a <=( (not A166)  and  A167 );
 a26115a <=( A170  and  a26114a );
 a26119a <=( (not A202)  and  (not A200) );
 a26120a <=( (not A199)  and  a26119a );
 a26121a <=( a26120a  and  a26115a );
 a26125a <=( A236  and  (not A233) );
 a26126a <=( A232  and  a26125a );
 a26130a <=( A269  and  A266 );
 a26131a <=( (not A265)  and  a26130a );
 a26132a <=( a26131a  and  a26126a );
 a26136a <=( (not A166)  and  A167 );
 a26137a <=( A170  and  a26136a );
 a26141a <=( (not A202)  and  (not A200) );
 a26142a <=( (not A199)  and  a26141a );
 a26143a <=( a26142a  and  a26137a );
 a26147a <=( A236  and  (not A233) );
 a26148a <=( A232  and  a26147a );
 a26152a <=( A269  and  (not A266) );
 a26153a <=( A265  and  a26152a );
 a26154a <=( a26153a  and  a26148a );
 a26158a <=( A166  and  (not A167) );
 a26159a <=( A170  and  a26158a );
 a26163a <=( (not A203)  and  (not A202) );
 a26164a <=( (not A201)  and  a26163a );
 a26165a <=( a26164a  and  a26159a );
 a26169a <=( A298  and  A234 );
 a26170a <=( A232  and  a26169a );
 a26174a <=( (not A301)  and  (not A300) );
 a26175a <=( A299  and  a26174a );
 a26176a <=( a26175a  and  a26170a );
 a26180a <=( A166  and  (not A167) );
 a26181a <=( A170  and  a26180a );
 a26185a <=( (not A203)  and  (not A202) );
 a26186a <=( (not A201)  and  a26185a );
 a26187a <=( a26186a  and  a26181a );
 a26191a <=( A298  and  A234 );
 a26192a <=( A233  and  a26191a );
 a26196a <=( (not A301)  and  (not A300) );
 a26197a <=( A299  and  a26196a );
 a26198a <=( a26197a  and  a26192a );
 a26202a <=( A166  and  (not A167) );
 a26203a <=( A170  and  a26202a );
 a26207a <=( (not A203)  and  (not A202) );
 a26208a <=( (not A201)  and  a26207a );
 a26209a <=( a26208a  and  a26203a );
 a26213a <=( A236  and  A233 );
 a26214a <=( (not A232)  and  a26213a );
 a26218a <=( (not A302)  and  (not A301) );
 a26219a <=( (not A300)  and  a26218a );
 a26220a <=( a26219a  and  a26214a );
 a26224a <=( A166  and  (not A167) );
 a26225a <=( A170  and  a26224a );
 a26229a <=( (not A203)  and  (not A202) );
 a26230a <=( (not A201)  and  a26229a );
 a26231a <=( a26230a  and  a26225a );
 a26235a <=( A236  and  A233 );
 a26236a <=( (not A232)  and  a26235a );
 a26240a <=( (not A301)  and  (not A299) );
 a26241a <=( (not A298)  and  a26240a );
 a26242a <=( a26241a  and  a26236a );
 a26246a <=( A166  and  (not A167) );
 a26247a <=( A170  and  a26246a );
 a26251a <=( (not A203)  and  (not A202) );
 a26252a <=( (not A201)  and  a26251a );
 a26253a <=( a26252a  and  a26247a );
 a26257a <=( A236  and  A233 );
 a26258a <=( (not A232)  and  a26257a );
 a26262a <=( A269  and  A266 );
 a26263a <=( (not A265)  and  a26262a );
 a26264a <=( a26263a  and  a26258a );
 a26268a <=( A166  and  (not A167) );
 a26269a <=( A170  and  a26268a );
 a26273a <=( (not A203)  and  (not A202) );
 a26274a <=( (not A201)  and  a26273a );
 a26275a <=( a26274a  and  a26269a );
 a26279a <=( A236  and  A233 );
 a26280a <=( (not A232)  and  a26279a );
 a26284a <=( A269  and  (not A266) );
 a26285a <=( A265  and  a26284a );
 a26286a <=( a26285a  and  a26280a );
 a26290a <=( A166  and  (not A167) );
 a26291a <=( A170  and  a26290a );
 a26295a <=( (not A203)  and  (not A202) );
 a26296a <=( (not A201)  and  a26295a );
 a26297a <=( a26296a  and  a26291a );
 a26301a <=( A236  and  (not A233) );
 a26302a <=( A232  and  a26301a );
 a26306a <=( (not A302)  and  (not A301) );
 a26307a <=( (not A300)  and  a26306a );
 a26308a <=( a26307a  and  a26302a );
 a26312a <=( A166  and  (not A167) );
 a26313a <=( A170  and  a26312a );
 a26317a <=( (not A203)  and  (not A202) );
 a26318a <=( (not A201)  and  a26317a );
 a26319a <=( a26318a  and  a26313a );
 a26323a <=( A236  and  (not A233) );
 a26324a <=( A232  and  a26323a );
 a26328a <=( (not A301)  and  (not A299) );
 a26329a <=( (not A298)  and  a26328a );
 a26330a <=( a26329a  and  a26324a );
 a26334a <=( A166  and  (not A167) );
 a26335a <=( A170  and  a26334a );
 a26339a <=( (not A203)  and  (not A202) );
 a26340a <=( (not A201)  and  a26339a );
 a26341a <=( a26340a  and  a26335a );
 a26345a <=( A236  and  (not A233) );
 a26346a <=( A232  and  a26345a );
 a26350a <=( A269  and  A266 );
 a26351a <=( (not A265)  and  a26350a );
 a26352a <=( a26351a  and  a26346a );
 a26356a <=( A166  and  (not A167) );
 a26357a <=( A170  and  a26356a );
 a26361a <=( (not A203)  and  (not A202) );
 a26362a <=( (not A201)  and  a26361a );
 a26363a <=( a26362a  and  a26357a );
 a26367a <=( A236  and  (not A233) );
 a26368a <=( A232  and  a26367a );
 a26372a <=( A269  and  (not A266) );
 a26373a <=( A265  and  a26372a );
 a26374a <=( a26373a  and  a26368a );
 a26378a <=( A166  and  (not A167) );
 a26379a <=( A170  and  a26378a );
 a26383a <=( (not A201)  and  A200 );
 a26384a <=( A199  and  a26383a );
 a26385a <=( a26384a  and  a26379a );
 a26389a <=( A298  and  A235 );
 a26390a <=( (not A202)  and  a26389a );
 a26394a <=( (not A301)  and  (not A300) );
 a26395a <=( A299  and  a26394a );
 a26396a <=( a26395a  and  a26390a );
 a26400a <=( A166  and  (not A167) );
 a26401a <=( A170  and  a26400a );
 a26405a <=( (not A201)  and  A200 );
 a26406a <=( A199  and  a26405a );
 a26407a <=( a26406a  and  a26401a );
 a26411a <=( A234  and  A232 );
 a26412a <=( (not A202)  and  a26411a );
 a26416a <=( (not A302)  and  (not A301) );
 a26417a <=( (not A300)  and  a26416a );
 a26418a <=( a26417a  and  a26412a );
 a26422a <=( A166  and  (not A167) );
 a26423a <=( A170  and  a26422a );
 a26427a <=( (not A201)  and  A200 );
 a26428a <=( A199  and  a26427a );
 a26429a <=( a26428a  and  a26423a );
 a26433a <=( A234  and  A232 );
 a26434a <=( (not A202)  and  a26433a );
 a26438a <=( (not A301)  and  (not A299) );
 a26439a <=( (not A298)  and  a26438a );
 a26440a <=( a26439a  and  a26434a );
 a26444a <=( A166  and  (not A167) );
 a26445a <=( A170  and  a26444a );
 a26449a <=( (not A201)  and  A200 );
 a26450a <=( A199  and  a26449a );
 a26451a <=( a26450a  and  a26445a );
 a26455a <=( A234  and  A232 );
 a26456a <=( (not A202)  and  a26455a );
 a26460a <=( A269  and  A266 );
 a26461a <=( (not A265)  and  a26460a );
 a26462a <=( a26461a  and  a26456a );
 a26466a <=( A166  and  (not A167) );
 a26467a <=( A170  and  a26466a );
 a26471a <=( (not A201)  and  A200 );
 a26472a <=( A199  and  a26471a );
 a26473a <=( a26472a  and  a26467a );
 a26477a <=( A234  and  A232 );
 a26478a <=( (not A202)  and  a26477a );
 a26482a <=( A269  and  (not A266) );
 a26483a <=( A265  and  a26482a );
 a26484a <=( a26483a  and  a26478a );
 a26488a <=( A166  and  (not A167) );
 a26489a <=( A170  and  a26488a );
 a26493a <=( (not A201)  and  A200 );
 a26494a <=( A199  and  a26493a );
 a26495a <=( a26494a  and  a26489a );
 a26499a <=( A234  and  A233 );
 a26500a <=( (not A202)  and  a26499a );
 a26504a <=( (not A302)  and  (not A301) );
 a26505a <=( (not A300)  and  a26504a );
 a26506a <=( a26505a  and  a26500a );
 a26510a <=( A166  and  (not A167) );
 a26511a <=( A170  and  a26510a );
 a26515a <=( (not A201)  and  A200 );
 a26516a <=( A199  and  a26515a );
 a26517a <=( a26516a  and  a26511a );
 a26521a <=( A234  and  A233 );
 a26522a <=( (not A202)  and  a26521a );
 a26526a <=( (not A301)  and  (not A299) );
 a26527a <=( (not A298)  and  a26526a );
 a26528a <=( a26527a  and  a26522a );
 a26532a <=( A166  and  (not A167) );
 a26533a <=( A170  and  a26532a );
 a26537a <=( (not A201)  and  A200 );
 a26538a <=( A199  and  a26537a );
 a26539a <=( a26538a  and  a26533a );
 a26543a <=( A234  and  A233 );
 a26544a <=( (not A202)  and  a26543a );
 a26548a <=( A269  and  A266 );
 a26549a <=( (not A265)  and  a26548a );
 a26550a <=( a26549a  and  a26544a );
 a26554a <=( A166  and  (not A167) );
 a26555a <=( A170  and  a26554a );
 a26559a <=( (not A201)  and  A200 );
 a26560a <=( A199  and  a26559a );
 a26561a <=( a26560a  and  a26555a );
 a26565a <=( A234  and  A233 );
 a26566a <=( (not A202)  and  a26565a );
 a26570a <=( A269  and  (not A266) );
 a26571a <=( A265  and  a26570a );
 a26572a <=( a26571a  and  a26566a );
 a26576a <=( A166  and  (not A167) );
 a26577a <=( A170  and  a26576a );
 a26581a <=( (not A201)  and  A200 );
 a26582a <=( A199  and  a26581a );
 a26583a <=( a26582a  and  a26577a );
 a26587a <=( A233  and  (not A232) );
 a26588a <=( (not A202)  and  a26587a );
 a26592a <=( A267  and  A265 );
 a26593a <=( A236  and  a26592a );
 a26594a <=( a26593a  and  a26588a );
 a26598a <=( A166  and  (not A167) );
 a26599a <=( A170  and  a26598a );
 a26603a <=( (not A201)  and  A200 );
 a26604a <=( A199  and  a26603a );
 a26605a <=( a26604a  and  a26599a );
 a26609a <=( A233  and  (not A232) );
 a26610a <=( (not A202)  and  a26609a );
 a26614a <=( A267  and  A266 );
 a26615a <=( A236  and  a26614a );
 a26616a <=( a26615a  and  a26610a );
 a26620a <=( A166  and  (not A167) );
 a26621a <=( A170  and  a26620a );
 a26625a <=( (not A201)  and  A200 );
 a26626a <=( A199  and  a26625a );
 a26627a <=( a26626a  and  a26621a );
 a26631a <=( (not A233)  and  A232 );
 a26632a <=( (not A202)  and  a26631a );
 a26636a <=( A267  and  A265 );
 a26637a <=( A236  and  a26636a );
 a26638a <=( a26637a  and  a26632a );
 a26642a <=( A166  and  (not A167) );
 a26643a <=( A170  and  a26642a );
 a26647a <=( (not A201)  and  A200 );
 a26648a <=( A199  and  a26647a );
 a26649a <=( a26648a  and  a26643a );
 a26653a <=( (not A233)  and  A232 );
 a26654a <=( (not A202)  and  a26653a );
 a26658a <=( A267  and  A266 );
 a26659a <=( A236  and  a26658a );
 a26660a <=( a26659a  and  a26654a );
 a26664a <=( A166  and  (not A167) );
 a26665a <=( A170  and  a26664a );
 a26669a <=( (not A202)  and  (not A200) );
 a26670a <=( (not A199)  and  a26669a );
 a26671a <=( a26670a  and  a26665a );
 a26675a <=( A298  and  A234 );
 a26676a <=( A232  and  a26675a );
 a26680a <=( (not A301)  and  (not A300) );
 a26681a <=( A299  and  a26680a );
 a26682a <=( a26681a  and  a26676a );
 a26686a <=( A166  and  (not A167) );
 a26687a <=( A170  and  a26686a );
 a26691a <=( (not A202)  and  (not A200) );
 a26692a <=( (not A199)  and  a26691a );
 a26693a <=( a26692a  and  a26687a );
 a26697a <=( A298  and  A234 );
 a26698a <=( A233  and  a26697a );
 a26702a <=( (not A301)  and  (not A300) );
 a26703a <=( A299  and  a26702a );
 a26704a <=( a26703a  and  a26698a );
 a26708a <=( A166  and  (not A167) );
 a26709a <=( A170  and  a26708a );
 a26713a <=( (not A202)  and  (not A200) );
 a26714a <=( (not A199)  and  a26713a );
 a26715a <=( a26714a  and  a26709a );
 a26719a <=( A236  and  A233 );
 a26720a <=( (not A232)  and  a26719a );
 a26724a <=( (not A302)  and  (not A301) );
 a26725a <=( (not A300)  and  a26724a );
 a26726a <=( a26725a  and  a26720a );
 a26730a <=( A166  and  (not A167) );
 a26731a <=( A170  and  a26730a );
 a26735a <=( (not A202)  and  (not A200) );
 a26736a <=( (not A199)  and  a26735a );
 a26737a <=( a26736a  and  a26731a );
 a26741a <=( A236  and  A233 );
 a26742a <=( (not A232)  and  a26741a );
 a26746a <=( (not A301)  and  (not A299) );
 a26747a <=( (not A298)  and  a26746a );
 a26748a <=( a26747a  and  a26742a );
 a26752a <=( A166  and  (not A167) );
 a26753a <=( A170  and  a26752a );
 a26757a <=( (not A202)  and  (not A200) );
 a26758a <=( (not A199)  and  a26757a );
 a26759a <=( a26758a  and  a26753a );
 a26763a <=( A236  and  A233 );
 a26764a <=( (not A232)  and  a26763a );
 a26768a <=( A269  and  A266 );
 a26769a <=( (not A265)  and  a26768a );
 a26770a <=( a26769a  and  a26764a );
 a26774a <=( A166  and  (not A167) );
 a26775a <=( A170  and  a26774a );
 a26779a <=( (not A202)  and  (not A200) );
 a26780a <=( (not A199)  and  a26779a );
 a26781a <=( a26780a  and  a26775a );
 a26785a <=( A236  and  A233 );
 a26786a <=( (not A232)  and  a26785a );
 a26790a <=( A269  and  (not A266) );
 a26791a <=( A265  and  a26790a );
 a26792a <=( a26791a  and  a26786a );
 a26796a <=( A166  and  (not A167) );
 a26797a <=( A170  and  a26796a );
 a26801a <=( (not A202)  and  (not A200) );
 a26802a <=( (not A199)  and  a26801a );
 a26803a <=( a26802a  and  a26797a );
 a26807a <=( A236  and  (not A233) );
 a26808a <=( A232  and  a26807a );
 a26812a <=( (not A302)  and  (not A301) );
 a26813a <=( (not A300)  and  a26812a );
 a26814a <=( a26813a  and  a26808a );
 a26818a <=( A166  and  (not A167) );
 a26819a <=( A170  and  a26818a );
 a26823a <=( (not A202)  and  (not A200) );
 a26824a <=( (not A199)  and  a26823a );
 a26825a <=( a26824a  and  a26819a );
 a26829a <=( A236  and  (not A233) );
 a26830a <=( A232  and  a26829a );
 a26834a <=( (not A301)  and  (not A299) );
 a26835a <=( (not A298)  and  a26834a );
 a26836a <=( a26835a  and  a26830a );
 a26840a <=( A166  and  (not A167) );
 a26841a <=( A170  and  a26840a );
 a26845a <=( (not A202)  and  (not A200) );
 a26846a <=( (not A199)  and  a26845a );
 a26847a <=( a26846a  and  a26841a );
 a26851a <=( A236  and  (not A233) );
 a26852a <=( A232  and  a26851a );
 a26856a <=( A269  and  A266 );
 a26857a <=( (not A265)  and  a26856a );
 a26858a <=( a26857a  and  a26852a );
 a26862a <=( A166  and  (not A167) );
 a26863a <=( A170  and  a26862a );
 a26867a <=( (not A202)  and  (not A200) );
 a26868a <=( (not A199)  and  a26867a );
 a26869a <=( a26868a  and  a26863a );
 a26873a <=( A236  and  (not A233) );
 a26874a <=( A232  and  a26873a );
 a26878a <=( A269  and  (not A266) );
 a26879a <=( A265  and  a26878a );
 a26880a <=( a26879a  and  a26874a );
 a26884a <=( (not A202)  and  (not A201) );
 a26885a <=( A169  and  a26884a );
 a26889a <=( (not A235)  and  (not A234) );
 a26890a <=( (not A203)  and  a26889a );
 a26891a <=( a26890a  and  a26885a );
 a26895a <=( (not A268)  and  (not A267) );
 a26896a <=( (not A236)  and  a26895a );
 a26900a <=( A300  and  A299 );
 a26901a <=( (not A269)  and  a26900a );
 a26902a <=( a26901a  and  a26896a );
 a26906a <=( (not A202)  and  (not A201) );
 a26907a <=( A169  and  a26906a );
 a26911a <=( (not A235)  and  (not A234) );
 a26912a <=( (not A203)  and  a26911a );
 a26913a <=( a26912a  and  a26907a );
 a26917a <=( (not A268)  and  (not A267) );
 a26918a <=( (not A236)  and  a26917a );
 a26922a <=( A300  and  A298 );
 a26923a <=( (not A269)  and  a26922a );
 a26924a <=( a26923a  and  a26918a );
 a26928a <=( (not A202)  and  (not A201) );
 a26929a <=( A169  and  a26928a );
 a26933a <=( (not A235)  and  (not A234) );
 a26934a <=( (not A203)  and  a26933a );
 a26935a <=( a26934a  and  a26929a );
 a26939a <=( A266  and  A265 );
 a26940a <=( (not A236)  and  a26939a );
 a26944a <=( A301  and  (not A268) );
 a26945a <=( (not A267)  and  a26944a );
 a26946a <=( a26945a  and  a26940a );
 a26950a <=( (not A202)  and  (not A201) );
 a26951a <=( A169  and  a26950a );
 a26955a <=( (not A235)  and  (not A234) );
 a26956a <=( (not A203)  and  a26955a );
 a26957a <=( a26956a  and  a26951a );
 a26961a <=( (not A266)  and  (not A265) );
 a26962a <=( (not A236)  and  a26961a );
 a26966a <=( A300  and  A299 );
 a26967a <=( (not A268)  and  a26966a );
 a26968a <=( a26967a  and  a26962a );
 a26972a <=( (not A202)  and  (not A201) );
 a26973a <=( A169  and  a26972a );
 a26977a <=( (not A235)  and  (not A234) );
 a26978a <=( (not A203)  and  a26977a );
 a26979a <=( a26978a  and  a26973a );
 a26983a <=( (not A266)  and  (not A265) );
 a26984a <=( (not A236)  and  a26983a );
 a26988a <=( A300  and  A298 );
 a26989a <=( (not A268)  and  a26988a );
 a26990a <=( a26989a  and  a26984a );
 a26994a <=( (not A202)  and  (not A201) );
 a26995a <=( A169  and  a26994a );
 a26999a <=( A233  and  A232 );
 a27000a <=( (not A203)  and  a26999a );
 a27001a <=( a27000a  and  a26995a );
 a27005a <=( (not A267)  and  (not A235) );
 a27006a <=( (not A234)  and  a27005a );
 a27010a <=( A301  and  (not A269) );
 a27011a <=( (not A268)  and  a27010a );
 a27012a <=( a27011a  and  a27006a );
 a27016a <=( (not A202)  and  (not A201) );
 a27017a <=( A169  and  a27016a );
 a27021a <=( A233  and  A232 );
 a27022a <=( (not A203)  and  a27021a );
 a27023a <=( a27022a  and  a27017a );
 a27027a <=( (not A265)  and  (not A235) );
 a27028a <=( (not A234)  and  a27027a );
 a27032a <=( A301  and  (not A268) );
 a27033a <=( (not A266)  and  a27032a );
 a27034a <=( a27033a  and  a27028a );
 a27038a <=( (not A202)  and  (not A201) );
 a27039a <=( A169  and  a27038a );
 a27043a <=( (not A233)  and  (not A232) );
 a27044a <=( (not A203)  and  a27043a );
 a27045a <=( a27044a  and  a27039a );
 a27049a <=( (not A268)  and  (not A267) );
 a27050a <=( (not A235)  and  a27049a );
 a27054a <=( A300  and  A299 );
 a27055a <=( (not A269)  and  a27054a );
 a27056a <=( a27055a  and  a27050a );
 a27060a <=( (not A202)  and  (not A201) );
 a27061a <=( A169  and  a27060a );
 a27065a <=( (not A233)  and  (not A232) );
 a27066a <=( (not A203)  and  a27065a );
 a27067a <=( a27066a  and  a27061a );
 a27071a <=( (not A268)  and  (not A267) );
 a27072a <=( (not A235)  and  a27071a );
 a27076a <=( A300  and  A298 );
 a27077a <=( (not A269)  and  a27076a );
 a27078a <=( a27077a  and  a27072a );
 a27082a <=( (not A202)  and  (not A201) );
 a27083a <=( A169  and  a27082a );
 a27087a <=( (not A233)  and  (not A232) );
 a27088a <=( (not A203)  and  a27087a );
 a27089a <=( a27088a  and  a27083a );
 a27093a <=( A266  and  A265 );
 a27094a <=( (not A235)  and  a27093a );
 a27098a <=( A301  and  (not A268) );
 a27099a <=( (not A267)  and  a27098a );
 a27100a <=( a27099a  and  a27094a );
 a27104a <=( (not A202)  and  (not A201) );
 a27105a <=( A169  and  a27104a );
 a27109a <=( (not A233)  and  (not A232) );
 a27110a <=( (not A203)  and  a27109a );
 a27111a <=( a27110a  and  a27105a );
 a27115a <=( (not A266)  and  (not A265) );
 a27116a <=( (not A235)  and  a27115a );
 a27120a <=( A300  and  A299 );
 a27121a <=( (not A268)  and  a27120a );
 a27122a <=( a27121a  and  a27116a );
 a27126a <=( (not A202)  and  (not A201) );
 a27127a <=( A169  and  a27126a );
 a27131a <=( (not A233)  and  (not A232) );
 a27132a <=( (not A203)  and  a27131a );
 a27133a <=( a27132a  and  a27127a );
 a27137a <=( (not A266)  and  (not A265) );
 a27138a <=( (not A235)  and  a27137a );
 a27142a <=( A300  and  A298 );
 a27143a <=( (not A268)  and  a27142a );
 a27144a <=( a27143a  and  a27138a );
 a27148a <=( A200  and  A199 );
 a27149a <=( A169  and  a27148a );
 a27153a <=( (not A234)  and  (not A202) );
 a27154a <=( (not A201)  and  a27153a );
 a27155a <=( a27154a  and  a27149a );
 a27159a <=( (not A267)  and  (not A236) );
 a27160a <=( (not A235)  and  a27159a );
 a27164a <=( A301  and  (not A269) );
 a27165a <=( (not A268)  and  a27164a );
 a27166a <=( a27165a  and  a27160a );
 a27170a <=( A200  and  A199 );
 a27171a <=( A169  and  a27170a );
 a27175a <=( (not A234)  and  (not A202) );
 a27176a <=( (not A201)  and  a27175a );
 a27177a <=( a27176a  and  a27171a );
 a27181a <=( (not A265)  and  (not A236) );
 a27182a <=( (not A235)  and  a27181a );
 a27186a <=( A301  and  (not A268) );
 a27187a <=( (not A266)  and  a27186a );
 a27188a <=( a27187a  and  a27182a );
 a27192a <=( A200  and  A199 );
 a27193a <=( A169  and  a27192a );
 a27197a <=( (not A232)  and  (not A202) );
 a27198a <=( (not A201)  and  a27197a );
 a27199a <=( a27198a  and  a27193a );
 a27203a <=( A298  and  A236 );
 a27204a <=( A233  and  a27203a );
 a27208a <=( (not A301)  and  (not A300) );
 a27209a <=( A299  and  a27208a );
 a27210a <=( a27209a  and  a27204a );
 a27214a <=( A200  and  A199 );
 a27215a <=( A169  and  a27214a );
 a27219a <=( A232  and  (not A202) );
 a27220a <=( (not A201)  and  a27219a );
 a27221a <=( a27220a  and  a27215a );
 a27225a <=( A298  and  A236 );
 a27226a <=( (not A233)  and  a27225a );
 a27230a <=( (not A301)  and  (not A300) );
 a27231a <=( A299  and  a27230a );
 a27232a <=( a27231a  and  a27226a );
 a27236a <=( A200  and  A199 );
 a27237a <=( A169  and  a27236a );
 a27241a <=( (not A232)  and  (not A202) );
 a27242a <=( (not A201)  and  a27241a );
 a27243a <=( a27242a  and  a27237a );
 a27247a <=( (not A267)  and  (not A235) );
 a27248a <=( (not A233)  and  a27247a );
 a27252a <=( A301  and  (not A269) );
 a27253a <=( (not A268)  and  a27252a );
 a27254a <=( a27253a  and  a27248a );
 a27258a <=( A200  and  A199 );
 a27259a <=( A169  and  a27258a );
 a27263a <=( (not A232)  and  (not A202) );
 a27264a <=( (not A201)  and  a27263a );
 a27265a <=( a27264a  and  a27259a );
 a27269a <=( (not A265)  and  (not A235) );
 a27270a <=( (not A233)  and  a27269a );
 a27274a <=( A301  and  (not A268) );
 a27275a <=( (not A266)  and  a27274a );
 a27276a <=( a27275a  and  a27270a );
 a27280a <=( (not A200)  and  (not A199) );
 a27281a <=( A169  and  a27280a );
 a27285a <=( (not A235)  and  (not A234) );
 a27286a <=( (not A202)  and  a27285a );
 a27287a <=( a27286a  and  a27281a );
 a27291a <=( (not A268)  and  (not A267) );
 a27292a <=( (not A236)  and  a27291a );
 a27296a <=( A300  and  A299 );
 a27297a <=( (not A269)  and  a27296a );
 a27298a <=( a27297a  and  a27292a );
 a27302a <=( (not A200)  and  (not A199) );
 a27303a <=( A169  and  a27302a );
 a27307a <=( (not A235)  and  (not A234) );
 a27308a <=( (not A202)  and  a27307a );
 a27309a <=( a27308a  and  a27303a );
 a27313a <=( (not A268)  and  (not A267) );
 a27314a <=( (not A236)  and  a27313a );
 a27318a <=( A300  and  A298 );
 a27319a <=( (not A269)  and  a27318a );
 a27320a <=( a27319a  and  a27314a );
 a27324a <=( (not A200)  and  (not A199) );
 a27325a <=( A169  and  a27324a );
 a27329a <=( (not A235)  and  (not A234) );
 a27330a <=( (not A202)  and  a27329a );
 a27331a <=( a27330a  and  a27325a );
 a27335a <=( A266  and  A265 );
 a27336a <=( (not A236)  and  a27335a );
 a27340a <=( A301  and  (not A268) );
 a27341a <=( (not A267)  and  a27340a );
 a27342a <=( a27341a  and  a27336a );
 a27346a <=( (not A200)  and  (not A199) );
 a27347a <=( A169  and  a27346a );
 a27351a <=( (not A235)  and  (not A234) );
 a27352a <=( (not A202)  and  a27351a );
 a27353a <=( a27352a  and  a27347a );
 a27357a <=( (not A266)  and  (not A265) );
 a27358a <=( (not A236)  and  a27357a );
 a27362a <=( A300  and  A299 );
 a27363a <=( (not A268)  and  a27362a );
 a27364a <=( a27363a  and  a27358a );
 a27368a <=( (not A200)  and  (not A199) );
 a27369a <=( A169  and  a27368a );
 a27373a <=( (not A235)  and  (not A234) );
 a27374a <=( (not A202)  and  a27373a );
 a27375a <=( a27374a  and  a27369a );
 a27379a <=( (not A266)  and  (not A265) );
 a27380a <=( (not A236)  and  a27379a );
 a27384a <=( A300  and  A298 );
 a27385a <=( (not A268)  and  a27384a );
 a27386a <=( a27385a  and  a27380a );
 a27390a <=( (not A200)  and  (not A199) );
 a27391a <=( A169  and  a27390a );
 a27395a <=( A233  and  A232 );
 a27396a <=( (not A202)  and  a27395a );
 a27397a <=( a27396a  and  a27391a );
 a27401a <=( (not A267)  and  (not A235) );
 a27402a <=( (not A234)  and  a27401a );
 a27406a <=( A301  and  (not A269) );
 a27407a <=( (not A268)  and  a27406a );
 a27408a <=( a27407a  and  a27402a );
 a27412a <=( (not A200)  and  (not A199) );
 a27413a <=( A169  and  a27412a );
 a27417a <=( A233  and  A232 );
 a27418a <=( (not A202)  and  a27417a );
 a27419a <=( a27418a  and  a27413a );
 a27423a <=( (not A265)  and  (not A235) );
 a27424a <=( (not A234)  and  a27423a );
 a27428a <=( A301  and  (not A268) );
 a27429a <=( (not A266)  and  a27428a );
 a27430a <=( a27429a  and  a27424a );
 a27434a <=( (not A200)  and  (not A199) );
 a27435a <=( A169  and  a27434a );
 a27439a <=( (not A233)  and  (not A232) );
 a27440a <=( (not A202)  and  a27439a );
 a27441a <=( a27440a  and  a27435a );
 a27445a <=( (not A268)  and  (not A267) );
 a27446a <=( (not A235)  and  a27445a );
 a27450a <=( A300  and  A299 );
 a27451a <=( (not A269)  and  a27450a );
 a27452a <=( a27451a  and  a27446a );
 a27456a <=( (not A200)  and  (not A199) );
 a27457a <=( A169  and  a27456a );
 a27461a <=( (not A233)  and  (not A232) );
 a27462a <=( (not A202)  and  a27461a );
 a27463a <=( a27462a  and  a27457a );
 a27467a <=( (not A268)  and  (not A267) );
 a27468a <=( (not A235)  and  a27467a );
 a27472a <=( A300  and  A298 );
 a27473a <=( (not A269)  and  a27472a );
 a27474a <=( a27473a  and  a27468a );
 a27478a <=( (not A200)  and  (not A199) );
 a27479a <=( A169  and  a27478a );
 a27483a <=( (not A233)  and  (not A232) );
 a27484a <=( (not A202)  and  a27483a );
 a27485a <=( a27484a  and  a27479a );
 a27489a <=( A266  and  A265 );
 a27490a <=( (not A235)  and  a27489a );
 a27494a <=( A301  and  (not A268) );
 a27495a <=( (not A267)  and  a27494a );
 a27496a <=( a27495a  and  a27490a );
 a27500a <=( (not A200)  and  (not A199) );
 a27501a <=( A169  and  a27500a );
 a27505a <=( (not A233)  and  (not A232) );
 a27506a <=( (not A202)  and  a27505a );
 a27507a <=( a27506a  and  a27501a );
 a27511a <=( (not A266)  and  (not A265) );
 a27512a <=( (not A235)  and  a27511a );
 a27516a <=( A300  and  A299 );
 a27517a <=( (not A268)  and  a27516a );
 a27518a <=( a27517a  and  a27512a );
 a27522a <=( (not A200)  and  (not A199) );
 a27523a <=( A169  and  a27522a );
 a27527a <=( (not A233)  and  (not A232) );
 a27528a <=( (not A202)  and  a27527a );
 a27529a <=( a27528a  and  a27523a );
 a27533a <=( (not A266)  and  (not A265) );
 a27534a <=( (not A235)  and  a27533a );
 a27538a <=( A300  and  A298 );
 a27539a <=( (not A268)  and  a27538a );
 a27540a <=( a27539a  and  a27534a );
 a27544a <=( (not A166)  and  (not A167) );
 a27545a <=( (not A169)  and  a27544a );
 a27549a <=( (not A235)  and  (not A234) );
 a27550a <=( A202  and  a27549a );
 a27551a <=( a27550a  and  a27545a );
 a27555a <=( (not A268)  and  (not A267) );
 a27556a <=( (not A236)  and  a27555a );
 a27560a <=( A300  and  A299 );
 a27561a <=( (not A269)  and  a27560a );
 a27562a <=( a27561a  and  a27556a );
 a27566a <=( (not A166)  and  (not A167) );
 a27567a <=( (not A169)  and  a27566a );
 a27571a <=( (not A235)  and  (not A234) );
 a27572a <=( A202  and  a27571a );
 a27573a <=( a27572a  and  a27567a );
 a27577a <=( (not A268)  and  (not A267) );
 a27578a <=( (not A236)  and  a27577a );
 a27582a <=( A300  and  A298 );
 a27583a <=( (not A269)  and  a27582a );
 a27584a <=( a27583a  and  a27578a );
 a27588a <=( (not A166)  and  (not A167) );
 a27589a <=( (not A169)  and  a27588a );
 a27593a <=( (not A235)  and  (not A234) );
 a27594a <=( A202  and  a27593a );
 a27595a <=( a27594a  and  a27589a );
 a27599a <=( A266  and  A265 );
 a27600a <=( (not A236)  and  a27599a );
 a27604a <=( A301  and  (not A268) );
 a27605a <=( (not A267)  and  a27604a );
 a27606a <=( a27605a  and  a27600a );
 a27610a <=( (not A166)  and  (not A167) );
 a27611a <=( (not A169)  and  a27610a );
 a27615a <=( (not A235)  and  (not A234) );
 a27616a <=( A202  and  a27615a );
 a27617a <=( a27616a  and  a27611a );
 a27621a <=( (not A266)  and  (not A265) );
 a27622a <=( (not A236)  and  a27621a );
 a27626a <=( A300  and  A299 );
 a27627a <=( (not A268)  and  a27626a );
 a27628a <=( a27627a  and  a27622a );
 a27632a <=( (not A166)  and  (not A167) );
 a27633a <=( (not A169)  and  a27632a );
 a27637a <=( (not A235)  and  (not A234) );
 a27638a <=( A202  and  a27637a );
 a27639a <=( a27638a  and  a27633a );
 a27643a <=( (not A266)  and  (not A265) );
 a27644a <=( (not A236)  and  a27643a );
 a27648a <=( A300  and  A298 );
 a27649a <=( (not A268)  and  a27648a );
 a27650a <=( a27649a  and  a27644a );
 a27654a <=( (not A166)  and  (not A167) );
 a27655a <=( (not A169)  and  a27654a );
 a27659a <=( A233  and  A232 );
 a27660a <=( A202  and  a27659a );
 a27661a <=( a27660a  and  a27655a );
 a27665a <=( (not A267)  and  (not A235) );
 a27666a <=( (not A234)  and  a27665a );
 a27670a <=( A301  and  (not A269) );
 a27671a <=( (not A268)  and  a27670a );
 a27672a <=( a27671a  and  a27666a );
 a27676a <=( (not A166)  and  (not A167) );
 a27677a <=( (not A169)  and  a27676a );
 a27681a <=( A233  and  A232 );
 a27682a <=( A202  and  a27681a );
 a27683a <=( a27682a  and  a27677a );
 a27687a <=( (not A265)  and  (not A235) );
 a27688a <=( (not A234)  and  a27687a );
 a27692a <=( A301  and  (not A268) );
 a27693a <=( (not A266)  and  a27692a );
 a27694a <=( a27693a  and  a27688a );
 a27698a <=( (not A166)  and  (not A167) );
 a27699a <=( (not A169)  and  a27698a );
 a27703a <=( (not A233)  and  (not A232) );
 a27704a <=( A202  and  a27703a );
 a27705a <=( a27704a  and  a27699a );
 a27709a <=( (not A268)  and  (not A267) );
 a27710a <=( (not A235)  and  a27709a );
 a27714a <=( A300  and  A299 );
 a27715a <=( (not A269)  and  a27714a );
 a27716a <=( a27715a  and  a27710a );
 a27720a <=( (not A166)  and  (not A167) );
 a27721a <=( (not A169)  and  a27720a );
 a27725a <=( (not A233)  and  (not A232) );
 a27726a <=( A202  and  a27725a );
 a27727a <=( a27726a  and  a27721a );
 a27731a <=( (not A268)  and  (not A267) );
 a27732a <=( (not A235)  and  a27731a );
 a27736a <=( A300  and  A298 );
 a27737a <=( (not A269)  and  a27736a );
 a27738a <=( a27737a  and  a27732a );
 a27742a <=( (not A166)  and  (not A167) );
 a27743a <=( (not A169)  and  a27742a );
 a27747a <=( (not A233)  and  (not A232) );
 a27748a <=( A202  and  a27747a );
 a27749a <=( a27748a  and  a27743a );
 a27753a <=( A266  and  A265 );
 a27754a <=( (not A235)  and  a27753a );
 a27758a <=( A301  and  (not A268) );
 a27759a <=( (not A267)  and  a27758a );
 a27760a <=( a27759a  and  a27754a );
 a27764a <=( (not A166)  and  (not A167) );
 a27765a <=( (not A169)  and  a27764a );
 a27769a <=( (not A233)  and  (not A232) );
 a27770a <=( A202  and  a27769a );
 a27771a <=( a27770a  and  a27765a );
 a27775a <=( (not A266)  and  (not A265) );
 a27776a <=( (not A235)  and  a27775a );
 a27780a <=( A300  and  A299 );
 a27781a <=( (not A268)  and  a27780a );
 a27782a <=( a27781a  and  a27776a );
 a27786a <=( (not A166)  and  (not A167) );
 a27787a <=( (not A169)  and  a27786a );
 a27791a <=( (not A233)  and  (not A232) );
 a27792a <=( A202  and  a27791a );
 a27793a <=( a27792a  and  a27787a );
 a27797a <=( (not A266)  and  (not A265) );
 a27798a <=( (not A235)  and  a27797a );
 a27802a <=( A300  and  A298 );
 a27803a <=( (not A268)  and  a27802a );
 a27804a <=( a27803a  and  a27798a );
 a27808a <=( (not A166)  and  (not A167) );
 a27809a <=( (not A169)  and  a27808a );
 a27813a <=( (not A234)  and  A201 );
 a27814a <=( A199  and  a27813a );
 a27815a <=( a27814a  and  a27809a );
 a27819a <=( (not A267)  and  (not A236) );
 a27820a <=( (not A235)  and  a27819a );
 a27824a <=( A301  and  (not A269) );
 a27825a <=( (not A268)  and  a27824a );
 a27826a <=( a27825a  and  a27820a );
 a27830a <=( (not A166)  and  (not A167) );
 a27831a <=( (not A169)  and  a27830a );
 a27835a <=( (not A234)  and  A201 );
 a27836a <=( A199  and  a27835a );
 a27837a <=( a27836a  and  a27831a );
 a27841a <=( (not A265)  and  (not A236) );
 a27842a <=( (not A235)  and  a27841a );
 a27846a <=( A301  and  (not A268) );
 a27847a <=( (not A266)  and  a27846a );
 a27848a <=( a27847a  and  a27842a );
 a27852a <=( (not A166)  and  (not A167) );
 a27853a <=( (not A169)  and  a27852a );
 a27857a <=( (not A232)  and  A201 );
 a27858a <=( A199  and  a27857a );
 a27859a <=( a27858a  and  a27853a );
 a27863a <=( A298  and  A236 );
 a27864a <=( A233  and  a27863a );
 a27868a <=( (not A301)  and  (not A300) );
 a27869a <=( A299  and  a27868a );
 a27870a <=( a27869a  and  a27864a );
 a27874a <=( (not A166)  and  (not A167) );
 a27875a <=( (not A169)  and  a27874a );
 a27879a <=( A232  and  A201 );
 a27880a <=( A199  and  a27879a );
 a27881a <=( a27880a  and  a27875a );
 a27885a <=( A298  and  A236 );
 a27886a <=( (not A233)  and  a27885a );
 a27890a <=( (not A301)  and  (not A300) );
 a27891a <=( A299  and  a27890a );
 a27892a <=( a27891a  and  a27886a );
 a27896a <=( (not A166)  and  (not A167) );
 a27897a <=( (not A169)  and  a27896a );
 a27901a <=( (not A232)  and  A201 );
 a27902a <=( A199  and  a27901a );
 a27903a <=( a27902a  and  a27897a );
 a27907a <=( (not A267)  and  (not A235) );
 a27908a <=( (not A233)  and  a27907a );
 a27912a <=( A301  and  (not A269) );
 a27913a <=( (not A268)  and  a27912a );
 a27914a <=( a27913a  and  a27908a );
 a27918a <=( (not A166)  and  (not A167) );
 a27919a <=( (not A169)  and  a27918a );
 a27923a <=( (not A232)  and  A201 );
 a27924a <=( A199  and  a27923a );
 a27925a <=( a27924a  and  a27919a );
 a27929a <=( (not A265)  and  (not A235) );
 a27930a <=( (not A233)  and  a27929a );
 a27934a <=( A301  and  (not A268) );
 a27935a <=( (not A266)  and  a27934a );
 a27936a <=( a27935a  and  a27930a );
 a27940a <=( (not A166)  and  (not A167) );
 a27941a <=( (not A169)  and  a27940a );
 a27945a <=( (not A234)  and  A201 );
 a27946a <=( A200  and  a27945a );
 a27947a <=( a27946a  and  a27941a );
 a27951a <=( (not A267)  and  (not A236) );
 a27952a <=( (not A235)  and  a27951a );
 a27956a <=( A301  and  (not A269) );
 a27957a <=( (not A268)  and  a27956a );
 a27958a <=( a27957a  and  a27952a );
 a27962a <=( (not A166)  and  (not A167) );
 a27963a <=( (not A169)  and  a27962a );
 a27967a <=( (not A234)  and  A201 );
 a27968a <=( A200  and  a27967a );
 a27969a <=( a27968a  and  a27963a );
 a27973a <=( (not A265)  and  (not A236) );
 a27974a <=( (not A235)  and  a27973a );
 a27978a <=( A301  and  (not A268) );
 a27979a <=( (not A266)  and  a27978a );
 a27980a <=( a27979a  and  a27974a );
 a27984a <=( (not A166)  and  (not A167) );
 a27985a <=( (not A169)  and  a27984a );
 a27989a <=( (not A232)  and  A201 );
 a27990a <=( A200  and  a27989a );
 a27991a <=( a27990a  and  a27985a );
 a27995a <=( A298  and  A236 );
 a27996a <=( A233  and  a27995a );
 a28000a <=( (not A301)  and  (not A300) );
 a28001a <=( A299  and  a28000a );
 a28002a <=( a28001a  and  a27996a );
 a28006a <=( (not A166)  and  (not A167) );
 a28007a <=( (not A169)  and  a28006a );
 a28011a <=( A232  and  A201 );
 a28012a <=( A200  and  a28011a );
 a28013a <=( a28012a  and  a28007a );
 a28017a <=( A298  and  A236 );
 a28018a <=( (not A233)  and  a28017a );
 a28022a <=( (not A301)  and  (not A300) );
 a28023a <=( A299  and  a28022a );
 a28024a <=( a28023a  and  a28018a );
 a28028a <=( (not A166)  and  (not A167) );
 a28029a <=( (not A169)  and  a28028a );
 a28033a <=( (not A232)  and  A201 );
 a28034a <=( A200  and  a28033a );
 a28035a <=( a28034a  and  a28029a );
 a28039a <=( (not A267)  and  (not A235) );
 a28040a <=( (not A233)  and  a28039a );
 a28044a <=( A301  and  (not A269) );
 a28045a <=( (not A268)  and  a28044a );
 a28046a <=( a28045a  and  a28040a );
 a28050a <=( (not A166)  and  (not A167) );
 a28051a <=( (not A169)  and  a28050a );
 a28055a <=( (not A232)  and  A201 );
 a28056a <=( A200  and  a28055a );
 a28057a <=( a28056a  and  a28051a );
 a28061a <=( (not A265)  and  (not A235) );
 a28062a <=( (not A233)  and  a28061a );
 a28066a <=( A301  and  (not A268) );
 a28067a <=( (not A266)  and  a28066a );
 a28068a <=( a28067a  and  a28062a );
 a28072a <=( (not A166)  and  (not A167) );
 a28073a <=( (not A169)  and  a28072a );
 a28077a <=( A203  and  A200 );
 a28078a <=( (not A199)  and  a28077a );
 a28079a <=( a28078a  and  a28073a );
 a28083a <=( A298  and  A234 );
 a28084a <=( A232  and  a28083a );
 a28088a <=( (not A301)  and  (not A300) );
 a28089a <=( A299  and  a28088a );
 a28090a <=( a28089a  and  a28084a );
 a28094a <=( (not A166)  and  (not A167) );
 a28095a <=( (not A169)  and  a28094a );
 a28099a <=( A203  and  A200 );
 a28100a <=( (not A199)  and  a28099a );
 a28101a <=( a28100a  and  a28095a );
 a28105a <=( A298  and  A234 );
 a28106a <=( A233  and  a28105a );
 a28110a <=( (not A301)  and  (not A300) );
 a28111a <=( A299  and  a28110a );
 a28112a <=( a28111a  and  a28106a );
 a28116a <=( (not A166)  and  (not A167) );
 a28117a <=( (not A169)  and  a28116a );
 a28121a <=( A203  and  A200 );
 a28122a <=( (not A199)  and  a28121a );
 a28123a <=( a28122a  and  a28117a );
 a28127a <=( A236  and  A233 );
 a28128a <=( (not A232)  and  a28127a );
 a28132a <=( (not A302)  and  (not A301) );
 a28133a <=( (not A300)  and  a28132a );
 a28134a <=( a28133a  and  a28128a );
 a28138a <=( (not A166)  and  (not A167) );
 a28139a <=( (not A169)  and  a28138a );
 a28143a <=( A203  and  A200 );
 a28144a <=( (not A199)  and  a28143a );
 a28145a <=( a28144a  and  a28139a );
 a28149a <=( A236  and  A233 );
 a28150a <=( (not A232)  and  a28149a );
 a28154a <=( (not A301)  and  (not A299) );
 a28155a <=( (not A298)  and  a28154a );
 a28156a <=( a28155a  and  a28150a );
 a28160a <=( (not A166)  and  (not A167) );
 a28161a <=( (not A169)  and  a28160a );
 a28165a <=( A203  and  A200 );
 a28166a <=( (not A199)  and  a28165a );
 a28167a <=( a28166a  and  a28161a );
 a28171a <=( A236  and  A233 );
 a28172a <=( (not A232)  and  a28171a );
 a28176a <=( A269  and  A266 );
 a28177a <=( (not A265)  and  a28176a );
 a28178a <=( a28177a  and  a28172a );
 a28182a <=( (not A166)  and  (not A167) );
 a28183a <=( (not A169)  and  a28182a );
 a28187a <=( A203  and  A200 );
 a28188a <=( (not A199)  and  a28187a );
 a28189a <=( a28188a  and  a28183a );
 a28193a <=( A236  and  A233 );
 a28194a <=( (not A232)  and  a28193a );
 a28198a <=( A269  and  (not A266) );
 a28199a <=( A265  and  a28198a );
 a28200a <=( a28199a  and  a28194a );
 a28204a <=( (not A166)  and  (not A167) );
 a28205a <=( (not A169)  and  a28204a );
 a28209a <=( A203  and  A200 );
 a28210a <=( (not A199)  and  a28209a );
 a28211a <=( a28210a  and  a28205a );
 a28215a <=( A236  and  (not A233) );
 a28216a <=( A232  and  a28215a );
 a28220a <=( (not A302)  and  (not A301) );
 a28221a <=( (not A300)  and  a28220a );
 a28222a <=( a28221a  and  a28216a );
 a28226a <=( (not A166)  and  (not A167) );
 a28227a <=( (not A169)  and  a28226a );
 a28231a <=( A203  and  A200 );
 a28232a <=( (not A199)  and  a28231a );
 a28233a <=( a28232a  and  a28227a );
 a28237a <=( A236  and  (not A233) );
 a28238a <=( A232  and  a28237a );
 a28242a <=( (not A301)  and  (not A299) );
 a28243a <=( (not A298)  and  a28242a );
 a28244a <=( a28243a  and  a28238a );
 a28248a <=( (not A166)  and  (not A167) );
 a28249a <=( (not A169)  and  a28248a );
 a28253a <=( A203  and  A200 );
 a28254a <=( (not A199)  and  a28253a );
 a28255a <=( a28254a  and  a28249a );
 a28259a <=( A236  and  (not A233) );
 a28260a <=( A232  and  a28259a );
 a28264a <=( A269  and  A266 );
 a28265a <=( (not A265)  and  a28264a );
 a28266a <=( a28265a  and  a28260a );
 a28270a <=( (not A166)  and  (not A167) );
 a28271a <=( (not A169)  and  a28270a );
 a28275a <=( A203  and  A200 );
 a28276a <=( (not A199)  and  a28275a );
 a28277a <=( a28276a  and  a28271a );
 a28281a <=( A236  and  (not A233) );
 a28282a <=( A232  and  a28281a );
 a28286a <=( A269  and  (not A266) );
 a28287a <=( A265  and  a28286a );
 a28288a <=( a28287a  and  a28282a );
 a28292a <=( (not A166)  and  (not A167) );
 a28293a <=( (not A169)  and  a28292a );
 a28297a <=( A203  and  (not A200) );
 a28298a <=( A199  and  a28297a );
 a28299a <=( a28298a  and  a28293a );
 a28303a <=( A298  and  A234 );
 a28304a <=( A232  and  a28303a );
 a28308a <=( (not A301)  and  (not A300) );
 a28309a <=( A299  and  a28308a );
 a28310a <=( a28309a  and  a28304a );
 a28314a <=( (not A166)  and  (not A167) );
 a28315a <=( (not A169)  and  a28314a );
 a28319a <=( A203  and  (not A200) );
 a28320a <=( A199  and  a28319a );
 a28321a <=( a28320a  and  a28315a );
 a28325a <=( A298  and  A234 );
 a28326a <=( A233  and  a28325a );
 a28330a <=( (not A301)  and  (not A300) );
 a28331a <=( A299  and  a28330a );
 a28332a <=( a28331a  and  a28326a );
 a28336a <=( (not A166)  and  (not A167) );
 a28337a <=( (not A169)  and  a28336a );
 a28341a <=( A203  and  (not A200) );
 a28342a <=( A199  and  a28341a );
 a28343a <=( a28342a  and  a28337a );
 a28347a <=( A236  and  A233 );
 a28348a <=( (not A232)  and  a28347a );
 a28352a <=( (not A302)  and  (not A301) );
 a28353a <=( (not A300)  and  a28352a );
 a28354a <=( a28353a  and  a28348a );
 a28358a <=( (not A166)  and  (not A167) );
 a28359a <=( (not A169)  and  a28358a );
 a28363a <=( A203  and  (not A200) );
 a28364a <=( A199  and  a28363a );
 a28365a <=( a28364a  and  a28359a );
 a28369a <=( A236  and  A233 );
 a28370a <=( (not A232)  and  a28369a );
 a28374a <=( (not A301)  and  (not A299) );
 a28375a <=( (not A298)  and  a28374a );
 a28376a <=( a28375a  and  a28370a );
 a28380a <=( (not A166)  and  (not A167) );
 a28381a <=( (not A169)  and  a28380a );
 a28385a <=( A203  and  (not A200) );
 a28386a <=( A199  and  a28385a );
 a28387a <=( a28386a  and  a28381a );
 a28391a <=( A236  and  A233 );
 a28392a <=( (not A232)  and  a28391a );
 a28396a <=( A269  and  A266 );
 a28397a <=( (not A265)  and  a28396a );
 a28398a <=( a28397a  and  a28392a );
 a28402a <=( (not A166)  and  (not A167) );
 a28403a <=( (not A169)  and  a28402a );
 a28407a <=( A203  and  (not A200) );
 a28408a <=( A199  and  a28407a );
 a28409a <=( a28408a  and  a28403a );
 a28413a <=( A236  and  A233 );
 a28414a <=( (not A232)  and  a28413a );
 a28418a <=( A269  and  (not A266) );
 a28419a <=( A265  and  a28418a );
 a28420a <=( a28419a  and  a28414a );
 a28424a <=( (not A166)  and  (not A167) );
 a28425a <=( (not A169)  and  a28424a );
 a28429a <=( A203  and  (not A200) );
 a28430a <=( A199  and  a28429a );
 a28431a <=( a28430a  and  a28425a );
 a28435a <=( A236  and  (not A233) );
 a28436a <=( A232  and  a28435a );
 a28440a <=( (not A302)  and  (not A301) );
 a28441a <=( (not A300)  and  a28440a );
 a28442a <=( a28441a  and  a28436a );
 a28446a <=( (not A166)  and  (not A167) );
 a28447a <=( (not A169)  and  a28446a );
 a28451a <=( A203  and  (not A200) );
 a28452a <=( A199  and  a28451a );
 a28453a <=( a28452a  and  a28447a );
 a28457a <=( A236  and  (not A233) );
 a28458a <=( A232  and  a28457a );
 a28462a <=( (not A301)  and  (not A299) );
 a28463a <=( (not A298)  and  a28462a );
 a28464a <=( a28463a  and  a28458a );
 a28468a <=( (not A166)  and  (not A167) );
 a28469a <=( (not A169)  and  a28468a );
 a28473a <=( A203  and  (not A200) );
 a28474a <=( A199  and  a28473a );
 a28475a <=( a28474a  and  a28469a );
 a28479a <=( A236  and  (not A233) );
 a28480a <=( A232  and  a28479a );
 a28484a <=( A269  and  A266 );
 a28485a <=( (not A265)  and  a28484a );
 a28486a <=( a28485a  and  a28480a );
 a28490a <=( (not A166)  and  (not A167) );
 a28491a <=( (not A169)  and  a28490a );
 a28495a <=( A203  and  (not A200) );
 a28496a <=( A199  and  a28495a );
 a28497a <=( a28496a  and  a28491a );
 a28501a <=( A236  and  (not A233) );
 a28502a <=( A232  and  a28501a );
 a28506a <=( A269  and  (not A266) );
 a28507a <=( A265  and  a28506a );
 a28508a <=( a28507a  and  a28502a );
 a28512a <=( A167  and  (not A168) );
 a28513a <=( (not A169)  and  a28512a );
 a28517a <=( (not A234)  and  A202 );
 a28518a <=( A166  and  a28517a );
 a28519a <=( a28518a  and  a28513a );
 a28523a <=( (not A267)  and  (not A236) );
 a28524a <=( (not A235)  and  a28523a );
 a28528a <=( A301  and  (not A269) );
 a28529a <=( (not A268)  and  a28528a );
 a28530a <=( a28529a  and  a28524a );
 a28534a <=( A167  and  (not A168) );
 a28535a <=( (not A169)  and  a28534a );
 a28539a <=( (not A234)  and  A202 );
 a28540a <=( A166  and  a28539a );
 a28541a <=( a28540a  and  a28535a );
 a28545a <=( (not A265)  and  (not A236) );
 a28546a <=( (not A235)  and  a28545a );
 a28550a <=( A301  and  (not A268) );
 a28551a <=( (not A266)  and  a28550a );
 a28552a <=( a28551a  and  a28546a );
 a28556a <=( A167  and  (not A168) );
 a28557a <=( (not A169)  and  a28556a );
 a28561a <=( (not A232)  and  A202 );
 a28562a <=( A166  and  a28561a );
 a28563a <=( a28562a  and  a28557a );
 a28567a <=( A298  and  A236 );
 a28568a <=( A233  and  a28567a );
 a28572a <=( (not A301)  and  (not A300) );
 a28573a <=( A299  and  a28572a );
 a28574a <=( a28573a  and  a28568a );
 a28578a <=( A167  and  (not A168) );
 a28579a <=( (not A169)  and  a28578a );
 a28583a <=( A232  and  A202 );
 a28584a <=( A166  and  a28583a );
 a28585a <=( a28584a  and  a28579a );
 a28589a <=( A298  and  A236 );
 a28590a <=( (not A233)  and  a28589a );
 a28594a <=( (not A301)  and  (not A300) );
 a28595a <=( A299  and  a28594a );
 a28596a <=( a28595a  and  a28590a );
 a28600a <=( A167  and  (not A168) );
 a28601a <=( (not A169)  and  a28600a );
 a28605a <=( (not A232)  and  A202 );
 a28606a <=( A166  and  a28605a );
 a28607a <=( a28606a  and  a28601a );
 a28611a <=( (not A267)  and  (not A235) );
 a28612a <=( (not A233)  and  a28611a );
 a28616a <=( A301  and  (not A269) );
 a28617a <=( (not A268)  and  a28616a );
 a28618a <=( a28617a  and  a28612a );
 a28622a <=( A167  and  (not A168) );
 a28623a <=( (not A169)  and  a28622a );
 a28627a <=( (not A232)  and  A202 );
 a28628a <=( A166  and  a28627a );
 a28629a <=( a28628a  and  a28623a );
 a28633a <=( (not A265)  and  (not A235) );
 a28634a <=( (not A233)  and  a28633a );
 a28638a <=( A301  and  (not A268) );
 a28639a <=( (not A266)  and  a28638a );
 a28640a <=( a28639a  and  a28634a );
 a28644a <=( A167  and  (not A168) );
 a28645a <=( (not A169)  and  a28644a );
 a28649a <=( A201  and  A199 );
 a28650a <=( A166  and  a28649a );
 a28651a <=( a28650a  and  a28645a );
 a28655a <=( A298  and  A234 );
 a28656a <=( A232  and  a28655a );
 a28660a <=( (not A301)  and  (not A300) );
 a28661a <=( A299  and  a28660a );
 a28662a <=( a28661a  and  a28656a );
 a28666a <=( A167  and  (not A168) );
 a28667a <=( (not A169)  and  a28666a );
 a28671a <=( A201  and  A199 );
 a28672a <=( A166  and  a28671a );
 a28673a <=( a28672a  and  a28667a );
 a28677a <=( A298  and  A234 );
 a28678a <=( A233  and  a28677a );
 a28682a <=( (not A301)  and  (not A300) );
 a28683a <=( A299  and  a28682a );
 a28684a <=( a28683a  and  a28678a );
 a28688a <=( A167  and  (not A168) );
 a28689a <=( (not A169)  and  a28688a );
 a28693a <=( A201  and  A199 );
 a28694a <=( A166  and  a28693a );
 a28695a <=( a28694a  and  a28689a );
 a28699a <=( A236  and  A233 );
 a28700a <=( (not A232)  and  a28699a );
 a28704a <=( (not A302)  and  (not A301) );
 a28705a <=( (not A300)  and  a28704a );
 a28706a <=( a28705a  and  a28700a );
 a28710a <=( A167  and  (not A168) );
 a28711a <=( (not A169)  and  a28710a );
 a28715a <=( A201  and  A199 );
 a28716a <=( A166  and  a28715a );
 a28717a <=( a28716a  and  a28711a );
 a28721a <=( A236  and  A233 );
 a28722a <=( (not A232)  and  a28721a );
 a28726a <=( (not A301)  and  (not A299) );
 a28727a <=( (not A298)  and  a28726a );
 a28728a <=( a28727a  and  a28722a );
 a28732a <=( A167  and  (not A168) );
 a28733a <=( (not A169)  and  a28732a );
 a28737a <=( A201  and  A199 );
 a28738a <=( A166  and  a28737a );
 a28739a <=( a28738a  and  a28733a );
 a28743a <=( A236  and  A233 );
 a28744a <=( (not A232)  and  a28743a );
 a28748a <=( A269  and  A266 );
 a28749a <=( (not A265)  and  a28748a );
 a28750a <=( a28749a  and  a28744a );
 a28754a <=( A167  and  (not A168) );
 a28755a <=( (not A169)  and  a28754a );
 a28759a <=( A201  and  A199 );
 a28760a <=( A166  and  a28759a );
 a28761a <=( a28760a  and  a28755a );
 a28765a <=( A236  and  A233 );
 a28766a <=( (not A232)  and  a28765a );
 a28770a <=( A269  and  (not A266) );
 a28771a <=( A265  and  a28770a );
 a28772a <=( a28771a  and  a28766a );
 a28776a <=( A167  and  (not A168) );
 a28777a <=( (not A169)  and  a28776a );
 a28781a <=( A201  and  A199 );
 a28782a <=( A166  and  a28781a );
 a28783a <=( a28782a  and  a28777a );
 a28787a <=( A236  and  (not A233) );
 a28788a <=( A232  and  a28787a );
 a28792a <=( (not A302)  and  (not A301) );
 a28793a <=( (not A300)  and  a28792a );
 a28794a <=( a28793a  and  a28788a );
 a28798a <=( A167  and  (not A168) );
 a28799a <=( (not A169)  and  a28798a );
 a28803a <=( A201  and  A199 );
 a28804a <=( A166  and  a28803a );
 a28805a <=( a28804a  and  a28799a );
 a28809a <=( A236  and  (not A233) );
 a28810a <=( A232  and  a28809a );
 a28814a <=( (not A301)  and  (not A299) );
 a28815a <=( (not A298)  and  a28814a );
 a28816a <=( a28815a  and  a28810a );
 a28820a <=( A167  and  (not A168) );
 a28821a <=( (not A169)  and  a28820a );
 a28825a <=( A201  and  A199 );
 a28826a <=( A166  and  a28825a );
 a28827a <=( a28826a  and  a28821a );
 a28831a <=( A236  and  (not A233) );
 a28832a <=( A232  and  a28831a );
 a28836a <=( A269  and  A266 );
 a28837a <=( (not A265)  and  a28836a );
 a28838a <=( a28837a  and  a28832a );
 a28842a <=( A167  and  (not A168) );
 a28843a <=( (not A169)  and  a28842a );
 a28847a <=( A201  and  A199 );
 a28848a <=( A166  and  a28847a );
 a28849a <=( a28848a  and  a28843a );
 a28853a <=( A236  and  (not A233) );
 a28854a <=( A232  and  a28853a );
 a28858a <=( A269  and  (not A266) );
 a28859a <=( A265  and  a28858a );
 a28860a <=( a28859a  and  a28854a );
 a28864a <=( A167  and  (not A168) );
 a28865a <=( (not A169)  and  a28864a );
 a28869a <=( A201  and  A200 );
 a28870a <=( A166  and  a28869a );
 a28871a <=( a28870a  and  a28865a );
 a28875a <=( A298  and  A234 );
 a28876a <=( A232  and  a28875a );
 a28880a <=( (not A301)  and  (not A300) );
 a28881a <=( A299  and  a28880a );
 a28882a <=( a28881a  and  a28876a );
 a28886a <=( A167  and  (not A168) );
 a28887a <=( (not A169)  and  a28886a );
 a28891a <=( A201  and  A200 );
 a28892a <=( A166  and  a28891a );
 a28893a <=( a28892a  and  a28887a );
 a28897a <=( A298  and  A234 );
 a28898a <=( A233  and  a28897a );
 a28902a <=( (not A301)  and  (not A300) );
 a28903a <=( A299  and  a28902a );
 a28904a <=( a28903a  and  a28898a );
 a28908a <=( A167  and  (not A168) );
 a28909a <=( (not A169)  and  a28908a );
 a28913a <=( A201  and  A200 );
 a28914a <=( A166  and  a28913a );
 a28915a <=( a28914a  and  a28909a );
 a28919a <=( A236  and  A233 );
 a28920a <=( (not A232)  and  a28919a );
 a28924a <=( (not A302)  and  (not A301) );
 a28925a <=( (not A300)  and  a28924a );
 a28926a <=( a28925a  and  a28920a );
 a28930a <=( A167  and  (not A168) );
 a28931a <=( (not A169)  and  a28930a );
 a28935a <=( A201  and  A200 );
 a28936a <=( A166  and  a28935a );
 a28937a <=( a28936a  and  a28931a );
 a28941a <=( A236  and  A233 );
 a28942a <=( (not A232)  and  a28941a );
 a28946a <=( (not A301)  and  (not A299) );
 a28947a <=( (not A298)  and  a28946a );
 a28948a <=( a28947a  and  a28942a );
 a28952a <=( A167  and  (not A168) );
 a28953a <=( (not A169)  and  a28952a );
 a28957a <=( A201  and  A200 );
 a28958a <=( A166  and  a28957a );
 a28959a <=( a28958a  and  a28953a );
 a28963a <=( A236  and  A233 );
 a28964a <=( (not A232)  and  a28963a );
 a28968a <=( A269  and  A266 );
 a28969a <=( (not A265)  and  a28968a );
 a28970a <=( a28969a  and  a28964a );
 a28974a <=( A167  and  (not A168) );
 a28975a <=( (not A169)  and  a28974a );
 a28979a <=( A201  and  A200 );
 a28980a <=( A166  and  a28979a );
 a28981a <=( a28980a  and  a28975a );
 a28985a <=( A236  and  A233 );
 a28986a <=( (not A232)  and  a28985a );
 a28990a <=( A269  and  (not A266) );
 a28991a <=( A265  and  a28990a );
 a28992a <=( a28991a  and  a28986a );
 a28996a <=( A167  and  (not A168) );
 a28997a <=( (not A169)  and  a28996a );
 a29001a <=( A201  and  A200 );
 a29002a <=( A166  and  a29001a );
 a29003a <=( a29002a  and  a28997a );
 a29007a <=( A236  and  (not A233) );
 a29008a <=( A232  and  a29007a );
 a29012a <=( (not A302)  and  (not A301) );
 a29013a <=( (not A300)  and  a29012a );
 a29014a <=( a29013a  and  a29008a );
 a29018a <=( A167  and  (not A168) );
 a29019a <=( (not A169)  and  a29018a );
 a29023a <=( A201  and  A200 );
 a29024a <=( A166  and  a29023a );
 a29025a <=( a29024a  and  a29019a );
 a29029a <=( A236  and  (not A233) );
 a29030a <=( A232  and  a29029a );
 a29034a <=( (not A301)  and  (not A299) );
 a29035a <=( (not A298)  and  a29034a );
 a29036a <=( a29035a  and  a29030a );
 a29040a <=( A167  and  (not A168) );
 a29041a <=( (not A169)  and  a29040a );
 a29045a <=( A201  and  A200 );
 a29046a <=( A166  and  a29045a );
 a29047a <=( a29046a  and  a29041a );
 a29051a <=( A236  and  (not A233) );
 a29052a <=( A232  and  a29051a );
 a29056a <=( A269  and  A266 );
 a29057a <=( (not A265)  and  a29056a );
 a29058a <=( a29057a  and  a29052a );
 a29062a <=( A167  and  (not A168) );
 a29063a <=( (not A169)  and  a29062a );
 a29067a <=( A201  and  A200 );
 a29068a <=( A166  and  a29067a );
 a29069a <=( a29068a  and  a29063a );
 a29073a <=( A236  and  (not A233) );
 a29074a <=( A232  and  a29073a );
 a29078a <=( A269  and  (not A266) );
 a29079a <=( A265  and  a29078a );
 a29080a <=( a29079a  and  a29074a );
 a29084a <=( A167  and  (not A168) );
 a29085a <=( (not A169)  and  a29084a );
 a29089a <=( A200  and  (not A199) );
 a29090a <=( A166  and  a29089a );
 a29091a <=( a29090a  and  a29085a );
 a29095a <=( A298  and  A235 );
 a29096a <=( A203  and  a29095a );
 a29100a <=( (not A301)  and  (not A300) );
 a29101a <=( A299  and  a29100a );
 a29102a <=( a29101a  and  a29096a );
 a29106a <=( A167  and  (not A168) );
 a29107a <=( (not A169)  and  a29106a );
 a29111a <=( A200  and  (not A199) );
 a29112a <=( A166  and  a29111a );
 a29113a <=( a29112a  and  a29107a );
 a29117a <=( A234  and  A232 );
 a29118a <=( A203  and  a29117a );
 a29122a <=( (not A302)  and  (not A301) );
 a29123a <=( (not A300)  and  a29122a );
 a29124a <=( a29123a  and  a29118a );
 a29128a <=( A167  and  (not A168) );
 a29129a <=( (not A169)  and  a29128a );
 a29133a <=( A200  and  (not A199) );
 a29134a <=( A166  and  a29133a );
 a29135a <=( a29134a  and  a29129a );
 a29139a <=( A234  and  A232 );
 a29140a <=( A203  and  a29139a );
 a29144a <=( (not A301)  and  (not A299) );
 a29145a <=( (not A298)  and  a29144a );
 a29146a <=( a29145a  and  a29140a );
 a29150a <=( A167  and  (not A168) );
 a29151a <=( (not A169)  and  a29150a );
 a29155a <=( A200  and  (not A199) );
 a29156a <=( A166  and  a29155a );
 a29157a <=( a29156a  and  a29151a );
 a29161a <=( A234  and  A232 );
 a29162a <=( A203  and  a29161a );
 a29166a <=( A269  and  A266 );
 a29167a <=( (not A265)  and  a29166a );
 a29168a <=( a29167a  and  a29162a );
 a29172a <=( A167  and  (not A168) );
 a29173a <=( (not A169)  and  a29172a );
 a29177a <=( A200  and  (not A199) );
 a29178a <=( A166  and  a29177a );
 a29179a <=( a29178a  and  a29173a );
 a29183a <=( A234  and  A232 );
 a29184a <=( A203  and  a29183a );
 a29188a <=( A269  and  (not A266) );
 a29189a <=( A265  and  a29188a );
 a29190a <=( a29189a  and  a29184a );
 a29194a <=( A167  and  (not A168) );
 a29195a <=( (not A169)  and  a29194a );
 a29199a <=( A200  and  (not A199) );
 a29200a <=( A166  and  a29199a );
 a29201a <=( a29200a  and  a29195a );
 a29205a <=( A234  and  A233 );
 a29206a <=( A203  and  a29205a );
 a29210a <=( (not A302)  and  (not A301) );
 a29211a <=( (not A300)  and  a29210a );
 a29212a <=( a29211a  and  a29206a );
 a29216a <=( A167  and  (not A168) );
 a29217a <=( (not A169)  and  a29216a );
 a29221a <=( A200  and  (not A199) );
 a29222a <=( A166  and  a29221a );
 a29223a <=( a29222a  and  a29217a );
 a29227a <=( A234  and  A233 );
 a29228a <=( A203  and  a29227a );
 a29232a <=( (not A301)  and  (not A299) );
 a29233a <=( (not A298)  and  a29232a );
 a29234a <=( a29233a  and  a29228a );
 a29238a <=( A167  and  (not A168) );
 a29239a <=( (not A169)  and  a29238a );
 a29243a <=( A200  and  (not A199) );
 a29244a <=( A166  and  a29243a );
 a29245a <=( a29244a  and  a29239a );
 a29249a <=( A234  and  A233 );
 a29250a <=( A203  and  a29249a );
 a29254a <=( A269  and  A266 );
 a29255a <=( (not A265)  and  a29254a );
 a29256a <=( a29255a  and  a29250a );
 a29260a <=( A167  and  (not A168) );
 a29261a <=( (not A169)  and  a29260a );
 a29265a <=( A200  and  (not A199) );
 a29266a <=( A166  and  a29265a );
 a29267a <=( a29266a  and  a29261a );
 a29271a <=( A234  and  A233 );
 a29272a <=( A203  and  a29271a );
 a29276a <=( A269  and  (not A266) );
 a29277a <=( A265  and  a29276a );
 a29278a <=( a29277a  and  a29272a );
 a29282a <=( A167  and  (not A168) );
 a29283a <=( (not A169)  and  a29282a );
 a29287a <=( A200  and  (not A199) );
 a29288a <=( A166  and  a29287a );
 a29289a <=( a29288a  and  a29283a );
 a29293a <=( A233  and  (not A232) );
 a29294a <=( A203  and  a29293a );
 a29298a <=( A267  and  A265 );
 a29299a <=( A236  and  a29298a );
 a29300a <=( a29299a  and  a29294a );
 a29304a <=( A167  and  (not A168) );
 a29305a <=( (not A169)  and  a29304a );
 a29309a <=( A200  and  (not A199) );
 a29310a <=( A166  and  a29309a );
 a29311a <=( a29310a  and  a29305a );
 a29315a <=( A233  and  (not A232) );
 a29316a <=( A203  and  a29315a );
 a29320a <=( A267  and  A266 );
 a29321a <=( A236  and  a29320a );
 a29322a <=( a29321a  and  a29316a );
 a29326a <=( A167  and  (not A168) );
 a29327a <=( (not A169)  and  a29326a );
 a29331a <=( A200  and  (not A199) );
 a29332a <=( A166  and  a29331a );
 a29333a <=( a29332a  and  a29327a );
 a29337a <=( (not A233)  and  A232 );
 a29338a <=( A203  and  a29337a );
 a29342a <=( A267  and  A265 );
 a29343a <=( A236  and  a29342a );
 a29344a <=( a29343a  and  a29338a );
 a29348a <=( A167  and  (not A168) );
 a29349a <=( (not A169)  and  a29348a );
 a29353a <=( A200  and  (not A199) );
 a29354a <=( A166  and  a29353a );
 a29355a <=( a29354a  and  a29349a );
 a29359a <=( (not A233)  and  A232 );
 a29360a <=( A203  and  a29359a );
 a29364a <=( A267  and  A266 );
 a29365a <=( A236  and  a29364a );
 a29366a <=( a29365a  and  a29360a );
 a29370a <=( A167  and  (not A168) );
 a29371a <=( (not A169)  and  a29370a );
 a29375a <=( (not A200)  and  A199 );
 a29376a <=( A166  and  a29375a );
 a29377a <=( a29376a  and  a29371a );
 a29381a <=( A298  and  A235 );
 a29382a <=( A203  and  a29381a );
 a29386a <=( (not A301)  and  (not A300) );
 a29387a <=( A299  and  a29386a );
 a29388a <=( a29387a  and  a29382a );
 a29392a <=( A167  and  (not A168) );
 a29393a <=( (not A169)  and  a29392a );
 a29397a <=( (not A200)  and  A199 );
 a29398a <=( A166  and  a29397a );
 a29399a <=( a29398a  and  a29393a );
 a29403a <=( A234  and  A232 );
 a29404a <=( A203  and  a29403a );
 a29408a <=( (not A302)  and  (not A301) );
 a29409a <=( (not A300)  and  a29408a );
 a29410a <=( a29409a  and  a29404a );
 a29414a <=( A167  and  (not A168) );
 a29415a <=( (not A169)  and  a29414a );
 a29419a <=( (not A200)  and  A199 );
 a29420a <=( A166  and  a29419a );
 a29421a <=( a29420a  and  a29415a );
 a29425a <=( A234  and  A232 );
 a29426a <=( A203  and  a29425a );
 a29430a <=( (not A301)  and  (not A299) );
 a29431a <=( (not A298)  and  a29430a );
 a29432a <=( a29431a  and  a29426a );
 a29436a <=( A167  and  (not A168) );
 a29437a <=( (not A169)  and  a29436a );
 a29441a <=( (not A200)  and  A199 );
 a29442a <=( A166  and  a29441a );
 a29443a <=( a29442a  and  a29437a );
 a29447a <=( A234  and  A232 );
 a29448a <=( A203  and  a29447a );
 a29452a <=( A269  and  A266 );
 a29453a <=( (not A265)  and  a29452a );
 a29454a <=( a29453a  and  a29448a );
 a29458a <=( A167  and  (not A168) );
 a29459a <=( (not A169)  and  a29458a );
 a29463a <=( (not A200)  and  A199 );
 a29464a <=( A166  and  a29463a );
 a29465a <=( a29464a  and  a29459a );
 a29469a <=( A234  and  A232 );
 a29470a <=( A203  and  a29469a );
 a29474a <=( A269  and  (not A266) );
 a29475a <=( A265  and  a29474a );
 a29476a <=( a29475a  and  a29470a );
 a29480a <=( A167  and  (not A168) );
 a29481a <=( (not A169)  and  a29480a );
 a29485a <=( (not A200)  and  A199 );
 a29486a <=( A166  and  a29485a );
 a29487a <=( a29486a  and  a29481a );
 a29491a <=( A234  and  A233 );
 a29492a <=( A203  and  a29491a );
 a29496a <=( (not A302)  and  (not A301) );
 a29497a <=( (not A300)  and  a29496a );
 a29498a <=( a29497a  and  a29492a );
 a29502a <=( A167  and  (not A168) );
 a29503a <=( (not A169)  and  a29502a );
 a29507a <=( (not A200)  and  A199 );
 a29508a <=( A166  and  a29507a );
 a29509a <=( a29508a  and  a29503a );
 a29513a <=( A234  and  A233 );
 a29514a <=( A203  and  a29513a );
 a29518a <=( (not A301)  and  (not A299) );
 a29519a <=( (not A298)  and  a29518a );
 a29520a <=( a29519a  and  a29514a );
 a29524a <=( A167  and  (not A168) );
 a29525a <=( (not A169)  and  a29524a );
 a29529a <=( (not A200)  and  A199 );
 a29530a <=( A166  and  a29529a );
 a29531a <=( a29530a  and  a29525a );
 a29535a <=( A234  and  A233 );
 a29536a <=( A203  and  a29535a );
 a29540a <=( A269  and  A266 );
 a29541a <=( (not A265)  and  a29540a );
 a29542a <=( a29541a  and  a29536a );
 a29546a <=( A167  and  (not A168) );
 a29547a <=( (not A169)  and  a29546a );
 a29551a <=( (not A200)  and  A199 );
 a29552a <=( A166  and  a29551a );
 a29553a <=( a29552a  and  a29547a );
 a29557a <=( A234  and  A233 );
 a29558a <=( A203  and  a29557a );
 a29562a <=( A269  and  (not A266) );
 a29563a <=( A265  and  a29562a );
 a29564a <=( a29563a  and  a29558a );
 a29568a <=( A167  and  (not A168) );
 a29569a <=( (not A169)  and  a29568a );
 a29573a <=( (not A200)  and  A199 );
 a29574a <=( A166  and  a29573a );
 a29575a <=( a29574a  and  a29569a );
 a29579a <=( A233  and  (not A232) );
 a29580a <=( A203  and  a29579a );
 a29584a <=( A267  and  A265 );
 a29585a <=( A236  and  a29584a );
 a29586a <=( a29585a  and  a29580a );
 a29590a <=( A167  and  (not A168) );
 a29591a <=( (not A169)  and  a29590a );
 a29595a <=( (not A200)  and  A199 );
 a29596a <=( A166  and  a29595a );
 a29597a <=( a29596a  and  a29591a );
 a29601a <=( A233  and  (not A232) );
 a29602a <=( A203  and  a29601a );
 a29606a <=( A267  and  A266 );
 a29607a <=( A236  and  a29606a );
 a29608a <=( a29607a  and  a29602a );
 a29612a <=( A167  and  (not A168) );
 a29613a <=( (not A169)  and  a29612a );
 a29617a <=( (not A200)  and  A199 );
 a29618a <=( A166  and  a29617a );
 a29619a <=( a29618a  and  a29613a );
 a29623a <=( (not A233)  and  A232 );
 a29624a <=( A203  and  a29623a );
 a29628a <=( A267  and  A265 );
 a29629a <=( A236  and  a29628a );
 a29630a <=( a29629a  and  a29624a );
 a29634a <=( A167  and  (not A168) );
 a29635a <=( (not A169)  and  a29634a );
 a29639a <=( (not A200)  and  A199 );
 a29640a <=( A166  and  a29639a );
 a29641a <=( a29640a  and  a29635a );
 a29645a <=( (not A233)  and  A232 );
 a29646a <=( A203  and  a29645a );
 a29650a <=( A267  and  A266 );
 a29651a <=( A236  and  a29650a );
 a29652a <=( a29651a  and  a29646a );
 a29656a <=( (not A168)  and  (not A169) );
 a29657a <=( (not A170)  and  a29656a );
 a29661a <=( (not A235)  and  (not A234) );
 a29662a <=( A202  and  a29661a );
 a29663a <=( a29662a  and  a29657a );
 a29667a <=( (not A268)  and  (not A267) );
 a29668a <=( (not A236)  and  a29667a );
 a29672a <=( A300  and  A299 );
 a29673a <=( (not A269)  and  a29672a );
 a29674a <=( a29673a  and  a29668a );
 a29678a <=( (not A168)  and  (not A169) );
 a29679a <=( (not A170)  and  a29678a );
 a29683a <=( (not A235)  and  (not A234) );
 a29684a <=( A202  and  a29683a );
 a29685a <=( a29684a  and  a29679a );
 a29689a <=( (not A268)  and  (not A267) );
 a29690a <=( (not A236)  and  a29689a );
 a29694a <=( A300  and  A298 );
 a29695a <=( (not A269)  and  a29694a );
 a29696a <=( a29695a  and  a29690a );
 a29700a <=( (not A168)  and  (not A169) );
 a29701a <=( (not A170)  and  a29700a );
 a29705a <=( (not A235)  and  (not A234) );
 a29706a <=( A202  and  a29705a );
 a29707a <=( a29706a  and  a29701a );
 a29711a <=( A266  and  A265 );
 a29712a <=( (not A236)  and  a29711a );
 a29716a <=( A301  and  (not A268) );
 a29717a <=( (not A267)  and  a29716a );
 a29718a <=( a29717a  and  a29712a );
 a29722a <=( (not A168)  and  (not A169) );
 a29723a <=( (not A170)  and  a29722a );
 a29727a <=( (not A235)  and  (not A234) );
 a29728a <=( A202  and  a29727a );
 a29729a <=( a29728a  and  a29723a );
 a29733a <=( (not A266)  and  (not A265) );
 a29734a <=( (not A236)  and  a29733a );
 a29738a <=( A300  and  A299 );
 a29739a <=( (not A268)  and  a29738a );
 a29740a <=( a29739a  and  a29734a );
 a29744a <=( (not A168)  and  (not A169) );
 a29745a <=( (not A170)  and  a29744a );
 a29749a <=( (not A235)  and  (not A234) );
 a29750a <=( A202  and  a29749a );
 a29751a <=( a29750a  and  a29745a );
 a29755a <=( (not A266)  and  (not A265) );
 a29756a <=( (not A236)  and  a29755a );
 a29760a <=( A300  and  A298 );
 a29761a <=( (not A268)  and  a29760a );
 a29762a <=( a29761a  and  a29756a );
 a29766a <=( (not A168)  and  (not A169) );
 a29767a <=( (not A170)  and  a29766a );
 a29771a <=( A233  and  A232 );
 a29772a <=( A202  and  a29771a );
 a29773a <=( a29772a  and  a29767a );
 a29777a <=( (not A267)  and  (not A235) );
 a29778a <=( (not A234)  and  a29777a );
 a29782a <=( A301  and  (not A269) );
 a29783a <=( (not A268)  and  a29782a );
 a29784a <=( a29783a  and  a29778a );
 a29788a <=( (not A168)  and  (not A169) );
 a29789a <=( (not A170)  and  a29788a );
 a29793a <=( A233  and  A232 );
 a29794a <=( A202  and  a29793a );
 a29795a <=( a29794a  and  a29789a );
 a29799a <=( (not A265)  and  (not A235) );
 a29800a <=( (not A234)  and  a29799a );
 a29804a <=( A301  and  (not A268) );
 a29805a <=( (not A266)  and  a29804a );
 a29806a <=( a29805a  and  a29800a );
 a29810a <=( (not A168)  and  (not A169) );
 a29811a <=( (not A170)  and  a29810a );
 a29815a <=( (not A233)  and  (not A232) );
 a29816a <=( A202  and  a29815a );
 a29817a <=( a29816a  and  a29811a );
 a29821a <=( (not A268)  and  (not A267) );
 a29822a <=( (not A235)  and  a29821a );
 a29826a <=( A300  and  A299 );
 a29827a <=( (not A269)  and  a29826a );
 a29828a <=( a29827a  and  a29822a );
 a29832a <=( (not A168)  and  (not A169) );
 a29833a <=( (not A170)  and  a29832a );
 a29837a <=( (not A233)  and  (not A232) );
 a29838a <=( A202  and  a29837a );
 a29839a <=( a29838a  and  a29833a );
 a29843a <=( (not A268)  and  (not A267) );
 a29844a <=( (not A235)  and  a29843a );
 a29848a <=( A300  and  A298 );
 a29849a <=( (not A269)  and  a29848a );
 a29850a <=( a29849a  and  a29844a );
 a29854a <=( (not A168)  and  (not A169) );
 a29855a <=( (not A170)  and  a29854a );
 a29859a <=( (not A233)  and  (not A232) );
 a29860a <=( A202  and  a29859a );
 a29861a <=( a29860a  and  a29855a );
 a29865a <=( A266  and  A265 );
 a29866a <=( (not A235)  and  a29865a );
 a29870a <=( A301  and  (not A268) );
 a29871a <=( (not A267)  and  a29870a );
 a29872a <=( a29871a  and  a29866a );
 a29876a <=( (not A168)  and  (not A169) );
 a29877a <=( (not A170)  and  a29876a );
 a29881a <=( (not A233)  and  (not A232) );
 a29882a <=( A202  and  a29881a );
 a29883a <=( a29882a  and  a29877a );
 a29887a <=( (not A266)  and  (not A265) );
 a29888a <=( (not A235)  and  a29887a );
 a29892a <=( A300  and  A299 );
 a29893a <=( (not A268)  and  a29892a );
 a29894a <=( a29893a  and  a29888a );
 a29898a <=( (not A168)  and  (not A169) );
 a29899a <=( (not A170)  and  a29898a );
 a29903a <=( (not A233)  and  (not A232) );
 a29904a <=( A202  and  a29903a );
 a29905a <=( a29904a  and  a29899a );
 a29909a <=( (not A266)  and  (not A265) );
 a29910a <=( (not A235)  and  a29909a );
 a29914a <=( A300  and  A298 );
 a29915a <=( (not A268)  and  a29914a );
 a29916a <=( a29915a  and  a29910a );
 a29920a <=( (not A168)  and  (not A169) );
 a29921a <=( (not A170)  and  a29920a );
 a29925a <=( (not A234)  and  A201 );
 a29926a <=( A199  and  a29925a );
 a29927a <=( a29926a  and  a29921a );
 a29931a <=( (not A267)  and  (not A236) );
 a29932a <=( (not A235)  and  a29931a );
 a29936a <=( A301  and  (not A269) );
 a29937a <=( (not A268)  and  a29936a );
 a29938a <=( a29937a  and  a29932a );
 a29942a <=( (not A168)  and  (not A169) );
 a29943a <=( (not A170)  and  a29942a );
 a29947a <=( (not A234)  and  A201 );
 a29948a <=( A199  and  a29947a );
 a29949a <=( a29948a  and  a29943a );
 a29953a <=( (not A265)  and  (not A236) );
 a29954a <=( (not A235)  and  a29953a );
 a29958a <=( A301  and  (not A268) );
 a29959a <=( (not A266)  and  a29958a );
 a29960a <=( a29959a  and  a29954a );
 a29964a <=( (not A168)  and  (not A169) );
 a29965a <=( (not A170)  and  a29964a );
 a29969a <=( (not A232)  and  A201 );
 a29970a <=( A199  and  a29969a );
 a29971a <=( a29970a  and  a29965a );
 a29975a <=( A298  and  A236 );
 a29976a <=( A233  and  a29975a );
 a29980a <=( (not A301)  and  (not A300) );
 a29981a <=( A299  and  a29980a );
 a29982a <=( a29981a  and  a29976a );
 a29986a <=( (not A168)  and  (not A169) );
 a29987a <=( (not A170)  and  a29986a );
 a29991a <=( A232  and  A201 );
 a29992a <=( A199  and  a29991a );
 a29993a <=( a29992a  and  a29987a );
 a29997a <=( A298  and  A236 );
 a29998a <=( (not A233)  and  a29997a );
 a30002a <=( (not A301)  and  (not A300) );
 a30003a <=( A299  and  a30002a );
 a30004a <=( a30003a  and  a29998a );
 a30008a <=( (not A168)  and  (not A169) );
 a30009a <=( (not A170)  and  a30008a );
 a30013a <=( (not A232)  and  A201 );
 a30014a <=( A199  and  a30013a );
 a30015a <=( a30014a  and  a30009a );
 a30019a <=( (not A267)  and  (not A235) );
 a30020a <=( (not A233)  and  a30019a );
 a30024a <=( A301  and  (not A269) );
 a30025a <=( (not A268)  and  a30024a );
 a30026a <=( a30025a  and  a30020a );
 a30030a <=( (not A168)  and  (not A169) );
 a30031a <=( (not A170)  and  a30030a );
 a30035a <=( (not A232)  and  A201 );
 a30036a <=( A199  and  a30035a );
 a30037a <=( a30036a  and  a30031a );
 a30041a <=( (not A265)  and  (not A235) );
 a30042a <=( (not A233)  and  a30041a );
 a30046a <=( A301  and  (not A268) );
 a30047a <=( (not A266)  and  a30046a );
 a30048a <=( a30047a  and  a30042a );
 a30052a <=( (not A168)  and  (not A169) );
 a30053a <=( (not A170)  and  a30052a );
 a30057a <=( (not A234)  and  A201 );
 a30058a <=( A200  and  a30057a );
 a30059a <=( a30058a  and  a30053a );
 a30063a <=( (not A267)  and  (not A236) );
 a30064a <=( (not A235)  and  a30063a );
 a30068a <=( A301  and  (not A269) );
 a30069a <=( (not A268)  and  a30068a );
 a30070a <=( a30069a  and  a30064a );
 a30074a <=( (not A168)  and  (not A169) );
 a30075a <=( (not A170)  and  a30074a );
 a30079a <=( (not A234)  and  A201 );
 a30080a <=( A200  and  a30079a );
 a30081a <=( a30080a  and  a30075a );
 a30085a <=( (not A265)  and  (not A236) );
 a30086a <=( (not A235)  and  a30085a );
 a30090a <=( A301  and  (not A268) );
 a30091a <=( (not A266)  and  a30090a );
 a30092a <=( a30091a  and  a30086a );
 a30096a <=( (not A168)  and  (not A169) );
 a30097a <=( (not A170)  and  a30096a );
 a30101a <=( (not A232)  and  A201 );
 a30102a <=( A200  and  a30101a );
 a30103a <=( a30102a  and  a30097a );
 a30107a <=( A298  and  A236 );
 a30108a <=( A233  and  a30107a );
 a30112a <=( (not A301)  and  (not A300) );
 a30113a <=( A299  and  a30112a );
 a30114a <=( a30113a  and  a30108a );
 a30118a <=( (not A168)  and  (not A169) );
 a30119a <=( (not A170)  and  a30118a );
 a30123a <=( A232  and  A201 );
 a30124a <=( A200  and  a30123a );
 a30125a <=( a30124a  and  a30119a );
 a30129a <=( A298  and  A236 );
 a30130a <=( (not A233)  and  a30129a );
 a30134a <=( (not A301)  and  (not A300) );
 a30135a <=( A299  and  a30134a );
 a30136a <=( a30135a  and  a30130a );
 a30140a <=( (not A168)  and  (not A169) );
 a30141a <=( (not A170)  and  a30140a );
 a30145a <=( (not A232)  and  A201 );
 a30146a <=( A200  and  a30145a );
 a30147a <=( a30146a  and  a30141a );
 a30151a <=( (not A267)  and  (not A235) );
 a30152a <=( (not A233)  and  a30151a );
 a30156a <=( A301  and  (not A269) );
 a30157a <=( (not A268)  and  a30156a );
 a30158a <=( a30157a  and  a30152a );
 a30162a <=( (not A168)  and  (not A169) );
 a30163a <=( (not A170)  and  a30162a );
 a30167a <=( (not A232)  and  A201 );
 a30168a <=( A200  and  a30167a );
 a30169a <=( a30168a  and  a30163a );
 a30173a <=( (not A265)  and  (not A235) );
 a30174a <=( (not A233)  and  a30173a );
 a30178a <=( A301  and  (not A268) );
 a30179a <=( (not A266)  and  a30178a );
 a30180a <=( a30179a  and  a30174a );
 a30184a <=( (not A168)  and  (not A169) );
 a30185a <=( (not A170)  and  a30184a );
 a30189a <=( A203  and  A200 );
 a30190a <=( (not A199)  and  a30189a );
 a30191a <=( a30190a  and  a30185a );
 a30195a <=( A298  and  A234 );
 a30196a <=( A232  and  a30195a );
 a30200a <=( (not A301)  and  (not A300) );
 a30201a <=( A299  and  a30200a );
 a30202a <=( a30201a  and  a30196a );
 a30206a <=( (not A168)  and  (not A169) );
 a30207a <=( (not A170)  and  a30206a );
 a30211a <=( A203  and  A200 );
 a30212a <=( (not A199)  and  a30211a );
 a30213a <=( a30212a  and  a30207a );
 a30217a <=( A298  and  A234 );
 a30218a <=( A233  and  a30217a );
 a30222a <=( (not A301)  and  (not A300) );
 a30223a <=( A299  and  a30222a );
 a30224a <=( a30223a  and  a30218a );
 a30228a <=( (not A168)  and  (not A169) );
 a30229a <=( (not A170)  and  a30228a );
 a30233a <=( A203  and  A200 );
 a30234a <=( (not A199)  and  a30233a );
 a30235a <=( a30234a  and  a30229a );
 a30239a <=( A236  and  A233 );
 a30240a <=( (not A232)  and  a30239a );
 a30244a <=( (not A302)  and  (not A301) );
 a30245a <=( (not A300)  and  a30244a );
 a30246a <=( a30245a  and  a30240a );
 a30250a <=( (not A168)  and  (not A169) );
 a30251a <=( (not A170)  and  a30250a );
 a30255a <=( A203  and  A200 );
 a30256a <=( (not A199)  and  a30255a );
 a30257a <=( a30256a  and  a30251a );
 a30261a <=( A236  and  A233 );
 a30262a <=( (not A232)  and  a30261a );
 a30266a <=( (not A301)  and  (not A299) );
 a30267a <=( (not A298)  and  a30266a );
 a30268a <=( a30267a  and  a30262a );
 a30272a <=( (not A168)  and  (not A169) );
 a30273a <=( (not A170)  and  a30272a );
 a30277a <=( A203  and  A200 );
 a30278a <=( (not A199)  and  a30277a );
 a30279a <=( a30278a  and  a30273a );
 a30283a <=( A236  and  A233 );
 a30284a <=( (not A232)  and  a30283a );
 a30288a <=( A269  and  A266 );
 a30289a <=( (not A265)  and  a30288a );
 a30290a <=( a30289a  and  a30284a );
 a30294a <=( (not A168)  and  (not A169) );
 a30295a <=( (not A170)  and  a30294a );
 a30299a <=( A203  and  A200 );
 a30300a <=( (not A199)  and  a30299a );
 a30301a <=( a30300a  and  a30295a );
 a30305a <=( A236  and  A233 );
 a30306a <=( (not A232)  and  a30305a );
 a30310a <=( A269  and  (not A266) );
 a30311a <=( A265  and  a30310a );
 a30312a <=( a30311a  and  a30306a );
 a30316a <=( (not A168)  and  (not A169) );
 a30317a <=( (not A170)  and  a30316a );
 a30321a <=( A203  and  A200 );
 a30322a <=( (not A199)  and  a30321a );
 a30323a <=( a30322a  and  a30317a );
 a30327a <=( A236  and  (not A233) );
 a30328a <=( A232  and  a30327a );
 a30332a <=( (not A302)  and  (not A301) );
 a30333a <=( (not A300)  and  a30332a );
 a30334a <=( a30333a  and  a30328a );
 a30338a <=( (not A168)  and  (not A169) );
 a30339a <=( (not A170)  and  a30338a );
 a30343a <=( A203  and  A200 );
 a30344a <=( (not A199)  and  a30343a );
 a30345a <=( a30344a  and  a30339a );
 a30349a <=( A236  and  (not A233) );
 a30350a <=( A232  and  a30349a );
 a30354a <=( (not A301)  and  (not A299) );
 a30355a <=( (not A298)  and  a30354a );
 a30356a <=( a30355a  and  a30350a );
 a30360a <=( (not A168)  and  (not A169) );
 a30361a <=( (not A170)  and  a30360a );
 a30365a <=( A203  and  A200 );
 a30366a <=( (not A199)  and  a30365a );
 a30367a <=( a30366a  and  a30361a );
 a30371a <=( A236  and  (not A233) );
 a30372a <=( A232  and  a30371a );
 a30376a <=( A269  and  A266 );
 a30377a <=( (not A265)  and  a30376a );
 a30378a <=( a30377a  and  a30372a );
 a30382a <=( (not A168)  and  (not A169) );
 a30383a <=( (not A170)  and  a30382a );
 a30387a <=( A203  and  A200 );
 a30388a <=( (not A199)  and  a30387a );
 a30389a <=( a30388a  and  a30383a );
 a30393a <=( A236  and  (not A233) );
 a30394a <=( A232  and  a30393a );
 a30398a <=( A269  and  (not A266) );
 a30399a <=( A265  and  a30398a );
 a30400a <=( a30399a  and  a30394a );
 a30404a <=( (not A168)  and  (not A169) );
 a30405a <=( (not A170)  and  a30404a );
 a30409a <=( A203  and  (not A200) );
 a30410a <=( A199  and  a30409a );
 a30411a <=( a30410a  and  a30405a );
 a30415a <=( A298  and  A234 );
 a30416a <=( A232  and  a30415a );
 a30420a <=( (not A301)  and  (not A300) );
 a30421a <=( A299  and  a30420a );
 a30422a <=( a30421a  and  a30416a );
 a30426a <=( (not A168)  and  (not A169) );
 a30427a <=( (not A170)  and  a30426a );
 a30431a <=( A203  and  (not A200) );
 a30432a <=( A199  and  a30431a );
 a30433a <=( a30432a  and  a30427a );
 a30437a <=( A298  and  A234 );
 a30438a <=( A233  and  a30437a );
 a30442a <=( (not A301)  and  (not A300) );
 a30443a <=( A299  and  a30442a );
 a30444a <=( a30443a  and  a30438a );
 a30448a <=( (not A168)  and  (not A169) );
 a30449a <=( (not A170)  and  a30448a );
 a30453a <=( A203  and  (not A200) );
 a30454a <=( A199  and  a30453a );
 a30455a <=( a30454a  and  a30449a );
 a30459a <=( A236  and  A233 );
 a30460a <=( (not A232)  and  a30459a );
 a30464a <=( (not A302)  and  (not A301) );
 a30465a <=( (not A300)  and  a30464a );
 a30466a <=( a30465a  and  a30460a );
 a30470a <=( (not A168)  and  (not A169) );
 a30471a <=( (not A170)  and  a30470a );
 a30475a <=( A203  and  (not A200) );
 a30476a <=( A199  and  a30475a );
 a30477a <=( a30476a  and  a30471a );
 a30481a <=( A236  and  A233 );
 a30482a <=( (not A232)  and  a30481a );
 a30486a <=( (not A301)  and  (not A299) );
 a30487a <=( (not A298)  and  a30486a );
 a30488a <=( a30487a  and  a30482a );
 a30492a <=( (not A168)  and  (not A169) );
 a30493a <=( (not A170)  and  a30492a );
 a30497a <=( A203  and  (not A200) );
 a30498a <=( A199  and  a30497a );
 a30499a <=( a30498a  and  a30493a );
 a30503a <=( A236  and  A233 );
 a30504a <=( (not A232)  and  a30503a );
 a30508a <=( A269  and  A266 );
 a30509a <=( (not A265)  and  a30508a );
 a30510a <=( a30509a  and  a30504a );
 a30514a <=( (not A168)  and  (not A169) );
 a30515a <=( (not A170)  and  a30514a );
 a30519a <=( A203  and  (not A200) );
 a30520a <=( A199  and  a30519a );
 a30521a <=( a30520a  and  a30515a );
 a30525a <=( A236  and  A233 );
 a30526a <=( (not A232)  and  a30525a );
 a30530a <=( A269  and  (not A266) );
 a30531a <=( A265  and  a30530a );
 a30532a <=( a30531a  and  a30526a );
 a30536a <=( (not A168)  and  (not A169) );
 a30537a <=( (not A170)  and  a30536a );
 a30541a <=( A203  and  (not A200) );
 a30542a <=( A199  and  a30541a );
 a30543a <=( a30542a  and  a30537a );
 a30547a <=( A236  and  (not A233) );
 a30548a <=( A232  and  a30547a );
 a30552a <=( (not A302)  and  (not A301) );
 a30553a <=( (not A300)  and  a30552a );
 a30554a <=( a30553a  and  a30548a );
 a30558a <=( (not A168)  and  (not A169) );
 a30559a <=( (not A170)  and  a30558a );
 a30563a <=( A203  and  (not A200) );
 a30564a <=( A199  and  a30563a );
 a30565a <=( a30564a  and  a30559a );
 a30569a <=( A236  and  (not A233) );
 a30570a <=( A232  and  a30569a );
 a30574a <=( (not A301)  and  (not A299) );
 a30575a <=( (not A298)  and  a30574a );
 a30576a <=( a30575a  and  a30570a );
 a30580a <=( (not A168)  and  (not A169) );
 a30581a <=( (not A170)  and  a30580a );
 a30585a <=( A203  and  (not A200) );
 a30586a <=( A199  and  a30585a );
 a30587a <=( a30586a  and  a30581a );
 a30591a <=( A236  and  (not A233) );
 a30592a <=( A232  and  a30591a );
 a30596a <=( A269  and  A266 );
 a30597a <=( (not A265)  and  a30596a );
 a30598a <=( a30597a  and  a30592a );
 a30602a <=( (not A168)  and  (not A169) );
 a30603a <=( (not A170)  and  a30602a );
 a30607a <=( A203  and  (not A200) );
 a30608a <=( A199  and  a30607a );
 a30609a <=( a30608a  and  a30603a );
 a30613a <=( A236  and  (not A233) );
 a30614a <=( A232  and  a30613a );
 a30618a <=( A269  and  (not A266) );
 a30619a <=( A265  and  a30618a );
 a30620a <=( a30619a  and  a30614a );
 a30624a <=( (not A201)  and  A166 );
 a30625a <=( A168  and  a30624a );
 a30629a <=( (not A234)  and  (not A203) );
 a30630a <=( (not A202)  and  a30629a );
 a30631a <=( a30630a  and  a30625a );
 a30635a <=( (not A267)  and  (not A236) );
 a30636a <=( (not A235)  and  a30635a );
 a30639a <=( (not A269)  and  (not A268) );
 a30642a <=( A300  and  A299 );
 a30643a <=( a30642a  and  a30639a );
 a30644a <=( a30643a  and  a30636a );
 a30648a <=( (not A201)  and  A166 );
 a30649a <=( A168  and  a30648a );
 a30653a <=( (not A234)  and  (not A203) );
 a30654a <=( (not A202)  and  a30653a );
 a30655a <=( a30654a  and  a30649a );
 a30659a <=( (not A267)  and  (not A236) );
 a30660a <=( (not A235)  and  a30659a );
 a30663a <=( (not A269)  and  (not A268) );
 a30666a <=( A300  and  A298 );
 a30667a <=( a30666a  and  a30663a );
 a30668a <=( a30667a  and  a30660a );
 a30672a <=( (not A201)  and  A166 );
 a30673a <=( A168  and  a30672a );
 a30677a <=( (not A234)  and  (not A203) );
 a30678a <=( (not A202)  and  a30677a );
 a30679a <=( a30678a  and  a30673a );
 a30683a <=( A265  and  (not A236) );
 a30684a <=( (not A235)  and  a30683a );
 a30687a <=( (not A267)  and  A266 );
 a30690a <=( A301  and  (not A268) );
 a30691a <=( a30690a  and  a30687a );
 a30692a <=( a30691a  and  a30684a );
 a30696a <=( (not A201)  and  A166 );
 a30697a <=( A168  and  a30696a );
 a30701a <=( (not A234)  and  (not A203) );
 a30702a <=( (not A202)  and  a30701a );
 a30703a <=( a30702a  and  a30697a );
 a30707a <=( (not A265)  and  (not A236) );
 a30708a <=( (not A235)  and  a30707a );
 a30711a <=( (not A268)  and  (not A266) );
 a30714a <=( A300  and  A299 );
 a30715a <=( a30714a  and  a30711a );
 a30716a <=( a30715a  and  a30708a );
 a30720a <=( (not A201)  and  A166 );
 a30721a <=( A168  and  a30720a );
 a30725a <=( (not A234)  and  (not A203) );
 a30726a <=( (not A202)  and  a30725a );
 a30727a <=( a30726a  and  a30721a );
 a30731a <=( (not A265)  and  (not A236) );
 a30732a <=( (not A235)  and  a30731a );
 a30735a <=( (not A268)  and  (not A266) );
 a30738a <=( A300  and  A298 );
 a30739a <=( a30738a  and  a30735a );
 a30740a <=( a30739a  and  a30732a );
 a30744a <=( (not A201)  and  A166 );
 a30745a <=( A168  and  a30744a );
 a30749a <=( A232  and  (not A203) );
 a30750a <=( (not A202)  and  a30749a );
 a30751a <=( a30750a  and  a30745a );
 a30755a <=( (not A235)  and  (not A234) );
 a30756a <=( A233  and  a30755a );
 a30759a <=( (not A268)  and  (not A267) );
 a30762a <=( A301  and  (not A269) );
 a30763a <=( a30762a  and  a30759a );
 a30764a <=( a30763a  and  a30756a );
 a30768a <=( (not A201)  and  A166 );
 a30769a <=( A168  and  a30768a );
 a30773a <=( A232  and  (not A203) );
 a30774a <=( (not A202)  and  a30773a );
 a30775a <=( a30774a  and  a30769a );
 a30779a <=( (not A235)  and  (not A234) );
 a30780a <=( A233  and  a30779a );
 a30783a <=( (not A266)  and  (not A265) );
 a30786a <=( A301  and  (not A268) );
 a30787a <=( a30786a  and  a30783a );
 a30788a <=( a30787a  and  a30780a );
 a30792a <=( (not A201)  and  A166 );
 a30793a <=( A168  and  a30792a );
 a30797a <=( (not A232)  and  (not A203) );
 a30798a <=( (not A202)  and  a30797a );
 a30799a <=( a30798a  and  a30793a );
 a30803a <=( (not A267)  and  (not A235) );
 a30804a <=( (not A233)  and  a30803a );
 a30807a <=( (not A269)  and  (not A268) );
 a30810a <=( A300  and  A299 );
 a30811a <=( a30810a  and  a30807a );
 a30812a <=( a30811a  and  a30804a );
 a30816a <=( (not A201)  and  A166 );
 a30817a <=( A168  and  a30816a );
 a30821a <=( (not A232)  and  (not A203) );
 a30822a <=( (not A202)  and  a30821a );
 a30823a <=( a30822a  and  a30817a );
 a30827a <=( (not A267)  and  (not A235) );
 a30828a <=( (not A233)  and  a30827a );
 a30831a <=( (not A269)  and  (not A268) );
 a30834a <=( A300  and  A298 );
 a30835a <=( a30834a  and  a30831a );
 a30836a <=( a30835a  and  a30828a );
 a30840a <=( (not A201)  and  A166 );
 a30841a <=( A168  and  a30840a );
 a30845a <=( (not A232)  and  (not A203) );
 a30846a <=( (not A202)  and  a30845a );
 a30847a <=( a30846a  and  a30841a );
 a30851a <=( A265  and  (not A235) );
 a30852a <=( (not A233)  and  a30851a );
 a30855a <=( (not A267)  and  A266 );
 a30858a <=( A301  and  (not A268) );
 a30859a <=( a30858a  and  a30855a );
 a30860a <=( a30859a  and  a30852a );
 a30864a <=( (not A201)  and  A166 );
 a30865a <=( A168  and  a30864a );
 a30869a <=( (not A232)  and  (not A203) );
 a30870a <=( (not A202)  and  a30869a );
 a30871a <=( a30870a  and  a30865a );
 a30875a <=( (not A265)  and  (not A235) );
 a30876a <=( (not A233)  and  a30875a );
 a30879a <=( (not A268)  and  (not A266) );
 a30882a <=( A300  and  A299 );
 a30883a <=( a30882a  and  a30879a );
 a30884a <=( a30883a  and  a30876a );
 a30888a <=( (not A201)  and  A166 );
 a30889a <=( A168  and  a30888a );
 a30893a <=( (not A232)  and  (not A203) );
 a30894a <=( (not A202)  and  a30893a );
 a30895a <=( a30894a  and  a30889a );
 a30899a <=( (not A265)  and  (not A235) );
 a30900a <=( (not A233)  and  a30899a );
 a30903a <=( (not A268)  and  (not A266) );
 a30906a <=( A300  and  A298 );
 a30907a <=( a30906a  and  a30903a );
 a30908a <=( a30907a  and  a30900a );
 a30912a <=( A199  and  A166 );
 a30913a <=( A168  and  a30912a );
 a30917a <=( (not A202)  and  (not A201) );
 a30918a <=( A200  and  a30917a );
 a30919a <=( a30918a  and  a30913a );
 a30923a <=( (not A236)  and  (not A235) );
 a30924a <=( (not A234)  and  a30923a );
 a30927a <=( (not A268)  and  (not A267) );
 a30930a <=( A301  and  (not A269) );
 a30931a <=( a30930a  and  a30927a );
 a30932a <=( a30931a  and  a30924a );
 a30936a <=( A199  and  A166 );
 a30937a <=( A168  and  a30936a );
 a30941a <=( (not A202)  and  (not A201) );
 a30942a <=( A200  and  a30941a );
 a30943a <=( a30942a  and  a30937a );
 a30947a <=( (not A236)  and  (not A235) );
 a30948a <=( (not A234)  and  a30947a );
 a30951a <=( (not A266)  and  (not A265) );
 a30954a <=( A301  and  (not A268) );
 a30955a <=( a30954a  and  a30951a );
 a30956a <=( a30955a  and  a30948a );
 a30960a <=( A199  and  A166 );
 a30961a <=( A168  and  a30960a );
 a30965a <=( (not A202)  and  (not A201) );
 a30966a <=( A200  and  a30965a );
 a30967a <=( a30966a  and  a30961a );
 a30971a <=( A236  and  A233 );
 a30972a <=( (not A232)  and  a30971a );
 a30975a <=( A299  and  A298 );
 a30978a <=( (not A301)  and  (not A300) );
 a30979a <=( a30978a  and  a30975a );
 a30980a <=( a30979a  and  a30972a );
 a30984a <=( A199  and  A166 );
 a30985a <=( A168  and  a30984a );
 a30989a <=( (not A202)  and  (not A201) );
 a30990a <=( A200  and  a30989a );
 a30991a <=( a30990a  and  a30985a );
 a30995a <=( A236  and  (not A233) );
 a30996a <=( A232  and  a30995a );
 a30999a <=( A299  and  A298 );
 a31002a <=( (not A301)  and  (not A300) );
 a31003a <=( a31002a  and  a30999a );
 a31004a <=( a31003a  and  a30996a );
 a31008a <=( A199  and  A166 );
 a31009a <=( A168  and  a31008a );
 a31013a <=( (not A202)  and  (not A201) );
 a31014a <=( A200  and  a31013a );
 a31015a <=( a31014a  and  a31009a );
 a31019a <=( (not A235)  and  (not A233) );
 a31020a <=( (not A232)  and  a31019a );
 a31023a <=( (not A268)  and  (not A267) );
 a31026a <=( A301  and  (not A269) );
 a31027a <=( a31026a  and  a31023a );
 a31028a <=( a31027a  and  a31020a );
 a31032a <=( A199  and  A166 );
 a31033a <=( A168  and  a31032a );
 a31037a <=( (not A202)  and  (not A201) );
 a31038a <=( A200  and  a31037a );
 a31039a <=( a31038a  and  a31033a );
 a31043a <=( (not A235)  and  (not A233) );
 a31044a <=( (not A232)  and  a31043a );
 a31047a <=( (not A266)  and  (not A265) );
 a31050a <=( A301  and  (not A268) );
 a31051a <=( a31050a  and  a31047a );
 a31052a <=( a31051a  and  a31044a );
 a31056a <=( (not A199)  and  A166 );
 a31057a <=( A168  and  a31056a );
 a31061a <=( (not A234)  and  (not A202) );
 a31062a <=( (not A200)  and  a31061a );
 a31063a <=( a31062a  and  a31057a );
 a31067a <=( (not A267)  and  (not A236) );
 a31068a <=( (not A235)  and  a31067a );
 a31071a <=( (not A269)  and  (not A268) );
 a31074a <=( A300  and  A299 );
 a31075a <=( a31074a  and  a31071a );
 a31076a <=( a31075a  and  a31068a );
 a31080a <=( (not A199)  and  A166 );
 a31081a <=( A168  and  a31080a );
 a31085a <=( (not A234)  and  (not A202) );
 a31086a <=( (not A200)  and  a31085a );
 a31087a <=( a31086a  and  a31081a );
 a31091a <=( (not A267)  and  (not A236) );
 a31092a <=( (not A235)  and  a31091a );
 a31095a <=( (not A269)  and  (not A268) );
 a31098a <=( A300  and  A298 );
 a31099a <=( a31098a  and  a31095a );
 a31100a <=( a31099a  and  a31092a );
 a31104a <=( (not A199)  and  A166 );
 a31105a <=( A168  and  a31104a );
 a31109a <=( (not A234)  and  (not A202) );
 a31110a <=( (not A200)  and  a31109a );
 a31111a <=( a31110a  and  a31105a );
 a31115a <=( A265  and  (not A236) );
 a31116a <=( (not A235)  and  a31115a );
 a31119a <=( (not A267)  and  A266 );
 a31122a <=( A301  and  (not A268) );
 a31123a <=( a31122a  and  a31119a );
 a31124a <=( a31123a  and  a31116a );
 a31128a <=( (not A199)  and  A166 );
 a31129a <=( A168  and  a31128a );
 a31133a <=( (not A234)  and  (not A202) );
 a31134a <=( (not A200)  and  a31133a );
 a31135a <=( a31134a  and  a31129a );
 a31139a <=( (not A265)  and  (not A236) );
 a31140a <=( (not A235)  and  a31139a );
 a31143a <=( (not A268)  and  (not A266) );
 a31146a <=( A300  and  A299 );
 a31147a <=( a31146a  and  a31143a );
 a31148a <=( a31147a  and  a31140a );
 a31152a <=( (not A199)  and  A166 );
 a31153a <=( A168  and  a31152a );
 a31157a <=( (not A234)  and  (not A202) );
 a31158a <=( (not A200)  and  a31157a );
 a31159a <=( a31158a  and  a31153a );
 a31163a <=( (not A265)  and  (not A236) );
 a31164a <=( (not A235)  and  a31163a );
 a31167a <=( (not A268)  and  (not A266) );
 a31170a <=( A300  and  A298 );
 a31171a <=( a31170a  and  a31167a );
 a31172a <=( a31171a  and  a31164a );
 a31176a <=( (not A199)  and  A166 );
 a31177a <=( A168  and  a31176a );
 a31181a <=( A232  and  (not A202) );
 a31182a <=( (not A200)  and  a31181a );
 a31183a <=( a31182a  and  a31177a );
 a31187a <=( (not A235)  and  (not A234) );
 a31188a <=( A233  and  a31187a );
 a31191a <=( (not A268)  and  (not A267) );
 a31194a <=( A301  and  (not A269) );
 a31195a <=( a31194a  and  a31191a );
 a31196a <=( a31195a  and  a31188a );
 a31200a <=( (not A199)  and  A166 );
 a31201a <=( A168  and  a31200a );
 a31205a <=( A232  and  (not A202) );
 a31206a <=( (not A200)  and  a31205a );
 a31207a <=( a31206a  and  a31201a );
 a31211a <=( (not A235)  and  (not A234) );
 a31212a <=( A233  and  a31211a );
 a31215a <=( (not A266)  and  (not A265) );
 a31218a <=( A301  and  (not A268) );
 a31219a <=( a31218a  and  a31215a );
 a31220a <=( a31219a  and  a31212a );
 a31224a <=( (not A199)  and  A166 );
 a31225a <=( A168  and  a31224a );
 a31229a <=( (not A232)  and  (not A202) );
 a31230a <=( (not A200)  and  a31229a );
 a31231a <=( a31230a  and  a31225a );
 a31235a <=( (not A267)  and  (not A235) );
 a31236a <=( (not A233)  and  a31235a );
 a31239a <=( (not A269)  and  (not A268) );
 a31242a <=( A300  and  A299 );
 a31243a <=( a31242a  and  a31239a );
 a31244a <=( a31243a  and  a31236a );
 a31248a <=( (not A199)  and  A166 );
 a31249a <=( A168  and  a31248a );
 a31253a <=( (not A232)  and  (not A202) );
 a31254a <=( (not A200)  and  a31253a );
 a31255a <=( a31254a  and  a31249a );
 a31259a <=( (not A267)  and  (not A235) );
 a31260a <=( (not A233)  and  a31259a );
 a31263a <=( (not A269)  and  (not A268) );
 a31266a <=( A300  and  A298 );
 a31267a <=( a31266a  and  a31263a );
 a31268a <=( a31267a  and  a31260a );
 a31272a <=( (not A199)  and  A166 );
 a31273a <=( A168  and  a31272a );
 a31277a <=( (not A232)  and  (not A202) );
 a31278a <=( (not A200)  and  a31277a );
 a31279a <=( a31278a  and  a31273a );
 a31283a <=( A265  and  (not A235) );
 a31284a <=( (not A233)  and  a31283a );
 a31287a <=( (not A267)  and  A266 );
 a31290a <=( A301  and  (not A268) );
 a31291a <=( a31290a  and  a31287a );
 a31292a <=( a31291a  and  a31284a );
 a31296a <=( (not A199)  and  A166 );
 a31297a <=( A168  and  a31296a );
 a31301a <=( (not A232)  and  (not A202) );
 a31302a <=( (not A200)  and  a31301a );
 a31303a <=( a31302a  and  a31297a );
 a31307a <=( (not A265)  and  (not A235) );
 a31308a <=( (not A233)  and  a31307a );
 a31311a <=( (not A268)  and  (not A266) );
 a31314a <=( A300  and  A299 );
 a31315a <=( a31314a  and  a31311a );
 a31316a <=( a31315a  and  a31308a );
 a31320a <=( (not A199)  and  A166 );
 a31321a <=( A168  and  a31320a );
 a31325a <=( (not A232)  and  (not A202) );
 a31326a <=( (not A200)  and  a31325a );
 a31327a <=( a31326a  and  a31321a );
 a31331a <=( (not A265)  and  (not A235) );
 a31332a <=( (not A233)  and  a31331a );
 a31335a <=( (not A268)  and  (not A266) );
 a31338a <=( A300  and  A298 );
 a31339a <=( a31338a  and  a31335a );
 a31340a <=( a31339a  and  a31332a );
 a31344a <=( (not A201)  and  A167 );
 a31345a <=( A168  and  a31344a );
 a31349a <=( (not A234)  and  (not A203) );
 a31350a <=( (not A202)  and  a31349a );
 a31351a <=( a31350a  and  a31345a );
 a31355a <=( (not A267)  and  (not A236) );
 a31356a <=( (not A235)  and  a31355a );
 a31359a <=( (not A269)  and  (not A268) );
 a31362a <=( A300  and  A299 );
 a31363a <=( a31362a  and  a31359a );
 a31364a <=( a31363a  and  a31356a );
 a31368a <=( (not A201)  and  A167 );
 a31369a <=( A168  and  a31368a );
 a31373a <=( (not A234)  and  (not A203) );
 a31374a <=( (not A202)  and  a31373a );
 a31375a <=( a31374a  and  a31369a );
 a31379a <=( (not A267)  and  (not A236) );
 a31380a <=( (not A235)  and  a31379a );
 a31383a <=( (not A269)  and  (not A268) );
 a31386a <=( A300  and  A298 );
 a31387a <=( a31386a  and  a31383a );
 a31388a <=( a31387a  and  a31380a );
 a31392a <=( (not A201)  and  A167 );
 a31393a <=( A168  and  a31392a );
 a31397a <=( (not A234)  and  (not A203) );
 a31398a <=( (not A202)  and  a31397a );
 a31399a <=( a31398a  and  a31393a );
 a31403a <=( A265  and  (not A236) );
 a31404a <=( (not A235)  and  a31403a );
 a31407a <=( (not A267)  and  A266 );
 a31410a <=( A301  and  (not A268) );
 a31411a <=( a31410a  and  a31407a );
 a31412a <=( a31411a  and  a31404a );
 a31416a <=( (not A201)  and  A167 );
 a31417a <=( A168  and  a31416a );
 a31421a <=( (not A234)  and  (not A203) );
 a31422a <=( (not A202)  and  a31421a );
 a31423a <=( a31422a  and  a31417a );
 a31427a <=( (not A265)  and  (not A236) );
 a31428a <=( (not A235)  and  a31427a );
 a31431a <=( (not A268)  and  (not A266) );
 a31434a <=( A300  and  A299 );
 a31435a <=( a31434a  and  a31431a );
 a31436a <=( a31435a  and  a31428a );
 a31440a <=( (not A201)  and  A167 );
 a31441a <=( A168  and  a31440a );
 a31445a <=( (not A234)  and  (not A203) );
 a31446a <=( (not A202)  and  a31445a );
 a31447a <=( a31446a  and  a31441a );
 a31451a <=( (not A265)  and  (not A236) );
 a31452a <=( (not A235)  and  a31451a );
 a31455a <=( (not A268)  and  (not A266) );
 a31458a <=( A300  and  A298 );
 a31459a <=( a31458a  and  a31455a );
 a31460a <=( a31459a  and  a31452a );
 a31464a <=( (not A201)  and  A167 );
 a31465a <=( A168  and  a31464a );
 a31469a <=( A232  and  (not A203) );
 a31470a <=( (not A202)  and  a31469a );
 a31471a <=( a31470a  and  a31465a );
 a31475a <=( (not A235)  and  (not A234) );
 a31476a <=( A233  and  a31475a );
 a31479a <=( (not A268)  and  (not A267) );
 a31482a <=( A301  and  (not A269) );
 a31483a <=( a31482a  and  a31479a );
 a31484a <=( a31483a  and  a31476a );
 a31488a <=( (not A201)  and  A167 );
 a31489a <=( A168  and  a31488a );
 a31493a <=( A232  and  (not A203) );
 a31494a <=( (not A202)  and  a31493a );
 a31495a <=( a31494a  and  a31489a );
 a31499a <=( (not A235)  and  (not A234) );
 a31500a <=( A233  and  a31499a );
 a31503a <=( (not A266)  and  (not A265) );
 a31506a <=( A301  and  (not A268) );
 a31507a <=( a31506a  and  a31503a );
 a31508a <=( a31507a  and  a31500a );
 a31512a <=( (not A201)  and  A167 );
 a31513a <=( A168  and  a31512a );
 a31517a <=( (not A232)  and  (not A203) );
 a31518a <=( (not A202)  and  a31517a );
 a31519a <=( a31518a  and  a31513a );
 a31523a <=( (not A267)  and  (not A235) );
 a31524a <=( (not A233)  and  a31523a );
 a31527a <=( (not A269)  and  (not A268) );
 a31530a <=( A300  and  A299 );
 a31531a <=( a31530a  and  a31527a );
 a31532a <=( a31531a  and  a31524a );
 a31536a <=( (not A201)  and  A167 );
 a31537a <=( A168  and  a31536a );
 a31541a <=( (not A232)  and  (not A203) );
 a31542a <=( (not A202)  and  a31541a );
 a31543a <=( a31542a  and  a31537a );
 a31547a <=( (not A267)  and  (not A235) );
 a31548a <=( (not A233)  and  a31547a );
 a31551a <=( (not A269)  and  (not A268) );
 a31554a <=( A300  and  A298 );
 a31555a <=( a31554a  and  a31551a );
 a31556a <=( a31555a  and  a31548a );
 a31560a <=( (not A201)  and  A167 );
 a31561a <=( A168  and  a31560a );
 a31565a <=( (not A232)  and  (not A203) );
 a31566a <=( (not A202)  and  a31565a );
 a31567a <=( a31566a  and  a31561a );
 a31571a <=( A265  and  (not A235) );
 a31572a <=( (not A233)  and  a31571a );
 a31575a <=( (not A267)  and  A266 );
 a31578a <=( A301  and  (not A268) );
 a31579a <=( a31578a  and  a31575a );
 a31580a <=( a31579a  and  a31572a );
 a31584a <=( (not A201)  and  A167 );
 a31585a <=( A168  and  a31584a );
 a31589a <=( (not A232)  and  (not A203) );
 a31590a <=( (not A202)  and  a31589a );
 a31591a <=( a31590a  and  a31585a );
 a31595a <=( (not A265)  and  (not A235) );
 a31596a <=( (not A233)  and  a31595a );
 a31599a <=( (not A268)  and  (not A266) );
 a31602a <=( A300  and  A299 );
 a31603a <=( a31602a  and  a31599a );
 a31604a <=( a31603a  and  a31596a );
 a31608a <=( (not A201)  and  A167 );
 a31609a <=( A168  and  a31608a );
 a31613a <=( (not A232)  and  (not A203) );
 a31614a <=( (not A202)  and  a31613a );
 a31615a <=( a31614a  and  a31609a );
 a31619a <=( (not A265)  and  (not A235) );
 a31620a <=( (not A233)  and  a31619a );
 a31623a <=( (not A268)  and  (not A266) );
 a31626a <=( A300  and  A298 );
 a31627a <=( a31626a  and  a31623a );
 a31628a <=( a31627a  and  a31620a );
 a31632a <=( A199  and  A167 );
 a31633a <=( A168  and  a31632a );
 a31637a <=( (not A202)  and  (not A201) );
 a31638a <=( A200  and  a31637a );
 a31639a <=( a31638a  and  a31633a );
 a31643a <=( (not A236)  and  (not A235) );
 a31644a <=( (not A234)  and  a31643a );
 a31647a <=( (not A268)  and  (not A267) );
 a31650a <=( A301  and  (not A269) );
 a31651a <=( a31650a  and  a31647a );
 a31652a <=( a31651a  and  a31644a );
 a31656a <=( A199  and  A167 );
 a31657a <=( A168  and  a31656a );
 a31661a <=( (not A202)  and  (not A201) );
 a31662a <=( A200  and  a31661a );
 a31663a <=( a31662a  and  a31657a );
 a31667a <=( (not A236)  and  (not A235) );
 a31668a <=( (not A234)  and  a31667a );
 a31671a <=( (not A266)  and  (not A265) );
 a31674a <=( A301  and  (not A268) );
 a31675a <=( a31674a  and  a31671a );
 a31676a <=( a31675a  and  a31668a );
 a31680a <=( A199  and  A167 );
 a31681a <=( A168  and  a31680a );
 a31685a <=( (not A202)  and  (not A201) );
 a31686a <=( A200  and  a31685a );
 a31687a <=( a31686a  and  a31681a );
 a31691a <=( A236  and  A233 );
 a31692a <=( (not A232)  and  a31691a );
 a31695a <=( A299  and  A298 );
 a31698a <=( (not A301)  and  (not A300) );
 a31699a <=( a31698a  and  a31695a );
 a31700a <=( a31699a  and  a31692a );
 a31704a <=( A199  and  A167 );
 a31705a <=( A168  and  a31704a );
 a31709a <=( (not A202)  and  (not A201) );
 a31710a <=( A200  and  a31709a );
 a31711a <=( a31710a  and  a31705a );
 a31715a <=( A236  and  (not A233) );
 a31716a <=( A232  and  a31715a );
 a31719a <=( A299  and  A298 );
 a31722a <=( (not A301)  and  (not A300) );
 a31723a <=( a31722a  and  a31719a );
 a31724a <=( a31723a  and  a31716a );
 a31728a <=( A199  and  A167 );
 a31729a <=( A168  and  a31728a );
 a31733a <=( (not A202)  and  (not A201) );
 a31734a <=( A200  and  a31733a );
 a31735a <=( a31734a  and  a31729a );
 a31739a <=( (not A235)  and  (not A233) );
 a31740a <=( (not A232)  and  a31739a );
 a31743a <=( (not A268)  and  (not A267) );
 a31746a <=( A301  and  (not A269) );
 a31747a <=( a31746a  and  a31743a );
 a31748a <=( a31747a  and  a31740a );
 a31752a <=( A199  and  A167 );
 a31753a <=( A168  and  a31752a );
 a31757a <=( (not A202)  and  (not A201) );
 a31758a <=( A200  and  a31757a );
 a31759a <=( a31758a  and  a31753a );
 a31763a <=( (not A235)  and  (not A233) );
 a31764a <=( (not A232)  and  a31763a );
 a31767a <=( (not A266)  and  (not A265) );
 a31770a <=( A301  and  (not A268) );
 a31771a <=( a31770a  and  a31767a );
 a31772a <=( a31771a  and  a31764a );
 a31776a <=( (not A199)  and  A167 );
 a31777a <=( A168  and  a31776a );
 a31781a <=( (not A234)  and  (not A202) );
 a31782a <=( (not A200)  and  a31781a );
 a31783a <=( a31782a  and  a31777a );
 a31787a <=( (not A267)  and  (not A236) );
 a31788a <=( (not A235)  and  a31787a );
 a31791a <=( (not A269)  and  (not A268) );
 a31794a <=( A300  and  A299 );
 a31795a <=( a31794a  and  a31791a );
 a31796a <=( a31795a  and  a31788a );
 a31800a <=( (not A199)  and  A167 );
 a31801a <=( A168  and  a31800a );
 a31805a <=( (not A234)  and  (not A202) );
 a31806a <=( (not A200)  and  a31805a );
 a31807a <=( a31806a  and  a31801a );
 a31811a <=( (not A267)  and  (not A236) );
 a31812a <=( (not A235)  and  a31811a );
 a31815a <=( (not A269)  and  (not A268) );
 a31818a <=( A300  and  A298 );
 a31819a <=( a31818a  and  a31815a );
 a31820a <=( a31819a  and  a31812a );
 a31824a <=( (not A199)  and  A167 );
 a31825a <=( A168  and  a31824a );
 a31829a <=( (not A234)  and  (not A202) );
 a31830a <=( (not A200)  and  a31829a );
 a31831a <=( a31830a  and  a31825a );
 a31835a <=( A265  and  (not A236) );
 a31836a <=( (not A235)  and  a31835a );
 a31839a <=( (not A267)  and  A266 );
 a31842a <=( A301  and  (not A268) );
 a31843a <=( a31842a  and  a31839a );
 a31844a <=( a31843a  and  a31836a );
 a31848a <=( (not A199)  and  A167 );
 a31849a <=( A168  and  a31848a );
 a31853a <=( (not A234)  and  (not A202) );
 a31854a <=( (not A200)  and  a31853a );
 a31855a <=( a31854a  and  a31849a );
 a31859a <=( (not A265)  and  (not A236) );
 a31860a <=( (not A235)  and  a31859a );
 a31863a <=( (not A268)  and  (not A266) );
 a31866a <=( A300  and  A299 );
 a31867a <=( a31866a  and  a31863a );
 a31868a <=( a31867a  and  a31860a );
 a31872a <=( (not A199)  and  A167 );
 a31873a <=( A168  and  a31872a );
 a31877a <=( (not A234)  and  (not A202) );
 a31878a <=( (not A200)  and  a31877a );
 a31879a <=( a31878a  and  a31873a );
 a31883a <=( (not A265)  and  (not A236) );
 a31884a <=( (not A235)  and  a31883a );
 a31887a <=( (not A268)  and  (not A266) );
 a31890a <=( A300  and  A298 );
 a31891a <=( a31890a  and  a31887a );
 a31892a <=( a31891a  and  a31884a );
 a31896a <=( (not A199)  and  A167 );
 a31897a <=( A168  and  a31896a );
 a31901a <=( A232  and  (not A202) );
 a31902a <=( (not A200)  and  a31901a );
 a31903a <=( a31902a  and  a31897a );
 a31907a <=( (not A235)  and  (not A234) );
 a31908a <=( A233  and  a31907a );
 a31911a <=( (not A268)  and  (not A267) );
 a31914a <=( A301  and  (not A269) );
 a31915a <=( a31914a  and  a31911a );
 a31916a <=( a31915a  and  a31908a );
 a31920a <=( (not A199)  and  A167 );
 a31921a <=( A168  and  a31920a );
 a31925a <=( A232  and  (not A202) );
 a31926a <=( (not A200)  and  a31925a );
 a31927a <=( a31926a  and  a31921a );
 a31931a <=( (not A235)  and  (not A234) );
 a31932a <=( A233  and  a31931a );
 a31935a <=( (not A266)  and  (not A265) );
 a31938a <=( A301  and  (not A268) );
 a31939a <=( a31938a  and  a31935a );
 a31940a <=( a31939a  and  a31932a );
 a31944a <=( (not A199)  and  A167 );
 a31945a <=( A168  and  a31944a );
 a31949a <=( (not A232)  and  (not A202) );
 a31950a <=( (not A200)  and  a31949a );
 a31951a <=( a31950a  and  a31945a );
 a31955a <=( (not A267)  and  (not A235) );
 a31956a <=( (not A233)  and  a31955a );
 a31959a <=( (not A269)  and  (not A268) );
 a31962a <=( A300  and  A299 );
 a31963a <=( a31962a  and  a31959a );
 a31964a <=( a31963a  and  a31956a );
 a31968a <=( (not A199)  and  A167 );
 a31969a <=( A168  and  a31968a );
 a31973a <=( (not A232)  and  (not A202) );
 a31974a <=( (not A200)  and  a31973a );
 a31975a <=( a31974a  and  a31969a );
 a31979a <=( (not A267)  and  (not A235) );
 a31980a <=( (not A233)  and  a31979a );
 a31983a <=( (not A269)  and  (not A268) );
 a31986a <=( A300  and  A298 );
 a31987a <=( a31986a  and  a31983a );
 a31988a <=( a31987a  and  a31980a );
 a31992a <=( (not A199)  and  A167 );
 a31993a <=( A168  and  a31992a );
 a31997a <=( (not A232)  and  (not A202) );
 a31998a <=( (not A200)  and  a31997a );
 a31999a <=( a31998a  and  a31993a );
 a32003a <=( A265  and  (not A235) );
 a32004a <=( (not A233)  and  a32003a );
 a32007a <=( (not A267)  and  A266 );
 a32010a <=( A301  and  (not A268) );
 a32011a <=( a32010a  and  a32007a );
 a32012a <=( a32011a  and  a32004a );
 a32016a <=( (not A199)  and  A167 );
 a32017a <=( A168  and  a32016a );
 a32021a <=( (not A232)  and  (not A202) );
 a32022a <=( (not A200)  and  a32021a );
 a32023a <=( a32022a  and  a32017a );
 a32027a <=( (not A265)  and  (not A235) );
 a32028a <=( (not A233)  and  a32027a );
 a32031a <=( (not A268)  and  (not A266) );
 a32034a <=( A300  and  A299 );
 a32035a <=( a32034a  and  a32031a );
 a32036a <=( a32035a  and  a32028a );
 a32040a <=( (not A199)  and  A167 );
 a32041a <=( A168  and  a32040a );
 a32045a <=( (not A232)  and  (not A202) );
 a32046a <=( (not A200)  and  a32045a );
 a32047a <=( a32046a  and  a32041a );
 a32051a <=( (not A265)  and  (not A235) );
 a32052a <=( (not A233)  and  a32051a );
 a32055a <=( (not A268)  and  (not A266) );
 a32058a <=( A300  and  A298 );
 a32059a <=( a32058a  and  a32055a );
 a32060a <=( a32059a  and  a32052a );
 a32064a <=( (not A166)  and  A167 );
 a32065a <=( A170  and  a32064a );
 a32069a <=( (not A203)  and  (not A202) );
 a32070a <=( (not A201)  and  a32069a );
 a32071a <=( a32070a  and  a32065a );
 a32075a <=( (not A236)  and  (not A235) );
 a32076a <=( (not A234)  and  a32075a );
 a32079a <=( (not A268)  and  (not A267) );
 a32082a <=( A301  and  (not A269) );
 a32083a <=( a32082a  and  a32079a );
 a32084a <=( a32083a  and  a32076a );
 a32088a <=( (not A166)  and  A167 );
 a32089a <=( A170  and  a32088a );
 a32093a <=( (not A203)  and  (not A202) );
 a32094a <=( (not A201)  and  a32093a );
 a32095a <=( a32094a  and  a32089a );
 a32099a <=( (not A236)  and  (not A235) );
 a32100a <=( (not A234)  and  a32099a );
 a32103a <=( (not A266)  and  (not A265) );
 a32106a <=( A301  and  (not A268) );
 a32107a <=( a32106a  and  a32103a );
 a32108a <=( a32107a  and  a32100a );
 a32112a <=( (not A166)  and  A167 );
 a32113a <=( A170  and  a32112a );
 a32117a <=( (not A203)  and  (not A202) );
 a32118a <=( (not A201)  and  a32117a );
 a32119a <=( a32118a  and  a32113a );
 a32123a <=( A236  and  A233 );
 a32124a <=( (not A232)  and  a32123a );
 a32127a <=( A299  and  A298 );
 a32130a <=( (not A301)  and  (not A300) );
 a32131a <=( a32130a  and  a32127a );
 a32132a <=( a32131a  and  a32124a );
 a32136a <=( (not A166)  and  A167 );
 a32137a <=( A170  and  a32136a );
 a32141a <=( (not A203)  and  (not A202) );
 a32142a <=( (not A201)  and  a32141a );
 a32143a <=( a32142a  and  a32137a );
 a32147a <=( A236  and  (not A233) );
 a32148a <=( A232  and  a32147a );
 a32151a <=( A299  and  A298 );
 a32154a <=( (not A301)  and  (not A300) );
 a32155a <=( a32154a  and  a32151a );
 a32156a <=( a32155a  and  a32148a );
 a32160a <=( (not A166)  and  A167 );
 a32161a <=( A170  and  a32160a );
 a32165a <=( (not A203)  and  (not A202) );
 a32166a <=( (not A201)  and  a32165a );
 a32167a <=( a32166a  and  a32161a );
 a32171a <=( (not A235)  and  (not A233) );
 a32172a <=( (not A232)  and  a32171a );
 a32175a <=( (not A268)  and  (not A267) );
 a32178a <=( A301  and  (not A269) );
 a32179a <=( a32178a  and  a32175a );
 a32180a <=( a32179a  and  a32172a );
 a32184a <=( (not A166)  and  A167 );
 a32185a <=( A170  and  a32184a );
 a32189a <=( (not A203)  and  (not A202) );
 a32190a <=( (not A201)  and  a32189a );
 a32191a <=( a32190a  and  a32185a );
 a32195a <=( (not A235)  and  (not A233) );
 a32196a <=( (not A232)  and  a32195a );
 a32199a <=( (not A266)  and  (not A265) );
 a32202a <=( A301  and  (not A268) );
 a32203a <=( a32202a  and  a32199a );
 a32204a <=( a32203a  and  a32196a );
 a32208a <=( (not A166)  and  A167 );
 a32209a <=( A170  and  a32208a );
 a32213a <=( (not A201)  and  A200 );
 a32214a <=( A199  and  a32213a );
 a32215a <=( a32214a  and  a32209a );
 a32219a <=( A234  and  A232 );
 a32220a <=( (not A202)  and  a32219a );
 a32223a <=( A299  and  A298 );
 a32226a <=( (not A301)  and  (not A300) );
 a32227a <=( a32226a  and  a32223a );
 a32228a <=( a32227a  and  a32220a );
 a32232a <=( (not A166)  and  A167 );
 a32233a <=( A170  and  a32232a );
 a32237a <=( (not A201)  and  A200 );
 a32238a <=( A199  and  a32237a );
 a32239a <=( a32238a  and  a32233a );
 a32243a <=( A234  and  A233 );
 a32244a <=( (not A202)  and  a32243a );
 a32247a <=( A299  and  A298 );
 a32250a <=( (not A301)  and  (not A300) );
 a32251a <=( a32250a  and  a32247a );
 a32252a <=( a32251a  and  a32244a );
 a32256a <=( (not A166)  and  A167 );
 a32257a <=( A170  and  a32256a );
 a32261a <=( (not A201)  and  A200 );
 a32262a <=( A199  and  a32261a );
 a32263a <=( a32262a  and  a32257a );
 a32267a <=( A233  and  (not A232) );
 a32268a <=( (not A202)  and  a32267a );
 a32271a <=( (not A300)  and  A236 );
 a32274a <=( (not A302)  and  (not A301) );
 a32275a <=( a32274a  and  a32271a );
 a32276a <=( a32275a  and  a32268a );
 a32280a <=( (not A166)  and  A167 );
 a32281a <=( A170  and  a32280a );
 a32285a <=( (not A201)  and  A200 );
 a32286a <=( A199  and  a32285a );
 a32287a <=( a32286a  and  a32281a );
 a32291a <=( A233  and  (not A232) );
 a32292a <=( (not A202)  and  a32291a );
 a32295a <=( (not A298)  and  A236 );
 a32298a <=( (not A301)  and  (not A299) );
 a32299a <=( a32298a  and  a32295a );
 a32300a <=( a32299a  and  a32292a );
 a32304a <=( (not A166)  and  A167 );
 a32305a <=( A170  and  a32304a );
 a32309a <=( (not A201)  and  A200 );
 a32310a <=( A199  and  a32309a );
 a32311a <=( a32310a  and  a32305a );
 a32315a <=( A233  and  (not A232) );
 a32316a <=( (not A202)  and  a32315a );
 a32319a <=( (not A265)  and  A236 );
 a32322a <=( A269  and  A266 );
 a32323a <=( a32322a  and  a32319a );
 a32324a <=( a32323a  and  a32316a );
 a32328a <=( (not A166)  and  A167 );
 a32329a <=( A170  and  a32328a );
 a32333a <=( (not A201)  and  A200 );
 a32334a <=( A199  and  a32333a );
 a32335a <=( a32334a  and  a32329a );
 a32339a <=( A233  and  (not A232) );
 a32340a <=( (not A202)  and  a32339a );
 a32343a <=( A265  and  A236 );
 a32346a <=( A269  and  (not A266) );
 a32347a <=( a32346a  and  a32343a );
 a32348a <=( a32347a  and  a32340a );
 a32352a <=( (not A166)  and  A167 );
 a32353a <=( A170  and  a32352a );
 a32357a <=( (not A201)  and  A200 );
 a32358a <=( A199  and  a32357a );
 a32359a <=( a32358a  and  a32353a );
 a32363a <=( (not A233)  and  A232 );
 a32364a <=( (not A202)  and  a32363a );
 a32367a <=( (not A300)  and  A236 );
 a32370a <=( (not A302)  and  (not A301) );
 a32371a <=( a32370a  and  a32367a );
 a32372a <=( a32371a  and  a32364a );
 a32376a <=( (not A166)  and  A167 );
 a32377a <=( A170  and  a32376a );
 a32381a <=( (not A201)  and  A200 );
 a32382a <=( A199  and  a32381a );
 a32383a <=( a32382a  and  a32377a );
 a32387a <=( (not A233)  and  A232 );
 a32388a <=( (not A202)  and  a32387a );
 a32391a <=( (not A298)  and  A236 );
 a32394a <=( (not A301)  and  (not A299) );
 a32395a <=( a32394a  and  a32391a );
 a32396a <=( a32395a  and  a32388a );
 a32400a <=( (not A166)  and  A167 );
 a32401a <=( A170  and  a32400a );
 a32405a <=( (not A201)  and  A200 );
 a32406a <=( A199  and  a32405a );
 a32407a <=( a32406a  and  a32401a );
 a32411a <=( (not A233)  and  A232 );
 a32412a <=( (not A202)  and  a32411a );
 a32415a <=( (not A265)  and  A236 );
 a32418a <=( A269  and  A266 );
 a32419a <=( a32418a  and  a32415a );
 a32420a <=( a32419a  and  a32412a );
 a32424a <=( (not A166)  and  A167 );
 a32425a <=( A170  and  a32424a );
 a32429a <=( (not A201)  and  A200 );
 a32430a <=( A199  and  a32429a );
 a32431a <=( a32430a  and  a32425a );
 a32435a <=( (not A233)  and  A232 );
 a32436a <=( (not A202)  and  a32435a );
 a32439a <=( A265  and  A236 );
 a32442a <=( A269  and  (not A266) );
 a32443a <=( a32442a  and  a32439a );
 a32444a <=( a32443a  and  a32436a );
 a32448a <=( (not A166)  and  A167 );
 a32449a <=( A170  and  a32448a );
 a32453a <=( (not A202)  and  (not A200) );
 a32454a <=( (not A199)  and  a32453a );
 a32455a <=( a32454a  and  a32449a );
 a32459a <=( (not A236)  and  (not A235) );
 a32460a <=( (not A234)  and  a32459a );
 a32463a <=( (not A268)  and  (not A267) );
 a32466a <=( A301  and  (not A269) );
 a32467a <=( a32466a  and  a32463a );
 a32468a <=( a32467a  and  a32460a );
 a32472a <=( (not A166)  and  A167 );
 a32473a <=( A170  and  a32472a );
 a32477a <=( (not A202)  and  (not A200) );
 a32478a <=( (not A199)  and  a32477a );
 a32479a <=( a32478a  and  a32473a );
 a32483a <=( (not A236)  and  (not A235) );
 a32484a <=( (not A234)  and  a32483a );
 a32487a <=( (not A266)  and  (not A265) );
 a32490a <=( A301  and  (not A268) );
 a32491a <=( a32490a  and  a32487a );
 a32492a <=( a32491a  and  a32484a );
 a32496a <=( (not A166)  and  A167 );
 a32497a <=( A170  and  a32496a );
 a32501a <=( (not A202)  and  (not A200) );
 a32502a <=( (not A199)  and  a32501a );
 a32503a <=( a32502a  and  a32497a );
 a32507a <=( A236  and  A233 );
 a32508a <=( (not A232)  and  a32507a );
 a32511a <=( A299  and  A298 );
 a32514a <=( (not A301)  and  (not A300) );
 a32515a <=( a32514a  and  a32511a );
 a32516a <=( a32515a  and  a32508a );
 a32520a <=( (not A166)  and  A167 );
 a32521a <=( A170  and  a32520a );
 a32525a <=( (not A202)  and  (not A200) );
 a32526a <=( (not A199)  and  a32525a );
 a32527a <=( a32526a  and  a32521a );
 a32531a <=( A236  and  (not A233) );
 a32532a <=( A232  and  a32531a );
 a32535a <=( A299  and  A298 );
 a32538a <=( (not A301)  and  (not A300) );
 a32539a <=( a32538a  and  a32535a );
 a32540a <=( a32539a  and  a32532a );
 a32544a <=( (not A166)  and  A167 );
 a32545a <=( A170  and  a32544a );
 a32549a <=( (not A202)  and  (not A200) );
 a32550a <=( (not A199)  and  a32549a );
 a32551a <=( a32550a  and  a32545a );
 a32555a <=( (not A235)  and  (not A233) );
 a32556a <=( (not A232)  and  a32555a );
 a32559a <=( (not A268)  and  (not A267) );
 a32562a <=( A301  and  (not A269) );
 a32563a <=( a32562a  and  a32559a );
 a32564a <=( a32563a  and  a32556a );
 a32568a <=( (not A166)  and  A167 );
 a32569a <=( A170  and  a32568a );
 a32573a <=( (not A202)  and  (not A200) );
 a32574a <=( (not A199)  and  a32573a );
 a32575a <=( a32574a  and  a32569a );
 a32579a <=( (not A235)  and  (not A233) );
 a32580a <=( (not A232)  and  a32579a );
 a32583a <=( (not A266)  and  (not A265) );
 a32586a <=( A301  and  (not A268) );
 a32587a <=( a32586a  and  a32583a );
 a32588a <=( a32587a  and  a32580a );
 a32592a <=( A166  and  (not A167) );
 a32593a <=( A170  and  a32592a );
 a32597a <=( (not A203)  and  (not A202) );
 a32598a <=( (not A201)  and  a32597a );
 a32599a <=( a32598a  and  a32593a );
 a32603a <=( (not A236)  and  (not A235) );
 a32604a <=( (not A234)  and  a32603a );
 a32607a <=( (not A268)  and  (not A267) );
 a32610a <=( A301  and  (not A269) );
 a32611a <=( a32610a  and  a32607a );
 a32612a <=( a32611a  and  a32604a );
 a32616a <=( A166  and  (not A167) );
 a32617a <=( A170  and  a32616a );
 a32621a <=( (not A203)  and  (not A202) );
 a32622a <=( (not A201)  and  a32621a );
 a32623a <=( a32622a  and  a32617a );
 a32627a <=( (not A236)  and  (not A235) );
 a32628a <=( (not A234)  and  a32627a );
 a32631a <=( (not A266)  and  (not A265) );
 a32634a <=( A301  and  (not A268) );
 a32635a <=( a32634a  and  a32631a );
 a32636a <=( a32635a  and  a32628a );
 a32640a <=( A166  and  (not A167) );
 a32641a <=( A170  and  a32640a );
 a32645a <=( (not A203)  and  (not A202) );
 a32646a <=( (not A201)  and  a32645a );
 a32647a <=( a32646a  and  a32641a );
 a32651a <=( A236  and  A233 );
 a32652a <=( (not A232)  and  a32651a );
 a32655a <=( A299  and  A298 );
 a32658a <=( (not A301)  and  (not A300) );
 a32659a <=( a32658a  and  a32655a );
 a32660a <=( a32659a  and  a32652a );
 a32664a <=( A166  and  (not A167) );
 a32665a <=( A170  and  a32664a );
 a32669a <=( (not A203)  and  (not A202) );
 a32670a <=( (not A201)  and  a32669a );
 a32671a <=( a32670a  and  a32665a );
 a32675a <=( A236  and  (not A233) );
 a32676a <=( A232  and  a32675a );
 a32679a <=( A299  and  A298 );
 a32682a <=( (not A301)  and  (not A300) );
 a32683a <=( a32682a  and  a32679a );
 a32684a <=( a32683a  and  a32676a );
 a32688a <=( A166  and  (not A167) );
 a32689a <=( A170  and  a32688a );
 a32693a <=( (not A203)  and  (not A202) );
 a32694a <=( (not A201)  and  a32693a );
 a32695a <=( a32694a  and  a32689a );
 a32699a <=( (not A235)  and  (not A233) );
 a32700a <=( (not A232)  and  a32699a );
 a32703a <=( (not A268)  and  (not A267) );
 a32706a <=( A301  and  (not A269) );
 a32707a <=( a32706a  and  a32703a );
 a32708a <=( a32707a  and  a32700a );
 a32712a <=( A166  and  (not A167) );
 a32713a <=( A170  and  a32712a );
 a32717a <=( (not A203)  and  (not A202) );
 a32718a <=( (not A201)  and  a32717a );
 a32719a <=( a32718a  and  a32713a );
 a32723a <=( (not A235)  and  (not A233) );
 a32724a <=( (not A232)  and  a32723a );
 a32727a <=( (not A266)  and  (not A265) );
 a32730a <=( A301  and  (not A268) );
 a32731a <=( a32730a  and  a32727a );
 a32732a <=( a32731a  and  a32724a );
 a32736a <=( A166  and  (not A167) );
 a32737a <=( A170  and  a32736a );
 a32741a <=( (not A201)  and  A200 );
 a32742a <=( A199  and  a32741a );
 a32743a <=( a32742a  and  a32737a );
 a32747a <=( A234  and  A232 );
 a32748a <=( (not A202)  and  a32747a );
 a32751a <=( A299  and  A298 );
 a32754a <=( (not A301)  and  (not A300) );
 a32755a <=( a32754a  and  a32751a );
 a32756a <=( a32755a  and  a32748a );
 a32760a <=( A166  and  (not A167) );
 a32761a <=( A170  and  a32760a );
 a32765a <=( (not A201)  and  A200 );
 a32766a <=( A199  and  a32765a );
 a32767a <=( a32766a  and  a32761a );
 a32771a <=( A234  and  A233 );
 a32772a <=( (not A202)  and  a32771a );
 a32775a <=( A299  and  A298 );
 a32778a <=( (not A301)  and  (not A300) );
 a32779a <=( a32778a  and  a32775a );
 a32780a <=( a32779a  and  a32772a );
 a32784a <=( A166  and  (not A167) );
 a32785a <=( A170  and  a32784a );
 a32789a <=( (not A201)  and  A200 );
 a32790a <=( A199  and  a32789a );
 a32791a <=( a32790a  and  a32785a );
 a32795a <=( A233  and  (not A232) );
 a32796a <=( (not A202)  and  a32795a );
 a32799a <=( (not A300)  and  A236 );
 a32802a <=( (not A302)  and  (not A301) );
 a32803a <=( a32802a  and  a32799a );
 a32804a <=( a32803a  and  a32796a );
 a32808a <=( A166  and  (not A167) );
 a32809a <=( A170  and  a32808a );
 a32813a <=( (not A201)  and  A200 );
 a32814a <=( A199  and  a32813a );
 a32815a <=( a32814a  and  a32809a );
 a32819a <=( A233  and  (not A232) );
 a32820a <=( (not A202)  and  a32819a );
 a32823a <=( (not A298)  and  A236 );
 a32826a <=( (not A301)  and  (not A299) );
 a32827a <=( a32826a  and  a32823a );
 a32828a <=( a32827a  and  a32820a );
 a32832a <=( A166  and  (not A167) );
 a32833a <=( A170  and  a32832a );
 a32837a <=( (not A201)  and  A200 );
 a32838a <=( A199  and  a32837a );
 a32839a <=( a32838a  and  a32833a );
 a32843a <=( A233  and  (not A232) );
 a32844a <=( (not A202)  and  a32843a );
 a32847a <=( (not A265)  and  A236 );
 a32850a <=( A269  and  A266 );
 a32851a <=( a32850a  and  a32847a );
 a32852a <=( a32851a  and  a32844a );
 a32856a <=( A166  and  (not A167) );
 a32857a <=( A170  and  a32856a );
 a32861a <=( (not A201)  and  A200 );
 a32862a <=( A199  and  a32861a );
 a32863a <=( a32862a  and  a32857a );
 a32867a <=( A233  and  (not A232) );
 a32868a <=( (not A202)  and  a32867a );
 a32871a <=( A265  and  A236 );
 a32874a <=( A269  and  (not A266) );
 a32875a <=( a32874a  and  a32871a );
 a32876a <=( a32875a  and  a32868a );
 a32880a <=( A166  and  (not A167) );
 a32881a <=( A170  and  a32880a );
 a32885a <=( (not A201)  and  A200 );
 a32886a <=( A199  and  a32885a );
 a32887a <=( a32886a  and  a32881a );
 a32891a <=( (not A233)  and  A232 );
 a32892a <=( (not A202)  and  a32891a );
 a32895a <=( (not A300)  and  A236 );
 a32898a <=( (not A302)  and  (not A301) );
 a32899a <=( a32898a  and  a32895a );
 a32900a <=( a32899a  and  a32892a );
 a32904a <=( A166  and  (not A167) );
 a32905a <=( A170  and  a32904a );
 a32909a <=( (not A201)  and  A200 );
 a32910a <=( A199  and  a32909a );
 a32911a <=( a32910a  and  a32905a );
 a32915a <=( (not A233)  and  A232 );
 a32916a <=( (not A202)  and  a32915a );
 a32919a <=( (not A298)  and  A236 );
 a32922a <=( (not A301)  and  (not A299) );
 a32923a <=( a32922a  and  a32919a );
 a32924a <=( a32923a  and  a32916a );
 a32928a <=( A166  and  (not A167) );
 a32929a <=( A170  and  a32928a );
 a32933a <=( (not A201)  and  A200 );
 a32934a <=( A199  and  a32933a );
 a32935a <=( a32934a  and  a32929a );
 a32939a <=( (not A233)  and  A232 );
 a32940a <=( (not A202)  and  a32939a );
 a32943a <=( (not A265)  and  A236 );
 a32946a <=( A269  and  A266 );
 a32947a <=( a32946a  and  a32943a );
 a32948a <=( a32947a  and  a32940a );
 a32952a <=( A166  and  (not A167) );
 a32953a <=( A170  and  a32952a );
 a32957a <=( (not A201)  and  A200 );
 a32958a <=( A199  and  a32957a );
 a32959a <=( a32958a  and  a32953a );
 a32963a <=( (not A233)  and  A232 );
 a32964a <=( (not A202)  and  a32963a );
 a32967a <=( A265  and  A236 );
 a32970a <=( A269  and  (not A266) );
 a32971a <=( a32970a  and  a32967a );
 a32972a <=( a32971a  and  a32964a );
 a32976a <=( A166  and  (not A167) );
 a32977a <=( A170  and  a32976a );
 a32981a <=( (not A202)  and  (not A200) );
 a32982a <=( (not A199)  and  a32981a );
 a32983a <=( a32982a  and  a32977a );
 a32987a <=( (not A236)  and  (not A235) );
 a32988a <=( (not A234)  and  a32987a );
 a32991a <=( (not A268)  and  (not A267) );
 a32994a <=( A301  and  (not A269) );
 a32995a <=( a32994a  and  a32991a );
 a32996a <=( a32995a  and  a32988a );
 a33000a <=( A166  and  (not A167) );
 a33001a <=( A170  and  a33000a );
 a33005a <=( (not A202)  and  (not A200) );
 a33006a <=( (not A199)  and  a33005a );
 a33007a <=( a33006a  and  a33001a );
 a33011a <=( (not A236)  and  (not A235) );
 a33012a <=( (not A234)  and  a33011a );
 a33015a <=( (not A266)  and  (not A265) );
 a33018a <=( A301  and  (not A268) );
 a33019a <=( a33018a  and  a33015a );
 a33020a <=( a33019a  and  a33012a );
 a33024a <=( A166  and  (not A167) );
 a33025a <=( A170  and  a33024a );
 a33029a <=( (not A202)  and  (not A200) );
 a33030a <=( (not A199)  and  a33029a );
 a33031a <=( a33030a  and  a33025a );
 a33035a <=( A236  and  A233 );
 a33036a <=( (not A232)  and  a33035a );
 a33039a <=( A299  and  A298 );
 a33042a <=( (not A301)  and  (not A300) );
 a33043a <=( a33042a  and  a33039a );
 a33044a <=( a33043a  and  a33036a );
 a33048a <=( A166  and  (not A167) );
 a33049a <=( A170  and  a33048a );
 a33053a <=( (not A202)  and  (not A200) );
 a33054a <=( (not A199)  and  a33053a );
 a33055a <=( a33054a  and  a33049a );
 a33059a <=( A236  and  (not A233) );
 a33060a <=( A232  and  a33059a );
 a33063a <=( A299  and  A298 );
 a33066a <=( (not A301)  and  (not A300) );
 a33067a <=( a33066a  and  a33063a );
 a33068a <=( a33067a  and  a33060a );
 a33072a <=( A166  and  (not A167) );
 a33073a <=( A170  and  a33072a );
 a33077a <=( (not A202)  and  (not A200) );
 a33078a <=( (not A199)  and  a33077a );
 a33079a <=( a33078a  and  a33073a );
 a33083a <=( (not A235)  and  (not A233) );
 a33084a <=( (not A232)  and  a33083a );
 a33087a <=( (not A268)  and  (not A267) );
 a33090a <=( A301  and  (not A269) );
 a33091a <=( a33090a  and  a33087a );
 a33092a <=( a33091a  and  a33084a );
 a33096a <=( A166  and  (not A167) );
 a33097a <=( A170  and  a33096a );
 a33101a <=( (not A202)  and  (not A200) );
 a33102a <=( (not A199)  and  a33101a );
 a33103a <=( a33102a  and  a33097a );
 a33107a <=( (not A235)  and  (not A233) );
 a33108a <=( (not A232)  and  a33107a );
 a33111a <=( (not A266)  and  (not A265) );
 a33114a <=( A301  and  (not A268) );
 a33115a <=( a33114a  and  a33111a );
 a33116a <=( a33115a  and  a33108a );
 a33120a <=( (not A202)  and  (not A201) );
 a33121a <=( A169  and  a33120a );
 a33125a <=( (not A235)  and  (not A234) );
 a33126a <=( (not A203)  and  a33125a );
 a33127a <=( a33126a  and  a33121a );
 a33131a <=( (not A268)  and  (not A267) );
 a33132a <=( (not A236)  and  a33131a );
 a33135a <=( A298  and  (not A269) );
 a33138a <=( A302  and  (not A299) );
 a33139a <=( a33138a  and  a33135a );
 a33140a <=( a33139a  and  a33132a );
 a33144a <=( (not A202)  and  (not A201) );
 a33145a <=( A169  and  a33144a );
 a33149a <=( (not A235)  and  (not A234) );
 a33150a <=( (not A203)  and  a33149a );
 a33151a <=( a33150a  and  a33145a );
 a33155a <=( (not A268)  and  (not A267) );
 a33156a <=( (not A236)  and  a33155a );
 a33159a <=( (not A298)  and  (not A269) );
 a33162a <=( A302  and  A299 );
 a33163a <=( a33162a  and  a33159a );
 a33164a <=( a33163a  and  a33156a );
 a33168a <=( (not A202)  and  (not A201) );
 a33169a <=( A169  and  a33168a );
 a33173a <=( (not A235)  and  (not A234) );
 a33174a <=( (not A203)  and  a33173a );
 a33175a <=( a33174a  and  a33169a );
 a33179a <=( A266  and  A265 );
 a33180a <=( (not A236)  and  a33179a );
 a33183a <=( (not A268)  and  (not A267) );
 a33186a <=( A300  and  A299 );
 a33187a <=( a33186a  and  a33183a );
 a33188a <=( a33187a  and  a33180a );
 a33192a <=( (not A202)  and  (not A201) );
 a33193a <=( A169  and  a33192a );
 a33197a <=( (not A235)  and  (not A234) );
 a33198a <=( (not A203)  and  a33197a );
 a33199a <=( a33198a  and  a33193a );
 a33203a <=( A266  and  A265 );
 a33204a <=( (not A236)  and  a33203a );
 a33207a <=( (not A268)  and  (not A267) );
 a33210a <=( A300  and  A298 );
 a33211a <=( a33210a  and  a33207a );
 a33212a <=( a33211a  and  a33204a );
 a33216a <=( (not A202)  and  (not A201) );
 a33217a <=( A169  and  a33216a );
 a33221a <=( (not A235)  and  (not A234) );
 a33222a <=( (not A203)  and  a33221a );
 a33223a <=( a33222a  and  a33217a );
 a33227a <=( (not A266)  and  (not A265) );
 a33228a <=( (not A236)  and  a33227a );
 a33231a <=( A298  and  (not A268) );
 a33234a <=( A302  and  (not A299) );
 a33235a <=( a33234a  and  a33231a );
 a33236a <=( a33235a  and  a33228a );
 a33240a <=( (not A202)  and  (not A201) );
 a33241a <=( A169  and  a33240a );
 a33245a <=( (not A235)  and  (not A234) );
 a33246a <=( (not A203)  and  a33245a );
 a33247a <=( a33246a  and  a33241a );
 a33251a <=( (not A266)  and  (not A265) );
 a33252a <=( (not A236)  and  a33251a );
 a33255a <=( (not A298)  and  (not A268) );
 a33258a <=( A302  and  A299 );
 a33259a <=( a33258a  and  a33255a );
 a33260a <=( a33259a  and  a33252a );
 a33264a <=( (not A202)  and  (not A201) );
 a33265a <=( A169  and  a33264a );
 a33269a <=( A233  and  A232 );
 a33270a <=( (not A203)  and  a33269a );
 a33271a <=( a33270a  and  a33265a );
 a33275a <=( (not A267)  and  (not A235) );
 a33276a <=( (not A234)  and  a33275a );
 a33279a <=( (not A269)  and  (not A268) );
 a33282a <=( A300  and  A299 );
 a33283a <=( a33282a  and  a33279a );
 a33284a <=( a33283a  and  a33276a );
 a33288a <=( (not A202)  and  (not A201) );
 a33289a <=( A169  and  a33288a );
 a33293a <=( A233  and  A232 );
 a33294a <=( (not A203)  and  a33293a );
 a33295a <=( a33294a  and  a33289a );
 a33299a <=( (not A267)  and  (not A235) );
 a33300a <=( (not A234)  and  a33299a );
 a33303a <=( (not A269)  and  (not A268) );
 a33306a <=( A300  and  A298 );
 a33307a <=( a33306a  and  a33303a );
 a33308a <=( a33307a  and  a33300a );
 a33312a <=( (not A202)  and  (not A201) );
 a33313a <=( A169  and  a33312a );
 a33317a <=( A233  and  A232 );
 a33318a <=( (not A203)  and  a33317a );
 a33319a <=( a33318a  and  a33313a );
 a33323a <=( A265  and  (not A235) );
 a33324a <=( (not A234)  and  a33323a );
 a33327a <=( (not A267)  and  A266 );
 a33330a <=( A301  and  (not A268) );
 a33331a <=( a33330a  and  a33327a );
 a33332a <=( a33331a  and  a33324a );
 a33336a <=( (not A202)  and  (not A201) );
 a33337a <=( A169  and  a33336a );
 a33341a <=( A233  and  A232 );
 a33342a <=( (not A203)  and  a33341a );
 a33343a <=( a33342a  and  a33337a );
 a33347a <=( (not A265)  and  (not A235) );
 a33348a <=( (not A234)  and  a33347a );
 a33351a <=( (not A268)  and  (not A266) );
 a33354a <=( A300  and  A299 );
 a33355a <=( a33354a  and  a33351a );
 a33356a <=( a33355a  and  a33348a );
 a33360a <=( (not A202)  and  (not A201) );
 a33361a <=( A169  and  a33360a );
 a33365a <=( A233  and  A232 );
 a33366a <=( (not A203)  and  a33365a );
 a33367a <=( a33366a  and  a33361a );
 a33371a <=( (not A265)  and  (not A235) );
 a33372a <=( (not A234)  and  a33371a );
 a33375a <=( (not A268)  and  (not A266) );
 a33378a <=( A300  and  A298 );
 a33379a <=( a33378a  and  a33375a );
 a33380a <=( a33379a  and  a33372a );
 a33384a <=( (not A202)  and  (not A201) );
 a33385a <=( A169  and  a33384a );
 a33389a <=( (not A233)  and  (not A232) );
 a33390a <=( (not A203)  and  a33389a );
 a33391a <=( a33390a  and  a33385a );
 a33395a <=( (not A268)  and  (not A267) );
 a33396a <=( (not A235)  and  a33395a );
 a33399a <=( A298  and  (not A269) );
 a33402a <=( A302  and  (not A299) );
 a33403a <=( a33402a  and  a33399a );
 a33404a <=( a33403a  and  a33396a );
 a33408a <=( (not A202)  and  (not A201) );
 a33409a <=( A169  and  a33408a );
 a33413a <=( (not A233)  and  (not A232) );
 a33414a <=( (not A203)  and  a33413a );
 a33415a <=( a33414a  and  a33409a );
 a33419a <=( (not A268)  and  (not A267) );
 a33420a <=( (not A235)  and  a33419a );
 a33423a <=( (not A298)  and  (not A269) );
 a33426a <=( A302  and  A299 );
 a33427a <=( a33426a  and  a33423a );
 a33428a <=( a33427a  and  a33420a );
 a33432a <=( (not A202)  and  (not A201) );
 a33433a <=( A169  and  a33432a );
 a33437a <=( (not A233)  and  (not A232) );
 a33438a <=( (not A203)  and  a33437a );
 a33439a <=( a33438a  and  a33433a );
 a33443a <=( A266  and  A265 );
 a33444a <=( (not A235)  and  a33443a );
 a33447a <=( (not A268)  and  (not A267) );
 a33450a <=( A300  and  A299 );
 a33451a <=( a33450a  and  a33447a );
 a33452a <=( a33451a  and  a33444a );
 a33456a <=( (not A202)  and  (not A201) );
 a33457a <=( A169  and  a33456a );
 a33461a <=( (not A233)  and  (not A232) );
 a33462a <=( (not A203)  and  a33461a );
 a33463a <=( a33462a  and  a33457a );
 a33467a <=( A266  and  A265 );
 a33468a <=( (not A235)  and  a33467a );
 a33471a <=( (not A268)  and  (not A267) );
 a33474a <=( A300  and  A298 );
 a33475a <=( a33474a  and  a33471a );
 a33476a <=( a33475a  and  a33468a );
 a33480a <=( (not A202)  and  (not A201) );
 a33481a <=( A169  and  a33480a );
 a33485a <=( (not A233)  and  (not A232) );
 a33486a <=( (not A203)  and  a33485a );
 a33487a <=( a33486a  and  a33481a );
 a33491a <=( (not A266)  and  (not A265) );
 a33492a <=( (not A235)  and  a33491a );
 a33495a <=( A298  and  (not A268) );
 a33498a <=( A302  and  (not A299) );
 a33499a <=( a33498a  and  a33495a );
 a33500a <=( a33499a  and  a33492a );
 a33504a <=( (not A202)  and  (not A201) );
 a33505a <=( A169  and  a33504a );
 a33509a <=( (not A233)  and  (not A232) );
 a33510a <=( (not A203)  and  a33509a );
 a33511a <=( a33510a  and  a33505a );
 a33515a <=( (not A266)  and  (not A265) );
 a33516a <=( (not A235)  and  a33515a );
 a33519a <=( (not A298)  and  (not A268) );
 a33522a <=( A302  and  A299 );
 a33523a <=( a33522a  and  a33519a );
 a33524a <=( a33523a  and  a33516a );
 a33528a <=( A200  and  A199 );
 a33529a <=( A169  and  a33528a );
 a33533a <=( (not A234)  and  (not A202) );
 a33534a <=( (not A201)  and  a33533a );
 a33535a <=( a33534a  and  a33529a );
 a33539a <=( (not A267)  and  (not A236) );
 a33540a <=( (not A235)  and  a33539a );
 a33543a <=( (not A269)  and  (not A268) );
 a33546a <=( A300  and  A299 );
 a33547a <=( a33546a  and  a33543a );
 a33548a <=( a33547a  and  a33540a );
 a33552a <=( A200  and  A199 );
 a33553a <=( A169  and  a33552a );
 a33557a <=( (not A234)  and  (not A202) );
 a33558a <=( (not A201)  and  a33557a );
 a33559a <=( a33558a  and  a33553a );
 a33563a <=( (not A267)  and  (not A236) );
 a33564a <=( (not A235)  and  a33563a );
 a33567a <=( (not A269)  and  (not A268) );
 a33570a <=( A300  and  A298 );
 a33571a <=( a33570a  and  a33567a );
 a33572a <=( a33571a  and  a33564a );
 a33576a <=( A200  and  A199 );
 a33577a <=( A169  and  a33576a );
 a33581a <=( (not A234)  and  (not A202) );
 a33582a <=( (not A201)  and  a33581a );
 a33583a <=( a33582a  and  a33577a );
 a33587a <=( A265  and  (not A236) );
 a33588a <=( (not A235)  and  a33587a );
 a33591a <=( (not A267)  and  A266 );
 a33594a <=( A301  and  (not A268) );
 a33595a <=( a33594a  and  a33591a );
 a33596a <=( a33595a  and  a33588a );
 a33600a <=( A200  and  A199 );
 a33601a <=( A169  and  a33600a );
 a33605a <=( (not A234)  and  (not A202) );
 a33606a <=( (not A201)  and  a33605a );
 a33607a <=( a33606a  and  a33601a );
 a33611a <=( (not A265)  and  (not A236) );
 a33612a <=( (not A235)  and  a33611a );
 a33615a <=( (not A268)  and  (not A266) );
 a33618a <=( A300  and  A299 );
 a33619a <=( a33618a  and  a33615a );
 a33620a <=( a33619a  and  a33612a );
 a33624a <=( A200  and  A199 );
 a33625a <=( A169  and  a33624a );
 a33629a <=( (not A234)  and  (not A202) );
 a33630a <=( (not A201)  and  a33629a );
 a33631a <=( a33630a  and  a33625a );
 a33635a <=( (not A265)  and  (not A236) );
 a33636a <=( (not A235)  and  a33635a );
 a33639a <=( (not A268)  and  (not A266) );
 a33642a <=( A300  and  A298 );
 a33643a <=( a33642a  and  a33639a );
 a33644a <=( a33643a  and  a33636a );
 a33648a <=( A200  and  A199 );
 a33649a <=( A169  and  a33648a );
 a33653a <=( A232  and  (not A202) );
 a33654a <=( (not A201)  and  a33653a );
 a33655a <=( a33654a  and  a33649a );
 a33659a <=( (not A235)  and  (not A234) );
 a33660a <=( A233  and  a33659a );
 a33663a <=( (not A268)  and  (not A267) );
 a33666a <=( A301  and  (not A269) );
 a33667a <=( a33666a  and  a33663a );
 a33668a <=( a33667a  and  a33660a );
 a33672a <=( A200  and  A199 );
 a33673a <=( A169  and  a33672a );
 a33677a <=( A232  and  (not A202) );
 a33678a <=( (not A201)  and  a33677a );
 a33679a <=( a33678a  and  a33673a );
 a33683a <=( (not A235)  and  (not A234) );
 a33684a <=( A233  and  a33683a );
 a33687a <=( (not A266)  and  (not A265) );
 a33690a <=( A301  and  (not A268) );
 a33691a <=( a33690a  and  a33687a );
 a33692a <=( a33691a  and  a33684a );
 a33696a <=( A200  and  A199 );
 a33697a <=( A169  and  a33696a );
 a33701a <=( (not A232)  and  (not A202) );
 a33702a <=( (not A201)  and  a33701a );
 a33703a <=( a33702a  and  a33697a );
 a33707a <=( (not A267)  and  (not A235) );
 a33708a <=( (not A233)  and  a33707a );
 a33711a <=( (not A269)  and  (not A268) );
 a33714a <=( A300  and  A299 );
 a33715a <=( a33714a  and  a33711a );
 a33716a <=( a33715a  and  a33708a );
 a33720a <=( A200  and  A199 );
 a33721a <=( A169  and  a33720a );
 a33725a <=( (not A232)  and  (not A202) );
 a33726a <=( (not A201)  and  a33725a );
 a33727a <=( a33726a  and  a33721a );
 a33731a <=( (not A267)  and  (not A235) );
 a33732a <=( (not A233)  and  a33731a );
 a33735a <=( (not A269)  and  (not A268) );
 a33738a <=( A300  and  A298 );
 a33739a <=( a33738a  and  a33735a );
 a33740a <=( a33739a  and  a33732a );
 a33744a <=( A200  and  A199 );
 a33745a <=( A169  and  a33744a );
 a33749a <=( (not A232)  and  (not A202) );
 a33750a <=( (not A201)  and  a33749a );
 a33751a <=( a33750a  and  a33745a );
 a33755a <=( A265  and  (not A235) );
 a33756a <=( (not A233)  and  a33755a );
 a33759a <=( (not A267)  and  A266 );
 a33762a <=( A301  and  (not A268) );
 a33763a <=( a33762a  and  a33759a );
 a33764a <=( a33763a  and  a33756a );
 a33768a <=( A200  and  A199 );
 a33769a <=( A169  and  a33768a );
 a33773a <=( (not A232)  and  (not A202) );
 a33774a <=( (not A201)  and  a33773a );
 a33775a <=( a33774a  and  a33769a );
 a33779a <=( (not A265)  and  (not A235) );
 a33780a <=( (not A233)  and  a33779a );
 a33783a <=( (not A268)  and  (not A266) );
 a33786a <=( A300  and  A299 );
 a33787a <=( a33786a  and  a33783a );
 a33788a <=( a33787a  and  a33780a );
 a33792a <=( A200  and  A199 );
 a33793a <=( A169  and  a33792a );
 a33797a <=( (not A232)  and  (not A202) );
 a33798a <=( (not A201)  and  a33797a );
 a33799a <=( a33798a  and  a33793a );
 a33803a <=( (not A265)  and  (not A235) );
 a33804a <=( (not A233)  and  a33803a );
 a33807a <=( (not A268)  and  (not A266) );
 a33810a <=( A300  and  A298 );
 a33811a <=( a33810a  and  a33807a );
 a33812a <=( a33811a  and  a33804a );
 a33816a <=( (not A200)  and  (not A199) );
 a33817a <=( A169  and  a33816a );
 a33821a <=( (not A235)  and  (not A234) );
 a33822a <=( (not A202)  and  a33821a );
 a33823a <=( a33822a  and  a33817a );
 a33827a <=( (not A268)  and  (not A267) );
 a33828a <=( (not A236)  and  a33827a );
 a33831a <=( A298  and  (not A269) );
 a33834a <=( A302  and  (not A299) );
 a33835a <=( a33834a  and  a33831a );
 a33836a <=( a33835a  and  a33828a );
 a33840a <=( (not A200)  and  (not A199) );
 a33841a <=( A169  and  a33840a );
 a33845a <=( (not A235)  and  (not A234) );
 a33846a <=( (not A202)  and  a33845a );
 a33847a <=( a33846a  and  a33841a );
 a33851a <=( (not A268)  and  (not A267) );
 a33852a <=( (not A236)  and  a33851a );
 a33855a <=( (not A298)  and  (not A269) );
 a33858a <=( A302  and  A299 );
 a33859a <=( a33858a  and  a33855a );
 a33860a <=( a33859a  and  a33852a );
 a33864a <=( (not A200)  and  (not A199) );
 a33865a <=( A169  and  a33864a );
 a33869a <=( (not A235)  and  (not A234) );
 a33870a <=( (not A202)  and  a33869a );
 a33871a <=( a33870a  and  a33865a );
 a33875a <=( A266  and  A265 );
 a33876a <=( (not A236)  and  a33875a );
 a33879a <=( (not A268)  and  (not A267) );
 a33882a <=( A300  and  A299 );
 a33883a <=( a33882a  and  a33879a );
 a33884a <=( a33883a  and  a33876a );
 a33888a <=( (not A200)  and  (not A199) );
 a33889a <=( A169  and  a33888a );
 a33893a <=( (not A235)  and  (not A234) );
 a33894a <=( (not A202)  and  a33893a );
 a33895a <=( a33894a  and  a33889a );
 a33899a <=( A266  and  A265 );
 a33900a <=( (not A236)  and  a33899a );
 a33903a <=( (not A268)  and  (not A267) );
 a33906a <=( A300  and  A298 );
 a33907a <=( a33906a  and  a33903a );
 a33908a <=( a33907a  and  a33900a );
 a33912a <=( (not A200)  and  (not A199) );
 a33913a <=( A169  and  a33912a );
 a33917a <=( (not A235)  and  (not A234) );
 a33918a <=( (not A202)  and  a33917a );
 a33919a <=( a33918a  and  a33913a );
 a33923a <=( (not A266)  and  (not A265) );
 a33924a <=( (not A236)  and  a33923a );
 a33927a <=( A298  and  (not A268) );
 a33930a <=( A302  and  (not A299) );
 a33931a <=( a33930a  and  a33927a );
 a33932a <=( a33931a  and  a33924a );
 a33936a <=( (not A200)  and  (not A199) );
 a33937a <=( A169  and  a33936a );
 a33941a <=( (not A235)  and  (not A234) );
 a33942a <=( (not A202)  and  a33941a );
 a33943a <=( a33942a  and  a33937a );
 a33947a <=( (not A266)  and  (not A265) );
 a33948a <=( (not A236)  and  a33947a );
 a33951a <=( (not A298)  and  (not A268) );
 a33954a <=( A302  and  A299 );
 a33955a <=( a33954a  and  a33951a );
 a33956a <=( a33955a  and  a33948a );
 a33960a <=( (not A200)  and  (not A199) );
 a33961a <=( A169  and  a33960a );
 a33965a <=( A233  and  A232 );
 a33966a <=( (not A202)  and  a33965a );
 a33967a <=( a33966a  and  a33961a );
 a33971a <=( (not A267)  and  (not A235) );
 a33972a <=( (not A234)  and  a33971a );
 a33975a <=( (not A269)  and  (not A268) );
 a33978a <=( A300  and  A299 );
 a33979a <=( a33978a  and  a33975a );
 a33980a <=( a33979a  and  a33972a );
 a33984a <=( (not A200)  and  (not A199) );
 a33985a <=( A169  and  a33984a );
 a33989a <=( A233  and  A232 );
 a33990a <=( (not A202)  and  a33989a );
 a33991a <=( a33990a  and  a33985a );
 a33995a <=( (not A267)  and  (not A235) );
 a33996a <=( (not A234)  and  a33995a );
 a33999a <=( (not A269)  and  (not A268) );
 a34002a <=( A300  and  A298 );
 a34003a <=( a34002a  and  a33999a );
 a34004a <=( a34003a  and  a33996a );
 a34008a <=( (not A200)  and  (not A199) );
 a34009a <=( A169  and  a34008a );
 a34013a <=( A233  and  A232 );
 a34014a <=( (not A202)  and  a34013a );
 a34015a <=( a34014a  and  a34009a );
 a34019a <=( A265  and  (not A235) );
 a34020a <=( (not A234)  and  a34019a );
 a34023a <=( (not A267)  and  A266 );
 a34026a <=( A301  and  (not A268) );
 a34027a <=( a34026a  and  a34023a );
 a34028a <=( a34027a  and  a34020a );
 a34032a <=( (not A200)  and  (not A199) );
 a34033a <=( A169  and  a34032a );
 a34037a <=( A233  and  A232 );
 a34038a <=( (not A202)  and  a34037a );
 a34039a <=( a34038a  and  a34033a );
 a34043a <=( (not A265)  and  (not A235) );
 a34044a <=( (not A234)  and  a34043a );
 a34047a <=( (not A268)  and  (not A266) );
 a34050a <=( A300  and  A299 );
 a34051a <=( a34050a  and  a34047a );
 a34052a <=( a34051a  and  a34044a );
 a34056a <=( (not A200)  and  (not A199) );
 a34057a <=( A169  and  a34056a );
 a34061a <=( A233  and  A232 );
 a34062a <=( (not A202)  and  a34061a );
 a34063a <=( a34062a  and  a34057a );
 a34067a <=( (not A265)  and  (not A235) );
 a34068a <=( (not A234)  and  a34067a );
 a34071a <=( (not A268)  and  (not A266) );
 a34074a <=( A300  and  A298 );
 a34075a <=( a34074a  and  a34071a );
 a34076a <=( a34075a  and  a34068a );
 a34080a <=( (not A200)  and  (not A199) );
 a34081a <=( A169  and  a34080a );
 a34085a <=( (not A233)  and  (not A232) );
 a34086a <=( (not A202)  and  a34085a );
 a34087a <=( a34086a  and  a34081a );
 a34091a <=( (not A268)  and  (not A267) );
 a34092a <=( (not A235)  and  a34091a );
 a34095a <=( A298  and  (not A269) );
 a34098a <=( A302  and  (not A299) );
 a34099a <=( a34098a  and  a34095a );
 a34100a <=( a34099a  and  a34092a );
 a34104a <=( (not A200)  and  (not A199) );
 a34105a <=( A169  and  a34104a );
 a34109a <=( (not A233)  and  (not A232) );
 a34110a <=( (not A202)  and  a34109a );
 a34111a <=( a34110a  and  a34105a );
 a34115a <=( (not A268)  and  (not A267) );
 a34116a <=( (not A235)  and  a34115a );
 a34119a <=( (not A298)  and  (not A269) );
 a34122a <=( A302  and  A299 );
 a34123a <=( a34122a  and  a34119a );
 a34124a <=( a34123a  and  a34116a );
 a34128a <=( (not A200)  and  (not A199) );
 a34129a <=( A169  and  a34128a );
 a34133a <=( (not A233)  and  (not A232) );
 a34134a <=( (not A202)  and  a34133a );
 a34135a <=( a34134a  and  a34129a );
 a34139a <=( A266  and  A265 );
 a34140a <=( (not A235)  and  a34139a );
 a34143a <=( (not A268)  and  (not A267) );
 a34146a <=( A300  and  A299 );
 a34147a <=( a34146a  and  a34143a );
 a34148a <=( a34147a  and  a34140a );
 a34152a <=( (not A200)  and  (not A199) );
 a34153a <=( A169  and  a34152a );
 a34157a <=( (not A233)  and  (not A232) );
 a34158a <=( (not A202)  and  a34157a );
 a34159a <=( a34158a  and  a34153a );
 a34163a <=( A266  and  A265 );
 a34164a <=( (not A235)  and  a34163a );
 a34167a <=( (not A268)  and  (not A267) );
 a34170a <=( A300  and  A298 );
 a34171a <=( a34170a  and  a34167a );
 a34172a <=( a34171a  and  a34164a );
 a34176a <=( (not A200)  and  (not A199) );
 a34177a <=( A169  and  a34176a );
 a34181a <=( (not A233)  and  (not A232) );
 a34182a <=( (not A202)  and  a34181a );
 a34183a <=( a34182a  and  a34177a );
 a34187a <=( (not A266)  and  (not A265) );
 a34188a <=( (not A235)  and  a34187a );
 a34191a <=( A298  and  (not A268) );
 a34194a <=( A302  and  (not A299) );
 a34195a <=( a34194a  and  a34191a );
 a34196a <=( a34195a  and  a34188a );
 a34200a <=( (not A200)  and  (not A199) );
 a34201a <=( A169  and  a34200a );
 a34205a <=( (not A233)  and  (not A232) );
 a34206a <=( (not A202)  and  a34205a );
 a34207a <=( a34206a  and  a34201a );
 a34211a <=( (not A266)  and  (not A265) );
 a34212a <=( (not A235)  and  a34211a );
 a34215a <=( (not A298)  and  (not A268) );
 a34218a <=( A302  and  A299 );
 a34219a <=( a34218a  and  a34215a );
 a34220a <=( a34219a  and  a34212a );
 a34224a <=( (not A166)  and  (not A167) );
 a34225a <=( (not A169)  and  a34224a );
 a34229a <=( (not A235)  and  (not A234) );
 a34230a <=( A202  and  a34229a );
 a34231a <=( a34230a  and  a34225a );
 a34235a <=( (not A268)  and  (not A267) );
 a34236a <=( (not A236)  and  a34235a );
 a34239a <=( A298  and  (not A269) );
 a34242a <=( A302  and  (not A299) );
 a34243a <=( a34242a  and  a34239a );
 a34244a <=( a34243a  and  a34236a );
 a34248a <=( (not A166)  and  (not A167) );
 a34249a <=( (not A169)  and  a34248a );
 a34253a <=( (not A235)  and  (not A234) );
 a34254a <=( A202  and  a34253a );
 a34255a <=( a34254a  and  a34249a );
 a34259a <=( (not A268)  and  (not A267) );
 a34260a <=( (not A236)  and  a34259a );
 a34263a <=( (not A298)  and  (not A269) );
 a34266a <=( A302  and  A299 );
 a34267a <=( a34266a  and  a34263a );
 a34268a <=( a34267a  and  a34260a );
 a34272a <=( (not A166)  and  (not A167) );
 a34273a <=( (not A169)  and  a34272a );
 a34277a <=( (not A235)  and  (not A234) );
 a34278a <=( A202  and  a34277a );
 a34279a <=( a34278a  and  a34273a );
 a34283a <=( A266  and  A265 );
 a34284a <=( (not A236)  and  a34283a );
 a34287a <=( (not A268)  and  (not A267) );
 a34290a <=( A300  and  A299 );
 a34291a <=( a34290a  and  a34287a );
 a34292a <=( a34291a  and  a34284a );
 a34296a <=( (not A166)  and  (not A167) );
 a34297a <=( (not A169)  and  a34296a );
 a34301a <=( (not A235)  and  (not A234) );
 a34302a <=( A202  and  a34301a );
 a34303a <=( a34302a  and  a34297a );
 a34307a <=( A266  and  A265 );
 a34308a <=( (not A236)  and  a34307a );
 a34311a <=( (not A268)  and  (not A267) );
 a34314a <=( A300  and  A298 );
 a34315a <=( a34314a  and  a34311a );
 a34316a <=( a34315a  and  a34308a );
 a34320a <=( (not A166)  and  (not A167) );
 a34321a <=( (not A169)  and  a34320a );
 a34325a <=( (not A235)  and  (not A234) );
 a34326a <=( A202  and  a34325a );
 a34327a <=( a34326a  and  a34321a );
 a34331a <=( (not A266)  and  (not A265) );
 a34332a <=( (not A236)  and  a34331a );
 a34335a <=( A298  and  (not A268) );
 a34338a <=( A302  and  (not A299) );
 a34339a <=( a34338a  and  a34335a );
 a34340a <=( a34339a  and  a34332a );
 a34344a <=( (not A166)  and  (not A167) );
 a34345a <=( (not A169)  and  a34344a );
 a34349a <=( (not A235)  and  (not A234) );
 a34350a <=( A202  and  a34349a );
 a34351a <=( a34350a  and  a34345a );
 a34355a <=( (not A266)  and  (not A265) );
 a34356a <=( (not A236)  and  a34355a );
 a34359a <=( (not A298)  and  (not A268) );
 a34362a <=( A302  and  A299 );
 a34363a <=( a34362a  and  a34359a );
 a34364a <=( a34363a  and  a34356a );
 a34368a <=( (not A166)  and  (not A167) );
 a34369a <=( (not A169)  and  a34368a );
 a34373a <=( A233  and  A232 );
 a34374a <=( A202  and  a34373a );
 a34375a <=( a34374a  and  a34369a );
 a34379a <=( (not A267)  and  (not A235) );
 a34380a <=( (not A234)  and  a34379a );
 a34383a <=( (not A269)  and  (not A268) );
 a34386a <=( A300  and  A299 );
 a34387a <=( a34386a  and  a34383a );
 a34388a <=( a34387a  and  a34380a );
 a34392a <=( (not A166)  and  (not A167) );
 a34393a <=( (not A169)  and  a34392a );
 a34397a <=( A233  and  A232 );
 a34398a <=( A202  and  a34397a );
 a34399a <=( a34398a  and  a34393a );
 a34403a <=( (not A267)  and  (not A235) );
 a34404a <=( (not A234)  and  a34403a );
 a34407a <=( (not A269)  and  (not A268) );
 a34410a <=( A300  and  A298 );
 a34411a <=( a34410a  and  a34407a );
 a34412a <=( a34411a  and  a34404a );
 a34416a <=( (not A166)  and  (not A167) );
 a34417a <=( (not A169)  and  a34416a );
 a34421a <=( A233  and  A232 );
 a34422a <=( A202  and  a34421a );
 a34423a <=( a34422a  and  a34417a );
 a34427a <=( A265  and  (not A235) );
 a34428a <=( (not A234)  and  a34427a );
 a34431a <=( (not A267)  and  A266 );
 a34434a <=( A301  and  (not A268) );
 a34435a <=( a34434a  and  a34431a );
 a34436a <=( a34435a  and  a34428a );
 a34440a <=( (not A166)  and  (not A167) );
 a34441a <=( (not A169)  and  a34440a );
 a34445a <=( A233  and  A232 );
 a34446a <=( A202  and  a34445a );
 a34447a <=( a34446a  and  a34441a );
 a34451a <=( (not A265)  and  (not A235) );
 a34452a <=( (not A234)  and  a34451a );
 a34455a <=( (not A268)  and  (not A266) );
 a34458a <=( A300  and  A299 );
 a34459a <=( a34458a  and  a34455a );
 a34460a <=( a34459a  and  a34452a );
 a34464a <=( (not A166)  and  (not A167) );
 a34465a <=( (not A169)  and  a34464a );
 a34469a <=( A233  and  A232 );
 a34470a <=( A202  and  a34469a );
 a34471a <=( a34470a  and  a34465a );
 a34475a <=( (not A265)  and  (not A235) );
 a34476a <=( (not A234)  and  a34475a );
 a34479a <=( (not A268)  and  (not A266) );
 a34482a <=( A300  and  A298 );
 a34483a <=( a34482a  and  a34479a );
 a34484a <=( a34483a  and  a34476a );
 a34488a <=( (not A166)  and  (not A167) );
 a34489a <=( (not A169)  and  a34488a );
 a34493a <=( (not A233)  and  (not A232) );
 a34494a <=( A202  and  a34493a );
 a34495a <=( a34494a  and  a34489a );
 a34499a <=( (not A268)  and  (not A267) );
 a34500a <=( (not A235)  and  a34499a );
 a34503a <=( A298  and  (not A269) );
 a34506a <=( A302  and  (not A299) );
 a34507a <=( a34506a  and  a34503a );
 a34508a <=( a34507a  and  a34500a );
 a34512a <=( (not A166)  and  (not A167) );
 a34513a <=( (not A169)  and  a34512a );
 a34517a <=( (not A233)  and  (not A232) );
 a34518a <=( A202  and  a34517a );
 a34519a <=( a34518a  and  a34513a );
 a34523a <=( (not A268)  and  (not A267) );
 a34524a <=( (not A235)  and  a34523a );
 a34527a <=( (not A298)  and  (not A269) );
 a34530a <=( A302  and  A299 );
 a34531a <=( a34530a  and  a34527a );
 a34532a <=( a34531a  and  a34524a );
 a34536a <=( (not A166)  and  (not A167) );
 a34537a <=( (not A169)  and  a34536a );
 a34541a <=( (not A233)  and  (not A232) );
 a34542a <=( A202  and  a34541a );
 a34543a <=( a34542a  and  a34537a );
 a34547a <=( A266  and  A265 );
 a34548a <=( (not A235)  and  a34547a );
 a34551a <=( (not A268)  and  (not A267) );
 a34554a <=( A300  and  A299 );
 a34555a <=( a34554a  and  a34551a );
 a34556a <=( a34555a  and  a34548a );
 a34560a <=( (not A166)  and  (not A167) );
 a34561a <=( (not A169)  and  a34560a );
 a34565a <=( (not A233)  and  (not A232) );
 a34566a <=( A202  and  a34565a );
 a34567a <=( a34566a  and  a34561a );
 a34571a <=( A266  and  A265 );
 a34572a <=( (not A235)  and  a34571a );
 a34575a <=( (not A268)  and  (not A267) );
 a34578a <=( A300  and  A298 );
 a34579a <=( a34578a  and  a34575a );
 a34580a <=( a34579a  and  a34572a );
 a34584a <=( (not A166)  and  (not A167) );
 a34585a <=( (not A169)  and  a34584a );
 a34589a <=( (not A233)  and  (not A232) );
 a34590a <=( A202  and  a34589a );
 a34591a <=( a34590a  and  a34585a );
 a34595a <=( (not A266)  and  (not A265) );
 a34596a <=( (not A235)  and  a34595a );
 a34599a <=( A298  and  (not A268) );
 a34602a <=( A302  and  (not A299) );
 a34603a <=( a34602a  and  a34599a );
 a34604a <=( a34603a  and  a34596a );
 a34608a <=( (not A166)  and  (not A167) );
 a34609a <=( (not A169)  and  a34608a );
 a34613a <=( (not A233)  and  (not A232) );
 a34614a <=( A202  and  a34613a );
 a34615a <=( a34614a  and  a34609a );
 a34619a <=( (not A266)  and  (not A265) );
 a34620a <=( (not A235)  and  a34619a );
 a34623a <=( (not A298)  and  (not A268) );
 a34626a <=( A302  and  A299 );
 a34627a <=( a34626a  and  a34623a );
 a34628a <=( a34627a  and  a34620a );
 a34632a <=( (not A166)  and  (not A167) );
 a34633a <=( (not A169)  and  a34632a );
 a34637a <=( (not A234)  and  A201 );
 a34638a <=( A199  and  a34637a );
 a34639a <=( a34638a  and  a34633a );
 a34643a <=( (not A267)  and  (not A236) );
 a34644a <=( (not A235)  and  a34643a );
 a34647a <=( (not A269)  and  (not A268) );
 a34650a <=( A300  and  A299 );
 a34651a <=( a34650a  and  a34647a );
 a34652a <=( a34651a  and  a34644a );
 a34656a <=( (not A166)  and  (not A167) );
 a34657a <=( (not A169)  and  a34656a );
 a34661a <=( (not A234)  and  A201 );
 a34662a <=( A199  and  a34661a );
 a34663a <=( a34662a  and  a34657a );
 a34667a <=( (not A267)  and  (not A236) );
 a34668a <=( (not A235)  and  a34667a );
 a34671a <=( (not A269)  and  (not A268) );
 a34674a <=( A300  and  A298 );
 a34675a <=( a34674a  and  a34671a );
 a34676a <=( a34675a  and  a34668a );
 a34680a <=( (not A166)  and  (not A167) );
 a34681a <=( (not A169)  and  a34680a );
 a34685a <=( (not A234)  and  A201 );
 a34686a <=( A199  and  a34685a );
 a34687a <=( a34686a  and  a34681a );
 a34691a <=( A265  and  (not A236) );
 a34692a <=( (not A235)  and  a34691a );
 a34695a <=( (not A267)  and  A266 );
 a34698a <=( A301  and  (not A268) );
 a34699a <=( a34698a  and  a34695a );
 a34700a <=( a34699a  and  a34692a );
 a34704a <=( (not A166)  and  (not A167) );
 a34705a <=( (not A169)  and  a34704a );
 a34709a <=( (not A234)  and  A201 );
 a34710a <=( A199  and  a34709a );
 a34711a <=( a34710a  and  a34705a );
 a34715a <=( (not A265)  and  (not A236) );
 a34716a <=( (not A235)  and  a34715a );
 a34719a <=( (not A268)  and  (not A266) );
 a34722a <=( A300  and  A299 );
 a34723a <=( a34722a  and  a34719a );
 a34724a <=( a34723a  and  a34716a );
 a34728a <=( (not A166)  and  (not A167) );
 a34729a <=( (not A169)  and  a34728a );
 a34733a <=( (not A234)  and  A201 );
 a34734a <=( A199  and  a34733a );
 a34735a <=( a34734a  and  a34729a );
 a34739a <=( (not A265)  and  (not A236) );
 a34740a <=( (not A235)  and  a34739a );
 a34743a <=( (not A268)  and  (not A266) );
 a34746a <=( A300  and  A298 );
 a34747a <=( a34746a  and  a34743a );
 a34748a <=( a34747a  and  a34740a );
 a34752a <=( (not A166)  and  (not A167) );
 a34753a <=( (not A169)  and  a34752a );
 a34757a <=( A232  and  A201 );
 a34758a <=( A199  and  a34757a );
 a34759a <=( a34758a  and  a34753a );
 a34763a <=( (not A235)  and  (not A234) );
 a34764a <=( A233  and  a34763a );
 a34767a <=( (not A268)  and  (not A267) );
 a34770a <=( A301  and  (not A269) );
 a34771a <=( a34770a  and  a34767a );
 a34772a <=( a34771a  and  a34764a );
 a34776a <=( (not A166)  and  (not A167) );
 a34777a <=( (not A169)  and  a34776a );
 a34781a <=( A232  and  A201 );
 a34782a <=( A199  and  a34781a );
 a34783a <=( a34782a  and  a34777a );
 a34787a <=( (not A235)  and  (not A234) );
 a34788a <=( A233  and  a34787a );
 a34791a <=( (not A266)  and  (not A265) );
 a34794a <=( A301  and  (not A268) );
 a34795a <=( a34794a  and  a34791a );
 a34796a <=( a34795a  and  a34788a );
 a34800a <=( (not A166)  and  (not A167) );
 a34801a <=( (not A169)  and  a34800a );
 a34805a <=( (not A232)  and  A201 );
 a34806a <=( A199  and  a34805a );
 a34807a <=( a34806a  and  a34801a );
 a34811a <=( (not A267)  and  (not A235) );
 a34812a <=( (not A233)  and  a34811a );
 a34815a <=( (not A269)  and  (not A268) );
 a34818a <=( A300  and  A299 );
 a34819a <=( a34818a  and  a34815a );
 a34820a <=( a34819a  and  a34812a );
 a34824a <=( (not A166)  and  (not A167) );
 a34825a <=( (not A169)  and  a34824a );
 a34829a <=( (not A232)  and  A201 );
 a34830a <=( A199  and  a34829a );
 a34831a <=( a34830a  and  a34825a );
 a34835a <=( (not A267)  and  (not A235) );
 a34836a <=( (not A233)  and  a34835a );
 a34839a <=( (not A269)  and  (not A268) );
 a34842a <=( A300  and  A298 );
 a34843a <=( a34842a  and  a34839a );
 a34844a <=( a34843a  and  a34836a );
 a34848a <=( (not A166)  and  (not A167) );
 a34849a <=( (not A169)  and  a34848a );
 a34853a <=( (not A232)  and  A201 );
 a34854a <=( A199  and  a34853a );
 a34855a <=( a34854a  and  a34849a );
 a34859a <=( A265  and  (not A235) );
 a34860a <=( (not A233)  and  a34859a );
 a34863a <=( (not A267)  and  A266 );
 a34866a <=( A301  and  (not A268) );
 a34867a <=( a34866a  and  a34863a );
 a34868a <=( a34867a  and  a34860a );
 a34872a <=( (not A166)  and  (not A167) );
 a34873a <=( (not A169)  and  a34872a );
 a34877a <=( (not A232)  and  A201 );
 a34878a <=( A199  and  a34877a );
 a34879a <=( a34878a  and  a34873a );
 a34883a <=( (not A265)  and  (not A235) );
 a34884a <=( (not A233)  and  a34883a );
 a34887a <=( (not A268)  and  (not A266) );
 a34890a <=( A300  and  A299 );
 a34891a <=( a34890a  and  a34887a );
 a34892a <=( a34891a  and  a34884a );
 a34896a <=( (not A166)  and  (not A167) );
 a34897a <=( (not A169)  and  a34896a );
 a34901a <=( (not A232)  and  A201 );
 a34902a <=( A199  and  a34901a );
 a34903a <=( a34902a  and  a34897a );
 a34907a <=( (not A265)  and  (not A235) );
 a34908a <=( (not A233)  and  a34907a );
 a34911a <=( (not A268)  and  (not A266) );
 a34914a <=( A300  and  A298 );
 a34915a <=( a34914a  and  a34911a );
 a34916a <=( a34915a  and  a34908a );
 a34920a <=( (not A166)  and  (not A167) );
 a34921a <=( (not A169)  and  a34920a );
 a34925a <=( (not A234)  and  A201 );
 a34926a <=( A200  and  a34925a );
 a34927a <=( a34926a  and  a34921a );
 a34931a <=( (not A267)  and  (not A236) );
 a34932a <=( (not A235)  and  a34931a );
 a34935a <=( (not A269)  and  (not A268) );
 a34938a <=( A300  and  A299 );
 a34939a <=( a34938a  and  a34935a );
 a34940a <=( a34939a  and  a34932a );
 a34944a <=( (not A166)  and  (not A167) );
 a34945a <=( (not A169)  and  a34944a );
 a34949a <=( (not A234)  and  A201 );
 a34950a <=( A200  and  a34949a );
 a34951a <=( a34950a  and  a34945a );
 a34955a <=( (not A267)  and  (not A236) );
 a34956a <=( (not A235)  and  a34955a );
 a34959a <=( (not A269)  and  (not A268) );
 a34962a <=( A300  and  A298 );
 a34963a <=( a34962a  and  a34959a );
 a34964a <=( a34963a  and  a34956a );
 a34968a <=( (not A166)  and  (not A167) );
 a34969a <=( (not A169)  and  a34968a );
 a34973a <=( (not A234)  and  A201 );
 a34974a <=( A200  and  a34973a );
 a34975a <=( a34974a  and  a34969a );
 a34979a <=( A265  and  (not A236) );
 a34980a <=( (not A235)  and  a34979a );
 a34983a <=( (not A267)  and  A266 );
 a34986a <=( A301  and  (not A268) );
 a34987a <=( a34986a  and  a34983a );
 a34988a <=( a34987a  and  a34980a );
 a34992a <=( (not A166)  and  (not A167) );
 a34993a <=( (not A169)  and  a34992a );
 a34997a <=( (not A234)  and  A201 );
 a34998a <=( A200  and  a34997a );
 a34999a <=( a34998a  and  a34993a );
 a35003a <=( (not A265)  and  (not A236) );
 a35004a <=( (not A235)  and  a35003a );
 a35007a <=( (not A268)  and  (not A266) );
 a35010a <=( A300  and  A299 );
 a35011a <=( a35010a  and  a35007a );
 a35012a <=( a35011a  and  a35004a );
 a35016a <=( (not A166)  and  (not A167) );
 a35017a <=( (not A169)  and  a35016a );
 a35021a <=( (not A234)  and  A201 );
 a35022a <=( A200  and  a35021a );
 a35023a <=( a35022a  and  a35017a );
 a35027a <=( (not A265)  and  (not A236) );
 a35028a <=( (not A235)  and  a35027a );
 a35031a <=( (not A268)  and  (not A266) );
 a35034a <=( A300  and  A298 );
 a35035a <=( a35034a  and  a35031a );
 a35036a <=( a35035a  and  a35028a );
 a35040a <=( (not A166)  and  (not A167) );
 a35041a <=( (not A169)  and  a35040a );
 a35045a <=( A232  and  A201 );
 a35046a <=( A200  and  a35045a );
 a35047a <=( a35046a  and  a35041a );
 a35051a <=( (not A235)  and  (not A234) );
 a35052a <=( A233  and  a35051a );
 a35055a <=( (not A268)  and  (not A267) );
 a35058a <=( A301  and  (not A269) );
 a35059a <=( a35058a  and  a35055a );
 a35060a <=( a35059a  and  a35052a );
 a35064a <=( (not A166)  and  (not A167) );
 a35065a <=( (not A169)  and  a35064a );
 a35069a <=( A232  and  A201 );
 a35070a <=( A200  and  a35069a );
 a35071a <=( a35070a  and  a35065a );
 a35075a <=( (not A235)  and  (not A234) );
 a35076a <=( A233  and  a35075a );
 a35079a <=( (not A266)  and  (not A265) );
 a35082a <=( A301  and  (not A268) );
 a35083a <=( a35082a  and  a35079a );
 a35084a <=( a35083a  and  a35076a );
 a35088a <=( (not A166)  and  (not A167) );
 a35089a <=( (not A169)  and  a35088a );
 a35093a <=( (not A232)  and  A201 );
 a35094a <=( A200  and  a35093a );
 a35095a <=( a35094a  and  a35089a );
 a35099a <=( (not A267)  and  (not A235) );
 a35100a <=( (not A233)  and  a35099a );
 a35103a <=( (not A269)  and  (not A268) );
 a35106a <=( A300  and  A299 );
 a35107a <=( a35106a  and  a35103a );
 a35108a <=( a35107a  and  a35100a );
 a35112a <=( (not A166)  and  (not A167) );
 a35113a <=( (not A169)  and  a35112a );
 a35117a <=( (not A232)  and  A201 );
 a35118a <=( A200  and  a35117a );
 a35119a <=( a35118a  and  a35113a );
 a35123a <=( (not A267)  and  (not A235) );
 a35124a <=( (not A233)  and  a35123a );
 a35127a <=( (not A269)  and  (not A268) );
 a35130a <=( A300  and  A298 );
 a35131a <=( a35130a  and  a35127a );
 a35132a <=( a35131a  and  a35124a );
 a35136a <=( (not A166)  and  (not A167) );
 a35137a <=( (not A169)  and  a35136a );
 a35141a <=( (not A232)  and  A201 );
 a35142a <=( A200  and  a35141a );
 a35143a <=( a35142a  and  a35137a );
 a35147a <=( A265  and  (not A235) );
 a35148a <=( (not A233)  and  a35147a );
 a35151a <=( (not A267)  and  A266 );
 a35154a <=( A301  and  (not A268) );
 a35155a <=( a35154a  and  a35151a );
 a35156a <=( a35155a  and  a35148a );
 a35160a <=( (not A166)  and  (not A167) );
 a35161a <=( (not A169)  and  a35160a );
 a35165a <=( (not A232)  and  A201 );
 a35166a <=( A200  and  a35165a );
 a35167a <=( a35166a  and  a35161a );
 a35171a <=( (not A265)  and  (not A235) );
 a35172a <=( (not A233)  and  a35171a );
 a35175a <=( (not A268)  and  (not A266) );
 a35178a <=( A300  and  A299 );
 a35179a <=( a35178a  and  a35175a );
 a35180a <=( a35179a  and  a35172a );
 a35184a <=( (not A166)  and  (not A167) );
 a35185a <=( (not A169)  and  a35184a );
 a35189a <=( (not A232)  and  A201 );
 a35190a <=( A200  and  a35189a );
 a35191a <=( a35190a  and  a35185a );
 a35195a <=( (not A265)  and  (not A235) );
 a35196a <=( (not A233)  and  a35195a );
 a35199a <=( (not A268)  and  (not A266) );
 a35202a <=( A300  and  A298 );
 a35203a <=( a35202a  and  a35199a );
 a35204a <=( a35203a  and  a35196a );
 a35208a <=( (not A166)  and  (not A167) );
 a35209a <=( (not A169)  and  a35208a );
 a35213a <=( A203  and  A200 );
 a35214a <=( (not A199)  and  a35213a );
 a35215a <=( a35214a  and  a35209a );
 a35219a <=( (not A236)  and  (not A235) );
 a35220a <=( (not A234)  and  a35219a );
 a35223a <=( (not A268)  and  (not A267) );
 a35226a <=( A301  and  (not A269) );
 a35227a <=( a35226a  and  a35223a );
 a35228a <=( a35227a  and  a35220a );
 a35232a <=( (not A166)  and  (not A167) );
 a35233a <=( (not A169)  and  a35232a );
 a35237a <=( A203  and  A200 );
 a35238a <=( (not A199)  and  a35237a );
 a35239a <=( a35238a  and  a35233a );
 a35243a <=( (not A236)  and  (not A235) );
 a35244a <=( (not A234)  and  a35243a );
 a35247a <=( (not A266)  and  (not A265) );
 a35250a <=( A301  and  (not A268) );
 a35251a <=( a35250a  and  a35247a );
 a35252a <=( a35251a  and  a35244a );
 a35256a <=( (not A166)  and  (not A167) );
 a35257a <=( (not A169)  and  a35256a );
 a35261a <=( A203  and  A200 );
 a35262a <=( (not A199)  and  a35261a );
 a35263a <=( a35262a  and  a35257a );
 a35267a <=( A236  and  A233 );
 a35268a <=( (not A232)  and  a35267a );
 a35271a <=( A299  and  A298 );
 a35274a <=( (not A301)  and  (not A300) );
 a35275a <=( a35274a  and  a35271a );
 a35276a <=( a35275a  and  a35268a );
 a35280a <=( (not A166)  and  (not A167) );
 a35281a <=( (not A169)  and  a35280a );
 a35285a <=( A203  and  A200 );
 a35286a <=( (not A199)  and  a35285a );
 a35287a <=( a35286a  and  a35281a );
 a35291a <=( A236  and  (not A233) );
 a35292a <=( A232  and  a35291a );
 a35295a <=( A299  and  A298 );
 a35298a <=( (not A301)  and  (not A300) );
 a35299a <=( a35298a  and  a35295a );
 a35300a <=( a35299a  and  a35292a );
 a35304a <=( (not A166)  and  (not A167) );
 a35305a <=( (not A169)  and  a35304a );
 a35309a <=( A203  and  A200 );
 a35310a <=( (not A199)  and  a35309a );
 a35311a <=( a35310a  and  a35305a );
 a35315a <=( (not A235)  and  (not A233) );
 a35316a <=( (not A232)  and  a35315a );
 a35319a <=( (not A268)  and  (not A267) );
 a35322a <=( A301  and  (not A269) );
 a35323a <=( a35322a  and  a35319a );
 a35324a <=( a35323a  and  a35316a );
 a35328a <=( (not A166)  and  (not A167) );
 a35329a <=( (not A169)  and  a35328a );
 a35333a <=( A203  and  A200 );
 a35334a <=( (not A199)  and  a35333a );
 a35335a <=( a35334a  and  a35329a );
 a35339a <=( (not A235)  and  (not A233) );
 a35340a <=( (not A232)  and  a35339a );
 a35343a <=( (not A266)  and  (not A265) );
 a35346a <=( A301  and  (not A268) );
 a35347a <=( a35346a  and  a35343a );
 a35348a <=( a35347a  and  a35340a );
 a35352a <=( (not A166)  and  (not A167) );
 a35353a <=( (not A169)  and  a35352a );
 a35357a <=( A203  and  (not A200) );
 a35358a <=( A199  and  a35357a );
 a35359a <=( a35358a  and  a35353a );
 a35363a <=( (not A236)  and  (not A235) );
 a35364a <=( (not A234)  and  a35363a );
 a35367a <=( (not A268)  and  (not A267) );
 a35370a <=( A301  and  (not A269) );
 a35371a <=( a35370a  and  a35367a );
 a35372a <=( a35371a  and  a35364a );
 a35376a <=( (not A166)  and  (not A167) );
 a35377a <=( (not A169)  and  a35376a );
 a35381a <=( A203  and  (not A200) );
 a35382a <=( A199  and  a35381a );
 a35383a <=( a35382a  and  a35377a );
 a35387a <=( (not A236)  and  (not A235) );
 a35388a <=( (not A234)  and  a35387a );
 a35391a <=( (not A266)  and  (not A265) );
 a35394a <=( A301  and  (not A268) );
 a35395a <=( a35394a  and  a35391a );
 a35396a <=( a35395a  and  a35388a );
 a35400a <=( (not A166)  and  (not A167) );
 a35401a <=( (not A169)  and  a35400a );
 a35405a <=( A203  and  (not A200) );
 a35406a <=( A199  and  a35405a );
 a35407a <=( a35406a  and  a35401a );
 a35411a <=( A236  and  A233 );
 a35412a <=( (not A232)  and  a35411a );
 a35415a <=( A299  and  A298 );
 a35418a <=( (not A301)  and  (not A300) );
 a35419a <=( a35418a  and  a35415a );
 a35420a <=( a35419a  and  a35412a );
 a35424a <=( (not A166)  and  (not A167) );
 a35425a <=( (not A169)  and  a35424a );
 a35429a <=( A203  and  (not A200) );
 a35430a <=( A199  and  a35429a );
 a35431a <=( a35430a  and  a35425a );
 a35435a <=( A236  and  (not A233) );
 a35436a <=( A232  and  a35435a );
 a35439a <=( A299  and  A298 );
 a35442a <=( (not A301)  and  (not A300) );
 a35443a <=( a35442a  and  a35439a );
 a35444a <=( a35443a  and  a35436a );
 a35448a <=( (not A166)  and  (not A167) );
 a35449a <=( (not A169)  and  a35448a );
 a35453a <=( A203  and  (not A200) );
 a35454a <=( A199  and  a35453a );
 a35455a <=( a35454a  and  a35449a );
 a35459a <=( (not A235)  and  (not A233) );
 a35460a <=( (not A232)  and  a35459a );
 a35463a <=( (not A268)  and  (not A267) );
 a35466a <=( A301  and  (not A269) );
 a35467a <=( a35466a  and  a35463a );
 a35468a <=( a35467a  and  a35460a );
 a35472a <=( (not A166)  and  (not A167) );
 a35473a <=( (not A169)  and  a35472a );
 a35477a <=( A203  and  (not A200) );
 a35478a <=( A199  and  a35477a );
 a35479a <=( a35478a  and  a35473a );
 a35483a <=( (not A235)  and  (not A233) );
 a35484a <=( (not A232)  and  a35483a );
 a35487a <=( (not A266)  and  (not A265) );
 a35490a <=( A301  and  (not A268) );
 a35491a <=( a35490a  and  a35487a );
 a35492a <=( a35491a  and  a35484a );
 a35496a <=( A167  and  (not A168) );
 a35497a <=( (not A169)  and  a35496a );
 a35501a <=( (not A234)  and  A202 );
 a35502a <=( A166  and  a35501a );
 a35503a <=( a35502a  and  a35497a );
 a35507a <=( (not A267)  and  (not A236) );
 a35508a <=( (not A235)  and  a35507a );
 a35511a <=( (not A269)  and  (not A268) );
 a35514a <=( A300  and  A299 );
 a35515a <=( a35514a  and  a35511a );
 a35516a <=( a35515a  and  a35508a );
 a35520a <=( A167  and  (not A168) );
 a35521a <=( (not A169)  and  a35520a );
 a35525a <=( (not A234)  and  A202 );
 a35526a <=( A166  and  a35525a );
 a35527a <=( a35526a  and  a35521a );
 a35531a <=( (not A267)  and  (not A236) );
 a35532a <=( (not A235)  and  a35531a );
 a35535a <=( (not A269)  and  (not A268) );
 a35538a <=( A300  and  A298 );
 a35539a <=( a35538a  and  a35535a );
 a35540a <=( a35539a  and  a35532a );
 a35544a <=( A167  and  (not A168) );
 a35545a <=( (not A169)  and  a35544a );
 a35549a <=( (not A234)  and  A202 );
 a35550a <=( A166  and  a35549a );
 a35551a <=( a35550a  and  a35545a );
 a35555a <=( A265  and  (not A236) );
 a35556a <=( (not A235)  and  a35555a );
 a35559a <=( (not A267)  and  A266 );
 a35562a <=( A301  and  (not A268) );
 a35563a <=( a35562a  and  a35559a );
 a35564a <=( a35563a  and  a35556a );
 a35568a <=( A167  and  (not A168) );
 a35569a <=( (not A169)  and  a35568a );
 a35573a <=( (not A234)  and  A202 );
 a35574a <=( A166  and  a35573a );
 a35575a <=( a35574a  and  a35569a );
 a35579a <=( (not A265)  and  (not A236) );
 a35580a <=( (not A235)  and  a35579a );
 a35583a <=( (not A268)  and  (not A266) );
 a35586a <=( A300  and  A299 );
 a35587a <=( a35586a  and  a35583a );
 a35588a <=( a35587a  and  a35580a );
 a35592a <=( A167  and  (not A168) );
 a35593a <=( (not A169)  and  a35592a );
 a35597a <=( (not A234)  and  A202 );
 a35598a <=( A166  and  a35597a );
 a35599a <=( a35598a  and  a35593a );
 a35603a <=( (not A265)  and  (not A236) );
 a35604a <=( (not A235)  and  a35603a );
 a35607a <=( (not A268)  and  (not A266) );
 a35610a <=( A300  and  A298 );
 a35611a <=( a35610a  and  a35607a );
 a35612a <=( a35611a  and  a35604a );
 a35616a <=( A167  and  (not A168) );
 a35617a <=( (not A169)  and  a35616a );
 a35621a <=( A232  and  A202 );
 a35622a <=( A166  and  a35621a );
 a35623a <=( a35622a  and  a35617a );
 a35627a <=( (not A235)  and  (not A234) );
 a35628a <=( A233  and  a35627a );
 a35631a <=( (not A268)  and  (not A267) );
 a35634a <=( A301  and  (not A269) );
 a35635a <=( a35634a  and  a35631a );
 a35636a <=( a35635a  and  a35628a );
 a35640a <=( A167  and  (not A168) );
 a35641a <=( (not A169)  and  a35640a );
 a35645a <=( A232  and  A202 );
 a35646a <=( A166  and  a35645a );
 a35647a <=( a35646a  and  a35641a );
 a35651a <=( (not A235)  and  (not A234) );
 a35652a <=( A233  and  a35651a );
 a35655a <=( (not A266)  and  (not A265) );
 a35658a <=( A301  and  (not A268) );
 a35659a <=( a35658a  and  a35655a );
 a35660a <=( a35659a  and  a35652a );
 a35664a <=( A167  and  (not A168) );
 a35665a <=( (not A169)  and  a35664a );
 a35669a <=( (not A232)  and  A202 );
 a35670a <=( A166  and  a35669a );
 a35671a <=( a35670a  and  a35665a );
 a35675a <=( (not A267)  and  (not A235) );
 a35676a <=( (not A233)  and  a35675a );
 a35679a <=( (not A269)  and  (not A268) );
 a35682a <=( A300  and  A299 );
 a35683a <=( a35682a  and  a35679a );
 a35684a <=( a35683a  and  a35676a );
 a35688a <=( A167  and  (not A168) );
 a35689a <=( (not A169)  and  a35688a );
 a35693a <=( (not A232)  and  A202 );
 a35694a <=( A166  and  a35693a );
 a35695a <=( a35694a  and  a35689a );
 a35699a <=( (not A267)  and  (not A235) );
 a35700a <=( (not A233)  and  a35699a );
 a35703a <=( (not A269)  and  (not A268) );
 a35706a <=( A300  and  A298 );
 a35707a <=( a35706a  and  a35703a );
 a35708a <=( a35707a  and  a35700a );
 a35712a <=( A167  and  (not A168) );
 a35713a <=( (not A169)  and  a35712a );
 a35717a <=( (not A232)  and  A202 );
 a35718a <=( A166  and  a35717a );
 a35719a <=( a35718a  and  a35713a );
 a35723a <=( A265  and  (not A235) );
 a35724a <=( (not A233)  and  a35723a );
 a35727a <=( (not A267)  and  A266 );
 a35730a <=( A301  and  (not A268) );
 a35731a <=( a35730a  and  a35727a );
 a35732a <=( a35731a  and  a35724a );
 a35736a <=( A167  and  (not A168) );
 a35737a <=( (not A169)  and  a35736a );
 a35741a <=( (not A232)  and  A202 );
 a35742a <=( A166  and  a35741a );
 a35743a <=( a35742a  and  a35737a );
 a35747a <=( (not A265)  and  (not A235) );
 a35748a <=( (not A233)  and  a35747a );
 a35751a <=( (not A268)  and  (not A266) );
 a35754a <=( A300  and  A299 );
 a35755a <=( a35754a  and  a35751a );
 a35756a <=( a35755a  and  a35748a );
 a35760a <=( A167  and  (not A168) );
 a35761a <=( (not A169)  and  a35760a );
 a35765a <=( (not A232)  and  A202 );
 a35766a <=( A166  and  a35765a );
 a35767a <=( a35766a  and  a35761a );
 a35771a <=( (not A265)  and  (not A235) );
 a35772a <=( (not A233)  and  a35771a );
 a35775a <=( (not A268)  and  (not A266) );
 a35778a <=( A300  and  A298 );
 a35779a <=( a35778a  and  a35775a );
 a35780a <=( a35779a  and  a35772a );
 a35784a <=( A167  and  (not A168) );
 a35785a <=( (not A169)  and  a35784a );
 a35789a <=( A201  and  A199 );
 a35790a <=( A166  and  a35789a );
 a35791a <=( a35790a  and  a35785a );
 a35795a <=( (not A236)  and  (not A235) );
 a35796a <=( (not A234)  and  a35795a );
 a35799a <=( (not A268)  and  (not A267) );
 a35802a <=( A301  and  (not A269) );
 a35803a <=( a35802a  and  a35799a );
 a35804a <=( a35803a  and  a35796a );
 a35808a <=( A167  and  (not A168) );
 a35809a <=( (not A169)  and  a35808a );
 a35813a <=( A201  and  A199 );
 a35814a <=( A166  and  a35813a );
 a35815a <=( a35814a  and  a35809a );
 a35819a <=( (not A236)  and  (not A235) );
 a35820a <=( (not A234)  and  a35819a );
 a35823a <=( (not A266)  and  (not A265) );
 a35826a <=( A301  and  (not A268) );
 a35827a <=( a35826a  and  a35823a );
 a35828a <=( a35827a  and  a35820a );
 a35832a <=( A167  and  (not A168) );
 a35833a <=( (not A169)  and  a35832a );
 a35837a <=( A201  and  A199 );
 a35838a <=( A166  and  a35837a );
 a35839a <=( a35838a  and  a35833a );
 a35843a <=( A236  and  A233 );
 a35844a <=( (not A232)  and  a35843a );
 a35847a <=( A299  and  A298 );
 a35850a <=( (not A301)  and  (not A300) );
 a35851a <=( a35850a  and  a35847a );
 a35852a <=( a35851a  and  a35844a );
 a35856a <=( A167  and  (not A168) );
 a35857a <=( (not A169)  and  a35856a );
 a35861a <=( A201  and  A199 );
 a35862a <=( A166  and  a35861a );
 a35863a <=( a35862a  and  a35857a );
 a35867a <=( A236  and  (not A233) );
 a35868a <=( A232  and  a35867a );
 a35871a <=( A299  and  A298 );
 a35874a <=( (not A301)  and  (not A300) );
 a35875a <=( a35874a  and  a35871a );
 a35876a <=( a35875a  and  a35868a );
 a35880a <=( A167  and  (not A168) );
 a35881a <=( (not A169)  and  a35880a );
 a35885a <=( A201  and  A199 );
 a35886a <=( A166  and  a35885a );
 a35887a <=( a35886a  and  a35881a );
 a35891a <=( (not A235)  and  (not A233) );
 a35892a <=( (not A232)  and  a35891a );
 a35895a <=( (not A268)  and  (not A267) );
 a35898a <=( A301  and  (not A269) );
 a35899a <=( a35898a  and  a35895a );
 a35900a <=( a35899a  and  a35892a );
 a35904a <=( A167  and  (not A168) );
 a35905a <=( (not A169)  and  a35904a );
 a35909a <=( A201  and  A199 );
 a35910a <=( A166  and  a35909a );
 a35911a <=( a35910a  and  a35905a );
 a35915a <=( (not A235)  and  (not A233) );
 a35916a <=( (not A232)  and  a35915a );
 a35919a <=( (not A266)  and  (not A265) );
 a35922a <=( A301  and  (not A268) );
 a35923a <=( a35922a  and  a35919a );
 a35924a <=( a35923a  and  a35916a );
 a35928a <=( A167  and  (not A168) );
 a35929a <=( (not A169)  and  a35928a );
 a35933a <=( A201  and  A200 );
 a35934a <=( A166  and  a35933a );
 a35935a <=( a35934a  and  a35929a );
 a35939a <=( (not A236)  and  (not A235) );
 a35940a <=( (not A234)  and  a35939a );
 a35943a <=( (not A268)  and  (not A267) );
 a35946a <=( A301  and  (not A269) );
 a35947a <=( a35946a  and  a35943a );
 a35948a <=( a35947a  and  a35940a );
 a35952a <=( A167  and  (not A168) );
 a35953a <=( (not A169)  and  a35952a );
 a35957a <=( A201  and  A200 );
 a35958a <=( A166  and  a35957a );
 a35959a <=( a35958a  and  a35953a );
 a35963a <=( (not A236)  and  (not A235) );
 a35964a <=( (not A234)  and  a35963a );
 a35967a <=( (not A266)  and  (not A265) );
 a35970a <=( A301  and  (not A268) );
 a35971a <=( a35970a  and  a35967a );
 a35972a <=( a35971a  and  a35964a );
 a35976a <=( A167  and  (not A168) );
 a35977a <=( (not A169)  and  a35976a );
 a35981a <=( A201  and  A200 );
 a35982a <=( A166  and  a35981a );
 a35983a <=( a35982a  and  a35977a );
 a35987a <=( A236  and  A233 );
 a35988a <=( (not A232)  and  a35987a );
 a35991a <=( A299  and  A298 );
 a35994a <=( (not A301)  and  (not A300) );
 a35995a <=( a35994a  and  a35991a );
 a35996a <=( a35995a  and  a35988a );
 a36000a <=( A167  and  (not A168) );
 a36001a <=( (not A169)  and  a36000a );
 a36005a <=( A201  and  A200 );
 a36006a <=( A166  and  a36005a );
 a36007a <=( a36006a  and  a36001a );
 a36011a <=( A236  and  (not A233) );
 a36012a <=( A232  and  a36011a );
 a36015a <=( A299  and  A298 );
 a36018a <=( (not A301)  and  (not A300) );
 a36019a <=( a36018a  and  a36015a );
 a36020a <=( a36019a  and  a36012a );
 a36024a <=( A167  and  (not A168) );
 a36025a <=( (not A169)  and  a36024a );
 a36029a <=( A201  and  A200 );
 a36030a <=( A166  and  a36029a );
 a36031a <=( a36030a  and  a36025a );
 a36035a <=( (not A235)  and  (not A233) );
 a36036a <=( (not A232)  and  a36035a );
 a36039a <=( (not A268)  and  (not A267) );
 a36042a <=( A301  and  (not A269) );
 a36043a <=( a36042a  and  a36039a );
 a36044a <=( a36043a  and  a36036a );
 a36048a <=( A167  and  (not A168) );
 a36049a <=( (not A169)  and  a36048a );
 a36053a <=( A201  and  A200 );
 a36054a <=( A166  and  a36053a );
 a36055a <=( a36054a  and  a36049a );
 a36059a <=( (not A235)  and  (not A233) );
 a36060a <=( (not A232)  and  a36059a );
 a36063a <=( (not A266)  and  (not A265) );
 a36066a <=( A301  and  (not A268) );
 a36067a <=( a36066a  and  a36063a );
 a36068a <=( a36067a  and  a36060a );
 a36072a <=( A167  and  (not A168) );
 a36073a <=( (not A169)  and  a36072a );
 a36077a <=( A200  and  (not A199) );
 a36078a <=( A166  and  a36077a );
 a36079a <=( a36078a  and  a36073a );
 a36083a <=( A234  and  A232 );
 a36084a <=( A203  and  a36083a );
 a36087a <=( A299  and  A298 );
 a36090a <=( (not A301)  and  (not A300) );
 a36091a <=( a36090a  and  a36087a );
 a36092a <=( a36091a  and  a36084a );
 a36096a <=( A167  and  (not A168) );
 a36097a <=( (not A169)  and  a36096a );
 a36101a <=( A200  and  (not A199) );
 a36102a <=( A166  and  a36101a );
 a36103a <=( a36102a  and  a36097a );
 a36107a <=( A234  and  A233 );
 a36108a <=( A203  and  a36107a );
 a36111a <=( A299  and  A298 );
 a36114a <=( (not A301)  and  (not A300) );
 a36115a <=( a36114a  and  a36111a );
 a36116a <=( a36115a  and  a36108a );
 a36120a <=( A167  and  (not A168) );
 a36121a <=( (not A169)  and  a36120a );
 a36125a <=( A200  and  (not A199) );
 a36126a <=( A166  and  a36125a );
 a36127a <=( a36126a  and  a36121a );
 a36131a <=( A233  and  (not A232) );
 a36132a <=( A203  and  a36131a );
 a36135a <=( (not A300)  and  A236 );
 a36138a <=( (not A302)  and  (not A301) );
 a36139a <=( a36138a  and  a36135a );
 a36140a <=( a36139a  and  a36132a );
 a36144a <=( A167  and  (not A168) );
 a36145a <=( (not A169)  and  a36144a );
 a36149a <=( A200  and  (not A199) );
 a36150a <=( A166  and  a36149a );
 a36151a <=( a36150a  and  a36145a );
 a36155a <=( A233  and  (not A232) );
 a36156a <=( A203  and  a36155a );
 a36159a <=( (not A298)  and  A236 );
 a36162a <=( (not A301)  and  (not A299) );
 a36163a <=( a36162a  and  a36159a );
 a36164a <=( a36163a  and  a36156a );
 a36168a <=( A167  and  (not A168) );
 a36169a <=( (not A169)  and  a36168a );
 a36173a <=( A200  and  (not A199) );
 a36174a <=( A166  and  a36173a );
 a36175a <=( a36174a  and  a36169a );
 a36179a <=( A233  and  (not A232) );
 a36180a <=( A203  and  a36179a );
 a36183a <=( (not A265)  and  A236 );
 a36186a <=( A269  and  A266 );
 a36187a <=( a36186a  and  a36183a );
 a36188a <=( a36187a  and  a36180a );
 a36192a <=( A167  and  (not A168) );
 a36193a <=( (not A169)  and  a36192a );
 a36197a <=( A200  and  (not A199) );
 a36198a <=( A166  and  a36197a );
 a36199a <=( a36198a  and  a36193a );
 a36203a <=( A233  and  (not A232) );
 a36204a <=( A203  and  a36203a );
 a36207a <=( A265  and  A236 );
 a36210a <=( A269  and  (not A266) );
 a36211a <=( a36210a  and  a36207a );
 a36212a <=( a36211a  and  a36204a );
 a36216a <=( A167  and  (not A168) );
 a36217a <=( (not A169)  and  a36216a );
 a36221a <=( A200  and  (not A199) );
 a36222a <=( A166  and  a36221a );
 a36223a <=( a36222a  and  a36217a );
 a36227a <=( (not A233)  and  A232 );
 a36228a <=( A203  and  a36227a );
 a36231a <=( (not A300)  and  A236 );
 a36234a <=( (not A302)  and  (not A301) );
 a36235a <=( a36234a  and  a36231a );
 a36236a <=( a36235a  and  a36228a );
 a36240a <=( A167  and  (not A168) );
 a36241a <=( (not A169)  and  a36240a );
 a36245a <=( A200  and  (not A199) );
 a36246a <=( A166  and  a36245a );
 a36247a <=( a36246a  and  a36241a );
 a36251a <=( (not A233)  and  A232 );
 a36252a <=( A203  and  a36251a );
 a36255a <=( (not A298)  and  A236 );
 a36258a <=( (not A301)  and  (not A299) );
 a36259a <=( a36258a  and  a36255a );
 a36260a <=( a36259a  and  a36252a );
 a36264a <=( A167  and  (not A168) );
 a36265a <=( (not A169)  and  a36264a );
 a36269a <=( A200  and  (not A199) );
 a36270a <=( A166  and  a36269a );
 a36271a <=( a36270a  and  a36265a );
 a36275a <=( (not A233)  and  A232 );
 a36276a <=( A203  and  a36275a );
 a36279a <=( (not A265)  and  A236 );
 a36282a <=( A269  and  A266 );
 a36283a <=( a36282a  and  a36279a );
 a36284a <=( a36283a  and  a36276a );
 a36288a <=( A167  and  (not A168) );
 a36289a <=( (not A169)  and  a36288a );
 a36293a <=( A200  and  (not A199) );
 a36294a <=( A166  and  a36293a );
 a36295a <=( a36294a  and  a36289a );
 a36299a <=( (not A233)  and  A232 );
 a36300a <=( A203  and  a36299a );
 a36303a <=( A265  and  A236 );
 a36306a <=( A269  and  (not A266) );
 a36307a <=( a36306a  and  a36303a );
 a36308a <=( a36307a  and  a36300a );
 a36312a <=( A167  and  (not A168) );
 a36313a <=( (not A169)  and  a36312a );
 a36317a <=( (not A200)  and  A199 );
 a36318a <=( A166  and  a36317a );
 a36319a <=( a36318a  and  a36313a );
 a36323a <=( A234  and  A232 );
 a36324a <=( A203  and  a36323a );
 a36327a <=( A299  and  A298 );
 a36330a <=( (not A301)  and  (not A300) );
 a36331a <=( a36330a  and  a36327a );
 a36332a <=( a36331a  and  a36324a );
 a36336a <=( A167  and  (not A168) );
 a36337a <=( (not A169)  and  a36336a );
 a36341a <=( (not A200)  and  A199 );
 a36342a <=( A166  and  a36341a );
 a36343a <=( a36342a  and  a36337a );
 a36347a <=( A234  and  A233 );
 a36348a <=( A203  and  a36347a );
 a36351a <=( A299  and  A298 );
 a36354a <=( (not A301)  and  (not A300) );
 a36355a <=( a36354a  and  a36351a );
 a36356a <=( a36355a  and  a36348a );
 a36360a <=( A167  and  (not A168) );
 a36361a <=( (not A169)  and  a36360a );
 a36365a <=( (not A200)  and  A199 );
 a36366a <=( A166  and  a36365a );
 a36367a <=( a36366a  and  a36361a );
 a36371a <=( A233  and  (not A232) );
 a36372a <=( A203  and  a36371a );
 a36375a <=( (not A300)  and  A236 );
 a36378a <=( (not A302)  and  (not A301) );
 a36379a <=( a36378a  and  a36375a );
 a36380a <=( a36379a  and  a36372a );
 a36384a <=( A167  and  (not A168) );
 a36385a <=( (not A169)  and  a36384a );
 a36389a <=( (not A200)  and  A199 );
 a36390a <=( A166  and  a36389a );
 a36391a <=( a36390a  and  a36385a );
 a36395a <=( A233  and  (not A232) );
 a36396a <=( A203  and  a36395a );
 a36399a <=( (not A298)  and  A236 );
 a36402a <=( (not A301)  and  (not A299) );
 a36403a <=( a36402a  and  a36399a );
 a36404a <=( a36403a  and  a36396a );
 a36408a <=( A167  and  (not A168) );
 a36409a <=( (not A169)  and  a36408a );
 a36413a <=( (not A200)  and  A199 );
 a36414a <=( A166  and  a36413a );
 a36415a <=( a36414a  and  a36409a );
 a36419a <=( A233  and  (not A232) );
 a36420a <=( A203  and  a36419a );
 a36423a <=( (not A265)  and  A236 );
 a36426a <=( A269  and  A266 );
 a36427a <=( a36426a  and  a36423a );
 a36428a <=( a36427a  and  a36420a );
 a36432a <=( A167  and  (not A168) );
 a36433a <=( (not A169)  and  a36432a );
 a36437a <=( (not A200)  and  A199 );
 a36438a <=( A166  and  a36437a );
 a36439a <=( a36438a  and  a36433a );
 a36443a <=( A233  and  (not A232) );
 a36444a <=( A203  and  a36443a );
 a36447a <=( A265  and  A236 );
 a36450a <=( A269  and  (not A266) );
 a36451a <=( a36450a  and  a36447a );
 a36452a <=( a36451a  and  a36444a );
 a36456a <=( A167  and  (not A168) );
 a36457a <=( (not A169)  and  a36456a );
 a36461a <=( (not A200)  and  A199 );
 a36462a <=( A166  and  a36461a );
 a36463a <=( a36462a  and  a36457a );
 a36467a <=( (not A233)  and  A232 );
 a36468a <=( A203  and  a36467a );
 a36471a <=( (not A300)  and  A236 );
 a36474a <=( (not A302)  and  (not A301) );
 a36475a <=( a36474a  and  a36471a );
 a36476a <=( a36475a  and  a36468a );
 a36480a <=( A167  and  (not A168) );
 a36481a <=( (not A169)  and  a36480a );
 a36485a <=( (not A200)  and  A199 );
 a36486a <=( A166  and  a36485a );
 a36487a <=( a36486a  and  a36481a );
 a36491a <=( (not A233)  and  A232 );
 a36492a <=( A203  and  a36491a );
 a36495a <=( (not A298)  and  A236 );
 a36498a <=( (not A301)  and  (not A299) );
 a36499a <=( a36498a  and  a36495a );
 a36500a <=( a36499a  and  a36492a );
 a36504a <=( A167  and  (not A168) );
 a36505a <=( (not A169)  and  a36504a );
 a36509a <=( (not A200)  and  A199 );
 a36510a <=( A166  and  a36509a );
 a36511a <=( a36510a  and  a36505a );
 a36515a <=( (not A233)  and  A232 );
 a36516a <=( A203  and  a36515a );
 a36519a <=( (not A265)  and  A236 );
 a36522a <=( A269  and  A266 );
 a36523a <=( a36522a  and  a36519a );
 a36524a <=( a36523a  and  a36516a );
 a36528a <=( A167  and  (not A168) );
 a36529a <=( (not A169)  and  a36528a );
 a36533a <=( (not A200)  and  A199 );
 a36534a <=( A166  and  a36533a );
 a36535a <=( a36534a  and  a36529a );
 a36539a <=( (not A233)  and  A232 );
 a36540a <=( A203  and  a36539a );
 a36543a <=( A265  and  A236 );
 a36546a <=( A269  and  (not A266) );
 a36547a <=( a36546a  and  a36543a );
 a36548a <=( a36547a  and  a36540a );
 a36552a <=( (not A168)  and  (not A169) );
 a36553a <=( (not A170)  and  a36552a );
 a36557a <=( (not A235)  and  (not A234) );
 a36558a <=( A202  and  a36557a );
 a36559a <=( a36558a  and  a36553a );
 a36563a <=( (not A268)  and  (not A267) );
 a36564a <=( (not A236)  and  a36563a );
 a36567a <=( A298  and  (not A269) );
 a36570a <=( A302  and  (not A299) );
 a36571a <=( a36570a  and  a36567a );
 a36572a <=( a36571a  and  a36564a );
 a36576a <=( (not A168)  and  (not A169) );
 a36577a <=( (not A170)  and  a36576a );
 a36581a <=( (not A235)  and  (not A234) );
 a36582a <=( A202  and  a36581a );
 a36583a <=( a36582a  and  a36577a );
 a36587a <=( (not A268)  and  (not A267) );
 a36588a <=( (not A236)  and  a36587a );
 a36591a <=( (not A298)  and  (not A269) );
 a36594a <=( A302  and  A299 );
 a36595a <=( a36594a  and  a36591a );
 a36596a <=( a36595a  and  a36588a );
 a36600a <=( (not A168)  and  (not A169) );
 a36601a <=( (not A170)  and  a36600a );
 a36605a <=( (not A235)  and  (not A234) );
 a36606a <=( A202  and  a36605a );
 a36607a <=( a36606a  and  a36601a );
 a36611a <=( A266  and  A265 );
 a36612a <=( (not A236)  and  a36611a );
 a36615a <=( (not A268)  and  (not A267) );
 a36618a <=( A300  and  A299 );
 a36619a <=( a36618a  and  a36615a );
 a36620a <=( a36619a  and  a36612a );
 a36624a <=( (not A168)  and  (not A169) );
 a36625a <=( (not A170)  and  a36624a );
 a36629a <=( (not A235)  and  (not A234) );
 a36630a <=( A202  and  a36629a );
 a36631a <=( a36630a  and  a36625a );
 a36635a <=( A266  and  A265 );
 a36636a <=( (not A236)  and  a36635a );
 a36639a <=( (not A268)  and  (not A267) );
 a36642a <=( A300  and  A298 );
 a36643a <=( a36642a  and  a36639a );
 a36644a <=( a36643a  and  a36636a );
 a36648a <=( (not A168)  and  (not A169) );
 a36649a <=( (not A170)  and  a36648a );
 a36653a <=( (not A235)  and  (not A234) );
 a36654a <=( A202  and  a36653a );
 a36655a <=( a36654a  and  a36649a );
 a36659a <=( (not A266)  and  (not A265) );
 a36660a <=( (not A236)  and  a36659a );
 a36663a <=( A298  and  (not A268) );
 a36666a <=( A302  and  (not A299) );
 a36667a <=( a36666a  and  a36663a );
 a36668a <=( a36667a  and  a36660a );
 a36672a <=( (not A168)  and  (not A169) );
 a36673a <=( (not A170)  and  a36672a );
 a36677a <=( (not A235)  and  (not A234) );
 a36678a <=( A202  and  a36677a );
 a36679a <=( a36678a  and  a36673a );
 a36683a <=( (not A266)  and  (not A265) );
 a36684a <=( (not A236)  and  a36683a );
 a36687a <=( (not A298)  and  (not A268) );
 a36690a <=( A302  and  A299 );
 a36691a <=( a36690a  and  a36687a );
 a36692a <=( a36691a  and  a36684a );
 a36696a <=( (not A168)  and  (not A169) );
 a36697a <=( (not A170)  and  a36696a );
 a36701a <=( A233  and  A232 );
 a36702a <=( A202  and  a36701a );
 a36703a <=( a36702a  and  a36697a );
 a36707a <=( (not A267)  and  (not A235) );
 a36708a <=( (not A234)  and  a36707a );
 a36711a <=( (not A269)  and  (not A268) );
 a36714a <=( A300  and  A299 );
 a36715a <=( a36714a  and  a36711a );
 a36716a <=( a36715a  and  a36708a );
 a36720a <=( (not A168)  and  (not A169) );
 a36721a <=( (not A170)  and  a36720a );
 a36725a <=( A233  and  A232 );
 a36726a <=( A202  and  a36725a );
 a36727a <=( a36726a  and  a36721a );
 a36731a <=( (not A267)  and  (not A235) );
 a36732a <=( (not A234)  and  a36731a );
 a36735a <=( (not A269)  and  (not A268) );
 a36738a <=( A300  and  A298 );
 a36739a <=( a36738a  and  a36735a );
 a36740a <=( a36739a  and  a36732a );
 a36744a <=( (not A168)  and  (not A169) );
 a36745a <=( (not A170)  and  a36744a );
 a36749a <=( A233  and  A232 );
 a36750a <=( A202  and  a36749a );
 a36751a <=( a36750a  and  a36745a );
 a36755a <=( A265  and  (not A235) );
 a36756a <=( (not A234)  and  a36755a );
 a36759a <=( (not A267)  and  A266 );
 a36762a <=( A301  and  (not A268) );
 a36763a <=( a36762a  and  a36759a );
 a36764a <=( a36763a  and  a36756a );
 a36768a <=( (not A168)  and  (not A169) );
 a36769a <=( (not A170)  and  a36768a );
 a36773a <=( A233  and  A232 );
 a36774a <=( A202  and  a36773a );
 a36775a <=( a36774a  and  a36769a );
 a36779a <=( (not A265)  and  (not A235) );
 a36780a <=( (not A234)  and  a36779a );
 a36783a <=( (not A268)  and  (not A266) );
 a36786a <=( A300  and  A299 );
 a36787a <=( a36786a  and  a36783a );
 a36788a <=( a36787a  and  a36780a );
 a36792a <=( (not A168)  and  (not A169) );
 a36793a <=( (not A170)  and  a36792a );
 a36797a <=( A233  and  A232 );
 a36798a <=( A202  and  a36797a );
 a36799a <=( a36798a  and  a36793a );
 a36803a <=( (not A265)  and  (not A235) );
 a36804a <=( (not A234)  and  a36803a );
 a36807a <=( (not A268)  and  (not A266) );
 a36810a <=( A300  and  A298 );
 a36811a <=( a36810a  and  a36807a );
 a36812a <=( a36811a  and  a36804a );
 a36816a <=( (not A168)  and  (not A169) );
 a36817a <=( (not A170)  and  a36816a );
 a36821a <=( (not A233)  and  (not A232) );
 a36822a <=( A202  and  a36821a );
 a36823a <=( a36822a  and  a36817a );
 a36827a <=( (not A268)  and  (not A267) );
 a36828a <=( (not A235)  and  a36827a );
 a36831a <=( A298  and  (not A269) );
 a36834a <=( A302  and  (not A299) );
 a36835a <=( a36834a  and  a36831a );
 a36836a <=( a36835a  and  a36828a );
 a36840a <=( (not A168)  and  (not A169) );
 a36841a <=( (not A170)  and  a36840a );
 a36845a <=( (not A233)  and  (not A232) );
 a36846a <=( A202  and  a36845a );
 a36847a <=( a36846a  and  a36841a );
 a36851a <=( (not A268)  and  (not A267) );
 a36852a <=( (not A235)  and  a36851a );
 a36855a <=( (not A298)  and  (not A269) );
 a36858a <=( A302  and  A299 );
 a36859a <=( a36858a  and  a36855a );
 a36860a <=( a36859a  and  a36852a );
 a36864a <=( (not A168)  and  (not A169) );
 a36865a <=( (not A170)  and  a36864a );
 a36869a <=( (not A233)  and  (not A232) );
 a36870a <=( A202  and  a36869a );
 a36871a <=( a36870a  and  a36865a );
 a36875a <=( A266  and  A265 );
 a36876a <=( (not A235)  and  a36875a );
 a36879a <=( (not A268)  and  (not A267) );
 a36882a <=( A300  and  A299 );
 a36883a <=( a36882a  and  a36879a );
 a36884a <=( a36883a  and  a36876a );
 a36888a <=( (not A168)  and  (not A169) );
 a36889a <=( (not A170)  and  a36888a );
 a36893a <=( (not A233)  and  (not A232) );
 a36894a <=( A202  and  a36893a );
 a36895a <=( a36894a  and  a36889a );
 a36899a <=( A266  and  A265 );
 a36900a <=( (not A235)  and  a36899a );
 a36903a <=( (not A268)  and  (not A267) );
 a36906a <=( A300  and  A298 );
 a36907a <=( a36906a  and  a36903a );
 a36908a <=( a36907a  and  a36900a );
 a36912a <=( (not A168)  and  (not A169) );
 a36913a <=( (not A170)  and  a36912a );
 a36917a <=( (not A233)  and  (not A232) );
 a36918a <=( A202  and  a36917a );
 a36919a <=( a36918a  and  a36913a );
 a36923a <=( (not A266)  and  (not A265) );
 a36924a <=( (not A235)  and  a36923a );
 a36927a <=( A298  and  (not A268) );
 a36930a <=( A302  and  (not A299) );
 a36931a <=( a36930a  and  a36927a );
 a36932a <=( a36931a  and  a36924a );
 a36936a <=( (not A168)  and  (not A169) );
 a36937a <=( (not A170)  and  a36936a );
 a36941a <=( (not A233)  and  (not A232) );
 a36942a <=( A202  and  a36941a );
 a36943a <=( a36942a  and  a36937a );
 a36947a <=( (not A266)  and  (not A265) );
 a36948a <=( (not A235)  and  a36947a );
 a36951a <=( (not A298)  and  (not A268) );
 a36954a <=( A302  and  A299 );
 a36955a <=( a36954a  and  a36951a );
 a36956a <=( a36955a  and  a36948a );
 a36960a <=( (not A168)  and  (not A169) );
 a36961a <=( (not A170)  and  a36960a );
 a36965a <=( (not A234)  and  A201 );
 a36966a <=( A199  and  a36965a );
 a36967a <=( a36966a  and  a36961a );
 a36971a <=( (not A267)  and  (not A236) );
 a36972a <=( (not A235)  and  a36971a );
 a36975a <=( (not A269)  and  (not A268) );
 a36978a <=( A300  and  A299 );
 a36979a <=( a36978a  and  a36975a );
 a36980a <=( a36979a  and  a36972a );
 a36984a <=( (not A168)  and  (not A169) );
 a36985a <=( (not A170)  and  a36984a );
 a36989a <=( (not A234)  and  A201 );
 a36990a <=( A199  and  a36989a );
 a36991a <=( a36990a  and  a36985a );
 a36995a <=( (not A267)  and  (not A236) );
 a36996a <=( (not A235)  and  a36995a );
 a36999a <=( (not A269)  and  (not A268) );
 a37002a <=( A300  and  A298 );
 a37003a <=( a37002a  and  a36999a );
 a37004a <=( a37003a  and  a36996a );
 a37008a <=( (not A168)  and  (not A169) );
 a37009a <=( (not A170)  and  a37008a );
 a37013a <=( (not A234)  and  A201 );
 a37014a <=( A199  and  a37013a );
 a37015a <=( a37014a  and  a37009a );
 a37019a <=( A265  and  (not A236) );
 a37020a <=( (not A235)  and  a37019a );
 a37023a <=( (not A267)  and  A266 );
 a37026a <=( A301  and  (not A268) );
 a37027a <=( a37026a  and  a37023a );
 a37028a <=( a37027a  and  a37020a );
 a37032a <=( (not A168)  and  (not A169) );
 a37033a <=( (not A170)  and  a37032a );
 a37037a <=( (not A234)  and  A201 );
 a37038a <=( A199  and  a37037a );
 a37039a <=( a37038a  and  a37033a );
 a37043a <=( (not A265)  and  (not A236) );
 a37044a <=( (not A235)  and  a37043a );
 a37047a <=( (not A268)  and  (not A266) );
 a37050a <=( A300  and  A299 );
 a37051a <=( a37050a  and  a37047a );
 a37052a <=( a37051a  and  a37044a );
 a37056a <=( (not A168)  and  (not A169) );
 a37057a <=( (not A170)  and  a37056a );
 a37061a <=( (not A234)  and  A201 );
 a37062a <=( A199  and  a37061a );
 a37063a <=( a37062a  and  a37057a );
 a37067a <=( (not A265)  and  (not A236) );
 a37068a <=( (not A235)  and  a37067a );
 a37071a <=( (not A268)  and  (not A266) );
 a37074a <=( A300  and  A298 );
 a37075a <=( a37074a  and  a37071a );
 a37076a <=( a37075a  and  a37068a );
 a37080a <=( (not A168)  and  (not A169) );
 a37081a <=( (not A170)  and  a37080a );
 a37085a <=( A232  and  A201 );
 a37086a <=( A199  and  a37085a );
 a37087a <=( a37086a  and  a37081a );
 a37091a <=( (not A235)  and  (not A234) );
 a37092a <=( A233  and  a37091a );
 a37095a <=( (not A268)  and  (not A267) );
 a37098a <=( A301  and  (not A269) );
 a37099a <=( a37098a  and  a37095a );
 a37100a <=( a37099a  and  a37092a );
 a37104a <=( (not A168)  and  (not A169) );
 a37105a <=( (not A170)  and  a37104a );
 a37109a <=( A232  and  A201 );
 a37110a <=( A199  and  a37109a );
 a37111a <=( a37110a  and  a37105a );
 a37115a <=( (not A235)  and  (not A234) );
 a37116a <=( A233  and  a37115a );
 a37119a <=( (not A266)  and  (not A265) );
 a37122a <=( A301  and  (not A268) );
 a37123a <=( a37122a  and  a37119a );
 a37124a <=( a37123a  and  a37116a );
 a37128a <=( (not A168)  and  (not A169) );
 a37129a <=( (not A170)  and  a37128a );
 a37133a <=( (not A232)  and  A201 );
 a37134a <=( A199  and  a37133a );
 a37135a <=( a37134a  and  a37129a );
 a37139a <=( (not A267)  and  (not A235) );
 a37140a <=( (not A233)  and  a37139a );
 a37143a <=( (not A269)  and  (not A268) );
 a37146a <=( A300  and  A299 );
 a37147a <=( a37146a  and  a37143a );
 a37148a <=( a37147a  and  a37140a );
 a37152a <=( (not A168)  and  (not A169) );
 a37153a <=( (not A170)  and  a37152a );
 a37157a <=( (not A232)  and  A201 );
 a37158a <=( A199  and  a37157a );
 a37159a <=( a37158a  and  a37153a );
 a37163a <=( (not A267)  and  (not A235) );
 a37164a <=( (not A233)  and  a37163a );
 a37167a <=( (not A269)  and  (not A268) );
 a37170a <=( A300  and  A298 );
 a37171a <=( a37170a  and  a37167a );
 a37172a <=( a37171a  and  a37164a );
 a37176a <=( (not A168)  and  (not A169) );
 a37177a <=( (not A170)  and  a37176a );
 a37181a <=( (not A232)  and  A201 );
 a37182a <=( A199  and  a37181a );
 a37183a <=( a37182a  and  a37177a );
 a37187a <=( A265  and  (not A235) );
 a37188a <=( (not A233)  and  a37187a );
 a37191a <=( (not A267)  and  A266 );
 a37194a <=( A301  and  (not A268) );
 a37195a <=( a37194a  and  a37191a );
 a37196a <=( a37195a  and  a37188a );
 a37200a <=( (not A168)  and  (not A169) );
 a37201a <=( (not A170)  and  a37200a );
 a37205a <=( (not A232)  and  A201 );
 a37206a <=( A199  and  a37205a );
 a37207a <=( a37206a  and  a37201a );
 a37211a <=( (not A265)  and  (not A235) );
 a37212a <=( (not A233)  and  a37211a );
 a37215a <=( (not A268)  and  (not A266) );
 a37218a <=( A300  and  A299 );
 a37219a <=( a37218a  and  a37215a );
 a37220a <=( a37219a  and  a37212a );
 a37224a <=( (not A168)  and  (not A169) );
 a37225a <=( (not A170)  and  a37224a );
 a37229a <=( (not A232)  and  A201 );
 a37230a <=( A199  and  a37229a );
 a37231a <=( a37230a  and  a37225a );
 a37235a <=( (not A265)  and  (not A235) );
 a37236a <=( (not A233)  and  a37235a );
 a37239a <=( (not A268)  and  (not A266) );
 a37242a <=( A300  and  A298 );
 a37243a <=( a37242a  and  a37239a );
 a37244a <=( a37243a  and  a37236a );
 a37248a <=( (not A168)  and  (not A169) );
 a37249a <=( (not A170)  and  a37248a );
 a37253a <=( (not A234)  and  A201 );
 a37254a <=( A200  and  a37253a );
 a37255a <=( a37254a  and  a37249a );
 a37259a <=( (not A267)  and  (not A236) );
 a37260a <=( (not A235)  and  a37259a );
 a37263a <=( (not A269)  and  (not A268) );
 a37266a <=( A300  and  A299 );
 a37267a <=( a37266a  and  a37263a );
 a37268a <=( a37267a  and  a37260a );
 a37272a <=( (not A168)  and  (not A169) );
 a37273a <=( (not A170)  and  a37272a );
 a37277a <=( (not A234)  and  A201 );
 a37278a <=( A200  and  a37277a );
 a37279a <=( a37278a  and  a37273a );
 a37283a <=( (not A267)  and  (not A236) );
 a37284a <=( (not A235)  and  a37283a );
 a37287a <=( (not A269)  and  (not A268) );
 a37290a <=( A300  and  A298 );
 a37291a <=( a37290a  and  a37287a );
 a37292a <=( a37291a  and  a37284a );
 a37296a <=( (not A168)  and  (not A169) );
 a37297a <=( (not A170)  and  a37296a );
 a37301a <=( (not A234)  and  A201 );
 a37302a <=( A200  and  a37301a );
 a37303a <=( a37302a  and  a37297a );
 a37307a <=( A265  and  (not A236) );
 a37308a <=( (not A235)  and  a37307a );
 a37311a <=( (not A267)  and  A266 );
 a37314a <=( A301  and  (not A268) );
 a37315a <=( a37314a  and  a37311a );
 a37316a <=( a37315a  and  a37308a );
 a37320a <=( (not A168)  and  (not A169) );
 a37321a <=( (not A170)  and  a37320a );
 a37325a <=( (not A234)  and  A201 );
 a37326a <=( A200  and  a37325a );
 a37327a <=( a37326a  and  a37321a );
 a37331a <=( (not A265)  and  (not A236) );
 a37332a <=( (not A235)  and  a37331a );
 a37335a <=( (not A268)  and  (not A266) );
 a37338a <=( A300  and  A299 );
 a37339a <=( a37338a  and  a37335a );
 a37340a <=( a37339a  and  a37332a );
 a37344a <=( (not A168)  and  (not A169) );
 a37345a <=( (not A170)  and  a37344a );
 a37349a <=( (not A234)  and  A201 );
 a37350a <=( A200  and  a37349a );
 a37351a <=( a37350a  and  a37345a );
 a37355a <=( (not A265)  and  (not A236) );
 a37356a <=( (not A235)  and  a37355a );
 a37359a <=( (not A268)  and  (not A266) );
 a37362a <=( A300  and  A298 );
 a37363a <=( a37362a  and  a37359a );
 a37364a <=( a37363a  and  a37356a );
 a37368a <=( (not A168)  and  (not A169) );
 a37369a <=( (not A170)  and  a37368a );
 a37373a <=( A232  and  A201 );
 a37374a <=( A200  and  a37373a );
 a37375a <=( a37374a  and  a37369a );
 a37379a <=( (not A235)  and  (not A234) );
 a37380a <=( A233  and  a37379a );
 a37383a <=( (not A268)  and  (not A267) );
 a37386a <=( A301  and  (not A269) );
 a37387a <=( a37386a  and  a37383a );
 a37388a <=( a37387a  and  a37380a );
 a37392a <=( (not A168)  and  (not A169) );
 a37393a <=( (not A170)  and  a37392a );
 a37397a <=( A232  and  A201 );
 a37398a <=( A200  and  a37397a );
 a37399a <=( a37398a  and  a37393a );
 a37403a <=( (not A235)  and  (not A234) );
 a37404a <=( A233  and  a37403a );
 a37407a <=( (not A266)  and  (not A265) );
 a37410a <=( A301  and  (not A268) );
 a37411a <=( a37410a  and  a37407a );
 a37412a <=( a37411a  and  a37404a );
 a37416a <=( (not A168)  and  (not A169) );
 a37417a <=( (not A170)  and  a37416a );
 a37421a <=( (not A232)  and  A201 );
 a37422a <=( A200  and  a37421a );
 a37423a <=( a37422a  and  a37417a );
 a37427a <=( (not A267)  and  (not A235) );
 a37428a <=( (not A233)  and  a37427a );
 a37431a <=( (not A269)  and  (not A268) );
 a37434a <=( A300  and  A299 );
 a37435a <=( a37434a  and  a37431a );
 a37436a <=( a37435a  and  a37428a );
 a37440a <=( (not A168)  and  (not A169) );
 a37441a <=( (not A170)  and  a37440a );
 a37445a <=( (not A232)  and  A201 );
 a37446a <=( A200  and  a37445a );
 a37447a <=( a37446a  and  a37441a );
 a37451a <=( (not A267)  and  (not A235) );
 a37452a <=( (not A233)  and  a37451a );
 a37455a <=( (not A269)  and  (not A268) );
 a37458a <=( A300  and  A298 );
 a37459a <=( a37458a  and  a37455a );
 a37460a <=( a37459a  and  a37452a );
 a37464a <=( (not A168)  and  (not A169) );
 a37465a <=( (not A170)  and  a37464a );
 a37469a <=( (not A232)  and  A201 );
 a37470a <=( A200  and  a37469a );
 a37471a <=( a37470a  and  a37465a );
 a37475a <=( A265  and  (not A235) );
 a37476a <=( (not A233)  and  a37475a );
 a37479a <=( (not A267)  and  A266 );
 a37482a <=( A301  and  (not A268) );
 a37483a <=( a37482a  and  a37479a );
 a37484a <=( a37483a  and  a37476a );
 a37488a <=( (not A168)  and  (not A169) );
 a37489a <=( (not A170)  and  a37488a );
 a37493a <=( (not A232)  and  A201 );
 a37494a <=( A200  and  a37493a );
 a37495a <=( a37494a  and  a37489a );
 a37499a <=( (not A265)  and  (not A235) );
 a37500a <=( (not A233)  and  a37499a );
 a37503a <=( (not A268)  and  (not A266) );
 a37506a <=( A300  and  A299 );
 a37507a <=( a37506a  and  a37503a );
 a37508a <=( a37507a  and  a37500a );
 a37512a <=( (not A168)  and  (not A169) );
 a37513a <=( (not A170)  and  a37512a );
 a37517a <=( (not A232)  and  A201 );
 a37518a <=( A200  and  a37517a );
 a37519a <=( a37518a  and  a37513a );
 a37523a <=( (not A265)  and  (not A235) );
 a37524a <=( (not A233)  and  a37523a );
 a37527a <=( (not A268)  and  (not A266) );
 a37530a <=( A300  and  A298 );
 a37531a <=( a37530a  and  a37527a );
 a37532a <=( a37531a  and  a37524a );
 a37536a <=( (not A168)  and  (not A169) );
 a37537a <=( (not A170)  and  a37536a );
 a37541a <=( A203  and  A200 );
 a37542a <=( (not A199)  and  a37541a );
 a37543a <=( a37542a  and  a37537a );
 a37547a <=( (not A236)  and  (not A235) );
 a37548a <=( (not A234)  and  a37547a );
 a37551a <=( (not A268)  and  (not A267) );
 a37554a <=( A301  and  (not A269) );
 a37555a <=( a37554a  and  a37551a );
 a37556a <=( a37555a  and  a37548a );
 a37560a <=( (not A168)  and  (not A169) );
 a37561a <=( (not A170)  and  a37560a );
 a37565a <=( A203  and  A200 );
 a37566a <=( (not A199)  and  a37565a );
 a37567a <=( a37566a  and  a37561a );
 a37571a <=( (not A236)  and  (not A235) );
 a37572a <=( (not A234)  and  a37571a );
 a37575a <=( (not A266)  and  (not A265) );
 a37578a <=( A301  and  (not A268) );
 a37579a <=( a37578a  and  a37575a );
 a37580a <=( a37579a  and  a37572a );
 a37584a <=( (not A168)  and  (not A169) );
 a37585a <=( (not A170)  and  a37584a );
 a37589a <=( A203  and  A200 );
 a37590a <=( (not A199)  and  a37589a );
 a37591a <=( a37590a  and  a37585a );
 a37595a <=( A236  and  A233 );
 a37596a <=( (not A232)  and  a37595a );
 a37599a <=( A299  and  A298 );
 a37602a <=( (not A301)  and  (not A300) );
 a37603a <=( a37602a  and  a37599a );
 a37604a <=( a37603a  and  a37596a );
 a37608a <=( (not A168)  and  (not A169) );
 a37609a <=( (not A170)  and  a37608a );
 a37613a <=( A203  and  A200 );
 a37614a <=( (not A199)  and  a37613a );
 a37615a <=( a37614a  and  a37609a );
 a37619a <=( A236  and  (not A233) );
 a37620a <=( A232  and  a37619a );
 a37623a <=( A299  and  A298 );
 a37626a <=( (not A301)  and  (not A300) );
 a37627a <=( a37626a  and  a37623a );
 a37628a <=( a37627a  and  a37620a );
 a37632a <=( (not A168)  and  (not A169) );
 a37633a <=( (not A170)  and  a37632a );
 a37637a <=( A203  and  A200 );
 a37638a <=( (not A199)  and  a37637a );
 a37639a <=( a37638a  and  a37633a );
 a37643a <=( (not A235)  and  (not A233) );
 a37644a <=( (not A232)  and  a37643a );
 a37647a <=( (not A268)  and  (not A267) );
 a37650a <=( A301  and  (not A269) );
 a37651a <=( a37650a  and  a37647a );
 a37652a <=( a37651a  and  a37644a );
 a37656a <=( (not A168)  and  (not A169) );
 a37657a <=( (not A170)  and  a37656a );
 a37661a <=( A203  and  A200 );
 a37662a <=( (not A199)  and  a37661a );
 a37663a <=( a37662a  and  a37657a );
 a37667a <=( (not A235)  and  (not A233) );
 a37668a <=( (not A232)  and  a37667a );
 a37671a <=( (not A266)  and  (not A265) );
 a37674a <=( A301  and  (not A268) );
 a37675a <=( a37674a  and  a37671a );
 a37676a <=( a37675a  and  a37668a );
 a37680a <=( (not A168)  and  (not A169) );
 a37681a <=( (not A170)  and  a37680a );
 a37685a <=( A203  and  (not A200) );
 a37686a <=( A199  and  a37685a );
 a37687a <=( a37686a  and  a37681a );
 a37691a <=( (not A236)  and  (not A235) );
 a37692a <=( (not A234)  and  a37691a );
 a37695a <=( (not A268)  and  (not A267) );
 a37698a <=( A301  and  (not A269) );
 a37699a <=( a37698a  and  a37695a );
 a37700a <=( a37699a  and  a37692a );
 a37704a <=( (not A168)  and  (not A169) );
 a37705a <=( (not A170)  and  a37704a );
 a37709a <=( A203  and  (not A200) );
 a37710a <=( A199  and  a37709a );
 a37711a <=( a37710a  and  a37705a );
 a37715a <=( (not A236)  and  (not A235) );
 a37716a <=( (not A234)  and  a37715a );
 a37719a <=( (not A266)  and  (not A265) );
 a37722a <=( A301  and  (not A268) );
 a37723a <=( a37722a  and  a37719a );
 a37724a <=( a37723a  and  a37716a );
 a37728a <=( (not A168)  and  (not A169) );
 a37729a <=( (not A170)  and  a37728a );
 a37733a <=( A203  and  (not A200) );
 a37734a <=( A199  and  a37733a );
 a37735a <=( a37734a  and  a37729a );
 a37739a <=( A236  and  A233 );
 a37740a <=( (not A232)  and  a37739a );
 a37743a <=( A299  and  A298 );
 a37746a <=( (not A301)  and  (not A300) );
 a37747a <=( a37746a  and  a37743a );
 a37748a <=( a37747a  and  a37740a );
 a37752a <=( (not A168)  and  (not A169) );
 a37753a <=( (not A170)  and  a37752a );
 a37757a <=( A203  and  (not A200) );
 a37758a <=( A199  and  a37757a );
 a37759a <=( a37758a  and  a37753a );
 a37763a <=( A236  and  (not A233) );
 a37764a <=( A232  and  a37763a );
 a37767a <=( A299  and  A298 );
 a37770a <=( (not A301)  and  (not A300) );
 a37771a <=( a37770a  and  a37767a );
 a37772a <=( a37771a  and  a37764a );
 a37776a <=( (not A168)  and  (not A169) );
 a37777a <=( (not A170)  and  a37776a );
 a37781a <=( A203  and  (not A200) );
 a37782a <=( A199  and  a37781a );
 a37783a <=( a37782a  and  a37777a );
 a37787a <=( (not A235)  and  (not A233) );
 a37788a <=( (not A232)  and  a37787a );
 a37791a <=( (not A268)  and  (not A267) );
 a37794a <=( A301  and  (not A269) );
 a37795a <=( a37794a  and  a37791a );
 a37796a <=( a37795a  and  a37788a );
 a37800a <=( (not A168)  and  (not A169) );
 a37801a <=( (not A170)  and  a37800a );
 a37805a <=( A203  and  (not A200) );
 a37806a <=( A199  and  a37805a );
 a37807a <=( a37806a  and  a37801a );
 a37811a <=( (not A235)  and  (not A233) );
 a37812a <=( (not A232)  and  a37811a );
 a37815a <=( (not A266)  and  (not A265) );
 a37818a <=( A301  and  (not A268) );
 a37819a <=( a37818a  and  a37815a );
 a37820a <=( a37819a  and  a37812a );
 a37824a <=( (not A201)  and  A166 );
 a37825a <=( A168  and  a37824a );
 a37828a <=( (not A203)  and  (not A202) );
 a37831a <=( (not A235)  and  (not A234) );
 a37832a <=( a37831a  and  a37828a );
 a37833a <=( a37832a  and  a37825a );
 a37837a <=( (not A268)  and  (not A267) );
 a37838a <=( (not A236)  and  a37837a );
 a37841a <=( A298  and  (not A269) );
 a37844a <=( A302  and  (not A299) );
 a37845a <=( a37844a  and  a37841a );
 a37846a <=( a37845a  and  a37838a );
 a37850a <=( (not A201)  and  A166 );
 a37851a <=( A168  and  a37850a );
 a37854a <=( (not A203)  and  (not A202) );
 a37857a <=( (not A235)  and  (not A234) );
 a37858a <=( a37857a  and  a37854a );
 a37859a <=( a37858a  and  a37851a );
 a37863a <=( (not A268)  and  (not A267) );
 a37864a <=( (not A236)  and  a37863a );
 a37867a <=( (not A298)  and  (not A269) );
 a37870a <=( A302  and  A299 );
 a37871a <=( a37870a  and  a37867a );
 a37872a <=( a37871a  and  a37864a );
 a37876a <=( (not A201)  and  A166 );
 a37877a <=( A168  and  a37876a );
 a37880a <=( (not A203)  and  (not A202) );
 a37883a <=( (not A235)  and  (not A234) );
 a37884a <=( a37883a  and  a37880a );
 a37885a <=( a37884a  and  a37877a );
 a37889a <=( A266  and  A265 );
 a37890a <=( (not A236)  and  a37889a );
 a37893a <=( (not A268)  and  (not A267) );
 a37896a <=( A300  and  A299 );
 a37897a <=( a37896a  and  a37893a );
 a37898a <=( a37897a  and  a37890a );
 a37902a <=( (not A201)  and  A166 );
 a37903a <=( A168  and  a37902a );
 a37906a <=( (not A203)  and  (not A202) );
 a37909a <=( (not A235)  and  (not A234) );
 a37910a <=( a37909a  and  a37906a );
 a37911a <=( a37910a  and  a37903a );
 a37915a <=( A266  and  A265 );
 a37916a <=( (not A236)  and  a37915a );
 a37919a <=( (not A268)  and  (not A267) );
 a37922a <=( A300  and  A298 );
 a37923a <=( a37922a  and  a37919a );
 a37924a <=( a37923a  and  a37916a );
 a37928a <=( (not A201)  and  A166 );
 a37929a <=( A168  and  a37928a );
 a37932a <=( (not A203)  and  (not A202) );
 a37935a <=( (not A235)  and  (not A234) );
 a37936a <=( a37935a  and  a37932a );
 a37937a <=( a37936a  and  a37929a );
 a37941a <=( (not A266)  and  (not A265) );
 a37942a <=( (not A236)  and  a37941a );
 a37945a <=( A298  and  (not A268) );
 a37948a <=( A302  and  (not A299) );
 a37949a <=( a37948a  and  a37945a );
 a37950a <=( a37949a  and  a37942a );
 a37954a <=( (not A201)  and  A166 );
 a37955a <=( A168  and  a37954a );
 a37958a <=( (not A203)  and  (not A202) );
 a37961a <=( (not A235)  and  (not A234) );
 a37962a <=( a37961a  and  a37958a );
 a37963a <=( a37962a  and  a37955a );
 a37967a <=( (not A266)  and  (not A265) );
 a37968a <=( (not A236)  and  a37967a );
 a37971a <=( (not A298)  and  (not A268) );
 a37974a <=( A302  and  A299 );
 a37975a <=( a37974a  and  a37971a );
 a37976a <=( a37975a  and  a37968a );
 a37980a <=( (not A201)  and  A166 );
 a37981a <=( A168  and  a37980a );
 a37984a <=( (not A203)  and  (not A202) );
 a37987a <=( A233  and  A232 );
 a37988a <=( a37987a  and  a37984a );
 a37989a <=( a37988a  and  a37981a );
 a37993a <=( (not A267)  and  (not A235) );
 a37994a <=( (not A234)  and  a37993a );
 a37997a <=( (not A269)  and  (not A268) );
 a38000a <=( A300  and  A299 );
 a38001a <=( a38000a  and  a37997a );
 a38002a <=( a38001a  and  a37994a );
 a38006a <=( (not A201)  and  A166 );
 a38007a <=( A168  and  a38006a );
 a38010a <=( (not A203)  and  (not A202) );
 a38013a <=( A233  and  A232 );
 a38014a <=( a38013a  and  a38010a );
 a38015a <=( a38014a  and  a38007a );
 a38019a <=( (not A267)  and  (not A235) );
 a38020a <=( (not A234)  and  a38019a );
 a38023a <=( (not A269)  and  (not A268) );
 a38026a <=( A300  and  A298 );
 a38027a <=( a38026a  and  a38023a );
 a38028a <=( a38027a  and  a38020a );
 a38032a <=( (not A201)  and  A166 );
 a38033a <=( A168  and  a38032a );
 a38036a <=( (not A203)  and  (not A202) );
 a38039a <=( A233  and  A232 );
 a38040a <=( a38039a  and  a38036a );
 a38041a <=( a38040a  and  a38033a );
 a38045a <=( A265  and  (not A235) );
 a38046a <=( (not A234)  and  a38045a );
 a38049a <=( (not A267)  and  A266 );
 a38052a <=( A301  and  (not A268) );
 a38053a <=( a38052a  and  a38049a );
 a38054a <=( a38053a  and  a38046a );
 a38058a <=( (not A201)  and  A166 );
 a38059a <=( A168  and  a38058a );
 a38062a <=( (not A203)  and  (not A202) );
 a38065a <=( A233  and  A232 );
 a38066a <=( a38065a  and  a38062a );
 a38067a <=( a38066a  and  a38059a );
 a38071a <=( (not A265)  and  (not A235) );
 a38072a <=( (not A234)  and  a38071a );
 a38075a <=( (not A268)  and  (not A266) );
 a38078a <=( A300  and  A299 );
 a38079a <=( a38078a  and  a38075a );
 a38080a <=( a38079a  and  a38072a );
 a38084a <=( (not A201)  and  A166 );
 a38085a <=( A168  and  a38084a );
 a38088a <=( (not A203)  and  (not A202) );
 a38091a <=( A233  and  A232 );
 a38092a <=( a38091a  and  a38088a );
 a38093a <=( a38092a  and  a38085a );
 a38097a <=( (not A265)  and  (not A235) );
 a38098a <=( (not A234)  and  a38097a );
 a38101a <=( (not A268)  and  (not A266) );
 a38104a <=( A300  and  A298 );
 a38105a <=( a38104a  and  a38101a );
 a38106a <=( a38105a  and  a38098a );
 a38110a <=( (not A201)  and  A166 );
 a38111a <=( A168  and  a38110a );
 a38114a <=( (not A203)  and  (not A202) );
 a38117a <=( (not A233)  and  (not A232) );
 a38118a <=( a38117a  and  a38114a );
 a38119a <=( a38118a  and  a38111a );
 a38123a <=( (not A268)  and  (not A267) );
 a38124a <=( (not A235)  and  a38123a );
 a38127a <=( A298  and  (not A269) );
 a38130a <=( A302  and  (not A299) );
 a38131a <=( a38130a  and  a38127a );
 a38132a <=( a38131a  and  a38124a );
 a38136a <=( (not A201)  and  A166 );
 a38137a <=( A168  and  a38136a );
 a38140a <=( (not A203)  and  (not A202) );
 a38143a <=( (not A233)  and  (not A232) );
 a38144a <=( a38143a  and  a38140a );
 a38145a <=( a38144a  and  a38137a );
 a38149a <=( (not A268)  and  (not A267) );
 a38150a <=( (not A235)  and  a38149a );
 a38153a <=( (not A298)  and  (not A269) );
 a38156a <=( A302  and  A299 );
 a38157a <=( a38156a  and  a38153a );
 a38158a <=( a38157a  and  a38150a );
 a38162a <=( (not A201)  and  A166 );
 a38163a <=( A168  and  a38162a );
 a38166a <=( (not A203)  and  (not A202) );
 a38169a <=( (not A233)  and  (not A232) );
 a38170a <=( a38169a  and  a38166a );
 a38171a <=( a38170a  and  a38163a );
 a38175a <=( A266  and  A265 );
 a38176a <=( (not A235)  and  a38175a );
 a38179a <=( (not A268)  and  (not A267) );
 a38182a <=( A300  and  A299 );
 a38183a <=( a38182a  and  a38179a );
 a38184a <=( a38183a  and  a38176a );
 a38188a <=( (not A201)  and  A166 );
 a38189a <=( A168  and  a38188a );
 a38192a <=( (not A203)  and  (not A202) );
 a38195a <=( (not A233)  and  (not A232) );
 a38196a <=( a38195a  and  a38192a );
 a38197a <=( a38196a  and  a38189a );
 a38201a <=( A266  and  A265 );
 a38202a <=( (not A235)  and  a38201a );
 a38205a <=( (not A268)  and  (not A267) );
 a38208a <=( A300  and  A298 );
 a38209a <=( a38208a  and  a38205a );
 a38210a <=( a38209a  and  a38202a );
 a38214a <=( (not A201)  and  A166 );
 a38215a <=( A168  and  a38214a );
 a38218a <=( (not A203)  and  (not A202) );
 a38221a <=( (not A233)  and  (not A232) );
 a38222a <=( a38221a  and  a38218a );
 a38223a <=( a38222a  and  a38215a );
 a38227a <=( (not A266)  and  (not A265) );
 a38228a <=( (not A235)  and  a38227a );
 a38231a <=( A298  and  (not A268) );
 a38234a <=( A302  and  (not A299) );
 a38235a <=( a38234a  and  a38231a );
 a38236a <=( a38235a  and  a38228a );
 a38240a <=( (not A201)  and  A166 );
 a38241a <=( A168  and  a38240a );
 a38244a <=( (not A203)  and  (not A202) );
 a38247a <=( (not A233)  and  (not A232) );
 a38248a <=( a38247a  and  a38244a );
 a38249a <=( a38248a  and  a38241a );
 a38253a <=( (not A266)  and  (not A265) );
 a38254a <=( (not A235)  and  a38253a );
 a38257a <=( (not A298)  and  (not A268) );
 a38260a <=( A302  and  A299 );
 a38261a <=( a38260a  and  a38257a );
 a38262a <=( a38261a  and  a38254a );
 a38266a <=( A199  and  A166 );
 a38267a <=( A168  and  a38266a );
 a38270a <=( (not A201)  and  A200 );
 a38273a <=( (not A234)  and  (not A202) );
 a38274a <=( a38273a  and  a38270a );
 a38275a <=( a38274a  and  a38267a );
 a38279a <=( (not A267)  and  (not A236) );
 a38280a <=( (not A235)  and  a38279a );
 a38283a <=( (not A269)  and  (not A268) );
 a38286a <=( A300  and  A299 );
 a38287a <=( a38286a  and  a38283a );
 a38288a <=( a38287a  and  a38280a );
 a38292a <=( A199  and  A166 );
 a38293a <=( A168  and  a38292a );
 a38296a <=( (not A201)  and  A200 );
 a38299a <=( (not A234)  and  (not A202) );
 a38300a <=( a38299a  and  a38296a );
 a38301a <=( a38300a  and  a38293a );
 a38305a <=( (not A267)  and  (not A236) );
 a38306a <=( (not A235)  and  a38305a );
 a38309a <=( (not A269)  and  (not A268) );
 a38312a <=( A300  and  A298 );
 a38313a <=( a38312a  and  a38309a );
 a38314a <=( a38313a  and  a38306a );
 a38318a <=( A199  and  A166 );
 a38319a <=( A168  and  a38318a );
 a38322a <=( (not A201)  and  A200 );
 a38325a <=( (not A234)  and  (not A202) );
 a38326a <=( a38325a  and  a38322a );
 a38327a <=( a38326a  and  a38319a );
 a38331a <=( A265  and  (not A236) );
 a38332a <=( (not A235)  and  a38331a );
 a38335a <=( (not A267)  and  A266 );
 a38338a <=( A301  and  (not A268) );
 a38339a <=( a38338a  and  a38335a );
 a38340a <=( a38339a  and  a38332a );
 a38344a <=( A199  and  A166 );
 a38345a <=( A168  and  a38344a );
 a38348a <=( (not A201)  and  A200 );
 a38351a <=( (not A234)  and  (not A202) );
 a38352a <=( a38351a  and  a38348a );
 a38353a <=( a38352a  and  a38345a );
 a38357a <=( (not A265)  and  (not A236) );
 a38358a <=( (not A235)  and  a38357a );
 a38361a <=( (not A268)  and  (not A266) );
 a38364a <=( A300  and  A299 );
 a38365a <=( a38364a  and  a38361a );
 a38366a <=( a38365a  and  a38358a );
 a38370a <=( A199  and  A166 );
 a38371a <=( A168  and  a38370a );
 a38374a <=( (not A201)  and  A200 );
 a38377a <=( (not A234)  and  (not A202) );
 a38378a <=( a38377a  and  a38374a );
 a38379a <=( a38378a  and  a38371a );
 a38383a <=( (not A265)  and  (not A236) );
 a38384a <=( (not A235)  and  a38383a );
 a38387a <=( (not A268)  and  (not A266) );
 a38390a <=( A300  and  A298 );
 a38391a <=( a38390a  and  a38387a );
 a38392a <=( a38391a  and  a38384a );
 a38396a <=( A199  and  A166 );
 a38397a <=( A168  and  a38396a );
 a38400a <=( (not A201)  and  A200 );
 a38403a <=( A232  and  (not A202) );
 a38404a <=( a38403a  and  a38400a );
 a38405a <=( a38404a  and  a38397a );
 a38409a <=( (not A235)  and  (not A234) );
 a38410a <=( A233  and  a38409a );
 a38413a <=( (not A268)  and  (not A267) );
 a38416a <=( A301  and  (not A269) );
 a38417a <=( a38416a  and  a38413a );
 a38418a <=( a38417a  and  a38410a );
 a38422a <=( A199  and  A166 );
 a38423a <=( A168  and  a38422a );
 a38426a <=( (not A201)  and  A200 );
 a38429a <=( A232  and  (not A202) );
 a38430a <=( a38429a  and  a38426a );
 a38431a <=( a38430a  and  a38423a );
 a38435a <=( (not A235)  and  (not A234) );
 a38436a <=( A233  and  a38435a );
 a38439a <=( (not A266)  and  (not A265) );
 a38442a <=( A301  and  (not A268) );
 a38443a <=( a38442a  and  a38439a );
 a38444a <=( a38443a  and  a38436a );
 a38448a <=( A199  and  A166 );
 a38449a <=( A168  and  a38448a );
 a38452a <=( (not A201)  and  A200 );
 a38455a <=( (not A232)  and  (not A202) );
 a38456a <=( a38455a  and  a38452a );
 a38457a <=( a38456a  and  a38449a );
 a38461a <=( (not A267)  and  (not A235) );
 a38462a <=( (not A233)  and  a38461a );
 a38465a <=( (not A269)  and  (not A268) );
 a38468a <=( A300  and  A299 );
 a38469a <=( a38468a  and  a38465a );
 a38470a <=( a38469a  and  a38462a );
 a38474a <=( A199  and  A166 );
 a38475a <=( A168  and  a38474a );
 a38478a <=( (not A201)  and  A200 );
 a38481a <=( (not A232)  and  (not A202) );
 a38482a <=( a38481a  and  a38478a );
 a38483a <=( a38482a  and  a38475a );
 a38487a <=( (not A267)  and  (not A235) );
 a38488a <=( (not A233)  and  a38487a );
 a38491a <=( (not A269)  and  (not A268) );
 a38494a <=( A300  and  A298 );
 a38495a <=( a38494a  and  a38491a );
 a38496a <=( a38495a  and  a38488a );
 a38500a <=( A199  and  A166 );
 a38501a <=( A168  and  a38500a );
 a38504a <=( (not A201)  and  A200 );
 a38507a <=( (not A232)  and  (not A202) );
 a38508a <=( a38507a  and  a38504a );
 a38509a <=( a38508a  and  a38501a );
 a38513a <=( A265  and  (not A235) );
 a38514a <=( (not A233)  and  a38513a );
 a38517a <=( (not A267)  and  A266 );
 a38520a <=( A301  and  (not A268) );
 a38521a <=( a38520a  and  a38517a );
 a38522a <=( a38521a  and  a38514a );
 a38526a <=( A199  and  A166 );
 a38527a <=( A168  and  a38526a );
 a38530a <=( (not A201)  and  A200 );
 a38533a <=( (not A232)  and  (not A202) );
 a38534a <=( a38533a  and  a38530a );
 a38535a <=( a38534a  and  a38527a );
 a38539a <=( (not A265)  and  (not A235) );
 a38540a <=( (not A233)  and  a38539a );
 a38543a <=( (not A268)  and  (not A266) );
 a38546a <=( A300  and  A299 );
 a38547a <=( a38546a  and  a38543a );
 a38548a <=( a38547a  and  a38540a );
 a38552a <=( A199  and  A166 );
 a38553a <=( A168  and  a38552a );
 a38556a <=( (not A201)  and  A200 );
 a38559a <=( (not A232)  and  (not A202) );
 a38560a <=( a38559a  and  a38556a );
 a38561a <=( a38560a  and  a38553a );
 a38565a <=( (not A265)  and  (not A235) );
 a38566a <=( (not A233)  and  a38565a );
 a38569a <=( (not A268)  and  (not A266) );
 a38572a <=( A300  and  A298 );
 a38573a <=( a38572a  and  a38569a );
 a38574a <=( a38573a  and  a38566a );
 a38578a <=( (not A199)  and  A166 );
 a38579a <=( A168  and  a38578a );
 a38582a <=( (not A202)  and  (not A200) );
 a38585a <=( (not A235)  and  (not A234) );
 a38586a <=( a38585a  and  a38582a );
 a38587a <=( a38586a  and  a38579a );
 a38591a <=( (not A268)  and  (not A267) );
 a38592a <=( (not A236)  and  a38591a );
 a38595a <=( A298  and  (not A269) );
 a38598a <=( A302  and  (not A299) );
 a38599a <=( a38598a  and  a38595a );
 a38600a <=( a38599a  and  a38592a );
 a38604a <=( (not A199)  and  A166 );
 a38605a <=( A168  and  a38604a );
 a38608a <=( (not A202)  and  (not A200) );
 a38611a <=( (not A235)  and  (not A234) );
 a38612a <=( a38611a  and  a38608a );
 a38613a <=( a38612a  and  a38605a );
 a38617a <=( (not A268)  and  (not A267) );
 a38618a <=( (not A236)  and  a38617a );
 a38621a <=( (not A298)  and  (not A269) );
 a38624a <=( A302  and  A299 );
 a38625a <=( a38624a  and  a38621a );
 a38626a <=( a38625a  and  a38618a );
 a38630a <=( (not A199)  and  A166 );
 a38631a <=( A168  and  a38630a );
 a38634a <=( (not A202)  and  (not A200) );
 a38637a <=( (not A235)  and  (not A234) );
 a38638a <=( a38637a  and  a38634a );
 a38639a <=( a38638a  and  a38631a );
 a38643a <=( A266  and  A265 );
 a38644a <=( (not A236)  and  a38643a );
 a38647a <=( (not A268)  and  (not A267) );
 a38650a <=( A300  and  A299 );
 a38651a <=( a38650a  and  a38647a );
 a38652a <=( a38651a  and  a38644a );
 a38656a <=( (not A199)  and  A166 );
 a38657a <=( A168  and  a38656a );
 a38660a <=( (not A202)  and  (not A200) );
 a38663a <=( (not A235)  and  (not A234) );
 a38664a <=( a38663a  and  a38660a );
 a38665a <=( a38664a  and  a38657a );
 a38669a <=( A266  and  A265 );
 a38670a <=( (not A236)  and  a38669a );
 a38673a <=( (not A268)  and  (not A267) );
 a38676a <=( A300  and  A298 );
 a38677a <=( a38676a  and  a38673a );
 a38678a <=( a38677a  and  a38670a );
 a38682a <=( (not A199)  and  A166 );
 a38683a <=( A168  and  a38682a );
 a38686a <=( (not A202)  and  (not A200) );
 a38689a <=( (not A235)  and  (not A234) );
 a38690a <=( a38689a  and  a38686a );
 a38691a <=( a38690a  and  a38683a );
 a38695a <=( (not A266)  and  (not A265) );
 a38696a <=( (not A236)  and  a38695a );
 a38699a <=( A298  and  (not A268) );
 a38702a <=( A302  and  (not A299) );
 a38703a <=( a38702a  and  a38699a );
 a38704a <=( a38703a  and  a38696a );
 a38708a <=( (not A199)  and  A166 );
 a38709a <=( A168  and  a38708a );
 a38712a <=( (not A202)  and  (not A200) );
 a38715a <=( (not A235)  and  (not A234) );
 a38716a <=( a38715a  and  a38712a );
 a38717a <=( a38716a  and  a38709a );
 a38721a <=( (not A266)  and  (not A265) );
 a38722a <=( (not A236)  and  a38721a );
 a38725a <=( (not A298)  and  (not A268) );
 a38728a <=( A302  and  A299 );
 a38729a <=( a38728a  and  a38725a );
 a38730a <=( a38729a  and  a38722a );
 a38734a <=( (not A199)  and  A166 );
 a38735a <=( A168  and  a38734a );
 a38738a <=( (not A202)  and  (not A200) );
 a38741a <=( A233  and  A232 );
 a38742a <=( a38741a  and  a38738a );
 a38743a <=( a38742a  and  a38735a );
 a38747a <=( (not A267)  and  (not A235) );
 a38748a <=( (not A234)  and  a38747a );
 a38751a <=( (not A269)  and  (not A268) );
 a38754a <=( A300  and  A299 );
 a38755a <=( a38754a  and  a38751a );
 a38756a <=( a38755a  and  a38748a );
 a38760a <=( (not A199)  and  A166 );
 a38761a <=( A168  and  a38760a );
 a38764a <=( (not A202)  and  (not A200) );
 a38767a <=( A233  and  A232 );
 a38768a <=( a38767a  and  a38764a );
 a38769a <=( a38768a  and  a38761a );
 a38773a <=( (not A267)  and  (not A235) );
 a38774a <=( (not A234)  and  a38773a );
 a38777a <=( (not A269)  and  (not A268) );
 a38780a <=( A300  and  A298 );
 a38781a <=( a38780a  and  a38777a );
 a38782a <=( a38781a  and  a38774a );
 a38786a <=( (not A199)  and  A166 );
 a38787a <=( A168  and  a38786a );
 a38790a <=( (not A202)  and  (not A200) );
 a38793a <=( A233  and  A232 );
 a38794a <=( a38793a  and  a38790a );
 a38795a <=( a38794a  and  a38787a );
 a38799a <=( A265  and  (not A235) );
 a38800a <=( (not A234)  and  a38799a );
 a38803a <=( (not A267)  and  A266 );
 a38806a <=( A301  and  (not A268) );
 a38807a <=( a38806a  and  a38803a );
 a38808a <=( a38807a  and  a38800a );
 a38812a <=( (not A199)  and  A166 );
 a38813a <=( A168  and  a38812a );
 a38816a <=( (not A202)  and  (not A200) );
 a38819a <=( A233  and  A232 );
 a38820a <=( a38819a  and  a38816a );
 a38821a <=( a38820a  and  a38813a );
 a38825a <=( (not A265)  and  (not A235) );
 a38826a <=( (not A234)  and  a38825a );
 a38829a <=( (not A268)  and  (not A266) );
 a38832a <=( A300  and  A299 );
 a38833a <=( a38832a  and  a38829a );
 a38834a <=( a38833a  and  a38826a );
 a38838a <=( (not A199)  and  A166 );
 a38839a <=( A168  and  a38838a );
 a38842a <=( (not A202)  and  (not A200) );
 a38845a <=( A233  and  A232 );
 a38846a <=( a38845a  and  a38842a );
 a38847a <=( a38846a  and  a38839a );
 a38851a <=( (not A265)  and  (not A235) );
 a38852a <=( (not A234)  and  a38851a );
 a38855a <=( (not A268)  and  (not A266) );
 a38858a <=( A300  and  A298 );
 a38859a <=( a38858a  and  a38855a );
 a38860a <=( a38859a  and  a38852a );
 a38864a <=( (not A199)  and  A166 );
 a38865a <=( A168  and  a38864a );
 a38868a <=( (not A202)  and  (not A200) );
 a38871a <=( (not A233)  and  (not A232) );
 a38872a <=( a38871a  and  a38868a );
 a38873a <=( a38872a  and  a38865a );
 a38877a <=( (not A268)  and  (not A267) );
 a38878a <=( (not A235)  and  a38877a );
 a38881a <=( A298  and  (not A269) );
 a38884a <=( A302  and  (not A299) );
 a38885a <=( a38884a  and  a38881a );
 a38886a <=( a38885a  and  a38878a );
 a38890a <=( (not A199)  and  A166 );
 a38891a <=( A168  and  a38890a );
 a38894a <=( (not A202)  and  (not A200) );
 a38897a <=( (not A233)  and  (not A232) );
 a38898a <=( a38897a  and  a38894a );
 a38899a <=( a38898a  and  a38891a );
 a38903a <=( (not A268)  and  (not A267) );
 a38904a <=( (not A235)  and  a38903a );
 a38907a <=( (not A298)  and  (not A269) );
 a38910a <=( A302  and  A299 );
 a38911a <=( a38910a  and  a38907a );
 a38912a <=( a38911a  and  a38904a );
 a38916a <=( (not A199)  and  A166 );
 a38917a <=( A168  and  a38916a );
 a38920a <=( (not A202)  and  (not A200) );
 a38923a <=( (not A233)  and  (not A232) );
 a38924a <=( a38923a  and  a38920a );
 a38925a <=( a38924a  and  a38917a );
 a38929a <=( A266  and  A265 );
 a38930a <=( (not A235)  and  a38929a );
 a38933a <=( (not A268)  and  (not A267) );
 a38936a <=( A300  and  A299 );
 a38937a <=( a38936a  and  a38933a );
 a38938a <=( a38937a  and  a38930a );
 a38942a <=( (not A199)  and  A166 );
 a38943a <=( A168  and  a38942a );
 a38946a <=( (not A202)  and  (not A200) );
 a38949a <=( (not A233)  and  (not A232) );
 a38950a <=( a38949a  and  a38946a );
 a38951a <=( a38950a  and  a38943a );
 a38955a <=( A266  and  A265 );
 a38956a <=( (not A235)  and  a38955a );
 a38959a <=( (not A268)  and  (not A267) );
 a38962a <=( A300  and  A298 );
 a38963a <=( a38962a  and  a38959a );
 a38964a <=( a38963a  and  a38956a );
 a38968a <=( (not A199)  and  A166 );
 a38969a <=( A168  and  a38968a );
 a38972a <=( (not A202)  and  (not A200) );
 a38975a <=( (not A233)  and  (not A232) );
 a38976a <=( a38975a  and  a38972a );
 a38977a <=( a38976a  and  a38969a );
 a38981a <=( (not A266)  and  (not A265) );
 a38982a <=( (not A235)  and  a38981a );
 a38985a <=( A298  and  (not A268) );
 a38988a <=( A302  and  (not A299) );
 a38989a <=( a38988a  and  a38985a );
 a38990a <=( a38989a  and  a38982a );
 a38994a <=( (not A199)  and  A166 );
 a38995a <=( A168  and  a38994a );
 a38998a <=( (not A202)  and  (not A200) );
 a39001a <=( (not A233)  and  (not A232) );
 a39002a <=( a39001a  and  a38998a );
 a39003a <=( a39002a  and  a38995a );
 a39007a <=( (not A266)  and  (not A265) );
 a39008a <=( (not A235)  and  a39007a );
 a39011a <=( (not A298)  and  (not A268) );
 a39014a <=( A302  and  A299 );
 a39015a <=( a39014a  and  a39011a );
 a39016a <=( a39015a  and  a39008a );
 a39020a <=( (not A201)  and  A167 );
 a39021a <=( A168  and  a39020a );
 a39024a <=( (not A203)  and  (not A202) );
 a39027a <=( (not A235)  and  (not A234) );
 a39028a <=( a39027a  and  a39024a );
 a39029a <=( a39028a  and  a39021a );
 a39033a <=( (not A268)  and  (not A267) );
 a39034a <=( (not A236)  and  a39033a );
 a39037a <=( A298  and  (not A269) );
 a39040a <=( A302  and  (not A299) );
 a39041a <=( a39040a  and  a39037a );
 a39042a <=( a39041a  and  a39034a );
 a39046a <=( (not A201)  and  A167 );
 a39047a <=( A168  and  a39046a );
 a39050a <=( (not A203)  and  (not A202) );
 a39053a <=( (not A235)  and  (not A234) );
 a39054a <=( a39053a  and  a39050a );
 a39055a <=( a39054a  and  a39047a );
 a39059a <=( (not A268)  and  (not A267) );
 a39060a <=( (not A236)  and  a39059a );
 a39063a <=( (not A298)  and  (not A269) );
 a39066a <=( A302  and  A299 );
 a39067a <=( a39066a  and  a39063a );
 a39068a <=( a39067a  and  a39060a );
 a39072a <=( (not A201)  and  A167 );
 a39073a <=( A168  and  a39072a );
 a39076a <=( (not A203)  and  (not A202) );
 a39079a <=( (not A235)  and  (not A234) );
 a39080a <=( a39079a  and  a39076a );
 a39081a <=( a39080a  and  a39073a );
 a39085a <=( A266  and  A265 );
 a39086a <=( (not A236)  and  a39085a );
 a39089a <=( (not A268)  and  (not A267) );
 a39092a <=( A300  and  A299 );
 a39093a <=( a39092a  and  a39089a );
 a39094a <=( a39093a  and  a39086a );
 a39098a <=( (not A201)  and  A167 );
 a39099a <=( A168  and  a39098a );
 a39102a <=( (not A203)  and  (not A202) );
 a39105a <=( (not A235)  and  (not A234) );
 a39106a <=( a39105a  and  a39102a );
 a39107a <=( a39106a  and  a39099a );
 a39111a <=( A266  and  A265 );
 a39112a <=( (not A236)  and  a39111a );
 a39115a <=( (not A268)  and  (not A267) );
 a39118a <=( A300  and  A298 );
 a39119a <=( a39118a  and  a39115a );
 a39120a <=( a39119a  and  a39112a );
 a39124a <=( (not A201)  and  A167 );
 a39125a <=( A168  and  a39124a );
 a39128a <=( (not A203)  and  (not A202) );
 a39131a <=( (not A235)  and  (not A234) );
 a39132a <=( a39131a  and  a39128a );
 a39133a <=( a39132a  and  a39125a );
 a39137a <=( (not A266)  and  (not A265) );
 a39138a <=( (not A236)  and  a39137a );
 a39141a <=( A298  and  (not A268) );
 a39144a <=( A302  and  (not A299) );
 a39145a <=( a39144a  and  a39141a );
 a39146a <=( a39145a  and  a39138a );
 a39150a <=( (not A201)  and  A167 );
 a39151a <=( A168  and  a39150a );
 a39154a <=( (not A203)  and  (not A202) );
 a39157a <=( (not A235)  and  (not A234) );
 a39158a <=( a39157a  and  a39154a );
 a39159a <=( a39158a  and  a39151a );
 a39163a <=( (not A266)  and  (not A265) );
 a39164a <=( (not A236)  and  a39163a );
 a39167a <=( (not A298)  and  (not A268) );
 a39170a <=( A302  and  A299 );
 a39171a <=( a39170a  and  a39167a );
 a39172a <=( a39171a  and  a39164a );
 a39176a <=( (not A201)  and  A167 );
 a39177a <=( A168  and  a39176a );
 a39180a <=( (not A203)  and  (not A202) );
 a39183a <=( A233  and  A232 );
 a39184a <=( a39183a  and  a39180a );
 a39185a <=( a39184a  and  a39177a );
 a39189a <=( (not A267)  and  (not A235) );
 a39190a <=( (not A234)  and  a39189a );
 a39193a <=( (not A269)  and  (not A268) );
 a39196a <=( A300  and  A299 );
 a39197a <=( a39196a  and  a39193a );
 a39198a <=( a39197a  and  a39190a );
 a39202a <=( (not A201)  and  A167 );
 a39203a <=( A168  and  a39202a );
 a39206a <=( (not A203)  and  (not A202) );
 a39209a <=( A233  and  A232 );
 a39210a <=( a39209a  and  a39206a );
 a39211a <=( a39210a  and  a39203a );
 a39215a <=( (not A267)  and  (not A235) );
 a39216a <=( (not A234)  and  a39215a );
 a39219a <=( (not A269)  and  (not A268) );
 a39222a <=( A300  and  A298 );
 a39223a <=( a39222a  and  a39219a );
 a39224a <=( a39223a  and  a39216a );
 a39228a <=( (not A201)  and  A167 );
 a39229a <=( A168  and  a39228a );
 a39232a <=( (not A203)  and  (not A202) );
 a39235a <=( A233  and  A232 );
 a39236a <=( a39235a  and  a39232a );
 a39237a <=( a39236a  and  a39229a );
 a39241a <=( A265  and  (not A235) );
 a39242a <=( (not A234)  and  a39241a );
 a39245a <=( (not A267)  and  A266 );
 a39248a <=( A301  and  (not A268) );
 a39249a <=( a39248a  and  a39245a );
 a39250a <=( a39249a  and  a39242a );
 a39254a <=( (not A201)  and  A167 );
 a39255a <=( A168  and  a39254a );
 a39258a <=( (not A203)  and  (not A202) );
 a39261a <=( A233  and  A232 );
 a39262a <=( a39261a  and  a39258a );
 a39263a <=( a39262a  and  a39255a );
 a39267a <=( (not A265)  and  (not A235) );
 a39268a <=( (not A234)  and  a39267a );
 a39271a <=( (not A268)  and  (not A266) );
 a39274a <=( A300  and  A299 );
 a39275a <=( a39274a  and  a39271a );
 a39276a <=( a39275a  and  a39268a );
 a39280a <=( (not A201)  and  A167 );
 a39281a <=( A168  and  a39280a );
 a39284a <=( (not A203)  and  (not A202) );
 a39287a <=( A233  and  A232 );
 a39288a <=( a39287a  and  a39284a );
 a39289a <=( a39288a  and  a39281a );
 a39293a <=( (not A265)  and  (not A235) );
 a39294a <=( (not A234)  and  a39293a );
 a39297a <=( (not A268)  and  (not A266) );
 a39300a <=( A300  and  A298 );
 a39301a <=( a39300a  and  a39297a );
 a39302a <=( a39301a  and  a39294a );
 a39306a <=( (not A201)  and  A167 );
 a39307a <=( A168  and  a39306a );
 a39310a <=( (not A203)  and  (not A202) );
 a39313a <=( (not A233)  and  (not A232) );
 a39314a <=( a39313a  and  a39310a );
 a39315a <=( a39314a  and  a39307a );
 a39319a <=( (not A268)  and  (not A267) );
 a39320a <=( (not A235)  and  a39319a );
 a39323a <=( A298  and  (not A269) );
 a39326a <=( A302  and  (not A299) );
 a39327a <=( a39326a  and  a39323a );
 a39328a <=( a39327a  and  a39320a );
 a39332a <=( (not A201)  and  A167 );
 a39333a <=( A168  and  a39332a );
 a39336a <=( (not A203)  and  (not A202) );
 a39339a <=( (not A233)  and  (not A232) );
 a39340a <=( a39339a  and  a39336a );
 a39341a <=( a39340a  and  a39333a );
 a39345a <=( (not A268)  and  (not A267) );
 a39346a <=( (not A235)  and  a39345a );
 a39349a <=( (not A298)  and  (not A269) );
 a39352a <=( A302  and  A299 );
 a39353a <=( a39352a  and  a39349a );
 a39354a <=( a39353a  and  a39346a );
 a39358a <=( (not A201)  and  A167 );
 a39359a <=( A168  and  a39358a );
 a39362a <=( (not A203)  and  (not A202) );
 a39365a <=( (not A233)  and  (not A232) );
 a39366a <=( a39365a  and  a39362a );
 a39367a <=( a39366a  and  a39359a );
 a39371a <=( A266  and  A265 );
 a39372a <=( (not A235)  and  a39371a );
 a39375a <=( (not A268)  and  (not A267) );
 a39378a <=( A300  and  A299 );
 a39379a <=( a39378a  and  a39375a );
 a39380a <=( a39379a  and  a39372a );
 a39384a <=( (not A201)  and  A167 );
 a39385a <=( A168  and  a39384a );
 a39388a <=( (not A203)  and  (not A202) );
 a39391a <=( (not A233)  and  (not A232) );
 a39392a <=( a39391a  and  a39388a );
 a39393a <=( a39392a  and  a39385a );
 a39397a <=( A266  and  A265 );
 a39398a <=( (not A235)  and  a39397a );
 a39401a <=( (not A268)  and  (not A267) );
 a39404a <=( A300  and  A298 );
 a39405a <=( a39404a  and  a39401a );
 a39406a <=( a39405a  and  a39398a );
 a39410a <=( (not A201)  and  A167 );
 a39411a <=( A168  and  a39410a );
 a39414a <=( (not A203)  and  (not A202) );
 a39417a <=( (not A233)  and  (not A232) );
 a39418a <=( a39417a  and  a39414a );
 a39419a <=( a39418a  and  a39411a );
 a39423a <=( (not A266)  and  (not A265) );
 a39424a <=( (not A235)  and  a39423a );
 a39427a <=( A298  and  (not A268) );
 a39430a <=( A302  and  (not A299) );
 a39431a <=( a39430a  and  a39427a );
 a39432a <=( a39431a  and  a39424a );
 a39436a <=( (not A201)  and  A167 );
 a39437a <=( A168  and  a39436a );
 a39440a <=( (not A203)  and  (not A202) );
 a39443a <=( (not A233)  and  (not A232) );
 a39444a <=( a39443a  and  a39440a );
 a39445a <=( a39444a  and  a39437a );
 a39449a <=( (not A266)  and  (not A265) );
 a39450a <=( (not A235)  and  a39449a );
 a39453a <=( (not A298)  and  (not A268) );
 a39456a <=( A302  and  A299 );
 a39457a <=( a39456a  and  a39453a );
 a39458a <=( a39457a  and  a39450a );
 a39462a <=( A199  and  A167 );
 a39463a <=( A168  and  a39462a );
 a39466a <=( (not A201)  and  A200 );
 a39469a <=( (not A234)  and  (not A202) );
 a39470a <=( a39469a  and  a39466a );
 a39471a <=( a39470a  and  a39463a );
 a39475a <=( (not A267)  and  (not A236) );
 a39476a <=( (not A235)  and  a39475a );
 a39479a <=( (not A269)  and  (not A268) );
 a39482a <=( A300  and  A299 );
 a39483a <=( a39482a  and  a39479a );
 a39484a <=( a39483a  and  a39476a );
 a39488a <=( A199  and  A167 );
 a39489a <=( A168  and  a39488a );
 a39492a <=( (not A201)  and  A200 );
 a39495a <=( (not A234)  and  (not A202) );
 a39496a <=( a39495a  and  a39492a );
 a39497a <=( a39496a  and  a39489a );
 a39501a <=( (not A267)  and  (not A236) );
 a39502a <=( (not A235)  and  a39501a );
 a39505a <=( (not A269)  and  (not A268) );
 a39508a <=( A300  and  A298 );
 a39509a <=( a39508a  and  a39505a );
 a39510a <=( a39509a  and  a39502a );
 a39514a <=( A199  and  A167 );
 a39515a <=( A168  and  a39514a );
 a39518a <=( (not A201)  and  A200 );
 a39521a <=( (not A234)  and  (not A202) );
 a39522a <=( a39521a  and  a39518a );
 a39523a <=( a39522a  and  a39515a );
 a39527a <=( A265  and  (not A236) );
 a39528a <=( (not A235)  and  a39527a );
 a39531a <=( (not A267)  and  A266 );
 a39534a <=( A301  and  (not A268) );
 a39535a <=( a39534a  and  a39531a );
 a39536a <=( a39535a  and  a39528a );
 a39540a <=( A199  and  A167 );
 a39541a <=( A168  and  a39540a );
 a39544a <=( (not A201)  and  A200 );
 a39547a <=( (not A234)  and  (not A202) );
 a39548a <=( a39547a  and  a39544a );
 a39549a <=( a39548a  and  a39541a );
 a39553a <=( (not A265)  and  (not A236) );
 a39554a <=( (not A235)  and  a39553a );
 a39557a <=( (not A268)  and  (not A266) );
 a39560a <=( A300  and  A299 );
 a39561a <=( a39560a  and  a39557a );
 a39562a <=( a39561a  and  a39554a );
 a39566a <=( A199  and  A167 );
 a39567a <=( A168  and  a39566a );
 a39570a <=( (not A201)  and  A200 );
 a39573a <=( (not A234)  and  (not A202) );
 a39574a <=( a39573a  and  a39570a );
 a39575a <=( a39574a  and  a39567a );
 a39579a <=( (not A265)  and  (not A236) );
 a39580a <=( (not A235)  and  a39579a );
 a39583a <=( (not A268)  and  (not A266) );
 a39586a <=( A300  and  A298 );
 a39587a <=( a39586a  and  a39583a );
 a39588a <=( a39587a  and  a39580a );
 a39592a <=( A199  and  A167 );
 a39593a <=( A168  and  a39592a );
 a39596a <=( (not A201)  and  A200 );
 a39599a <=( A232  and  (not A202) );
 a39600a <=( a39599a  and  a39596a );
 a39601a <=( a39600a  and  a39593a );
 a39605a <=( (not A235)  and  (not A234) );
 a39606a <=( A233  and  a39605a );
 a39609a <=( (not A268)  and  (not A267) );
 a39612a <=( A301  and  (not A269) );
 a39613a <=( a39612a  and  a39609a );
 a39614a <=( a39613a  and  a39606a );
 a39618a <=( A199  and  A167 );
 a39619a <=( A168  and  a39618a );
 a39622a <=( (not A201)  and  A200 );
 a39625a <=( A232  and  (not A202) );
 a39626a <=( a39625a  and  a39622a );
 a39627a <=( a39626a  and  a39619a );
 a39631a <=( (not A235)  and  (not A234) );
 a39632a <=( A233  and  a39631a );
 a39635a <=( (not A266)  and  (not A265) );
 a39638a <=( A301  and  (not A268) );
 a39639a <=( a39638a  and  a39635a );
 a39640a <=( a39639a  and  a39632a );
 a39644a <=( A199  and  A167 );
 a39645a <=( A168  and  a39644a );
 a39648a <=( (not A201)  and  A200 );
 a39651a <=( (not A232)  and  (not A202) );
 a39652a <=( a39651a  and  a39648a );
 a39653a <=( a39652a  and  a39645a );
 a39657a <=( (not A267)  and  (not A235) );
 a39658a <=( (not A233)  and  a39657a );
 a39661a <=( (not A269)  and  (not A268) );
 a39664a <=( A300  and  A299 );
 a39665a <=( a39664a  and  a39661a );
 a39666a <=( a39665a  and  a39658a );
 a39670a <=( A199  and  A167 );
 a39671a <=( A168  and  a39670a );
 a39674a <=( (not A201)  and  A200 );
 a39677a <=( (not A232)  and  (not A202) );
 a39678a <=( a39677a  and  a39674a );
 a39679a <=( a39678a  and  a39671a );
 a39683a <=( (not A267)  and  (not A235) );
 a39684a <=( (not A233)  and  a39683a );
 a39687a <=( (not A269)  and  (not A268) );
 a39690a <=( A300  and  A298 );
 a39691a <=( a39690a  and  a39687a );
 a39692a <=( a39691a  and  a39684a );
 a39696a <=( A199  and  A167 );
 a39697a <=( A168  and  a39696a );
 a39700a <=( (not A201)  and  A200 );
 a39703a <=( (not A232)  and  (not A202) );
 a39704a <=( a39703a  and  a39700a );
 a39705a <=( a39704a  and  a39697a );
 a39709a <=( A265  and  (not A235) );
 a39710a <=( (not A233)  and  a39709a );
 a39713a <=( (not A267)  and  A266 );
 a39716a <=( A301  and  (not A268) );
 a39717a <=( a39716a  and  a39713a );
 a39718a <=( a39717a  and  a39710a );
 a39722a <=( A199  and  A167 );
 a39723a <=( A168  and  a39722a );
 a39726a <=( (not A201)  and  A200 );
 a39729a <=( (not A232)  and  (not A202) );
 a39730a <=( a39729a  and  a39726a );
 a39731a <=( a39730a  and  a39723a );
 a39735a <=( (not A265)  and  (not A235) );
 a39736a <=( (not A233)  and  a39735a );
 a39739a <=( (not A268)  and  (not A266) );
 a39742a <=( A300  and  A299 );
 a39743a <=( a39742a  and  a39739a );
 a39744a <=( a39743a  and  a39736a );
 a39748a <=( A199  and  A167 );
 a39749a <=( A168  and  a39748a );
 a39752a <=( (not A201)  and  A200 );
 a39755a <=( (not A232)  and  (not A202) );
 a39756a <=( a39755a  and  a39752a );
 a39757a <=( a39756a  and  a39749a );
 a39761a <=( (not A265)  and  (not A235) );
 a39762a <=( (not A233)  and  a39761a );
 a39765a <=( (not A268)  and  (not A266) );
 a39768a <=( A300  and  A298 );
 a39769a <=( a39768a  and  a39765a );
 a39770a <=( a39769a  and  a39762a );
 a39774a <=( (not A199)  and  A167 );
 a39775a <=( A168  and  a39774a );
 a39778a <=( (not A202)  and  (not A200) );
 a39781a <=( (not A235)  and  (not A234) );
 a39782a <=( a39781a  and  a39778a );
 a39783a <=( a39782a  and  a39775a );
 a39787a <=( (not A268)  and  (not A267) );
 a39788a <=( (not A236)  and  a39787a );
 a39791a <=( A298  and  (not A269) );
 a39794a <=( A302  and  (not A299) );
 a39795a <=( a39794a  and  a39791a );
 a39796a <=( a39795a  and  a39788a );
 a39800a <=( (not A199)  and  A167 );
 a39801a <=( A168  and  a39800a );
 a39804a <=( (not A202)  and  (not A200) );
 a39807a <=( (not A235)  and  (not A234) );
 a39808a <=( a39807a  and  a39804a );
 a39809a <=( a39808a  and  a39801a );
 a39813a <=( (not A268)  and  (not A267) );
 a39814a <=( (not A236)  and  a39813a );
 a39817a <=( (not A298)  and  (not A269) );
 a39820a <=( A302  and  A299 );
 a39821a <=( a39820a  and  a39817a );
 a39822a <=( a39821a  and  a39814a );
 a39826a <=( (not A199)  and  A167 );
 a39827a <=( A168  and  a39826a );
 a39830a <=( (not A202)  and  (not A200) );
 a39833a <=( (not A235)  and  (not A234) );
 a39834a <=( a39833a  and  a39830a );
 a39835a <=( a39834a  and  a39827a );
 a39839a <=( A266  and  A265 );
 a39840a <=( (not A236)  and  a39839a );
 a39843a <=( (not A268)  and  (not A267) );
 a39846a <=( A300  and  A299 );
 a39847a <=( a39846a  and  a39843a );
 a39848a <=( a39847a  and  a39840a );
 a39852a <=( (not A199)  and  A167 );
 a39853a <=( A168  and  a39852a );
 a39856a <=( (not A202)  and  (not A200) );
 a39859a <=( (not A235)  and  (not A234) );
 a39860a <=( a39859a  and  a39856a );
 a39861a <=( a39860a  and  a39853a );
 a39865a <=( A266  and  A265 );
 a39866a <=( (not A236)  and  a39865a );
 a39869a <=( (not A268)  and  (not A267) );
 a39872a <=( A300  and  A298 );
 a39873a <=( a39872a  and  a39869a );
 a39874a <=( a39873a  and  a39866a );
 a39878a <=( (not A199)  and  A167 );
 a39879a <=( A168  and  a39878a );
 a39882a <=( (not A202)  and  (not A200) );
 a39885a <=( (not A235)  and  (not A234) );
 a39886a <=( a39885a  and  a39882a );
 a39887a <=( a39886a  and  a39879a );
 a39891a <=( (not A266)  and  (not A265) );
 a39892a <=( (not A236)  and  a39891a );
 a39895a <=( A298  and  (not A268) );
 a39898a <=( A302  and  (not A299) );
 a39899a <=( a39898a  and  a39895a );
 a39900a <=( a39899a  and  a39892a );
 a39904a <=( (not A199)  and  A167 );
 a39905a <=( A168  and  a39904a );
 a39908a <=( (not A202)  and  (not A200) );
 a39911a <=( (not A235)  and  (not A234) );
 a39912a <=( a39911a  and  a39908a );
 a39913a <=( a39912a  and  a39905a );
 a39917a <=( (not A266)  and  (not A265) );
 a39918a <=( (not A236)  and  a39917a );
 a39921a <=( (not A298)  and  (not A268) );
 a39924a <=( A302  and  A299 );
 a39925a <=( a39924a  and  a39921a );
 a39926a <=( a39925a  and  a39918a );
 a39930a <=( (not A199)  and  A167 );
 a39931a <=( A168  and  a39930a );
 a39934a <=( (not A202)  and  (not A200) );
 a39937a <=( A233  and  A232 );
 a39938a <=( a39937a  and  a39934a );
 a39939a <=( a39938a  and  a39931a );
 a39943a <=( (not A267)  and  (not A235) );
 a39944a <=( (not A234)  and  a39943a );
 a39947a <=( (not A269)  and  (not A268) );
 a39950a <=( A300  and  A299 );
 a39951a <=( a39950a  and  a39947a );
 a39952a <=( a39951a  and  a39944a );
 a39956a <=( (not A199)  and  A167 );
 a39957a <=( A168  and  a39956a );
 a39960a <=( (not A202)  and  (not A200) );
 a39963a <=( A233  and  A232 );
 a39964a <=( a39963a  and  a39960a );
 a39965a <=( a39964a  and  a39957a );
 a39969a <=( (not A267)  and  (not A235) );
 a39970a <=( (not A234)  and  a39969a );
 a39973a <=( (not A269)  and  (not A268) );
 a39976a <=( A300  and  A298 );
 a39977a <=( a39976a  and  a39973a );
 a39978a <=( a39977a  and  a39970a );
 a39982a <=( (not A199)  and  A167 );
 a39983a <=( A168  and  a39982a );
 a39986a <=( (not A202)  and  (not A200) );
 a39989a <=( A233  and  A232 );
 a39990a <=( a39989a  and  a39986a );
 a39991a <=( a39990a  and  a39983a );
 a39995a <=( A265  and  (not A235) );
 a39996a <=( (not A234)  and  a39995a );
 a39999a <=( (not A267)  and  A266 );
 a40002a <=( A301  and  (not A268) );
 a40003a <=( a40002a  and  a39999a );
 a40004a <=( a40003a  and  a39996a );
 a40008a <=( (not A199)  and  A167 );
 a40009a <=( A168  and  a40008a );
 a40012a <=( (not A202)  and  (not A200) );
 a40015a <=( A233  and  A232 );
 a40016a <=( a40015a  and  a40012a );
 a40017a <=( a40016a  and  a40009a );
 a40021a <=( (not A265)  and  (not A235) );
 a40022a <=( (not A234)  and  a40021a );
 a40025a <=( (not A268)  and  (not A266) );
 a40028a <=( A300  and  A299 );
 a40029a <=( a40028a  and  a40025a );
 a40030a <=( a40029a  and  a40022a );
 a40034a <=( (not A199)  and  A167 );
 a40035a <=( A168  and  a40034a );
 a40038a <=( (not A202)  and  (not A200) );
 a40041a <=( A233  and  A232 );
 a40042a <=( a40041a  and  a40038a );
 a40043a <=( a40042a  and  a40035a );
 a40047a <=( (not A265)  and  (not A235) );
 a40048a <=( (not A234)  and  a40047a );
 a40051a <=( (not A268)  and  (not A266) );
 a40054a <=( A300  and  A298 );
 a40055a <=( a40054a  and  a40051a );
 a40056a <=( a40055a  and  a40048a );
 a40060a <=( (not A199)  and  A167 );
 a40061a <=( A168  and  a40060a );
 a40064a <=( (not A202)  and  (not A200) );
 a40067a <=( (not A233)  and  (not A232) );
 a40068a <=( a40067a  and  a40064a );
 a40069a <=( a40068a  and  a40061a );
 a40073a <=( (not A268)  and  (not A267) );
 a40074a <=( (not A235)  and  a40073a );
 a40077a <=( A298  and  (not A269) );
 a40080a <=( A302  and  (not A299) );
 a40081a <=( a40080a  and  a40077a );
 a40082a <=( a40081a  and  a40074a );
 a40086a <=( (not A199)  and  A167 );
 a40087a <=( A168  and  a40086a );
 a40090a <=( (not A202)  and  (not A200) );
 a40093a <=( (not A233)  and  (not A232) );
 a40094a <=( a40093a  and  a40090a );
 a40095a <=( a40094a  and  a40087a );
 a40099a <=( (not A268)  and  (not A267) );
 a40100a <=( (not A235)  and  a40099a );
 a40103a <=( (not A298)  and  (not A269) );
 a40106a <=( A302  and  A299 );
 a40107a <=( a40106a  and  a40103a );
 a40108a <=( a40107a  and  a40100a );
 a40112a <=( (not A199)  and  A167 );
 a40113a <=( A168  and  a40112a );
 a40116a <=( (not A202)  and  (not A200) );
 a40119a <=( (not A233)  and  (not A232) );
 a40120a <=( a40119a  and  a40116a );
 a40121a <=( a40120a  and  a40113a );
 a40125a <=( A266  and  A265 );
 a40126a <=( (not A235)  and  a40125a );
 a40129a <=( (not A268)  and  (not A267) );
 a40132a <=( A300  and  A299 );
 a40133a <=( a40132a  and  a40129a );
 a40134a <=( a40133a  and  a40126a );
 a40138a <=( (not A199)  and  A167 );
 a40139a <=( A168  and  a40138a );
 a40142a <=( (not A202)  and  (not A200) );
 a40145a <=( (not A233)  and  (not A232) );
 a40146a <=( a40145a  and  a40142a );
 a40147a <=( a40146a  and  a40139a );
 a40151a <=( A266  and  A265 );
 a40152a <=( (not A235)  and  a40151a );
 a40155a <=( (not A268)  and  (not A267) );
 a40158a <=( A300  and  A298 );
 a40159a <=( a40158a  and  a40155a );
 a40160a <=( a40159a  and  a40152a );
 a40164a <=( (not A199)  and  A167 );
 a40165a <=( A168  and  a40164a );
 a40168a <=( (not A202)  and  (not A200) );
 a40171a <=( (not A233)  and  (not A232) );
 a40172a <=( a40171a  and  a40168a );
 a40173a <=( a40172a  and  a40165a );
 a40177a <=( (not A266)  and  (not A265) );
 a40178a <=( (not A235)  and  a40177a );
 a40181a <=( A298  and  (not A268) );
 a40184a <=( A302  and  (not A299) );
 a40185a <=( a40184a  and  a40181a );
 a40186a <=( a40185a  and  a40178a );
 a40190a <=( (not A199)  and  A167 );
 a40191a <=( A168  and  a40190a );
 a40194a <=( (not A202)  and  (not A200) );
 a40197a <=( (not A233)  and  (not A232) );
 a40198a <=( a40197a  and  a40194a );
 a40199a <=( a40198a  and  a40191a );
 a40203a <=( (not A266)  and  (not A265) );
 a40204a <=( (not A235)  and  a40203a );
 a40207a <=( (not A298)  and  (not A268) );
 a40210a <=( A302  and  A299 );
 a40211a <=( a40210a  and  a40207a );
 a40212a <=( a40211a  and  a40204a );
 a40216a <=( (not A166)  and  A167 );
 a40217a <=( A170  and  a40216a );
 a40220a <=( (not A202)  and  (not A201) );
 a40223a <=( (not A234)  and  (not A203) );
 a40224a <=( a40223a  and  a40220a );
 a40225a <=( a40224a  and  a40217a );
 a40229a <=( (not A267)  and  (not A236) );
 a40230a <=( (not A235)  and  a40229a );
 a40233a <=( (not A269)  and  (not A268) );
 a40236a <=( A300  and  A299 );
 a40237a <=( a40236a  and  a40233a );
 a40238a <=( a40237a  and  a40230a );
 a40242a <=( (not A166)  and  A167 );
 a40243a <=( A170  and  a40242a );
 a40246a <=( (not A202)  and  (not A201) );
 a40249a <=( (not A234)  and  (not A203) );
 a40250a <=( a40249a  and  a40246a );
 a40251a <=( a40250a  and  a40243a );
 a40255a <=( (not A267)  and  (not A236) );
 a40256a <=( (not A235)  and  a40255a );
 a40259a <=( (not A269)  and  (not A268) );
 a40262a <=( A300  and  A298 );
 a40263a <=( a40262a  and  a40259a );
 a40264a <=( a40263a  and  a40256a );
 a40268a <=( (not A166)  and  A167 );
 a40269a <=( A170  and  a40268a );
 a40272a <=( (not A202)  and  (not A201) );
 a40275a <=( (not A234)  and  (not A203) );
 a40276a <=( a40275a  and  a40272a );
 a40277a <=( a40276a  and  a40269a );
 a40281a <=( A265  and  (not A236) );
 a40282a <=( (not A235)  and  a40281a );
 a40285a <=( (not A267)  and  A266 );
 a40288a <=( A301  and  (not A268) );
 a40289a <=( a40288a  and  a40285a );
 a40290a <=( a40289a  and  a40282a );
 a40294a <=( (not A166)  and  A167 );
 a40295a <=( A170  and  a40294a );
 a40298a <=( (not A202)  and  (not A201) );
 a40301a <=( (not A234)  and  (not A203) );
 a40302a <=( a40301a  and  a40298a );
 a40303a <=( a40302a  and  a40295a );
 a40307a <=( (not A265)  and  (not A236) );
 a40308a <=( (not A235)  and  a40307a );
 a40311a <=( (not A268)  and  (not A266) );
 a40314a <=( A300  and  A299 );
 a40315a <=( a40314a  and  a40311a );
 a40316a <=( a40315a  and  a40308a );
 a40320a <=( (not A166)  and  A167 );
 a40321a <=( A170  and  a40320a );
 a40324a <=( (not A202)  and  (not A201) );
 a40327a <=( (not A234)  and  (not A203) );
 a40328a <=( a40327a  and  a40324a );
 a40329a <=( a40328a  and  a40321a );
 a40333a <=( (not A265)  and  (not A236) );
 a40334a <=( (not A235)  and  a40333a );
 a40337a <=( (not A268)  and  (not A266) );
 a40340a <=( A300  and  A298 );
 a40341a <=( a40340a  and  a40337a );
 a40342a <=( a40341a  and  a40334a );
 a40346a <=( (not A166)  and  A167 );
 a40347a <=( A170  and  a40346a );
 a40350a <=( (not A202)  and  (not A201) );
 a40353a <=( A232  and  (not A203) );
 a40354a <=( a40353a  and  a40350a );
 a40355a <=( a40354a  and  a40347a );
 a40359a <=( (not A235)  and  (not A234) );
 a40360a <=( A233  and  a40359a );
 a40363a <=( (not A268)  and  (not A267) );
 a40366a <=( A301  and  (not A269) );
 a40367a <=( a40366a  and  a40363a );
 a40368a <=( a40367a  and  a40360a );
 a40372a <=( (not A166)  and  A167 );
 a40373a <=( A170  and  a40372a );
 a40376a <=( (not A202)  and  (not A201) );
 a40379a <=( A232  and  (not A203) );
 a40380a <=( a40379a  and  a40376a );
 a40381a <=( a40380a  and  a40373a );
 a40385a <=( (not A235)  and  (not A234) );
 a40386a <=( A233  and  a40385a );
 a40389a <=( (not A266)  and  (not A265) );
 a40392a <=( A301  and  (not A268) );
 a40393a <=( a40392a  and  a40389a );
 a40394a <=( a40393a  and  a40386a );
 a40398a <=( (not A166)  and  A167 );
 a40399a <=( A170  and  a40398a );
 a40402a <=( (not A202)  and  (not A201) );
 a40405a <=( (not A232)  and  (not A203) );
 a40406a <=( a40405a  and  a40402a );
 a40407a <=( a40406a  and  a40399a );
 a40411a <=( (not A267)  and  (not A235) );
 a40412a <=( (not A233)  and  a40411a );
 a40415a <=( (not A269)  and  (not A268) );
 a40418a <=( A300  and  A299 );
 a40419a <=( a40418a  and  a40415a );
 a40420a <=( a40419a  and  a40412a );
 a40424a <=( (not A166)  and  A167 );
 a40425a <=( A170  and  a40424a );
 a40428a <=( (not A202)  and  (not A201) );
 a40431a <=( (not A232)  and  (not A203) );
 a40432a <=( a40431a  and  a40428a );
 a40433a <=( a40432a  and  a40425a );
 a40437a <=( (not A267)  and  (not A235) );
 a40438a <=( (not A233)  and  a40437a );
 a40441a <=( (not A269)  and  (not A268) );
 a40444a <=( A300  and  A298 );
 a40445a <=( a40444a  and  a40441a );
 a40446a <=( a40445a  and  a40438a );
 a40450a <=( (not A166)  and  A167 );
 a40451a <=( A170  and  a40450a );
 a40454a <=( (not A202)  and  (not A201) );
 a40457a <=( (not A232)  and  (not A203) );
 a40458a <=( a40457a  and  a40454a );
 a40459a <=( a40458a  and  a40451a );
 a40463a <=( A265  and  (not A235) );
 a40464a <=( (not A233)  and  a40463a );
 a40467a <=( (not A267)  and  A266 );
 a40470a <=( A301  and  (not A268) );
 a40471a <=( a40470a  and  a40467a );
 a40472a <=( a40471a  and  a40464a );
 a40476a <=( (not A166)  and  A167 );
 a40477a <=( A170  and  a40476a );
 a40480a <=( (not A202)  and  (not A201) );
 a40483a <=( (not A232)  and  (not A203) );
 a40484a <=( a40483a  and  a40480a );
 a40485a <=( a40484a  and  a40477a );
 a40489a <=( (not A265)  and  (not A235) );
 a40490a <=( (not A233)  and  a40489a );
 a40493a <=( (not A268)  and  (not A266) );
 a40496a <=( A300  and  A299 );
 a40497a <=( a40496a  and  a40493a );
 a40498a <=( a40497a  and  a40490a );
 a40502a <=( (not A166)  and  A167 );
 a40503a <=( A170  and  a40502a );
 a40506a <=( (not A202)  and  (not A201) );
 a40509a <=( (not A232)  and  (not A203) );
 a40510a <=( a40509a  and  a40506a );
 a40511a <=( a40510a  and  a40503a );
 a40515a <=( (not A265)  and  (not A235) );
 a40516a <=( (not A233)  and  a40515a );
 a40519a <=( (not A268)  and  (not A266) );
 a40522a <=( A300  and  A298 );
 a40523a <=( a40522a  and  a40519a );
 a40524a <=( a40523a  and  a40516a );
 a40528a <=( (not A166)  and  A167 );
 a40529a <=( A170  and  a40528a );
 a40532a <=( A200  and  A199 );
 a40535a <=( (not A202)  and  (not A201) );
 a40536a <=( a40535a  and  a40532a );
 a40537a <=( a40536a  and  a40529a );
 a40541a <=( (not A236)  and  (not A235) );
 a40542a <=( (not A234)  and  a40541a );
 a40545a <=( (not A268)  and  (not A267) );
 a40548a <=( A301  and  (not A269) );
 a40549a <=( a40548a  and  a40545a );
 a40550a <=( a40549a  and  a40542a );
 a40554a <=( (not A166)  and  A167 );
 a40555a <=( A170  and  a40554a );
 a40558a <=( A200  and  A199 );
 a40561a <=( (not A202)  and  (not A201) );
 a40562a <=( a40561a  and  a40558a );
 a40563a <=( a40562a  and  a40555a );
 a40567a <=( (not A236)  and  (not A235) );
 a40568a <=( (not A234)  and  a40567a );
 a40571a <=( (not A266)  and  (not A265) );
 a40574a <=( A301  and  (not A268) );
 a40575a <=( a40574a  and  a40571a );
 a40576a <=( a40575a  and  a40568a );
 a40580a <=( (not A166)  and  A167 );
 a40581a <=( A170  and  a40580a );
 a40584a <=( A200  and  A199 );
 a40587a <=( (not A202)  and  (not A201) );
 a40588a <=( a40587a  and  a40584a );
 a40589a <=( a40588a  and  a40581a );
 a40593a <=( A236  and  A233 );
 a40594a <=( (not A232)  and  a40593a );
 a40597a <=( A299  and  A298 );
 a40600a <=( (not A301)  and  (not A300) );
 a40601a <=( a40600a  and  a40597a );
 a40602a <=( a40601a  and  a40594a );
 a40606a <=( (not A166)  and  A167 );
 a40607a <=( A170  and  a40606a );
 a40610a <=( A200  and  A199 );
 a40613a <=( (not A202)  and  (not A201) );
 a40614a <=( a40613a  and  a40610a );
 a40615a <=( a40614a  and  a40607a );
 a40619a <=( A236  and  (not A233) );
 a40620a <=( A232  and  a40619a );
 a40623a <=( A299  and  A298 );
 a40626a <=( (not A301)  and  (not A300) );
 a40627a <=( a40626a  and  a40623a );
 a40628a <=( a40627a  and  a40620a );
 a40632a <=( (not A166)  and  A167 );
 a40633a <=( A170  and  a40632a );
 a40636a <=( A200  and  A199 );
 a40639a <=( (not A202)  and  (not A201) );
 a40640a <=( a40639a  and  a40636a );
 a40641a <=( a40640a  and  a40633a );
 a40645a <=( (not A235)  and  (not A233) );
 a40646a <=( (not A232)  and  a40645a );
 a40649a <=( (not A268)  and  (not A267) );
 a40652a <=( A301  and  (not A269) );
 a40653a <=( a40652a  and  a40649a );
 a40654a <=( a40653a  and  a40646a );
 a40658a <=( (not A166)  and  A167 );
 a40659a <=( A170  and  a40658a );
 a40662a <=( A200  and  A199 );
 a40665a <=( (not A202)  and  (not A201) );
 a40666a <=( a40665a  and  a40662a );
 a40667a <=( a40666a  and  a40659a );
 a40671a <=( (not A235)  and  (not A233) );
 a40672a <=( (not A232)  and  a40671a );
 a40675a <=( (not A266)  and  (not A265) );
 a40678a <=( A301  and  (not A268) );
 a40679a <=( a40678a  and  a40675a );
 a40680a <=( a40679a  and  a40672a );
 a40684a <=( (not A166)  and  A167 );
 a40685a <=( A170  and  a40684a );
 a40688a <=( (not A200)  and  (not A199) );
 a40691a <=( (not A234)  and  (not A202) );
 a40692a <=( a40691a  and  a40688a );
 a40693a <=( a40692a  and  a40685a );
 a40697a <=( (not A267)  and  (not A236) );
 a40698a <=( (not A235)  and  a40697a );
 a40701a <=( (not A269)  and  (not A268) );
 a40704a <=( A300  and  A299 );
 a40705a <=( a40704a  and  a40701a );
 a40706a <=( a40705a  and  a40698a );
 a40710a <=( (not A166)  and  A167 );
 a40711a <=( A170  and  a40710a );
 a40714a <=( (not A200)  and  (not A199) );
 a40717a <=( (not A234)  and  (not A202) );
 a40718a <=( a40717a  and  a40714a );
 a40719a <=( a40718a  and  a40711a );
 a40723a <=( (not A267)  and  (not A236) );
 a40724a <=( (not A235)  and  a40723a );
 a40727a <=( (not A269)  and  (not A268) );
 a40730a <=( A300  and  A298 );
 a40731a <=( a40730a  and  a40727a );
 a40732a <=( a40731a  and  a40724a );
 a40736a <=( (not A166)  and  A167 );
 a40737a <=( A170  and  a40736a );
 a40740a <=( (not A200)  and  (not A199) );
 a40743a <=( (not A234)  and  (not A202) );
 a40744a <=( a40743a  and  a40740a );
 a40745a <=( a40744a  and  a40737a );
 a40749a <=( A265  and  (not A236) );
 a40750a <=( (not A235)  and  a40749a );
 a40753a <=( (not A267)  and  A266 );
 a40756a <=( A301  and  (not A268) );
 a40757a <=( a40756a  and  a40753a );
 a40758a <=( a40757a  and  a40750a );
 a40762a <=( (not A166)  and  A167 );
 a40763a <=( A170  and  a40762a );
 a40766a <=( (not A200)  and  (not A199) );
 a40769a <=( (not A234)  and  (not A202) );
 a40770a <=( a40769a  and  a40766a );
 a40771a <=( a40770a  and  a40763a );
 a40775a <=( (not A265)  and  (not A236) );
 a40776a <=( (not A235)  and  a40775a );
 a40779a <=( (not A268)  and  (not A266) );
 a40782a <=( A300  and  A299 );
 a40783a <=( a40782a  and  a40779a );
 a40784a <=( a40783a  and  a40776a );
 a40788a <=( (not A166)  and  A167 );
 a40789a <=( A170  and  a40788a );
 a40792a <=( (not A200)  and  (not A199) );
 a40795a <=( (not A234)  and  (not A202) );
 a40796a <=( a40795a  and  a40792a );
 a40797a <=( a40796a  and  a40789a );
 a40801a <=( (not A265)  and  (not A236) );
 a40802a <=( (not A235)  and  a40801a );
 a40805a <=( (not A268)  and  (not A266) );
 a40808a <=( A300  and  A298 );
 a40809a <=( a40808a  and  a40805a );
 a40810a <=( a40809a  and  a40802a );
 a40814a <=( (not A166)  and  A167 );
 a40815a <=( A170  and  a40814a );
 a40818a <=( (not A200)  and  (not A199) );
 a40821a <=( A232  and  (not A202) );
 a40822a <=( a40821a  and  a40818a );
 a40823a <=( a40822a  and  a40815a );
 a40827a <=( (not A235)  and  (not A234) );
 a40828a <=( A233  and  a40827a );
 a40831a <=( (not A268)  and  (not A267) );
 a40834a <=( A301  and  (not A269) );
 a40835a <=( a40834a  and  a40831a );
 a40836a <=( a40835a  and  a40828a );
 a40840a <=( (not A166)  and  A167 );
 a40841a <=( A170  and  a40840a );
 a40844a <=( (not A200)  and  (not A199) );
 a40847a <=( A232  and  (not A202) );
 a40848a <=( a40847a  and  a40844a );
 a40849a <=( a40848a  and  a40841a );
 a40853a <=( (not A235)  and  (not A234) );
 a40854a <=( A233  and  a40853a );
 a40857a <=( (not A266)  and  (not A265) );
 a40860a <=( A301  and  (not A268) );
 a40861a <=( a40860a  and  a40857a );
 a40862a <=( a40861a  and  a40854a );
 a40866a <=( (not A166)  and  A167 );
 a40867a <=( A170  and  a40866a );
 a40870a <=( (not A200)  and  (not A199) );
 a40873a <=( (not A232)  and  (not A202) );
 a40874a <=( a40873a  and  a40870a );
 a40875a <=( a40874a  and  a40867a );
 a40879a <=( (not A267)  and  (not A235) );
 a40880a <=( (not A233)  and  a40879a );
 a40883a <=( (not A269)  and  (not A268) );
 a40886a <=( A300  and  A299 );
 a40887a <=( a40886a  and  a40883a );
 a40888a <=( a40887a  and  a40880a );
 a40892a <=( (not A166)  and  A167 );
 a40893a <=( A170  and  a40892a );
 a40896a <=( (not A200)  and  (not A199) );
 a40899a <=( (not A232)  and  (not A202) );
 a40900a <=( a40899a  and  a40896a );
 a40901a <=( a40900a  and  a40893a );
 a40905a <=( (not A267)  and  (not A235) );
 a40906a <=( (not A233)  and  a40905a );
 a40909a <=( (not A269)  and  (not A268) );
 a40912a <=( A300  and  A298 );
 a40913a <=( a40912a  and  a40909a );
 a40914a <=( a40913a  and  a40906a );
 a40918a <=( (not A166)  and  A167 );
 a40919a <=( A170  and  a40918a );
 a40922a <=( (not A200)  and  (not A199) );
 a40925a <=( (not A232)  and  (not A202) );
 a40926a <=( a40925a  and  a40922a );
 a40927a <=( a40926a  and  a40919a );
 a40931a <=( A265  and  (not A235) );
 a40932a <=( (not A233)  and  a40931a );
 a40935a <=( (not A267)  and  A266 );
 a40938a <=( A301  and  (not A268) );
 a40939a <=( a40938a  and  a40935a );
 a40940a <=( a40939a  and  a40932a );
 a40944a <=( (not A166)  and  A167 );
 a40945a <=( A170  and  a40944a );
 a40948a <=( (not A200)  and  (not A199) );
 a40951a <=( (not A232)  and  (not A202) );
 a40952a <=( a40951a  and  a40948a );
 a40953a <=( a40952a  and  a40945a );
 a40957a <=( (not A265)  and  (not A235) );
 a40958a <=( (not A233)  and  a40957a );
 a40961a <=( (not A268)  and  (not A266) );
 a40964a <=( A300  and  A299 );
 a40965a <=( a40964a  and  a40961a );
 a40966a <=( a40965a  and  a40958a );
 a40970a <=( (not A166)  and  A167 );
 a40971a <=( A170  and  a40970a );
 a40974a <=( (not A200)  and  (not A199) );
 a40977a <=( (not A232)  and  (not A202) );
 a40978a <=( a40977a  and  a40974a );
 a40979a <=( a40978a  and  a40971a );
 a40983a <=( (not A265)  and  (not A235) );
 a40984a <=( (not A233)  and  a40983a );
 a40987a <=( (not A268)  and  (not A266) );
 a40990a <=( A300  and  A298 );
 a40991a <=( a40990a  and  a40987a );
 a40992a <=( a40991a  and  a40984a );
 a40996a <=( A166  and  (not A167) );
 a40997a <=( A170  and  a40996a );
 a41000a <=( (not A202)  and  (not A201) );
 a41003a <=( (not A234)  and  (not A203) );
 a41004a <=( a41003a  and  a41000a );
 a41005a <=( a41004a  and  a40997a );
 a41009a <=( (not A267)  and  (not A236) );
 a41010a <=( (not A235)  and  a41009a );
 a41013a <=( (not A269)  and  (not A268) );
 a41016a <=( A300  and  A299 );
 a41017a <=( a41016a  and  a41013a );
 a41018a <=( a41017a  and  a41010a );
 a41022a <=( A166  and  (not A167) );
 a41023a <=( A170  and  a41022a );
 a41026a <=( (not A202)  and  (not A201) );
 a41029a <=( (not A234)  and  (not A203) );
 a41030a <=( a41029a  and  a41026a );
 a41031a <=( a41030a  and  a41023a );
 a41035a <=( (not A267)  and  (not A236) );
 a41036a <=( (not A235)  and  a41035a );
 a41039a <=( (not A269)  and  (not A268) );
 a41042a <=( A300  and  A298 );
 a41043a <=( a41042a  and  a41039a );
 a41044a <=( a41043a  and  a41036a );
 a41048a <=( A166  and  (not A167) );
 a41049a <=( A170  and  a41048a );
 a41052a <=( (not A202)  and  (not A201) );
 a41055a <=( (not A234)  and  (not A203) );
 a41056a <=( a41055a  and  a41052a );
 a41057a <=( a41056a  and  a41049a );
 a41061a <=( A265  and  (not A236) );
 a41062a <=( (not A235)  and  a41061a );
 a41065a <=( (not A267)  and  A266 );
 a41068a <=( A301  and  (not A268) );
 a41069a <=( a41068a  and  a41065a );
 a41070a <=( a41069a  and  a41062a );
 a41074a <=( A166  and  (not A167) );
 a41075a <=( A170  and  a41074a );
 a41078a <=( (not A202)  and  (not A201) );
 a41081a <=( (not A234)  and  (not A203) );
 a41082a <=( a41081a  and  a41078a );
 a41083a <=( a41082a  and  a41075a );
 a41087a <=( (not A265)  and  (not A236) );
 a41088a <=( (not A235)  and  a41087a );
 a41091a <=( (not A268)  and  (not A266) );
 a41094a <=( A300  and  A299 );
 a41095a <=( a41094a  and  a41091a );
 a41096a <=( a41095a  and  a41088a );
 a41100a <=( A166  and  (not A167) );
 a41101a <=( A170  and  a41100a );
 a41104a <=( (not A202)  and  (not A201) );
 a41107a <=( (not A234)  and  (not A203) );
 a41108a <=( a41107a  and  a41104a );
 a41109a <=( a41108a  and  a41101a );
 a41113a <=( (not A265)  and  (not A236) );
 a41114a <=( (not A235)  and  a41113a );
 a41117a <=( (not A268)  and  (not A266) );
 a41120a <=( A300  and  A298 );
 a41121a <=( a41120a  and  a41117a );
 a41122a <=( a41121a  and  a41114a );
 a41126a <=( A166  and  (not A167) );
 a41127a <=( A170  and  a41126a );
 a41130a <=( (not A202)  and  (not A201) );
 a41133a <=( A232  and  (not A203) );
 a41134a <=( a41133a  and  a41130a );
 a41135a <=( a41134a  and  a41127a );
 a41139a <=( (not A235)  and  (not A234) );
 a41140a <=( A233  and  a41139a );
 a41143a <=( (not A268)  and  (not A267) );
 a41146a <=( A301  and  (not A269) );
 a41147a <=( a41146a  and  a41143a );
 a41148a <=( a41147a  and  a41140a );
 a41152a <=( A166  and  (not A167) );
 a41153a <=( A170  and  a41152a );
 a41156a <=( (not A202)  and  (not A201) );
 a41159a <=( A232  and  (not A203) );
 a41160a <=( a41159a  and  a41156a );
 a41161a <=( a41160a  and  a41153a );
 a41165a <=( (not A235)  and  (not A234) );
 a41166a <=( A233  and  a41165a );
 a41169a <=( (not A266)  and  (not A265) );
 a41172a <=( A301  and  (not A268) );
 a41173a <=( a41172a  and  a41169a );
 a41174a <=( a41173a  and  a41166a );
 a41178a <=( A166  and  (not A167) );
 a41179a <=( A170  and  a41178a );
 a41182a <=( (not A202)  and  (not A201) );
 a41185a <=( (not A232)  and  (not A203) );
 a41186a <=( a41185a  and  a41182a );
 a41187a <=( a41186a  and  a41179a );
 a41191a <=( (not A267)  and  (not A235) );
 a41192a <=( (not A233)  and  a41191a );
 a41195a <=( (not A269)  and  (not A268) );
 a41198a <=( A300  and  A299 );
 a41199a <=( a41198a  and  a41195a );
 a41200a <=( a41199a  and  a41192a );
 a41204a <=( A166  and  (not A167) );
 a41205a <=( A170  and  a41204a );
 a41208a <=( (not A202)  and  (not A201) );
 a41211a <=( (not A232)  and  (not A203) );
 a41212a <=( a41211a  and  a41208a );
 a41213a <=( a41212a  and  a41205a );
 a41217a <=( (not A267)  and  (not A235) );
 a41218a <=( (not A233)  and  a41217a );
 a41221a <=( (not A269)  and  (not A268) );
 a41224a <=( A300  and  A298 );
 a41225a <=( a41224a  and  a41221a );
 a41226a <=( a41225a  and  a41218a );
 a41230a <=( A166  and  (not A167) );
 a41231a <=( A170  and  a41230a );
 a41234a <=( (not A202)  and  (not A201) );
 a41237a <=( (not A232)  and  (not A203) );
 a41238a <=( a41237a  and  a41234a );
 a41239a <=( a41238a  and  a41231a );
 a41243a <=( A265  and  (not A235) );
 a41244a <=( (not A233)  and  a41243a );
 a41247a <=( (not A267)  and  A266 );
 a41250a <=( A301  and  (not A268) );
 a41251a <=( a41250a  and  a41247a );
 a41252a <=( a41251a  and  a41244a );
 a41256a <=( A166  and  (not A167) );
 a41257a <=( A170  and  a41256a );
 a41260a <=( (not A202)  and  (not A201) );
 a41263a <=( (not A232)  and  (not A203) );
 a41264a <=( a41263a  and  a41260a );
 a41265a <=( a41264a  and  a41257a );
 a41269a <=( (not A265)  and  (not A235) );
 a41270a <=( (not A233)  and  a41269a );
 a41273a <=( (not A268)  and  (not A266) );
 a41276a <=( A300  and  A299 );
 a41277a <=( a41276a  and  a41273a );
 a41278a <=( a41277a  and  a41270a );
 a41282a <=( A166  and  (not A167) );
 a41283a <=( A170  and  a41282a );
 a41286a <=( (not A202)  and  (not A201) );
 a41289a <=( (not A232)  and  (not A203) );
 a41290a <=( a41289a  and  a41286a );
 a41291a <=( a41290a  and  a41283a );
 a41295a <=( (not A265)  and  (not A235) );
 a41296a <=( (not A233)  and  a41295a );
 a41299a <=( (not A268)  and  (not A266) );
 a41302a <=( A300  and  A298 );
 a41303a <=( a41302a  and  a41299a );
 a41304a <=( a41303a  and  a41296a );
 a41308a <=( A166  and  (not A167) );
 a41309a <=( A170  and  a41308a );
 a41312a <=( A200  and  A199 );
 a41315a <=( (not A202)  and  (not A201) );
 a41316a <=( a41315a  and  a41312a );
 a41317a <=( a41316a  and  a41309a );
 a41321a <=( (not A236)  and  (not A235) );
 a41322a <=( (not A234)  and  a41321a );
 a41325a <=( (not A268)  and  (not A267) );
 a41328a <=( A301  and  (not A269) );
 a41329a <=( a41328a  and  a41325a );
 a41330a <=( a41329a  and  a41322a );
 a41334a <=( A166  and  (not A167) );
 a41335a <=( A170  and  a41334a );
 a41338a <=( A200  and  A199 );
 a41341a <=( (not A202)  and  (not A201) );
 a41342a <=( a41341a  and  a41338a );
 a41343a <=( a41342a  and  a41335a );
 a41347a <=( (not A236)  and  (not A235) );
 a41348a <=( (not A234)  and  a41347a );
 a41351a <=( (not A266)  and  (not A265) );
 a41354a <=( A301  and  (not A268) );
 a41355a <=( a41354a  and  a41351a );
 a41356a <=( a41355a  and  a41348a );
 a41360a <=( A166  and  (not A167) );
 a41361a <=( A170  and  a41360a );
 a41364a <=( A200  and  A199 );
 a41367a <=( (not A202)  and  (not A201) );
 a41368a <=( a41367a  and  a41364a );
 a41369a <=( a41368a  and  a41361a );
 a41373a <=( A236  and  A233 );
 a41374a <=( (not A232)  and  a41373a );
 a41377a <=( A299  and  A298 );
 a41380a <=( (not A301)  and  (not A300) );
 a41381a <=( a41380a  and  a41377a );
 a41382a <=( a41381a  and  a41374a );
 a41386a <=( A166  and  (not A167) );
 a41387a <=( A170  and  a41386a );
 a41390a <=( A200  and  A199 );
 a41393a <=( (not A202)  and  (not A201) );
 a41394a <=( a41393a  and  a41390a );
 a41395a <=( a41394a  and  a41387a );
 a41399a <=( A236  and  (not A233) );
 a41400a <=( A232  and  a41399a );
 a41403a <=( A299  and  A298 );
 a41406a <=( (not A301)  and  (not A300) );
 a41407a <=( a41406a  and  a41403a );
 a41408a <=( a41407a  and  a41400a );
 a41412a <=( A166  and  (not A167) );
 a41413a <=( A170  and  a41412a );
 a41416a <=( A200  and  A199 );
 a41419a <=( (not A202)  and  (not A201) );
 a41420a <=( a41419a  and  a41416a );
 a41421a <=( a41420a  and  a41413a );
 a41425a <=( (not A235)  and  (not A233) );
 a41426a <=( (not A232)  and  a41425a );
 a41429a <=( (not A268)  and  (not A267) );
 a41432a <=( A301  and  (not A269) );
 a41433a <=( a41432a  and  a41429a );
 a41434a <=( a41433a  and  a41426a );
 a41438a <=( A166  and  (not A167) );
 a41439a <=( A170  and  a41438a );
 a41442a <=( A200  and  A199 );
 a41445a <=( (not A202)  and  (not A201) );
 a41446a <=( a41445a  and  a41442a );
 a41447a <=( a41446a  and  a41439a );
 a41451a <=( (not A235)  and  (not A233) );
 a41452a <=( (not A232)  and  a41451a );
 a41455a <=( (not A266)  and  (not A265) );
 a41458a <=( A301  and  (not A268) );
 a41459a <=( a41458a  and  a41455a );
 a41460a <=( a41459a  and  a41452a );
 a41464a <=( A166  and  (not A167) );
 a41465a <=( A170  and  a41464a );
 a41468a <=( (not A200)  and  (not A199) );
 a41471a <=( (not A234)  and  (not A202) );
 a41472a <=( a41471a  and  a41468a );
 a41473a <=( a41472a  and  a41465a );
 a41477a <=( (not A267)  and  (not A236) );
 a41478a <=( (not A235)  and  a41477a );
 a41481a <=( (not A269)  and  (not A268) );
 a41484a <=( A300  and  A299 );
 a41485a <=( a41484a  and  a41481a );
 a41486a <=( a41485a  and  a41478a );
 a41490a <=( A166  and  (not A167) );
 a41491a <=( A170  and  a41490a );
 a41494a <=( (not A200)  and  (not A199) );
 a41497a <=( (not A234)  and  (not A202) );
 a41498a <=( a41497a  and  a41494a );
 a41499a <=( a41498a  and  a41491a );
 a41503a <=( (not A267)  and  (not A236) );
 a41504a <=( (not A235)  and  a41503a );
 a41507a <=( (not A269)  and  (not A268) );
 a41510a <=( A300  and  A298 );
 a41511a <=( a41510a  and  a41507a );
 a41512a <=( a41511a  and  a41504a );
 a41516a <=( A166  and  (not A167) );
 a41517a <=( A170  and  a41516a );
 a41520a <=( (not A200)  and  (not A199) );
 a41523a <=( (not A234)  and  (not A202) );
 a41524a <=( a41523a  and  a41520a );
 a41525a <=( a41524a  and  a41517a );
 a41529a <=( A265  and  (not A236) );
 a41530a <=( (not A235)  and  a41529a );
 a41533a <=( (not A267)  and  A266 );
 a41536a <=( A301  and  (not A268) );
 a41537a <=( a41536a  and  a41533a );
 a41538a <=( a41537a  and  a41530a );
 a41542a <=( A166  and  (not A167) );
 a41543a <=( A170  and  a41542a );
 a41546a <=( (not A200)  and  (not A199) );
 a41549a <=( (not A234)  and  (not A202) );
 a41550a <=( a41549a  and  a41546a );
 a41551a <=( a41550a  and  a41543a );
 a41555a <=( (not A265)  and  (not A236) );
 a41556a <=( (not A235)  and  a41555a );
 a41559a <=( (not A268)  and  (not A266) );
 a41562a <=( A300  and  A299 );
 a41563a <=( a41562a  and  a41559a );
 a41564a <=( a41563a  and  a41556a );
 a41568a <=( A166  and  (not A167) );
 a41569a <=( A170  and  a41568a );
 a41572a <=( (not A200)  and  (not A199) );
 a41575a <=( (not A234)  and  (not A202) );
 a41576a <=( a41575a  and  a41572a );
 a41577a <=( a41576a  and  a41569a );
 a41581a <=( (not A265)  and  (not A236) );
 a41582a <=( (not A235)  and  a41581a );
 a41585a <=( (not A268)  and  (not A266) );
 a41588a <=( A300  and  A298 );
 a41589a <=( a41588a  and  a41585a );
 a41590a <=( a41589a  and  a41582a );
 a41594a <=( A166  and  (not A167) );
 a41595a <=( A170  and  a41594a );
 a41598a <=( (not A200)  and  (not A199) );
 a41601a <=( A232  and  (not A202) );
 a41602a <=( a41601a  and  a41598a );
 a41603a <=( a41602a  and  a41595a );
 a41607a <=( (not A235)  and  (not A234) );
 a41608a <=( A233  and  a41607a );
 a41611a <=( (not A268)  and  (not A267) );
 a41614a <=( A301  and  (not A269) );
 a41615a <=( a41614a  and  a41611a );
 a41616a <=( a41615a  and  a41608a );
 a41620a <=( A166  and  (not A167) );
 a41621a <=( A170  and  a41620a );
 a41624a <=( (not A200)  and  (not A199) );
 a41627a <=( A232  and  (not A202) );
 a41628a <=( a41627a  and  a41624a );
 a41629a <=( a41628a  and  a41621a );
 a41633a <=( (not A235)  and  (not A234) );
 a41634a <=( A233  and  a41633a );
 a41637a <=( (not A266)  and  (not A265) );
 a41640a <=( A301  and  (not A268) );
 a41641a <=( a41640a  and  a41637a );
 a41642a <=( a41641a  and  a41634a );
 a41646a <=( A166  and  (not A167) );
 a41647a <=( A170  and  a41646a );
 a41650a <=( (not A200)  and  (not A199) );
 a41653a <=( (not A232)  and  (not A202) );
 a41654a <=( a41653a  and  a41650a );
 a41655a <=( a41654a  and  a41647a );
 a41659a <=( (not A267)  and  (not A235) );
 a41660a <=( (not A233)  and  a41659a );
 a41663a <=( (not A269)  and  (not A268) );
 a41666a <=( A300  and  A299 );
 a41667a <=( a41666a  and  a41663a );
 a41668a <=( a41667a  and  a41660a );
 a41672a <=( A166  and  (not A167) );
 a41673a <=( A170  and  a41672a );
 a41676a <=( (not A200)  and  (not A199) );
 a41679a <=( (not A232)  and  (not A202) );
 a41680a <=( a41679a  and  a41676a );
 a41681a <=( a41680a  and  a41673a );
 a41685a <=( (not A267)  and  (not A235) );
 a41686a <=( (not A233)  and  a41685a );
 a41689a <=( (not A269)  and  (not A268) );
 a41692a <=( A300  and  A298 );
 a41693a <=( a41692a  and  a41689a );
 a41694a <=( a41693a  and  a41686a );
 a41698a <=( A166  and  (not A167) );
 a41699a <=( A170  and  a41698a );
 a41702a <=( (not A200)  and  (not A199) );
 a41705a <=( (not A232)  and  (not A202) );
 a41706a <=( a41705a  and  a41702a );
 a41707a <=( a41706a  and  a41699a );
 a41711a <=( A265  and  (not A235) );
 a41712a <=( (not A233)  and  a41711a );
 a41715a <=( (not A267)  and  A266 );
 a41718a <=( A301  and  (not A268) );
 a41719a <=( a41718a  and  a41715a );
 a41720a <=( a41719a  and  a41712a );
 a41724a <=( A166  and  (not A167) );
 a41725a <=( A170  and  a41724a );
 a41728a <=( (not A200)  and  (not A199) );
 a41731a <=( (not A232)  and  (not A202) );
 a41732a <=( a41731a  and  a41728a );
 a41733a <=( a41732a  and  a41725a );
 a41737a <=( (not A265)  and  (not A235) );
 a41738a <=( (not A233)  and  a41737a );
 a41741a <=( (not A268)  and  (not A266) );
 a41744a <=( A300  and  A299 );
 a41745a <=( a41744a  and  a41741a );
 a41746a <=( a41745a  and  a41738a );
 a41750a <=( A166  and  (not A167) );
 a41751a <=( A170  and  a41750a );
 a41754a <=( (not A200)  and  (not A199) );
 a41757a <=( (not A232)  and  (not A202) );
 a41758a <=( a41757a  and  a41754a );
 a41759a <=( a41758a  and  a41751a );
 a41763a <=( (not A265)  and  (not A235) );
 a41764a <=( (not A233)  and  a41763a );
 a41767a <=( (not A268)  and  (not A266) );
 a41770a <=( A300  and  A298 );
 a41771a <=( a41770a  and  a41767a );
 a41772a <=( a41771a  and  a41764a );
 a41776a <=( (not A202)  and  (not A201) );
 a41777a <=( A169  and  a41776a );
 a41780a <=( (not A234)  and  (not A203) );
 a41783a <=( (not A236)  and  (not A235) );
 a41784a <=( a41783a  and  a41780a );
 a41785a <=( a41784a  and  a41777a );
 a41789a <=( (not A267)  and  A266 );
 a41790a <=( A265  and  a41789a );
 a41793a <=( A298  and  (not A268) );
 a41796a <=( A302  and  (not A299) );
 a41797a <=( a41796a  and  a41793a );
 a41798a <=( a41797a  and  a41790a );
 a41802a <=( (not A202)  and  (not A201) );
 a41803a <=( A169  and  a41802a );
 a41806a <=( (not A234)  and  (not A203) );
 a41809a <=( (not A236)  and  (not A235) );
 a41810a <=( a41809a  and  a41806a );
 a41811a <=( a41810a  and  a41803a );
 a41815a <=( (not A267)  and  A266 );
 a41816a <=( A265  and  a41815a );
 a41819a <=( (not A298)  and  (not A268) );
 a41822a <=( A302  and  A299 );
 a41823a <=( a41822a  and  a41819a );
 a41824a <=( a41823a  and  a41816a );
 a41828a <=( (not A202)  and  (not A201) );
 a41829a <=( A169  and  a41828a );
 a41832a <=( A232  and  (not A203) );
 a41835a <=( (not A234)  and  A233 );
 a41836a <=( a41835a  and  a41832a );
 a41837a <=( a41836a  and  a41829a );
 a41841a <=( (not A268)  and  (not A267) );
 a41842a <=( (not A235)  and  a41841a );
 a41845a <=( A298  and  (not A269) );
 a41848a <=( A302  and  (not A299) );
 a41849a <=( a41848a  and  a41845a );
 a41850a <=( a41849a  and  a41842a );
 a41854a <=( (not A202)  and  (not A201) );
 a41855a <=( A169  and  a41854a );
 a41858a <=( A232  and  (not A203) );
 a41861a <=( (not A234)  and  A233 );
 a41862a <=( a41861a  and  a41858a );
 a41863a <=( a41862a  and  a41855a );
 a41867a <=( (not A268)  and  (not A267) );
 a41868a <=( (not A235)  and  a41867a );
 a41871a <=( (not A298)  and  (not A269) );
 a41874a <=( A302  and  A299 );
 a41875a <=( a41874a  and  a41871a );
 a41876a <=( a41875a  and  a41868a );
 a41880a <=( (not A202)  and  (not A201) );
 a41881a <=( A169  and  a41880a );
 a41884a <=( A232  and  (not A203) );
 a41887a <=( (not A234)  and  A233 );
 a41888a <=( a41887a  and  a41884a );
 a41889a <=( a41888a  and  a41881a );
 a41893a <=( A266  and  A265 );
 a41894a <=( (not A235)  and  a41893a );
 a41897a <=( (not A268)  and  (not A267) );
 a41900a <=( A300  and  A299 );
 a41901a <=( a41900a  and  a41897a );
 a41902a <=( a41901a  and  a41894a );
 a41906a <=( (not A202)  and  (not A201) );
 a41907a <=( A169  and  a41906a );
 a41910a <=( A232  and  (not A203) );
 a41913a <=( (not A234)  and  A233 );
 a41914a <=( a41913a  and  a41910a );
 a41915a <=( a41914a  and  a41907a );
 a41919a <=( A266  and  A265 );
 a41920a <=( (not A235)  and  a41919a );
 a41923a <=( (not A268)  and  (not A267) );
 a41926a <=( A300  and  A298 );
 a41927a <=( a41926a  and  a41923a );
 a41928a <=( a41927a  and  a41920a );
 a41932a <=( (not A202)  and  (not A201) );
 a41933a <=( A169  and  a41932a );
 a41936a <=( A232  and  (not A203) );
 a41939a <=( (not A234)  and  A233 );
 a41940a <=( a41939a  and  a41936a );
 a41941a <=( a41940a  and  a41933a );
 a41945a <=( (not A266)  and  (not A265) );
 a41946a <=( (not A235)  and  a41945a );
 a41949a <=( A298  and  (not A268) );
 a41952a <=( A302  and  (not A299) );
 a41953a <=( a41952a  and  a41949a );
 a41954a <=( a41953a  and  a41946a );
 a41958a <=( (not A202)  and  (not A201) );
 a41959a <=( A169  and  a41958a );
 a41962a <=( A232  and  (not A203) );
 a41965a <=( (not A234)  and  A233 );
 a41966a <=( a41965a  and  a41962a );
 a41967a <=( a41966a  and  a41959a );
 a41971a <=( (not A266)  and  (not A265) );
 a41972a <=( (not A235)  and  a41971a );
 a41975a <=( (not A298)  and  (not A268) );
 a41978a <=( A302  and  A299 );
 a41979a <=( a41978a  and  a41975a );
 a41980a <=( a41979a  and  a41972a );
 a41984a <=( (not A202)  and  (not A201) );
 a41985a <=( A169  and  a41984a );
 a41988a <=( (not A232)  and  (not A203) );
 a41991a <=( (not A235)  and  (not A233) );
 a41992a <=( a41991a  and  a41988a );
 a41993a <=( a41992a  and  a41985a );
 a41997a <=( (not A267)  and  A266 );
 a41998a <=( A265  and  a41997a );
 a42001a <=( A298  and  (not A268) );
 a42004a <=( A302  and  (not A299) );
 a42005a <=( a42004a  and  a42001a );
 a42006a <=( a42005a  and  a41998a );
 a42010a <=( (not A202)  and  (not A201) );
 a42011a <=( A169  and  a42010a );
 a42014a <=( (not A232)  and  (not A203) );
 a42017a <=( (not A235)  and  (not A233) );
 a42018a <=( a42017a  and  a42014a );
 a42019a <=( a42018a  and  a42011a );
 a42023a <=( (not A267)  and  A266 );
 a42024a <=( A265  and  a42023a );
 a42027a <=( (not A298)  and  (not A268) );
 a42030a <=( A302  and  A299 );
 a42031a <=( a42030a  and  a42027a );
 a42032a <=( a42031a  and  a42024a );
 a42036a <=( A200  and  A199 );
 a42037a <=( A169  and  a42036a );
 a42040a <=( (not A202)  and  (not A201) );
 a42043a <=( (not A235)  and  (not A234) );
 a42044a <=( a42043a  and  a42040a );
 a42045a <=( a42044a  and  a42037a );
 a42049a <=( (not A268)  and  (not A267) );
 a42050a <=( (not A236)  and  a42049a );
 a42053a <=( A298  and  (not A269) );
 a42056a <=( A302  and  (not A299) );
 a42057a <=( a42056a  and  a42053a );
 a42058a <=( a42057a  and  a42050a );
 a42062a <=( A200  and  A199 );
 a42063a <=( A169  and  a42062a );
 a42066a <=( (not A202)  and  (not A201) );
 a42069a <=( (not A235)  and  (not A234) );
 a42070a <=( a42069a  and  a42066a );
 a42071a <=( a42070a  and  a42063a );
 a42075a <=( (not A268)  and  (not A267) );
 a42076a <=( (not A236)  and  a42075a );
 a42079a <=( (not A298)  and  (not A269) );
 a42082a <=( A302  and  A299 );
 a42083a <=( a42082a  and  a42079a );
 a42084a <=( a42083a  and  a42076a );
 a42088a <=( A200  and  A199 );
 a42089a <=( A169  and  a42088a );
 a42092a <=( (not A202)  and  (not A201) );
 a42095a <=( (not A235)  and  (not A234) );
 a42096a <=( a42095a  and  a42092a );
 a42097a <=( a42096a  and  a42089a );
 a42101a <=( A266  and  A265 );
 a42102a <=( (not A236)  and  a42101a );
 a42105a <=( (not A268)  and  (not A267) );
 a42108a <=( A300  and  A299 );
 a42109a <=( a42108a  and  a42105a );
 a42110a <=( a42109a  and  a42102a );
 a42114a <=( A200  and  A199 );
 a42115a <=( A169  and  a42114a );
 a42118a <=( (not A202)  and  (not A201) );
 a42121a <=( (not A235)  and  (not A234) );
 a42122a <=( a42121a  and  a42118a );
 a42123a <=( a42122a  and  a42115a );
 a42127a <=( A266  and  A265 );
 a42128a <=( (not A236)  and  a42127a );
 a42131a <=( (not A268)  and  (not A267) );
 a42134a <=( A300  and  A298 );
 a42135a <=( a42134a  and  a42131a );
 a42136a <=( a42135a  and  a42128a );
 a42140a <=( A200  and  A199 );
 a42141a <=( A169  and  a42140a );
 a42144a <=( (not A202)  and  (not A201) );
 a42147a <=( (not A235)  and  (not A234) );
 a42148a <=( a42147a  and  a42144a );
 a42149a <=( a42148a  and  a42141a );
 a42153a <=( (not A266)  and  (not A265) );
 a42154a <=( (not A236)  and  a42153a );
 a42157a <=( A298  and  (not A268) );
 a42160a <=( A302  and  (not A299) );
 a42161a <=( a42160a  and  a42157a );
 a42162a <=( a42161a  and  a42154a );
 a42166a <=( A200  and  A199 );
 a42167a <=( A169  and  a42166a );
 a42170a <=( (not A202)  and  (not A201) );
 a42173a <=( (not A235)  and  (not A234) );
 a42174a <=( a42173a  and  a42170a );
 a42175a <=( a42174a  and  a42167a );
 a42179a <=( (not A266)  and  (not A265) );
 a42180a <=( (not A236)  and  a42179a );
 a42183a <=( (not A298)  and  (not A268) );
 a42186a <=( A302  and  A299 );
 a42187a <=( a42186a  and  a42183a );
 a42188a <=( a42187a  and  a42180a );
 a42192a <=( A200  and  A199 );
 a42193a <=( A169  and  a42192a );
 a42196a <=( (not A202)  and  (not A201) );
 a42199a <=( A233  and  A232 );
 a42200a <=( a42199a  and  a42196a );
 a42201a <=( a42200a  and  a42193a );
 a42205a <=( (not A267)  and  (not A235) );
 a42206a <=( (not A234)  and  a42205a );
 a42209a <=( (not A269)  and  (not A268) );
 a42212a <=( A300  and  A299 );
 a42213a <=( a42212a  and  a42209a );
 a42214a <=( a42213a  and  a42206a );
 a42218a <=( A200  and  A199 );
 a42219a <=( A169  and  a42218a );
 a42222a <=( (not A202)  and  (not A201) );
 a42225a <=( A233  and  A232 );
 a42226a <=( a42225a  and  a42222a );
 a42227a <=( a42226a  and  a42219a );
 a42231a <=( (not A267)  and  (not A235) );
 a42232a <=( (not A234)  and  a42231a );
 a42235a <=( (not A269)  and  (not A268) );
 a42238a <=( A300  and  A298 );
 a42239a <=( a42238a  and  a42235a );
 a42240a <=( a42239a  and  a42232a );
 a42244a <=( A200  and  A199 );
 a42245a <=( A169  and  a42244a );
 a42248a <=( (not A202)  and  (not A201) );
 a42251a <=( A233  and  A232 );
 a42252a <=( a42251a  and  a42248a );
 a42253a <=( a42252a  and  a42245a );
 a42257a <=( A265  and  (not A235) );
 a42258a <=( (not A234)  and  a42257a );
 a42261a <=( (not A267)  and  A266 );
 a42264a <=( A301  and  (not A268) );
 a42265a <=( a42264a  and  a42261a );
 a42266a <=( a42265a  and  a42258a );
 a42270a <=( A200  and  A199 );
 a42271a <=( A169  and  a42270a );
 a42274a <=( (not A202)  and  (not A201) );
 a42277a <=( A233  and  A232 );
 a42278a <=( a42277a  and  a42274a );
 a42279a <=( a42278a  and  a42271a );
 a42283a <=( (not A265)  and  (not A235) );
 a42284a <=( (not A234)  and  a42283a );
 a42287a <=( (not A268)  and  (not A266) );
 a42290a <=( A300  and  A299 );
 a42291a <=( a42290a  and  a42287a );
 a42292a <=( a42291a  and  a42284a );
 a42296a <=( A200  and  A199 );
 a42297a <=( A169  and  a42296a );
 a42300a <=( (not A202)  and  (not A201) );
 a42303a <=( A233  and  A232 );
 a42304a <=( a42303a  and  a42300a );
 a42305a <=( a42304a  and  a42297a );
 a42309a <=( (not A265)  and  (not A235) );
 a42310a <=( (not A234)  and  a42309a );
 a42313a <=( (not A268)  and  (not A266) );
 a42316a <=( A300  and  A298 );
 a42317a <=( a42316a  and  a42313a );
 a42318a <=( a42317a  and  a42310a );
 a42322a <=( A200  and  A199 );
 a42323a <=( A169  and  a42322a );
 a42326a <=( (not A202)  and  (not A201) );
 a42329a <=( (not A233)  and  (not A232) );
 a42330a <=( a42329a  and  a42326a );
 a42331a <=( a42330a  and  a42323a );
 a42335a <=( (not A268)  and  (not A267) );
 a42336a <=( (not A235)  and  a42335a );
 a42339a <=( A298  and  (not A269) );
 a42342a <=( A302  and  (not A299) );
 a42343a <=( a42342a  and  a42339a );
 a42344a <=( a42343a  and  a42336a );
 a42348a <=( A200  and  A199 );
 a42349a <=( A169  and  a42348a );
 a42352a <=( (not A202)  and  (not A201) );
 a42355a <=( (not A233)  and  (not A232) );
 a42356a <=( a42355a  and  a42352a );
 a42357a <=( a42356a  and  a42349a );
 a42361a <=( (not A268)  and  (not A267) );
 a42362a <=( (not A235)  and  a42361a );
 a42365a <=( (not A298)  and  (not A269) );
 a42368a <=( A302  and  A299 );
 a42369a <=( a42368a  and  a42365a );
 a42370a <=( a42369a  and  a42362a );
 a42374a <=( A200  and  A199 );
 a42375a <=( A169  and  a42374a );
 a42378a <=( (not A202)  and  (not A201) );
 a42381a <=( (not A233)  and  (not A232) );
 a42382a <=( a42381a  and  a42378a );
 a42383a <=( a42382a  and  a42375a );
 a42387a <=( A266  and  A265 );
 a42388a <=( (not A235)  and  a42387a );
 a42391a <=( (not A268)  and  (not A267) );
 a42394a <=( A300  and  A299 );
 a42395a <=( a42394a  and  a42391a );
 a42396a <=( a42395a  and  a42388a );
 a42400a <=( A200  and  A199 );
 a42401a <=( A169  and  a42400a );
 a42404a <=( (not A202)  and  (not A201) );
 a42407a <=( (not A233)  and  (not A232) );
 a42408a <=( a42407a  and  a42404a );
 a42409a <=( a42408a  and  a42401a );
 a42413a <=( A266  and  A265 );
 a42414a <=( (not A235)  and  a42413a );
 a42417a <=( (not A268)  and  (not A267) );
 a42420a <=( A300  and  A298 );
 a42421a <=( a42420a  and  a42417a );
 a42422a <=( a42421a  and  a42414a );
 a42426a <=( A200  and  A199 );
 a42427a <=( A169  and  a42426a );
 a42430a <=( (not A202)  and  (not A201) );
 a42433a <=( (not A233)  and  (not A232) );
 a42434a <=( a42433a  and  a42430a );
 a42435a <=( a42434a  and  a42427a );
 a42439a <=( (not A266)  and  (not A265) );
 a42440a <=( (not A235)  and  a42439a );
 a42443a <=( A298  and  (not A268) );
 a42446a <=( A302  and  (not A299) );
 a42447a <=( a42446a  and  a42443a );
 a42448a <=( a42447a  and  a42440a );
 a42452a <=( A200  and  A199 );
 a42453a <=( A169  and  a42452a );
 a42456a <=( (not A202)  and  (not A201) );
 a42459a <=( (not A233)  and  (not A232) );
 a42460a <=( a42459a  and  a42456a );
 a42461a <=( a42460a  and  a42453a );
 a42465a <=( (not A266)  and  (not A265) );
 a42466a <=( (not A235)  and  a42465a );
 a42469a <=( (not A298)  and  (not A268) );
 a42472a <=( A302  and  A299 );
 a42473a <=( a42472a  and  a42469a );
 a42474a <=( a42473a  and  a42466a );
 a42478a <=( (not A200)  and  (not A199) );
 a42479a <=( A169  and  a42478a );
 a42482a <=( (not A234)  and  (not A202) );
 a42485a <=( (not A236)  and  (not A235) );
 a42486a <=( a42485a  and  a42482a );
 a42487a <=( a42486a  and  a42479a );
 a42491a <=( (not A267)  and  A266 );
 a42492a <=( A265  and  a42491a );
 a42495a <=( A298  and  (not A268) );
 a42498a <=( A302  and  (not A299) );
 a42499a <=( a42498a  and  a42495a );
 a42500a <=( a42499a  and  a42492a );
 a42504a <=( (not A200)  and  (not A199) );
 a42505a <=( A169  and  a42504a );
 a42508a <=( (not A234)  and  (not A202) );
 a42511a <=( (not A236)  and  (not A235) );
 a42512a <=( a42511a  and  a42508a );
 a42513a <=( a42512a  and  a42505a );
 a42517a <=( (not A267)  and  A266 );
 a42518a <=( A265  and  a42517a );
 a42521a <=( (not A298)  and  (not A268) );
 a42524a <=( A302  and  A299 );
 a42525a <=( a42524a  and  a42521a );
 a42526a <=( a42525a  and  a42518a );
 a42530a <=( (not A200)  and  (not A199) );
 a42531a <=( A169  and  a42530a );
 a42534a <=( A232  and  (not A202) );
 a42537a <=( (not A234)  and  A233 );
 a42538a <=( a42537a  and  a42534a );
 a42539a <=( a42538a  and  a42531a );
 a42543a <=( (not A268)  and  (not A267) );
 a42544a <=( (not A235)  and  a42543a );
 a42547a <=( A298  and  (not A269) );
 a42550a <=( A302  and  (not A299) );
 a42551a <=( a42550a  and  a42547a );
 a42552a <=( a42551a  and  a42544a );
 a42556a <=( (not A200)  and  (not A199) );
 a42557a <=( A169  and  a42556a );
 a42560a <=( A232  and  (not A202) );
 a42563a <=( (not A234)  and  A233 );
 a42564a <=( a42563a  and  a42560a );
 a42565a <=( a42564a  and  a42557a );
 a42569a <=( (not A268)  and  (not A267) );
 a42570a <=( (not A235)  and  a42569a );
 a42573a <=( (not A298)  and  (not A269) );
 a42576a <=( A302  and  A299 );
 a42577a <=( a42576a  and  a42573a );
 a42578a <=( a42577a  and  a42570a );
 a42582a <=( (not A200)  and  (not A199) );
 a42583a <=( A169  and  a42582a );
 a42586a <=( A232  and  (not A202) );
 a42589a <=( (not A234)  and  A233 );
 a42590a <=( a42589a  and  a42586a );
 a42591a <=( a42590a  and  a42583a );
 a42595a <=( A266  and  A265 );
 a42596a <=( (not A235)  and  a42595a );
 a42599a <=( (not A268)  and  (not A267) );
 a42602a <=( A300  and  A299 );
 a42603a <=( a42602a  and  a42599a );
 a42604a <=( a42603a  and  a42596a );
 a42608a <=( (not A200)  and  (not A199) );
 a42609a <=( A169  and  a42608a );
 a42612a <=( A232  and  (not A202) );
 a42615a <=( (not A234)  and  A233 );
 a42616a <=( a42615a  and  a42612a );
 a42617a <=( a42616a  and  a42609a );
 a42621a <=( A266  and  A265 );
 a42622a <=( (not A235)  and  a42621a );
 a42625a <=( (not A268)  and  (not A267) );
 a42628a <=( A300  and  A298 );
 a42629a <=( a42628a  and  a42625a );
 a42630a <=( a42629a  and  a42622a );
 a42634a <=( (not A200)  and  (not A199) );
 a42635a <=( A169  and  a42634a );
 a42638a <=( A232  and  (not A202) );
 a42641a <=( (not A234)  and  A233 );
 a42642a <=( a42641a  and  a42638a );
 a42643a <=( a42642a  and  a42635a );
 a42647a <=( (not A266)  and  (not A265) );
 a42648a <=( (not A235)  and  a42647a );
 a42651a <=( A298  and  (not A268) );
 a42654a <=( A302  and  (not A299) );
 a42655a <=( a42654a  and  a42651a );
 a42656a <=( a42655a  and  a42648a );
 a42660a <=( (not A200)  and  (not A199) );
 a42661a <=( A169  and  a42660a );
 a42664a <=( A232  and  (not A202) );
 a42667a <=( (not A234)  and  A233 );
 a42668a <=( a42667a  and  a42664a );
 a42669a <=( a42668a  and  a42661a );
 a42673a <=( (not A266)  and  (not A265) );
 a42674a <=( (not A235)  and  a42673a );
 a42677a <=( (not A298)  and  (not A268) );
 a42680a <=( A302  and  A299 );
 a42681a <=( a42680a  and  a42677a );
 a42682a <=( a42681a  and  a42674a );
 a42686a <=( (not A200)  and  (not A199) );
 a42687a <=( A169  and  a42686a );
 a42690a <=( (not A232)  and  (not A202) );
 a42693a <=( (not A235)  and  (not A233) );
 a42694a <=( a42693a  and  a42690a );
 a42695a <=( a42694a  and  a42687a );
 a42699a <=( (not A267)  and  A266 );
 a42700a <=( A265  and  a42699a );
 a42703a <=( A298  and  (not A268) );
 a42706a <=( A302  and  (not A299) );
 a42707a <=( a42706a  and  a42703a );
 a42708a <=( a42707a  and  a42700a );
 a42712a <=( (not A200)  and  (not A199) );
 a42713a <=( A169  and  a42712a );
 a42716a <=( (not A232)  and  (not A202) );
 a42719a <=( (not A235)  and  (not A233) );
 a42720a <=( a42719a  and  a42716a );
 a42721a <=( a42720a  and  a42713a );
 a42725a <=( (not A267)  and  A266 );
 a42726a <=( A265  and  a42725a );
 a42729a <=( (not A298)  and  (not A268) );
 a42732a <=( A302  and  A299 );
 a42733a <=( a42732a  and  a42729a );
 a42734a <=( a42733a  and  a42726a );
 a42738a <=( (not A166)  and  (not A167) );
 a42739a <=( (not A169)  and  a42738a );
 a42742a <=( (not A234)  and  A202 );
 a42745a <=( (not A236)  and  (not A235) );
 a42746a <=( a42745a  and  a42742a );
 a42747a <=( a42746a  and  a42739a );
 a42751a <=( (not A267)  and  A266 );
 a42752a <=( A265  and  a42751a );
 a42755a <=( A298  and  (not A268) );
 a42758a <=( A302  and  (not A299) );
 a42759a <=( a42758a  and  a42755a );
 a42760a <=( a42759a  and  a42752a );
 a42764a <=( (not A166)  and  (not A167) );
 a42765a <=( (not A169)  and  a42764a );
 a42768a <=( (not A234)  and  A202 );
 a42771a <=( (not A236)  and  (not A235) );
 a42772a <=( a42771a  and  a42768a );
 a42773a <=( a42772a  and  a42765a );
 a42777a <=( (not A267)  and  A266 );
 a42778a <=( A265  and  a42777a );
 a42781a <=( (not A298)  and  (not A268) );
 a42784a <=( A302  and  A299 );
 a42785a <=( a42784a  and  a42781a );
 a42786a <=( a42785a  and  a42778a );
 a42790a <=( (not A166)  and  (not A167) );
 a42791a <=( (not A169)  and  a42790a );
 a42794a <=( A232  and  A202 );
 a42797a <=( (not A234)  and  A233 );
 a42798a <=( a42797a  and  a42794a );
 a42799a <=( a42798a  and  a42791a );
 a42803a <=( (not A268)  and  (not A267) );
 a42804a <=( (not A235)  and  a42803a );
 a42807a <=( A298  and  (not A269) );
 a42810a <=( A302  and  (not A299) );
 a42811a <=( a42810a  and  a42807a );
 a42812a <=( a42811a  and  a42804a );
 a42816a <=( (not A166)  and  (not A167) );
 a42817a <=( (not A169)  and  a42816a );
 a42820a <=( A232  and  A202 );
 a42823a <=( (not A234)  and  A233 );
 a42824a <=( a42823a  and  a42820a );
 a42825a <=( a42824a  and  a42817a );
 a42829a <=( (not A268)  and  (not A267) );
 a42830a <=( (not A235)  and  a42829a );
 a42833a <=( (not A298)  and  (not A269) );
 a42836a <=( A302  and  A299 );
 a42837a <=( a42836a  and  a42833a );
 a42838a <=( a42837a  and  a42830a );
 a42842a <=( (not A166)  and  (not A167) );
 a42843a <=( (not A169)  and  a42842a );
 a42846a <=( A232  and  A202 );
 a42849a <=( (not A234)  and  A233 );
 a42850a <=( a42849a  and  a42846a );
 a42851a <=( a42850a  and  a42843a );
 a42855a <=( A266  and  A265 );
 a42856a <=( (not A235)  and  a42855a );
 a42859a <=( (not A268)  and  (not A267) );
 a42862a <=( A300  and  A299 );
 a42863a <=( a42862a  and  a42859a );
 a42864a <=( a42863a  and  a42856a );
 a42868a <=( (not A166)  and  (not A167) );
 a42869a <=( (not A169)  and  a42868a );
 a42872a <=( A232  and  A202 );
 a42875a <=( (not A234)  and  A233 );
 a42876a <=( a42875a  and  a42872a );
 a42877a <=( a42876a  and  a42869a );
 a42881a <=( A266  and  A265 );
 a42882a <=( (not A235)  and  a42881a );
 a42885a <=( (not A268)  and  (not A267) );
 a42888a <=( A300  and  A298 );
 a42889a <=( a42888a  and  a42885a );
 a42890a <=( a42889a  and  a42882a );
 a42894a <=( (not A166)  and  (not A167) );
 a42895a <=( (not A169)  and  a42894a );
 a42898a <=( A232  and  A202 );
 a42901a <=( (not A234)  and  A233 );
 a42902a <=( a42901a  and  a42898a );
 a42903a <=( a42902a  and  a42895a );
 a42907a <=( (not A266)  and  (not A265) );
 a42908a <=( (not A235)  and  a42907a );
 a42911a <=( A298  and  (not A268) );
 a42914a <=( A302  and  (not A299) );
 a42915a <=( a42914a  and  a42911a );
 a42916a <=( a42915a  and  a42908a );
 a42920a <=( (not A166)  and  (not A167) );
 a42921a <=( (not A169)  and  a42920a );
 a42924a <=( A232  and  A202 );
 a42927a <=( (not A234)  and  A233 );
 a42928a <=( a42927a  and  a42924a );
 a42929a <=( a42928a  and  a42921a );
 a42933a <=( (not A266)  and  (not A265) );
 a42934a <=( (not A235)  and  a42933a );
 a42937a <=( (not A298)  and  (not A268) );
 a42940a <=( A302  and  A299 );
 a42941a <=( a42940a  and  a42937a );
 a42942a <=( a42941a  and  a42934a );
 a42946a <=( (not A166)  and  (not A167) );
 a42947a <=( (not A169)  and  a42946a );
 a42950a <=( (not A232)  and  A202 );
 a42953a <=( (not A235)  and  (not A233) );
 a42954a <=( a42953a  and  a42950a );
 a42955a <=( a42954a  and  a42947a );
 a42959a <=( (not A267)  and  A266 );
 a42960a <=( A265  and  a42959a );
 a42963a <=( A298  and  (not A268) );
 a42966a <=( A302  and  (not A299) );
 a42967a <=( a42966a  and  a42963a );
 a42968a <=( a42967a  and  a42960a );
 a42972a <=( (not A166)  and  (not A167) );
 a42973a <=( (not A169)  and  a42972a );
 a42976a <=( (not A232)  and  A202 );
 a42979a <=( (not A235)  and  (not A233) );
 a42980a <=( a42979a  and  a42976a );
 a42981a <=( a42980a  and  a42973a );
 a42985a <=( (not A267)  and  A266 );
 a42986a <=( A265  and  a42985a );
 a42989a <=( (not A298)  and  (not A268) );
 a42992a <=( A302  and  A299 );
 a42993a <=( a42992a  and  a42989a );
 a42994a <=( a42993a  and  a42986a );
 a42998a <=( (not A166)  and  (not A167) );
 a42999a <=( (not A169)  and  a42998a );
 a43002a <=( A201  and  A199 );
 a43005a <=( (not A235)  and  (not A234) );
 a43006a <=( a43005a  and  a43002a );
 a43007a <=( a43006a  and  a42999a );
 a43011a <=( (not A268)  and  (not A267) );
 a43012a <=( (not A236)  and  a43011a );
 a43015a <=( A298  and  (not A269) );
 a43018a <=( A302  and  (not A299) );
 a43019a <=( a43018a  and  a43015a );
 a43020a <=( a43019a  and  a43012a );
 a43024a <=( (not A166)  and  (not A167) );
 a43025a <=( (not A169)  and  a43024a );
 a43028a <=( A201  and  A199 );
 a43031a <=( (not A235)  and  (not A234) );
 a43032a <=( a43031a  and  a43028a );
 a43033a <=( a43032a  and  a43025a );
 a43037a <=( (not A268)  and  (not A267) );
 a43038a <=( (not A236)  and  a43037a );
 a43041a <=( (not A298)  and  (not A269) );
 a43044a <=( A302  and  A299 );
 a43045a <=( a43044a  and  a43041a );
 a43046a <=( a43045a  and  a43038a );
 a43050a <=( (not A166)  and  (not A167) );
 a43051a <=( (not A169)  and  a43050a );
 a43054a <=( A201  and  A199 );
 a43057a <=( (not A235)  and  (not A234) );
 a43058a <=( a43057a  and  a43054a );
 a43059a <=( a43058a  and  a43051a );
 a43063a <=( A266  and  A265 );
 a43064a <=( (not A236)  and  a43063a );
 a43067a <=( (not A268)  and  (not A267) );
 a43070a <=( A300  and  A299 );
 a43071a <=( a43070a  and  a43067a );
 a43072a <=( a43071a  and  a43064a );
 a43076a <=( (not A166)  and  (not A167) );
 a43077a <=( (not A169)  and  a43076a );
 a43080a <=( A201  and  A199 );
 a43083a <=( (not A235)  and  (not A234) );
 a43084a <=( a43083a  and  a43080a );
 a43085a <=( a43084a  and  a43077a );
 a43089a <=( A266  and  A265 );
 a43090a <=( (not A236)  and  a43089a );
 a43093a <=( (not A268)  and  (not A267) );
 a43096a <=( A300  and  A298 );
 a43097a <=( a43096a  and  a43093a );
 a43098a <=( a43097a  and  a43090a );
 a43102a <=( (not A166)  and  (not A167) );
 a43103a <=( (not A169)  and  a43102a );
 a43106a <=( A201  and  A199 );
 a43109a <=( (not A235)  and  (not A234) );
 a43110a <=( a43109a  and  a43106a );
 a43111a <=( a43110a  and  a43103a );
 a43115a <=( (not A266)  and  (not A265) );
 a43116a <=( (not A236)  and  a43115a );
 a43119a <=( A298  and  (not A268) );
 a43122a <=( A302  and  (not A299) );
 a43123a <=( a43122a  and  a43119a );
 a43124a <=( a43123a  and  a43116a );
 a43128a <=( (not A166)  and  (not A167) );
 a43129a <=( (not A169)  and  a43128a );
 a43132a <=( A201  and  A199 );
 a43135a <=( (not A235)  and  (not A234) );
 a43136a <=( a43135a  and  a43132a );
 a43137a <=( a43136a  and  a43129a );
 a43141a <=( (not A266)  and  (not A265) );
 a43142a <=( (not A236)  and  a43141a );
 a43145a <=( (not A298)  and  (not A268) );
 a43148a <=( A302  and  A299 );
 a43149a <=( a43148a  and  a43145a );
 a43150a <=( a43149a  and  a43142a );
 a43154a <=( (not A166)  and  (not A167) );
 a43155a <=( (not A169)  and  a43154a );
 a43158a <=( A201  and  A199 );
 a43161a <=( A233  and  A232 );
 a43162a <=( a43161a  and  a43158a );
 a43163a <=( a43162a  and  a43155a );
 a43167a <=( (not A267)  and  (not A235) );
 a43168a <=( (not A234)  and  a43167a );
 a43171a <=( (not A269)  and  (not A268) );
 a43174a <=( A300  and  A299 );
 a43175a <=( a43174a  and  a43171a );
 a43176a <=( a43175a  and  a43168a );
 a43180a <=( (not A166)  and  (not A167) );
 a43181a <=( (not A169)  and  a43180a );
 a43184a <=( A201  and  A199 );
 a43187a <=( A233  and  A232 );
 a43188a <=( a43187a  and  a43184a );
 a43189a <=( a43188a  and  a43181a );
 a43193a <=( (not A267)  and  (not A235) );
 a43194a <=( (not A234)  and  a43193a );
 a43197a <=( (not A269)  and  (not A268) );
 a43200a <=( A300  and  A298 );
 a43201a <=( a43200a  and  a43197a );
 a43202a <=( a43201a  and  a43194a );
 a43206a <=( (not A166)  and  (not A167) );
 a43207a <=( (not A169)  and  a43206a );
 a43210a <=( A201  and  A199 );
 a43213a <=( A233  and  A232 );
 a43214a <=( a43213a  and  a43210a );
 a43215a <=( a43214a  and  a43207a );
 a43219a <=( A265  and  (not A235) );
 a43220a <=( (not A234)  and  a43219a );
 a43223a <=( (not A267)  and  A266 );
 a43226a <=( A301  and  (not A268) );
 a43227a <=( a43226a  and  a43223a );
 a43228a <=( a43227a  and  a43220a );
 a43232a <=( (not A166)  and  (not A167) );
 a43233a <=( (not A169)  and  a43232a );
 a43236a <=( A201  and  A199 );
 a43239a <=( A233  and  A232 );
 a43240a <=( a43239a  and  a43236a );
 a43241a <=( a43240a  and  a43233a );
 a43245a <=( (not A265)  and  (not A235) );
 a43246a <=( (not A234)  and  a43245a );
 a43249a <=( (not A268)  and  (not A266) );
 a43252a <=( A300  and  A299 );
 a43253a <=( a43252a  and  a43249a );
 a43254a <=( a43253a  and  a43246a );
 a43258a <=( (not A166)  and  (not A167) );
 a43259a <=( (not A169)  and  a43258a );
 a43262a <=( A201  and  A199 );
 a43265a <=( A233  and  A232 );
 a43266a <=( a43265a  and  a43262a );
 a43267a <=( a43266a  and  a43259a );
 a43271a <=( (not A265)  and  (not A235) );
 a43272a <=( (not A234)  and  a43271a );
 a43275a <=( (not A268)  and  (not A266) );
 a43278a <=( A300  and  A298 );
 a43279a <=( a43278a  and  a43275a );
 a43280a <=( a43279a  and  a43272a );
 a43284a <=( (not A166)  and  (not A167) );
 a43285a <=( (not A169)  and  a43284a );
 a43288a <=( A201  and  A199 );
 a43291a <=( (not A233)  and  (not A232) );
 a43292a <=( a43291a  and  a43288a );
 a43293a <=( a43292a  and  a43285a );
 a43297a <=( (not A268)  and  (not A267) );
 a43298a <=( (not A235)  and  a43297a );
 a43301a <=( A298  and  (not A269) );
 a43304a <=( A302  and  (not A299) );
 a43305a <=( a43304a  and  a43301a );
 a43306a <=( a43305a  and  a43298a );
 a43310a <=( (not A166)  and  (not A167) );
 a43311a <=( (not A169)  and  a43310a );
 a43314a <=( A201  and  A199 );
 a43317a <=( (not A233)  and  (not A232) );
 a43318a <=( a43317a  and  a43314a );
 a43319a <=( a43318a  and  a43311a );
 a43323a <=( (not A268)  and  (not A267) );
 a43324a <=( (not A235)  and  a43323a );
 a43327a <=( (not A298)  and  (not A269) );
 a43330a <=( A302  and  A299 );
 a43331a <=( a43330a  and  a43327a );
 a43332a <=( a43331a  and  a43324a );
 a43336a <=( (not A166)  and  (not A167) );
 a43337a <=( (not A169)  and  a43336a );
 a43340a <=( A201  and  A199 );
 a43343a <=( (not A233)  and  (not A232) );
 a43344a <=( a43343a  and  a43340a );
 a43345a <=( a43344a  and  a43337a );
 a43349a <=( A266  and  A265 );
 a43350a <=( (not A235)  and  a43349a );
 a43353a <=( (not A268)  and  (not A267) );
 a43356a <=( A300  and  A299 );
 a43357a <=( a43356a  and  a43353a );
 a43358a <=( a43357a  and  a43350a );
 a43362a <=( (not A166)  and  (not A167) );
 a43363a <=( (not A169)  and  a43362a );
 a43366a <=( A201  and  A199 );
 a43369a <=( (not A233)  and  (not A232) );
 a43370a <=( a43369a  and  a43366a );
 a43371a <=( a43370a  and  a43363a );
 a43375a <=( A266  and  A265 );
 a43376a <=( (not A235)  and  a43375a );
 a43379a <=( (not A268)  and  (not A267) );
 a43382a <=( A300  and  A298 );
 a43383a <=( a43382a  and  a43379a );
 a43384a <=( a43383a  and  a43376a );
 a43388a <=( (not A166)  and  (not A167) );
 a43389a <=( (not A169)  and  a43388a );
 a43392a <=( A201  and  A199 );
 a43395a <=( (not A233)  and  (not A232) );
 a43396a <=( a43395a  and  a43392a );
 a43397a <=( a43396a  and  a43389a );
 a43401a <=( (not A266)  and  (not A265) );
 a43402a <=( (not A235)  and  a43401a );
 a43405a <=( A298  and  (not A268) );
 a43408a <=( A302  and  (not A299) );
 a43409a <=( a43408a  and  a43405a );
 a43410a <=( a43409a  and  a43402a );
 a43414a <=( (not A166)  and  (not A167) );
 a43415a <=( (not A169)  and  a43414a );
 a43418a <=( A201  and  A199 );
 a43421a <=( (not A233)  and  (not A232) );
 a43422a <=( a43421a  and  a43418a );
 a43423a <=( a43422a  and  a43415a );
 a43427a <=( (not A266)  and  (not A265) );
 a43428a <=( (not A235)  and  a43427a );
 a43431a <=( (not A298)  and  (not A268) );
 a43434a <=( A302  and  A299 );
 a43435a <=( a43434a  and  a43431a );
 a43436a <=( a43435a  and  a43428a );
 a43440a <=( (not A166)  and  (not A167) );
 a43441a <=( (not A169)  and  a43440a );
 a43444a <=( A201  and  A200 );
 a43447a <=( (not A235)  and  (not A234) );
 a43448a <=( a43447a  and  a43444a );
 a43449a <=( a43448a  and  a43441a );
 a43453a <=( (not A268)  and  (not A267) );
 a43454a <=( (not A236)  and  a43453a );
 a43457a <=( A298  and  (not A269) );
 a43460a <=( A302  and  (not A299) );
 a43461a <=( a43460a  and  a43457a );
 a43462a <=( a43461a  and  a43454a );
 a43466a <=( (not A166)  and  (not A167) );
 a43467a <=( (not A169)  and  a43466a );
 a43470a <=( A201  and  A200 );
 a43473a <=( (not A235)  and  (not A234) );
 a43474a <=( a43473a  and  a43470a );
 a43475a <=( a43474a  and  a43467a );
 a43479a <=( (not A268)  and  (not A267) );
 a43480a <=( (not A236)  and  a43479a );
 a43483a <=( (not A298)  and  (not A269) );
 a43486a <=( A302  and  A299 );
 a43487a <=( a43486a  and  a43483a );
 a43488a <=( a43487a  and  a43480a );
 a43492a <=( (not A166)  and  (not A167) );
 a43493a <=( (not A169)  and  a43492a );
 a43496a <=( A201  and  A200 );
 a43499a <=( (not A235)  and  (not A234) );
 a43500a <=( a43499a  and  a43496a );
 a43501a <=( a43500a  and  a43493a );
 a43505a <=( A266  and  A265 );
 a43506a <=( (not A236)  and  a43505a );
 a43509a <=( (not A268)  and  (not A267) );
 a43512a <=( A300  and  A299 );
 a43513a <=( a43512a  and  a43509a );
 a43514a <=( a43513a  and  a43506a );
 a43518a <=( (not A166)  and  (not A167) );
 a43519a <=( (not A169)  and  a43518a );
 a43522a <=( A201  and  A200 );
 a43525a <=( (not A235)  and  (not A234) );
 a43526a <=( a43525a  and  a43522a );
 a43527a <=( a43526a  and  a43519a );
 a43531a <=( A266  and  A265 );
 a43532a <=( (not A236)  and  a43531a );
 a43535a <=( (not A268)  and  (not A267) );
 a43538a <=( A300  and  A298 );
 a43539a <=( a43538a  and  a43535a );
 a43540a <=( a43539a  and  a43532a );
 a43544a <=( (not A166)  and  (not A167) );
 a43545a <=( (not A169)  and  a43544a );
 a43548a <=( A201  and  A200 );
 a43551a <=( (not A235)  and  (not A234) );
 a43552a <=( a43551a  and  a43548a );
 a43553a <=( a43552a  and  a43545a );
 a43557a <=( (not A266)  and  (not A265) );
 a43558a <=( (not A236)  and  a43557a );
 a43561a <=( A298  and  (not A268) );
 a43564a <=( A302  and  (not A299) );
 a43565a <=( a43564a  and  a43561a );
 a43566a <=( a43565a  and  a43558a );
 a43570a <=( (not A166)  and  (not A167) );
 a43571a <=( (not A169)  and  a43570a );
 a43574a <=( A201  and  A200 );
 a43577a <=( (not A235)  and  (not A234) );
 a43578a <=( a43577a  and  a43574a );
 a43579a <=( a43578a  and  a43571a );
 a43583a <=( (not A266)  and  (not A265) );
 a43584a <=( (not A236)  and  a43583a );
 a43587a <=( (not A298)  and  (not A268) );
 a43590a <=( A302  and  A299 );
 a43591a <=( a43590a  and  a43587a );
 a43592a <=( a43591a  and  a43584a );
 a43596a <=( (not A166)  and  (not A167) );
 a43597a <=( (not A169)  and  a43596a );
 a43600a <=( A201  and  A200 );
 a43603a <=( A233  and  A232 );
 a43604a <=( a43603a  and  a43600a );
 a43605a <=( a43604a  and  a43597a );
 a43609a <=( (not A267)  and  (not A235) );
 a43610a <=( (not A234)  and  a43609a );
 a43613a <=( (not A269)  and  (not A268) );
 a43616a <=( A300  and  A299 );
 a43617a <=( a43616a  and  a43613a );
 a43618a <=( a43617a  and  a43610a );
 a43622a <=( (not A166)  and  (not A167) );
 a43623a <=( (not A169)  and  a43622a );
 a43626a <=( A201  and  A200 );
 a43629a <=( A233  and  A232 );
 a43630a <=( a43629a  and  a43626a );
 a43631a <=( a43630a  and  a43623a );
 a43635a <=( (not A267)  and  (not A235) );
 a43636a <=( (not A234)  and  a43635a );
 a43639a <=( (not A269)  and  (not A268) );
 a43642a <=( A300  and  A298 );
 a43643a <=( a43642a  and  a43639a );
 a43644a <=( a43643a  and  a43636a );
 a43648a <=( (not A166)  and  (not A167) );
 a43649a <=( (not A169)  and  a43648a );
 a43652a <=( A201  and  A200 );
 a43655a <=( A233  and  A232 );
 a43656a <=( a43655a  and  a43652a );
 a43657a <=( a43656a  and  a43649a );
 a43661a <=( A265  and  (not A235) );
 a43662a <=( (not A234)  and  a43661a );
 a43665a <=( (not A267)  and  A266 );
 a43668a <=( A301  and  (not A268) );
 a43669a <=( a43668a  and  a43665a );
 a43670a <=( a43669a  and  a43662a );
 a43674a <=( (not A166)  and  (not A167) );
 a43675a <=( (not A169)  and  a43674a );
 a43678a <=( A201  and  A200 );
 a43681a <=( A233  and  A232 );
 a43682a <=( a43681a  and  a43678a );
 a43683a <=( a43682a  and  a43675a );
 a43687a <=( (not A265)  and  (not A235) );
 a43688a <=( (not A234)  and  a43687a );
 a43691a <=( (not A268)  and  (not A266) );
 a43694a <=( A300  and  A299 );
 a43695a <=( a43694a  and  a43691a );
 a43696a <=( a43695a  and  a43688a );
 a43700a <=( (not A166)  and  (not A167) );
 a43701a <=( (not A169)  and  a43700a );
 a43704a <=( A201  and  A200 );
 a43707a <=( A233  and  A232 );
 a43708a <=( a43707a  and  a43704a );
 a43709a <=( a43708a  and  a43701a );
 a43713a <=( (not A265)  and  (not A235) );
 a43714a <=( (not A234)  and  a43713a );
 a43717a <=( (not A268)  and  (not A266) );
 a43720a <=( A300  and  A298 );
 a43721a <=( a43720a  and  a43717a );
 a43722a <=( a43721a  and  a43714a );
 a43726a <=( (not A166)  and  (not A167) );
 a43727a <=( (not A169)  and  a43726a );
 a43730a <=( A201  and  A200 );
 a43733a <=( (not A233)  and  (not A232) );
 a43734a <=( a43733a  and  a43730a );
 a43735a <=( a43734a  and  a43727a );
 a43739a <=( (not A268)  and  (not A267) );
 a43740a <=( (not A235)  and  a43739a );
 a43743a <=( A298  and  (not A269) );
 a43746a <=( A302  and  (not A299) );
 a43747a <=( a43746a  and  a43743a );
 a43748a <=( a43747a  and  a43740a );
 a43752a <=( (not A166)  and  (not A167) );
 a43753a <=( (not A169)  and  a43752a );
 a43756a <=( A201  and  A200 );
 a43759a <=( (not A233)  and  (not A232) );
 a43760a <=( a43759a  and  a43756a );
 a43761a <=( a43760a  and  a43753a );
 a43765a <=( (not A268)  and  (not A267) );
 a43766a <=( (not A235)  and  a43765a );
 a43769a <=( (not A298)  and  (not A269) );
 a43772a <=( A302  and  A299 );
 a43773a <=( a43772a  and  a43769a );
 a43774a <=( a43773a  and  a43766a );
 a43778a <=( (not A166)  and  (not A167) );
 a43779a <=( (not A169)  and  a43778a );
 a43782a <=( A201  and  A200 );
 a43785a <=( (not A233)  and  (not A232) );
 a43786a <=( a43785a  and  a43782a );
 a43787a <=( a43786a  and  a43779a );
 a43791a <=( A266  and  A265 );
 a43792a <=( (not A235)  and  a43791a );
 a43795a <=( (not A268)  and  (not A267) );
 a43798a <=( A300  and  A299 );
 a43799a <=( a43798a  and  a43795a );
 a43800a <=( a43799a  and  a43792a );
 a43804a <=( (not A166)  and  (not A167) );
 a43805a <=( (not A169)  and  a43804a );
 a43808a <=( A201  and  A200 );
 a43811a <=( (not A233)  and  (not A232) );
 a43812a <=( a43811a  and  a43808a );
 a43813a <=( a43812a  and  a43805a );
 a43817a <=( A266  and  A265 );
 a43818a <=( (not A235)  and  a43817a );
 a43821a <=( (not A268)  and  (not A267) );
 a43824a <=( A300  and  A298 );
 a43825a <=( a43824a  and  a43821a );
 a43826a <=( a43825a  and  a43818a );
 a43830a <=( (not A166)  and  (not A167) );
 a43831a <=( (not A169)  and  a43830a );
 a43834a <=( A201  and  A200 );
 a43837a <=( (not A233)  and  (not A232) );
 a43838a <=( a43837a  and  a43834a );
 a43839a <=( a43838a  and  a43831a );
 a43843a <=( (not A266)  and  (not A265) );
 a43844a <=( (not A235)  and  a43843a );
 a43847a <=( A298  and  (not A268) );
 a43850a <=( A302  and  (not A299) );
 a43851a <=( a43850a  and  a43847a );
 a43852a <=( a43851a  and  a43844a );
 a43856a <=( (not A166)  and  (not A167) );
 a43857a <=( (not A169)  and  a43856a );
 a43860a <=( A201  and  A200 );
 a43863a <=( (not A233)  and  (not A232) );
 a43864a <=( a43863a  and  a43860a );
 a43865a <=( a43864a  and  a43857a );
 a43869a <=( (not A266)  and  (not A265) );
 a43870a <=( (not A235)  and  a43869a );
 a43873a <=( (not A298)  and  (not A268) );
 a43876a <=( A302  and  A299 );
 a43877a <=( a43876a  and  a43873a );
 a43878a <=( a43877a  and  a43870a );
 a43882a <=( (not A166)  and  (not A167) );
 a43883a <=( (not A169)  and  a43882a );
 a43886a <=( A200  and  (not A199) );
 a43889a <=( (not A234)  and  A203 );
 a43890a <=( a43889a  and  a43886a );
 a43891a <=( a43890a  and  a43883a );
 a43895a <=( (not A267)  and  (not A236) );
 a43896a <=( (not A235)  and  a43895a );
 a43899a <=( (not A269)  and  (not A268) );
 a43902a <=( A300  and  A299 );
 a43903a <=( a43902a  and  a43899a );
 a43904a <=( a43903a  and  a43896a );
 a43908a <=( (not A166)  and  (not A167) );
 a43909a <=( (not A169)  and  a43908a );
 a43912a <=( A200  and  (not A199) );
 a43915a <=( (not A234)  and  A203 );
 a43916a <=( a43915a  and  a43912a );
 a43917a <=( a43916a  and  a43909a );
 a43921a <=( (not A267)  and  (not A236) );
 a43922a <=( (not A235)  and  a43921a );
 a43925a <=( (not A269)  and  (not A268) );
 a43928a <=( A300  and  A298 );
 a43929a <=( a43928a  and  a43925a );
 a43930a <=( a43929a  and  a43922a );
 a43934a <=( (not A166)  and  (not A167) );
 a43935a <=( (not A169)  and  a43934a );
 a43938a <=( A200  and  (not A199) );
 a43941a <=( (not A234)  and  A203 );
 a43942a <=( a43941a  and  a43938a );
 a43943a <=( a43942a  and  a43935a );
 a43947a <=( A265  and  (not A236) );
 a43948a <=( (not A235)  and  a43947a );
 a43951a <=( (not A267)  and  A266 );
 a43954a <=( A301  and  (not A268) );
 a43955a <=( a43954a  and  a43951a );
 a43956a <=( a43955a  and  a43948a );
 a43960a <=( (not A166)  and  (not A167) );
 a43961a <=( (not A169)  and  a43960a );
 a43964a <=( A200  and  (not A199) );
 a43967a <=( (not A234)  and  A203 );
 a43968a <=( a43967a  and  a43964a );
 a43969a <=( a43968a  and  a43961a );
 a43973a <=( (not A265)  and  (not A236) );
 a43974a <=( (not A235)  and  a43973a );
 a43977a <=( (not A268)  and  (not A266) );
 a43980a <=( A300  and  A299 );
 a43981a <=( a43980a  and  a43977a );
 a43982a <=( a43981a  and  a43974a );
 a43986a <=( (not A166)  and  (not A167) );
 a43987a <=( (not A169)  and  a43986a );
 a43990a <=( A200  and  (not A199) );
 a43993a <=( (not A234)  and  A203 );
 a43994a <=( a43993a  and  a43990a );
 a43995a <=( a43994a  and  a43987a );
 a43999a <=( (not A265)  and  (not A236) );
 a44000a <=( (not A235)  and  a43999a );
 a44003a <=( (not A268)  and  (not A266) );
 a44006a <=( A300  and  A298 );
 a44007a <=( a44006a  and  a44003a );
 a44008a <=( a44007a  and  a44000a );
 a44012a <=( (not A166)  and  (not A167) );
 a44013a <=( (not A169)  and  a44012a );
 a44016a <=( A200  and  (not A199) );
 a44019a <=( A232  and  A203 );
 a44020a <=( a44019a  and  a44016a );
 a44021a <=( a44020a  and  a44013a );
 a44025a <=( (not A235)  and  (not A234) );
 a44026a <=( A233  and  a44025a );
 a44029a <=( (not A268)  and  (not A267) );
 a44032a <=( A301  and  (not A269) );
 a44033a <=( a44032a  and  a44029a );
 a44034a <=( a44033a  and  a44026a );
 a44038a <=( (not A166)  and  (not A167) );
 a44039a <=( (not A169)  and  a44038a );
 a44042a <=( A200  and  (not A199) );
 a44045a <=( A232  and  A203 );
 a44046a <=( a44045a  and  a44042a );
 a44047a <=( a44046a  and  a44039a );
 a44051a <=( (not A235)  and  (not A234) );
 a44052a <=( A233  and  a44051a );
 a44055a <=( (not A266)  and  (not A265) );
 a44058a <=( A301  and  (not A268) );
 a44059a <=( a44058a  and  a44055a );
 a44060a <=( a44059a  and  a44052a );
 a44064a <=( (not A166)  and  (not A167) );
 a44065a <=( (not A169)  and  a44064a );
 a44068a <=( A200  and  (not A199) );
 a44071a <=( (not A232)  and  A203 );
 a44072a <=( a44071a  and  a44068a );
 a44073a <=( a44072a  and  a44065a );
 a44077a <=( (not A267)  and  (not A235) );
 a44078a <=( (not A233)  and  a44077a );
 a44081a <=( (not A269)  and  (not A268) );
 a44084a <=( A300  and  A299 );
 a44085a <=( a44084a  and  a44081a );
 a44086a <=( a44085a  and  a44078a );
 a44090a <=( (not A166)  and  (not A167) );
 a44091a <=( (not A169)  and  a44090a );
 a44094a <=( A200  and  (not A199) );
 a44097a <=( (not A232)  and  A203 );
 a44098a <=( a44097a  and  a44094a );
 a44099a <=( a44098a  and  a44091a );
 a44103a <=( (not A267)  and  (not A235) );
 a44104a <=( (not A233)  and  a44103a );
 a44107a <=( (not A269)  and  (not A268) );
 a44110a <=( A300  and  A298 );
 a44111a <=( a44110a  and  a44107a );
 a44112a <=( a44111a  and  a44104a );
 a44116a <=( (not A166)  and  (not A167) );
 a44117a <=( (not A169)  and  a44116a );
 a44120a <=( A200  and  (not A199) );
 a44123a <=( (not A232)  and  A203 );
 a44124a <=( a44123a  and  a44120a );
 a44125a <=( a44124a  and  a44117a );
 a44129a <=( A265  and  (not A235) );
 a44130a <=( (not A233)  and  a44129a );
 a44133a <=( (not A267)  and  A266 );
 a44136a <=( A301  and  (not A268) );
 a44137a <=( a44136a  and  a44133a );
 a44138a <=( a44137a  and  a44130a );
 a44142a <=( (not A166)  and  (not A167) );
 a44143a <=( (not A169)  and  a44142a );
 a44146a <=( A200  and  (not A199) );
 a44149a <=( (not A232)  and  A203 );
 a44150a <=( a44149a  and  a44146a );
 a44151a <=( a44150a  and  a44143a );
 a44155a <=( (not A265)  and  (not A235) );
 a44156a <=( (not A233)  and  a44155a );
 a44159a <=( (not A268)  and  (not A266) );
 a44162a <=( A300  and  A299 );
 a44163a <=( a44162a  and  a44159a );
 a44164a <=( a44163a  and  a44156a );
 a44168a <=( (not A166)  and  (not A167) );
 a44169a <=( (not A169)  and  a44168a );
 a44172a <=( A200  and  (not A199) );
 a44175a <=( (not A232)  and  A203 );
 a44176a <=( a44175a  and  a44172a );
 a44177a <=( a44176a  and  a44169a );
 a44181a <=( (not A265)  and  (not A235) );
 a44182a <=( (not A233)  and  a44181a );
 a44185a <=( (not A268)  and  (not A266) );
 a44188a <=( A300  and  A298 );
 a44189a <=( a44188a  and  a44185a );
 a44190a <=( a44189a  and  a44182a );
 a44194a <=( (not A166)  and  (not A167) );
 a44195a <=( (not A169)  and  a44194a );
 a44198a <=( (not A200)  and  A199 );
 a44201a <=( (not A234)  and  A203 );
 a44202a <=( a44201a  and  a44198a );
 a44203a <=( a44202a  and  a44195a );
 a44207a <=( (not A267)  and  (not A236) );
 a44208a <=( (not A235)  and  a44207a );
 a44211a <=( (not A269)  and  (not A268) );
 a44214a <=( A300  and  A299 );
 a44215a <=( a44214a  and  a44211a );
 a44216a <=( a44215a  and  a44208a );
 a44220a <=( (not A166)  and  (not A167) );
 a44221a <=( (not A169)  and  a44220a );
 a44224a <=( (not A200)  and  A199 );
 a44227a <=( (not A234)  and  A203 );
 a44228a <=( a44227a  and  a44224a );
 a44229a <=( a44228a  and  a44221a );
 a44233a <=( (not A267)  and  (not A236) );
 a44234a <=( (not A235)  and  a44233a );
 a44237a <=( (not A269)  and  (not A268) );
 a44240a <=( A300  and  A298 );
 a44241a <=( a44240a  and  a44237a );
 a44242a <=( a44241a  and  a44234a );
 a44246a <=( (not A166)  and  (not A167) );
 a44247a <=( (not A169)  and  a44246a );
 a44250a <=( (not A200)  and  A199 );
 a44253a <=( (not A234)  and  A203 );
 a44254a <=( a44253a  and  a44250a );
 a44255a <=( a44254a  and  a44247a );
 a44259a <=( A265  and  (not A236) );
 a44260a <=( (not A235)  and  a44259a );
 a44263a <=( (not A267)  and  A266 );
 a44266a <=( A301  and  (not A268) );
 a44267a <=( a44266a  and  a44263a );
 a44268a <=( a44267a  and  a44260a );
 a44272a <=( (not A166)  and  (not A167) );
 a44273a <=( (not A169)  and  a44272a );
 a44276a <=( (not A200)  and  A199 );
 a44279a <=( (not A234)  and  A203 );
 a44280a <=( a44279a  and  a44276a );
 a44281a <=( a44280a  and  a44273a );
 a44285a <=( (not A265)  and  (not A236) );
 a44286a <=( (not A235)  and  a44285a );
 a44289a <=( (not A268)  and  (not A266) );
 a44292a <=( A300  and  A299 );
 a44293a <=( a44292a  and  a44289a );
 a44294a <=( a44293a  and  a44286a );
 a44298a <=( (not A166)  and  (not A167) );
 a44299a <=( (not A169)  and  a44298a );
 a44302a <=( (not A200)  and  A199 );
 a44305a <=( (not A234)  and  A203 );
 a44306a <=( a44305a  and  a44302a );
 a44307a <=( a44306a  and  a44299a );
 a44311a <=( (not A265)  and  (not A236) );
 a44312a <=( (not A235)  and  a44311a );
 a44315a <=( (not A268)  and  (not A266) );
 a44318a <=( A300  and  A298 );
 a44319a <=( a44318a  and  a44315a );
 a44320a <=( a44319a  and  a44312a );
 a44324a <=( (not A166)  and  (not A167) );
 a44325a <=( (not A169)  and  a44324a );
 a44328a <=( (not A200)  and  A199 );
 a44331a <=( A232  and  A203 );
 a44332a <=( a44331a  and  a44328a );
 a44333a <=( a44332a  and  a44325a );
 a44337a <=( (not A235)  and  (not A234) );
 a44338a <=( A233  and  a44337a );
 a44341a <=( (not A268)  and  (not A267) );
 a44344a <=( A301  and  (not A269) );
 a44345a <=( a44344a  and  a44341a );
 a44346a <=( a44345a  and  a44338a );
 a44350a <=( (not A166)  and  (not A167) );
 a44351a <=( (not A169)  and  a44350a );
 a44354a <=( (not A200)  and  A199 );
 a44357a <=( A232  and  A203 );
 a44358a <=( a44357a  and  a44354a );
 a44359a <=( a44358a  and  a44351a );
 a44363a <=( (not A235)  and  (not A234) );
 a44364a <=( A233  and  a44363a );
 a44367a <=( (not A266)  and  (not A265) );
 a44370a <=( A301  and  (not A268) );
 a44371a <=( a44370a  and  a44367a );
 a44372a <=( a44371a  and  a44364a );
 a44376a <=( (not A166)  and  (not A167) );
 a44377a <=( (not A169)  and  a44376a );
 a44380a <=( (not A200)  and  A199 );
 a44383a <=( (not A232)  and  A203 );
 a44384a <=( a44383a  and  a44380a );
 a44385a <=( a44384a  and  a44377a );
 a44389a <=( (not A267)  and  (not A235) );
 a44390a <=( (not A233)  and  a44389a );
 a44393a <=( (not A269)  and  (not A268) );
 a44396a <=( A300  and  A299 );
 a44397a <=( a44396a  and  a44393a );
 a44398a <=( a44397a  and  a44390a );
 a44402a <=( (not A166)  and  (not A167) );
 a44403a <=( (not A169)  and  a44402a );
 a44406a <=( (not A200)  and  A199 );
 a44409a <=( (not A232)  and  A203 );
 a44410a <=( a44409a  and  a44406a );
 a44411a <=( a44410a  and  a44403a );
 a44415a <=( (not A267)  and  (not A235) );
 a44416a <=( (not A233)  and  a44415a );
 a44419a <=( (not A269)  and  (not A268) );
 a44422a <=( A300  and  A298 );
 a44423a <=( a44422a  and  a44419a );
 a44424a <=( a44423a  and  a44416a );
 a44428a <=( (not A166)  and  (not A167) );
 a44429a <=( (not A169)  and  a44428a );
 a44432a <=( (not A200)  and  A199 );
 a44435a <=( (not A232)  and  A203 );
 a44436a <=( a44435a  and  a44432a );
 a44437a <=( a44436a  and  a44429a );
 a44441a <=( A265  and  (not A235) );
 a44442a <=( (not A233)  and  a44441a );
 a44445a <=( (not A267)  and  A266 );
 a44448a <=( A301  and  (not A268) );
 a44449a <=( a44448a  and  a44445a );
 a44450a <=( a44449a  and  a44442a );
 a44454a <=( (not A166)  and  (not A167) );
 a44455a <=( (not A169)  and  a44454a );
 a44458a <=( (not A200)  and  A199 );
 a44461a <=( (not A232)  and  A203 );
 a44462a <=( a44461a  and  a44458a );
 a44463a <=( a44462a  and  a44455a );
 a44467a <=( (not A265)  and  (not A235) );
 a44468a <=( (not A233)  and  a44467a );
 a44471a <=( (not A268)  and  (not A266) );
 a44474a <=( A300  and  A299 );
 a44475a <=( a44474a  and  a44471a );
 a44476a <=( a44475a  and  a44468a );
 a44480a <=( (not A166)  and  (not A167) );
 a44481a <=( (not A169)  and  a44480a );
 a44484a <=( (not A200)  and  A199 );
 a44487a <=( (not A232)  and  A203 );
 a44488a <=( a44487a  and  a44484a );
 a44489a <=( a44488a  and  a44481a );
 a44493a <=( (not A265)  and  (not A235) );
 a44494a <=( (not A233)  and  a44493a );
 a44497a <=( (not A268)  and  (not A266) );
 a44500a <=( A300  and  A298 );
 a44501a <=( a44500a  and  a44497a );
 a44502a <=( a44501a  and  a44494a );
 a44506a <=( A167  and  (not A168) );
 a44507a <=( (not A169)  and  a44506a );
 a44510a <=( A202  and  A166 );
 a44513a <=( (not A235)  and  (not A234) );
 a44514a <=( a44513a  and  a44510a );
 a44515a <=( a44514a  and  a44507a );
 a44519a <=( (not A268)  and  (not A267) );
 a44520a <=( (not A236)  and  a44519a );
 a44523a <=( A298  and  (not A269) );
 a44526a <=( A302  and  (not A299) );
 a44527a <=( a44526a  and  a44523a );
 a44528a <=( a44527a  and  a44520a );
 a44532a <=( A167  and  (not A168) );
 a44533a <=( (not A169)  and  a44532a );
 a44536a <=( A202  and  A166 );
 a44539a <=( (not A235)  and  (not A234) );
 a44540a <=( a44539a  and  a44536a );
 a44541a <=( a44540a  and  a44533a );
 a44545a <=( (not A268)  and  (not A267) );
 a44546a <=( (not A236)  and  a44545a );
 a44549a <=( (not A298)  and  (not A269) );
 a44552a <=( A302  and  A299 );
 a44553a <=( a44552a  and  a44549a );
 a44554a <=( a44553a  and  a44546a );
 a44558a <=( A167  and  (not A168) );
 a44559a <=( (not A169)  and  a44558a );
 a44562a <=( A202  and  A166 );
 a44565a <=( (not A235)  and  (not A234) );
 a44566a <=( a44565a  and  a44562a );
 a44567a <=( a44566a  and  a44559a );
 a44571a <=( A266  and  A265 );
 a44572a <=( (not A236)  and  a44571a );
 a44575a <=( (not A268)  and  (not A267) );
 a44578a <=( A300  and  A299 );
 a44579a <=( a44578a  and  a44575a );
 a44580a <=( a44579a  and  a44572a );
 a44584a <=( A167  and  (not A168) );
 a44585a <=( (not A169)  and  a44584a );
 a44588a <=( A202  and  A166 );
 a44591a <=( (not A235)  and  (not A234) );
 a44592a <=( a44591a  and  a44588a );
 a44593a <=( a44592a  and  a44585a );
 a44597a <=( A266  and  A265 );
 a44598a <=( (not A236)  and  a44597a );
 a44601a <=( (not A268)  and  (not A267) );
 a44604a <=( A300  and  A298 );
 a44605a <=( a44604a  and  a44601a );
 a44606a <=( a44605a  and  a44598a );
 a44610a <=( A167  and  (not A168) );
 a44611a <=( (not A169)  and  a44610a );
 a44614a <=( A202  and  A166 );
 a44617a <=( (not A235)  and  (not A234) );
 a44618a <=( a44617a  and  a44614a );
 a44619a <=( a44618a  and  a44611a );
 a44623a <=( (not A266)  and  (not A265) );
 a44624a <=( (not A236)  and  a44623a );
 a44627a <=( A298  and  (not A268) );
 a44630a <=( A302  and  (not A299) );
 a44631a <=( a44630a  and  a44627a );
 a44632a <=( a44631a  and  a44624a );
 a44636a <=( A167  and  (not A168) );
 a44637a <=( (not A169)  and  a44636a );
 a44640a <=( A202  and  A166 );
 a44643a <=( (not A235)  and  (not A234) );
 a44644a <=( a44643a  and  a44640a );
 a44645a <=( a44644a  and  a44637a );
 a44649a <=( (not A266)  and  (not A265) );
 a44650a <=( (not A236)  and  a44649a );
 a44653a <=( (not A298)  and  (not A268) );
 a44656a <=( A302  and  A299 );
 a44657a <=( a44656a  and  a44653a );
 a44658a <=( a44657a  and  a44650a );
 a44662a <=( A167  and  (not A168) );
 a44663a <=( (not A169)  and  a44662a );
 a44666a <=( A202  and  A166 );
 a44669a <=( A233  and  A232 );
 a44670a <=( a44669a  and  a44666a );
 a44671a <=( a44670a  and  a44663a );
 a44675a <=( (not A267)  and  (not A235) );
 a44676a <=( (not A234)  and  a44675a );
 a44679a <=( (not A269)  and  (not A268) );
 a44682a <=( A300  and  A299 );
 a44683a <=( a44682a  and  a44679a );
 a44684a <=( a44683a  and  a44676a );
 a44688a <=( A167  and  (not A168) );
 a44689a <=( (not A169)  and  a44688a );
 a44692a <=( A202  and  A166 );
 a44695a <=( A233  and  A232 );
 a44696a <=( a44695a  and  a44692a );
 a44697a <=( a44696a  and  a44689a );
 a44701a <=( (not A267)  and  (not A235) );
 a44702a <=( (not A234)  and  a44701a );
 a44705a <=( (not A269)  and  (not A268) );
 a44708a <=( A300  and  A298 );
 a44709a <=( a44708a  and  a44705a );
 a44710a <=( a44709a  and  a44702a );
 a44714a <=( A167  and  (not A168) );
 a44715a <=( (not A169)  and  a44714a );
 a44718a <=( A202  and  A166 );
 a44721a <=( A233  and  A232 );
 a44722a <=( a44721a  and  a44718a );
 a44723a <=( a44722a  and  a44715a );
 a44727a <=( A265  and  (not A235) );
 a44728a <=( (not A234)  and  a44727a );
 a44731a <=( (not A267)  and  A266 );
 a44734a <=( A301  and  (not A268) );
 a44735a <=( a44734a  and  a44731a );
 a44736a <=( a44735a  and  a44728a );
 a44740a <=( A167  and  (not A168) );
 a44741a <=( (not A169)  and  a44740a );
 a44744a <=( A202  and  A166 );
 a44747a <=( A233  and  A232 );
 a44748a <=( a44747a  and  a44744a );
 a44749a <=( a44748a  and  a44741a );
 a44753a <=( (not A265)  and  (not A235) );
 a44754a <=( (not A234)  and  a44753a );
 a44757a <=( (not A268)  and  (not A266) );
 a44760a <=( A300  and  A299 );
 a44761a <=( a44760a  and  a44757a );
 a44762a <=( a44761a  and  a44754a );
 a44766a <=( A167  and  (not A168) );
 a44767a <=( (not A169)  and  a44766a );
 a44770a <=( A202  and  A166 );
 a44773a <=( A233  and  A232 );
 a44774a <=( a44773a  and  a44770a );
 a44775a <=( a44774a  and  a44767a );
 a44779a <=( (not A265)  and  (not A235) );
 a44780a <=( (not A234)  and  a44779a );
 a44783a <=( (not A268)  and  (not A266) );
 a44786a <=( A300  and  A298 );
 a44787a <=( a44786a  and  a44783a );
 a44788a <=( a44787a  and  a44780a );
 a44792a <=( A167  and  (not A168) );
 a44793a <=( (not A169)  and  a44792a );
 a44796a <=( A202  and  A166 );
 a44799a <=( (not A233)  and  (not A232) );
 a44800a <=( a44799a  and  a44796a );
 a44801a <=( a44800a  and  a44793a );
 a44805a <=( (not A268)  and  (not A267) );
 a44806a <=( (not A235)  and  a44805a );
 a44809a <=( A298  and  (not A269) );
 a44812a <=( A302  and  (not A299) );
 a44813a <=( a44812a  and  a44809a );
 a44814a <=( a44813a  and  a44806a );
 a44818a <=( A167  and  (not A168) );
 a44819a <=( (not A169)  and  a44818a );
 a44822a <=( A202  and  A166 );
 a44825a <=( (not A233)  and  (not A232) );
 a44826a <=( a44825a  and  a44822a );
 a44827a <=( a44826a  and  a44819a );
 a44831a <=( (not A268)  and  (not A267) );
 a44832a <=( (not A235)  and  a44831a );
 a44835a <=( (not A298)  and  (not A269) );
 a44838a <=( A302  and  A299 );
 a44839a <=( a44838a  and  a44835a );
 a44840a <=( a44839a  and  a44832a );
 a44844a <=( A167  and  (not A168) );
 a44845a <=( (not A169)  and  a44844a );
 a44848a <=( A202  and  A166 );
 a44851a <=( (not A233)  and  (not A232) );
 a44852a <=( a44851a  and  a44848a );
 a44853a <=( a44852a  and  a44845a );
 a44857a <=( A266  and  A265 );
 a44858a <=( (not A235)  and  a44857a );
 a44861a <=( (not A268)  and  (not A267) );
 a44864a <=( A300  and  A299 );
 a44865a <=( a44864a  and  a44861a );
 a44866a <=( a44865a  and  a44858a );
 a44870a <=( A167  and  (not A168) );
 a44871a <=( (not A169)  and  a44870a );
 a44874a <=( A202  and  A166 );
 a44877a <=( (not A233)  and  (not A232) );
 a44878a <=( a44877a  and  a44874a );
 a44879a <=( a44878a  and  a44871a );
 a44883a <=( A266  and  A265 );
 a44884a <=( (not A235)  and  a44883a );
 a44887a <=( (not A268)  and  (not A267) );
 a44890a <=( A300  and  A298 );
 a44891a <=( a44890a  and  a44887a );
 a44892a <=( a44891a  and  a44884a );
 a44896a <=( A167  and  (not A168) );
 a44897a <=( (not A169)  and  a44896a );
 a44900a <=( A202  and  A166 );
 a44903a <=( (not A233)  and  (not A232) );
 a44904a <=( a44903a  and  a44900a );
 a44905a <=( a44904a  and  a44897a );
 a44909a <=( (not A266)  and  (not A265) );
 a44910a <=( (not A235)  and  a44909a );
 a44913a <=( A298  and  (not A268) );
 a44916a <=( A302  and  (not A299) );
 a44917a <=( a44916a  and  a44913a );
 a44918a <=( a44917a  and  a44910a );
 a44922a <=( A167  and  (not A168) );
 a44923a <=( (not A169)  and  a44922a );
 a44926a <=( A202  and  A166 );
 a44929a <=( (not A233)  and  (not A232) );
 a44930a <=( a44929a  and  a44926a );
 a44931a <=( a44930a  and  a44923a );
 a44935a <=( (not A266)  and  (not A265) );
 a44936a <=( (not A235)  and  a44935a );
 a44939a <=( (not A298)  and  (not A268) );
 a44942a <=( A302  and  A299 );
 a44943a <=( a44942a  and  a44939a );
 a44944a <=( a44943a  and  a44936a );
 a44948a <=( A167  and  (not A168) );
 a44949a <=( (not A169)  and  a44948a );
 a44952a <=( A199  and  A166 );
 a44955a <=( (not A234)  and  A201 );
 a44956a <=( a44955a  and  a44952a );
 a44957a <=( a44956a  and  a44949a );
 a44961a <=( (not A267)  and  (not A236) );
 a44962a <=( (not A235)  and  a44961a );
 a44965a <=( (not A269)  and  (not A268) );
 a44968a <=( A300  and  A299 );
 a44969a <=( a44968a  and  a44965a );
 a44970a <=( a44969a  and  a44962a );
 a44974a <=( A167  and  (not A168) );
 a44975a <=( (not A169)  and  a44974a );
 a44978a <=( A199  and  A166 );
 a44981a <=( (not A234)  and  A201 );
 a44982a <=( a44981a  and  a44978a );
 a44983a <=( a44982a  and  a44975a );
 a44987a <=( (not A267)  and  (not A236) );
 a44988a <=( (not A235)  and  a44987a );
 a44991a <=( (not A269)  and  (not A268) );
 a44994a <=( A300  and  A298 );
 a44995a <=( a44994a  and  a44991a );
 a44996a <=( a44995a  and  a44988a );
 a45000a <=( A167  and  (not A168) );
 a45001a <=( (not A169)  and  a45000a );
 a45004a <=( A199  and  A166 );
 a45007a <=( (not A234)  and  A201 );
 a45008a <=( a45007a  and  a45004a );
 a45009a <=( a45008a  and  a45001a );
 a45013a <=( A265  and  (not A236) );
 a45014a <=( (not A235)  and  a45013a );
 a45017a <=( (not A267)  and  A266 );
 a45020a <=( A301  and  (not A268) );
 a45021a <=( a45020a  and  a45017a );
 a45022a <=( a45021a  and  a45014a );
 a45026a <=( A167  and  (not A168) );
 a45027a <=( (not A169)  and  a45026a );
 a45030a <=( A199  and  A166 );
 a45033a <=( (not A234)  and  A201 );
 a45034a <=( a45033a  and  a45030a );
 a45035a <=( a45034a  and  a45027a );
 a45039a <=( (not A265)  and  (not A236) );
 a45040a <=( (not A235)  and  a45039a );
 a45043a <=( (not A268)  and  (not A266) );
 a45046a <=( A300  and  A299 );
 a45047a <=( a45046a  and  a45043a );
 a45048a <=( a45047a  and  a45040a );
 a45052a <=( A167  and  (not A168) );
 a45053a <=( (not A169)  and  a45052a );
 a45056a <=( A199  and  A166 );
 a45059a <=( (not A234)  and  A201 );
 a45060a <=( a45059a  and  a45056a );
 a45061a <=( a45060a  and  a45053a );
 a45065a <=( (not A265)  and  (not A236) );
 a45066a <=( (not A235)  and  a45065a );
 a45069a <=( (not A268)  and  (not A266) );
 a45072a <=( A300  and  A298 );
 a45073a <=( a45072a  and  a45069a );
 a45074a <=( a45073a  and  a45066a );
 a45078a <=( A167  and  (not A168) );
 a45079a <=( (not A169)  and  a45078a );
 a45082a <=( A199  and  A166 );
 a45085a <=( A232  and  A201 );
 a45086a <=( a45085a  and  a45082a );
 a45087a <=( a45086a  and  a45079a );
 a45091a <=( (not A235)  and  (not A234) );
 a45092a <=( A233  and  a45091a );
 a45095a <=( (not A268)  and  (not A267) );
 a45098a <=( A301  and  (not A269) );
 a45099a <=( a45098a  and  a45095a );
 a45100a <=( a45099a  and  a45092a );
 a45104a <=( A167  and  (not A168) );
 a45105a <=( (not A169)  and  a45104a );
 a45108a <=( A199  and  A166 );
 a45111a <=( A232  and  A201 );
 a45112a <=( a45111a  and  a45108a );
 a45113a <=( a45112a  and  a45105a );
 a45117a <=( (not A235)  and  (not A234) );
 a45118a <=( A233  and  a45117a );
 a45121a <=( (not A266)  and  (not A265) );
 a45124a <=( A301  and  (not A268) );
 a45125a <=( a45124a  and  a45121a );
 a45126a <=( a45125a  and  a45118a );
 a45130a <=( A167  and  (not A168) );
 a45131a <=( (not A169)  and  a45130a );
 a45134a <=( A199  and  A166 );
 a45137a <=( (not A232)  and  A201 );
 a45138a <=( a45137a  and  a45134a );
 a45139a <=( a45138a  and  a45131a );
 a45143a <=( (not A267)  and  (not A235) );
 a45144a <=( (not A233)  and  a45143a );
 a45147a <=( (not A269)  and  (not A268) );
 a45150a <=( A300  and  A299 );
 a45151a <=( a45150a  and  a45147a );
 a45152a <=( a45151a  and  a45144a );
 a45156a <=( A167  and  (not A168) );
 a45157a <=( (not A169)  and  a45156a );
 a45160a <=( A199  and  A166 );
 a45163a <=( (not A232)  and  A201 );
 a45164a <=( a45163a  and  a45160a );
 a45165a <=( a45164a  and  a45157a );
 a45169a <=( (not A267)  and  (not A235) );
 a45170a <=( (not A233)  and  a45169a );
 a45173a <=( (not A269)  and  (not A268) );
 a45176a <=( A300  and  A298 );
 a45177a <=( a45176a  and  a45173a );
 a45178a <=( a45177a  and  a45170a );
 a45182a <=( A167  and  (not A168) );
 a45183a <=( (not A169)  and  a45182a );
 a45186a <=( A199  and  A166 );
 a45189a <=( (not A232)  and  A201 );
 a45190a <=( a45189a  and  a45186a );
 a45191a <=( a45190a  and  a45183a );
 a45195a <=( A265  and  (not A235) );
 a45196a <=( (not A233)  and  a45195a );
 a45199a <=( (not A267)  and  A266 );
 a45202a <=( A301  and  (not A268) );
 a45203a <=( a45202a  and  a45199a );
 a45204a <=( a45203a  and  a45196a );
 a45208a <=( A167  and  (not A168) );
 a45209a <=( (not A169)  and  a45208a );
 a45212a <=( A199  and  A166 );
 a45215a <=( (not A232)  and  A201 );
 a45216a <=( a45215a  and  a45212a );
 a45217a <=( a45216a  and  a45209a );
 a45221a <=( (not A265)  and  (not A235) );
 a45222a <=( (not A233)  and  a45221a );
 a45225a <=( (not A268)  and  (not A266) );
 a45228a <=( A300  and  A299 );
 a45229a <=( a45228a  and  a45225a );
 a45230a <=( a45229a  and  a45222a );
 a45234a <=( A167  and  (not A168) );
 a45235a <=( (not A169)  and  a45234a );
 a45238a <=( A199  and  A166 );
 a45241a <=( (not A232)  and  A201 );
 a45242a <=( a45241a  and  a45238a );
 a45243a <=( a45242a  and  a45235a );
 a45247a <=( (not A265)  and  (not A235) );
 a45248a <=( (not A233)  and  a45247a );
 a45251a <=( (not A268)  and  (not A266) );
 a45254a <=( A300  and  A298 );
 a45255a <=( a45254a  and  a45251a );
 a45256a <=( a45255a  and  a45248a );
 a45260a <=( A167  and  (not A168) );
 a45261a <=( (not A169)  and  a45260a );
 a45264a <=( A200  and  A166 );
 a45267a <=( (not A234)  and  A201 );
 a45268a <=( a45267a  and  a45264a );
 a45269a <=( a45268a  and  a45261a );
 a45273a <=( (not A267)  and  (not A236) );
 a45274a <=( (not A235)  and  a45273a );
 a45277a <=( (not A269)  and  (not A268) );
 a45280a <=( A300  and  A299 );
 a45281a <=( a45280a  and  a45277a );
 a45282a <=( a45281a  and  a45274a );
 a45286a <=( A167  and  (not A168) );
 a45287a <=( (not A169)  and  a45286a );
 a45290a <=( A200  and  A166 );
 a45293a <=( (not A234)  and  A201 );
 a45294a <=( a45293a  and  a45290a );
 a45295a <=( a45294a  and  a45287a );
 a45299a <=( (not A267)  and  (not A236) );
 a45300a <=( (not A235)  and  a45299a );
 a45303a <=( (not A269)  and  (not A268) );
 a45306a <=( A300  and  A298 );
 a45307a <=( a45306a  and  a45303a );
 a45308a <=( a45307a  and  a45300a );
 a45312a <=( A167  and  (not A168) );
 a45313a <=( (not A169)  and  a45312a );
 a45316a <=( A200  and  A166 );
 a45319a <=( (not A234)  and  A201 );
 a45320a <=( a45319a  and  a45316a );
 a45321a <=( a45320a  and  a45313a );
 a45325a <=( A265  and  (not A236) );
 a45326a <=( (not A235)  and  a45325a );
 a45329a <=( (not A267)  and  A266 );
 a45332a <=( A301  and  (not A268) );
 a45333a <=( a45332a  and  a45329a );
 a45334a <=( a45333a  and  a45326a );
 a45338a <=( A167  and  (not A168) );
 a45339a <=( (not A169)  and  a45338a );
 a45342a <=( A200  and  A166 );
 a45345a <=( (not A234)  and  A201 );
 a45346a <=( a45345a  and  a45342a );
 a45347a <=( a45346a  and  a45339a );
 a45351a <=( (not A265)  and  (not A236) );
 a45352a <=( (not A235)  and  a45351a );
 a45355a <=( (not A268)  and  (not A266) );
 a45358a <=( A300  and  A299 );
 a45359a <=( a45358a  and  a45355a );
 a45360a <=( a45359a  and  a45352a );
 a45364a <=( A167  and  (not A168) );
 a45365a <=( (not A169)  and  a45364a );
 a45368a <=( A200  and  A166 );
 a45371a <=( (not A234)  and  A201 );
 a45372a <=( a45371a  and  a45368a );
 a45373a <=( a45372a  and  a45365a );
 a45377a <=( (not A265)  and  (not A236) );
 a45378a <=( (not A235)  and  a45377a );
 a45381a <=( (not A268)  and  (not A266) );
 a45384a <=( A300  and  A298 );
 a45385a <=( a45384a  and  a45381a );
 a45386a <=( a45385a  and  a45378a );
 a45390a <=( A167  and  (not A168) );
 a45391a <=( (not A169)  and  a45390a );
 a45394a <=( A200  and  A166 );
 a45397a <=( A232  and  A201 );
 a45398a <=( a45397a  and  a45394a );
 a45399a <=( a45398a  and  a45391a );
 a45403a <=( (not A235)  and  (not A234) );
 a45404a <=( A233  and  a45403a );
 a45407a <=( (not A268)  and  (not A267) );
 a45410a <=( A301  and  (not A269) );
 a45411a <=( a45410a  and  a45407a );
 a45412a <=( a45411a  and  a45404a );
 a45416a <=( A167  and  (not A168) );
 a45417a <=( (not A169)  and  a45416a );
 a45420a <=( A200  and  A166 );
 a45423a <=( A232  and  A201 );
 a45424a <=( a45423a  and  a45420a );
 a45425a <=( a45424a  and  a45417a );
 a45429a <=( (not A235)  and  (not A234) );
 a45430a <=( A233  and  a45429a );
 a45433a <=( (not A266)  and  (not A265) );
 a45436a <=( A301  and  (not A268) );
 a45437a <=( a45436a  and  a45433a );
 a45438a <=( a45437a  and  a45430a );
 a45442a <=( A167  and  (not A168) );
 a45443a <=( (not A169)  and  a45442a );
 a45446a <=( A200  and  A166 );
 a45449a <=( (not A232)  and  A201 );
 a45450a <=( a45449a  and  a45446a );
 a45451a <=( a45450a  and  a45443a );
 a45455a <=( (not A267)  and  (not A235) );
 a45456a <=( (not A233)  and  a45455a );
 a45459a <=( (not A269)  and  (not A268) );
 a45462a <=( A300  and  A299 );
 a45463a <=( a45462a  and  a45459a );
 a45464a <=( a45463a  and  a45456a );
 a45468a <=( A167  and  (not A168) );
 a45469a <=( (not A169)  and  a45468a );
 a45472a <=( A200  and  A166 );
 a45475a <=( (not A232)  and  A201 );
 a45476a <=( a45475a  and  a45472a );
 a45477a <=( a45476a  and  a45469a );
 a45481a <=( (not A267)  and  (not A235) );
 a45482a <=( (not A233)  and  a45481a );
 a45485a <=( (not A269)  and  (not A268) );
 a45488a <=( A300  and  A298 );
 a45489a <=( a45488a  and  a45485a );
 a45490a <=( a45489a  and  a45482a );
 a45494a <=( A167  and  (not A168) );
 a45495a <=( (not A169)  and  a45494a );
 a45498a <=( A200  and  A166 );
 a45501a <=( (not A232)  and  A201 );
 a45502a <=( a45501a  and  a45498a );
 a45503a <=( a45502a  and  a45495a );
 a45507a <=( A265  and  (not A235) );
 a45508a <=( (not A233)  and  a45507a );
 a45511a <=( (not A267)  and  A266 );
 a45514a <=( A301  and  (not A268) );
 a45515a <=( a45514a  and  a45511a );
 a45516a <=( a45515a  and  a45508a );
 a45520a <=( A167  and  (not A168) );
 a45521a <=( (not A169)  and  a45520a );
 a45524a <=( A200  and  A166 );
 a45527a <=( (not A232)  and  A201 );
 a45528a <=( a45527a  and  a45524a );
 a45529a <=( a45528a  and  a45521a );
 a45533a <=( (not A265)  and  (not A235) );
 a45534a <=( (not A233)  and  a45533a );
 a45537a <=( (not A268)  and  (not A266) );
 a45540a <=( A300  and  A299 );
 a45541a <=( a45540a  and  a45537a );
 a45542a <=( a45541a  and  a45534a );
 a45546a <=( A167  and  (not A168) );
 a45547a <=( (not A169)  and  a45546a );
 a45550a <=( A200  and  A166 );
 a45553a <=( (not A232)  and  A201 );
 a45554a <=( a45553a  and  a45550a );
 a45555a <=( a45554a  and  a45547a );
 a45559a <=( (not A265)  and  (not A235) );
 a45560a <=( (not A233)  and  a45559a );
 a45563a <=( (not A268)  and  (not A266) );
 a45566a <=( A300  and  A298 );
 a45567a <=( a45566a  and  a45563a );
 a45568a <=( a45567a  and  a45560a );
 a45572a <=( A167  and  (not A168) );
 a45573a <=( (not A169)  and  a45572a );
 a45576a <=( (not A199)  and  A166 );
 a45579a <=( A203  and  A200 );
 a45580a <=( a45579a  and  a45576a );
 a45581a <=( a45580a  and  a45573a );
 a45585a <=( (not A236)  and  (not A235) );
 a45586a <=( (not A234)  and  a45585a );
 a45589a <=( (not A268)  and  (not A267) );
 a45592a <=( A301  and  (not A269) );
 a45593a <=( a45592a  and  a45589a );
 a45594a <=( a45593a  and  a45586a );
 a45598a <=( A167  and  (not A168) );
 a45599a <=( (not A169)  and  a45598a );
 a45602a <=( (not A199)  and  A166 );
 a45605a <=( A203  and  A200 );
 a45606a <=( a45605a  and  a45602a );
 a45607a <=( a45606a  and  a45599a );
 a45611a <=( (not A236)  and  (not A235) );
 a45612a <=( (not A234)  and  a45611a );
 a45615a <=( (not A266)  and  (not A265) );
 a45618a <=( A301  and  (not A268) );
 a45619a <=( a45618a  and  a45615a );
 a45620a <=( a45619a  and  a45612a );
 a45624a <=( A167  and  (not A168) );
 a45625a <=( (not A169)  and  a45624a );
 a45628a <=( (not A199)  and  A166 );
 a45631a <=( A203  and  A200 );
 a45632a <=( a45631a  and  a45628a );
 a45633a <=( a45632a  and  a45625a );
 a45637a <=( A236  and  A233 );
 a45638a <=( (not A232)  and  a45637a );
 a45641a <=( A299  and  A298 );
 a45644a <=( (not A301)  and  (not A300) );
 a45645a <=( a45644a  and  a45641a );
 a45646a <=( a45645a  and  a45638a );
 a45650a <=( A167  and  (not A168) );
 a45651a <=( (not A169)  and  a45650a );
 a45654a <=( (not A199)  and  A166 );
 a45657a <=( A203  and  A200 );
 a45658a <=( a45657a  and  a45654a );
 a45659a <=( a45658a  and  a45651a );
 a45663a <=( A236  and  (not A233) );
 a45664a <=( A232  and  a45663a );
 a45667a <=( A299  and  A298 );
 a45670a <=( (not A301)  and  (not A300) );
 a45671a <=( a45670a  and  a45667a );
 a45672a <=( a45671a  and  a45664a );
 a45676a <=( A167  and  (not A168) );
 a45677a <=( (not A169)  and  a45676a );
 a45680a <=( (not A199)  and  A166 );
 a45683a <=( A203  and  A200 );
 a45684a <=( a45683a  and  a45680a );
 a45685a <=( a45684a  and  a45677a );
 a45689a <=( (not A235)  and  (not A233) );
 a45690a <=( (not A232)  and  a45689a );
 a45693a <=( (not A268)  and  (not A267) );
 a45696a <=( A301  and  (not A269) );
 a45697a <=( a45696a  and  a45693a );
 a45698a <=( a45697a  and  a45690a );
 a45702a <=( A167  and  (not A168) );
 a45703a <=( (not A169)  and  a45702a );
 a45706a <=( (not A199)  and  A166 );
 a45709a <=( A203  and  A200 );
 a45710a <=( a45709a  and  a45706a );
 a45711a <=( a45710a  and  a45703a );
 a45715a <=( (not A235)  and  (not A233) );
 a45716a <=( (not A232)  and  a45715a );
 a45719a <=( (not A266)  and  (not A265) );
 a45722a <=( A301  and  (not A268) );
 a45723a <=( a45722a  and  a45719a );
 a45724a <=( a45723a  and  a45716a );
 a45728a <=( A167  and  (not A168) );
 a45729a <=( (not A169)  and  a45728a );
 a45732a <=( A199  and  A166 );
 a45735a <=( A203  and  (not A200) );
 a45736a <=( a45735a  and  a45732a );
 a45737a <=( a45736a  and  a45729a );
 a45741a <=( (not A236)  and  (not A235) );
 a45742a <=( (not A234)  and  a45741a );
 a45745a <=( (not A268)  and  (not A267) );
 a45748a <=( A301  and  (not A269) );
 a45749a <=( a45748a  and  a45745a );
 a45750a <=( a45749a  and  a45742a );
 a45754a <=( A167  and  (not A168) );
 a45755a <=( (not A169)  and  a45754a );
 a45758a <=( A199  and  A166 );
 a45761a <=( A203  and  (not A200) );
 a45762a <=( a45761a  and  a45758a );
 a45763a <=( a45762a  and  a45755a );
 a45767a <=( (not A236)  and  (not A235) );
 a45768a <=( (not A234)  and  a45767a );
 a45771a <=( (not A266)  and  (not A265) );
 a45774a <=( A301  and  (not A268) );
 a45775a <=( a45774a  and  a45771a );
 a45776a <=( a45775a  and  a45768a );
 a45780a <=( A167  and  (not A168) );
 a45781a <=( (not A169)  and  a45780a );
 a45784a <=( A199  and  A166 );
 a45787a <=( A203  and  (not A200) );
 a45788a <=( a45787a  and  a45784a );
 a45789a <=( a45788a  and  a45781a );
 a45793a <=( A236  and  A233 );
 a45794a <=( (not A232)  and  a45793a );
 a45797a <=( A299  and  A298 );
 a45800a <=( (not A301)  and  (not A300) );
 a45801a <=( a45800a  and  a45797a );
 a45802a <=( a45801a  and  a45794a );
 a45806a <=( A167  and  (not A168) );
 a45807a <=( (not A169)  and  a45806a );
 a45810a <=( A199  and  A166 );
 a45813a <=( A203  and  (not A200) );
 a45814a <=( a45813a  and  a45810a );
 a45815a <=( a45814a  and  a45807a );
 a45819a <=( A236  and  (not A233) );
 a45820a <=( A232  and  a45819a );
 a45823a <=( A299  and  A298 );
 a45826a <=( (not A301)  and  (not A300) );
 a45827a <=( a45826a  and  a45823a );
 a45828a <=( a45827a  and  a45820a );
 a45832a <=( A167  and  (not A168) );
 a45833a <=( (not A169)  and  a45832a );
 a45836a <=( A199  and  A166 );
 a45839a <=( A203  and  (not A200) );
 a45840a <=( a45839a  and  a45836a );
 a45841a <=( a45840a  and  a45833a );
 a45845a <=( (not A235)  and  (not A233) );
 a45846a <=( (not A232)  and  a45845a );
 a45849a <=( (not A268)  and  (not A267) );
 a45852a <=( A301  and  (not A269) );
 a45853a <=( a45852a  and  a45849a );
 a45854a <=( a45853a  and  a45846a );
 a45858a <=( A167  and  (not A168) );
 a45859a <=( (not A169)  and  a45858a );
 a45862a <=( A199  and  A166 );
 a45865a <=( A203  and  (not A200) );
 a45866a <=( a45865a  and  a45862a );
 a45867a <=( a45866a  and  a45859a );
 a45871a <=( (not A235)  and  (not A233) );
 a45872a <=( (not A232)  and  a45871a );
 a45875a <=( (not A266)  and  (not A265) );
 a45878a <=( A301  and  (not A268) );
 a45879a <=( a45878a  and  a45875a );
 a45880a <=( a45879a  and  a45872a );
 a45884a <=( (not A168)  and  (not A169) );
 a45885a <=( (not A170)  and  a45884a );
 a45888a <=( (not A234)  and  A202 );
 a45891a <=( (not A236)  and  (not A235) );
 a45892a <=( a45891a  and  a45888a );
 a45893a <=( a45892a  and  a45885a );
 a45897a <=( (not A267)  and  A266 );
 a45898a <=( A265  and  a45897a );
 a45901a <=( A298  and  (not A268) );
 a45904a <=( A302  and  (not A299) );
 a45905a <=( a45904a  and  a45901a );
 a45906a <=( a45905a  and  a45898a );
 a45910a <=( (not A168)  and  (not A169) );
 a45911a <=( (not A170)  and  a45910a );
 a45914a <=( (not A234)  and  A202 );
 a45917a <=( (not A236)  and  (not A235) );
 a45918a <=( a45917a  and  a45914a );
 a45919a <=( a45918a  and  a45911a );
 a45923a <=( (not A267)  and  A266 );
 a45924a <=( A265  and  a45923a );
 a45927a <=( (not A298)  and  (not A268) );
 a45930a <=( A302  and  A299 );
 a45931a <=( a45930a  and  a45927a );
 a45932a <=( a45931a  and  a45924a );
 a45936a <=( (not A168)  and  (not A169) );
 a45937a <=( (not A170)  and  a45936a );
 a45940a <=( A232  and  A202 );
 a45943a <=( (not A234)  and  A233 );
 a45944a <=( a45943a  and  a45940a );
 a45945a <=( a45944a  and  a45937a );
 a45949a <=( (not A268)  and  (not A267) );
 a45950a <=( (not A235)  and  a45949a );
 a45953a <=( A298  and  (not A269) );
 a45956a <=( A302  and  (not A299) );
 a45957a <=( a45956a  and  a45953a );
 a45958a <=( a45957a  and  a45950a );
 a45962a <=( (not A168)  and  (not A169) );
 a45963a <=( (not A170)  and  a45962a );
 a45966a <=( A232  and  A202 );
 a45969a <=( (not A234)  and  A233 );
 a45970a <=( a45969a  and  a45966a );
 a45971a <=( a45970a  and  a45963a );
 a45975a <=( (not A268)  and  (not A267) );
 a45976a <=( (not A235)  and  a45975a );
 a45979a <=( (not A298)  and  (not A269) );
 a45982a <=( A302  and  A299 );
 a45983a <=( a45982a  and  a45979a );
 a45984a <=( a45983a  and  a45976a );
 a45988a <=( (not A168)  and  (not A169) );
 a45989a <=( (not A170)  and  a45988a );
 a45992a <=( A232  and  A202 );
 a45995a <=( (not A234)  and  A233 );
 a45996a <=( a45995a  and  a45992a );
 a45997a <=( a45996a  and  a45989a );
 a46001a <=( A266  and  A265 );
 a46002a <=( (not A235)  and  a46001a );
 a46005a <=( (not A268)  and  (not A267) );
 a46008a <=( A300  and  A299 );
 a46009a <=( a46008a  and  a46005a );
 a46010a <=( a46009a  and  a46002a );
 a46014a <=( (not A168)  and  (not A169) );
 a46015a <=( (not A170)  and  a46014a );
 a46018a <=( A232  and  A202 );
 a46021a <=( (not A234)  and  A233 );
 a46022a <=( a46021a  and  a46018a );
 a46023a <=( a46022a  and  a46015a );
 a46027a <=( A266  and  A265 );
 a46028a <=( (not A235)  and  a46027a );
 a46031a <=( (not A268)  and  (not A267) );
 a46034a <=( A300  and  A298 );
 a46035a <=( a46034a  and  a46031a );
 a46036a <=( a46035a  and  a46028a );
 a46040a <=( (not A168)  and  (not A169) );
 a46041a <=( (not A170)  and  a46040a );
 a46044a <=( A232  and  A202 );
 a46047a <=( (not A234)  and  A233 );
 a46048a <=( a46047a  and  a46044a );
 a46049a <=( a46048a  and  a46041a );
 a46053a <=( (not A266)  and  (not A265) );
 a46054a <=( (not A235)  and  a46053a );
 a46057a <=( A298  and  (not A268) );
 a46060a <=( A302  and  (not A299) );
 a46061a <=( a46060a  and  a46057a );
 a46062a <=( a46061a  and  a46054a );
 a46066a <=( (not A168)  and  (not A169) );
 a46067a <=( (not A170)  and  a46066a );
 a46070a <=( A232  and  A202 );
 a46073a <=( (not A234)  and  A233 );
 a46074a <=( a46073a  and  a46070a );
 a46075a <=( a46074a  and  a46067a );
 a46079a <=( (not A266)  and  (not A265) );
 a46080a <=( (not A235)  and  a46079a );
 a46083a <=( (not A298)  and  (not A268) );
 a46086a <=( A302  and  A299 );
 a46087a <=( a46086a  and  a46083a );
 a46088a <=( a46087a  and  a46080a );
 a46092a <=( (not A168)  and  (not A169) );
 a46093a <=( (not A170)  and  a46092a );
 a46096a <=( (not A232)  and  A202 );
 a46099a <=( (not A235)  and  (not A233) );
 a46100a <=( a46099a  and  a46096a );
 a46101a <=( a46100a  and  a46093a );
 a46105a <=( (not A267)  and  A266 );
 a46106a <=( A265  and  a46105a );
 a46109a <=( A298  and  (not A268) );
 a46112a <=( A302  and  (not A299) );
 a46113a <=( a46112a  and  a46109a );
 a46114a <=( a46113a  and  a46106a );
 a46118a <=( (not A168)  and  (not A169) );
 a46119a <=( (not A170)  and  a46118a );
 a46122a <=( (not A232)  and  A202 );
 a46125a <=( (not A235)  and  (not A233) );
 a46126a <=( a46125a  and  a46122a );
 a46127a <=( a46126a  and  a46119a );
 a46131a <=( (not A267)  and  A266 );
 a46132a <=( A265  and  a46131a );
 a46135a <=( (not A298)  and  (not A268) );
 a46138a <=( A302  and  A299 );
 a46139a <=( a46138a  and  a46135a );
 a46140a <=( a46139a  and  a46132a );
 a46144a <=( (not A168)  and  (not A169) );
 a46145a <=( (not A170)  and  a46144a );
 a46148a <=( A201  and  A199 );
 a46151a <=( (not A235)  and  (not A234) );
 a46152a <=( a46151a  and  a46148a );
 a46153a <=( a46152a  and  a46145a );
 a46157a <=( (not A268)  and  (not A267) );
 a46158a <=( (not A236)  and  a46157a );
 a46161a <=( A298  and  (not A269) );
 a46164a <=( A302  and  (not A299) );
 a46165a <=( a46164a  and  a46161a );
 a46166a <=( a46165a  and  a46158a );
 a46170a <=( (not A168)  and  (not A169) );
 a46171a <=( (not A170)  and  a46170a );
 a46174a <=( A201  and  A199 );
 a46177a <=( (not A235)  and  (not A234) );
 a46178a <=( a46177a  and  a46174a );
 a46179a <=( a46178a  and  a46171a );
 a46183a <=( (not A268)  and  (not A267) );
 a46184a <=( (not A236)  and  a46183a );
 a46187a <=( (not A298)  and  (not A269) );
 a46190a <=( A302  and  A299 );
 a46191a <=( a46190a  and  a46187a );
 a46192a <=( a46191a  and  a46184a );
 a46196a <=( (not A168)  and  (not A169) );
 a46197a <=( (not A170)  and  a46196a );
 a46200a <=( A201  and  A199 );
 a46203a <=( (not A235)  and  (not A234) );
 a46204a <=( a46203a  and  a46200a );
 a46205a <=( a46204a  and  a46197a );
 a46209a <=( A266  and  A265 );
 a46210a <=( (not A236)  and  a46209a );
 a46213a <=( (not A268)  and  (not A267) );
 a46216a <=( A300  and  A299 );
 a46217a <=( a46216a  and  a46213a );
 a46218a <=( a46217a  and  a46210a );
 a46222a <=( (not A168)  and  (not A169) );
 a46223a <=( (not A170)  and  a46222a );
 a46226a <=( A201  and  A199 );
 a46229a <=( (not A235)  and  (not A234) );
 a46230a <=( a46229a  and  a46226a );
 a46231a <=( a46230a  and  a46223a );
 a46235a <=( A266  and  A265 );
 a46236a <=( (not A236)  and  a46235a );
 a46239a <=( (not A268)  and  (not A267) );
 a46242a <=( A300  and  A298 );
 a46243a <=( a46242a  and  a46239a );
 a46244a <=( a46243a  and  a46236a );
 a46248a <=( (not A168)  and  (not A169) );
 a46249a <=( (not A170)  and  a46248a );
 a46252a <=( A201  and  A199 );
 a46255a <=( (not A235)  and  (not A234) );
 a46256a <=( a46255a  and  a46252a );
 a46257a <=( a46256a  and  a46249a );
 a46261a <=( (not A266)  and  (not A265) );
 a46262a <=( (not A236)  and  a46261a );
 a46265a <=( A298  and  (not A268) );
 a46268a <=( A302  and  (not A299) );
 a46269a <=( a46268a  and  a46265a );
 a46270a <=( a46269a  and  a46262a );
 a46274a <=( (not A168)  and  (not A169) );
 a46275a <=( (not A170)  and  a46274a );
 a46278a <=( A201  and  A199 );
 a46281a <=( (not A235)  and  (not A234) );
 a46282a <=( a46281a  and  a46278a );
 a46283a <=( a46282a  and  a46275a );
 a46287a <=( (not A266)  and  (not A265) );
 a46288a <=( (not A236)  and  a46287a );
 a46291a <=( (not A298)  and  (not A268) );
 a46294a <=( A302  and  A299 );
 a46295a <=( a46294a  and  a46291a );
 a46296a <=( a46295a  and  a46288a );
 a46300a <=( (not A168)  and  (not A169) );
 a46301a <=( (not A170)  and  a46300a );
 a46304a <=( A201  and  A199 );
 a46307a <=( A233  and  A232 );
 a46308a <=( a46307a  and  a46304a );
 a46309a <=( a46308a  and  a46301a );
 a46313a <=( (not A267)  and  (not A235) );
 a46314a <=( (not A234)  and  a46313a );
 a46317a <=( (not A269)  and  (not A268) );
 a46320a <=( A300  and  A299 );
 a46321a <=( a46320a  and  a46317a );
 a46322a <=( a46321a  and  a46314a );
 a46326a <=( (not A168)  and  (not A169) );
 a46327a <=( (not A170)  and  a46326a );
 a46330a <=( A201  and  A199 );
 a46333a <=( A233  and  A232 );
 a46334a <=( a46333a  and  a46330a );
 a46335a <=( a46334a  and  a46327a );
 a46339a <=( (not A267)  and  (not A235) );
 a46340a <=( (not A234)  and  a46339a );
 a46343a <=( (not A269)  and  (not A268) );
 a46346a <=( A300  and  A298 );
 a46347a <=( a46346a  and  a46343a );
 a46348a <=( a46347a  and  a46340a );
 a46352a <=( (not A168)  and  (not A169) );
 a46353a <=( (not A170)  and  a46352a );
 a46356a <=( A201  and  A199 );
 a46359a <=( A233  and  A232 );
 a46360a <=( a46359a  and  a46356a );
 a46361a <=( a46360a  and  a46353a );
 a46365a <=( A265  and  (not A235) );
 a46366a <=( (not A234)  and  a46365a );
 a46369a <=( (not A267)  and  A266 );
 a46372a <=( A301  and  (not A268) );
 a46373a <=( a46372a  and  a46369a );
 a46374a <=( a46373a  and  a46366a );
 a46378a <=( (not A168)  and  (not A169) );
 a46379a <=( (not A170)  and  a46378a );
 a46382a <=( A201  and  A199 );
 a46385a <=( A233  and  A232 );
 a46386a <=( a46385a  and  a46382a );
 a46387a <=( a46386a  and  a46379a );
 a46391a <=( (not A265)  and  (not A235) );
 a46392a <=( (not A234)  and  a46391a );
 a46395a <=( (not A268)  and  (not A266) );
 a46398a <=( A300  and  A299 );
 a46399a <=( a46398a  and  a46395a );
 a46400a <=( a46399a  and  a46392a );
 a46404a <=( (not A168)  and  (not A169) );
 a46405a <=( (not A170)  and  a46404a );
 a46408a <=( A201  and  A199 );
 a46411a <=( A233  and  A232 );
 a46412a <=( a46411a  and  a46408a );
 a46413a <=( a46412a  and  a46405a );
 a46417a <=( (not A265)  and  (not A235) );
 a46418a <=( (not A234)  and  a46417a );
 a46421a <=( (not A268)  and  (not A266) );
 a46424a <=( A300  and  A298 );
 a46425a <=( a46424a  and  a46421a );
 a46426a <=( a46425a  and  a46418a );
 a46430a <=( (not A168)  and  (not A169) );
 a46431a <=( (not A170)  and  a46430a );
 a46434a <=( A201  and  A199 );
 a46437a <=( (not A233)  and  (not A232) );
 a46438a <=( a46437a  and  a46434a );
 a46439a <=( a46438a  and  a46431a );
 a46443a <=( (not A268)  and  (not A267) );
 a46444a <=( (not A235)  and  a46443a );
 a46447a <=( A298  and  (not A269) );
 a46450a <=( A302  and  (not A299) );
 a46451a <=( a46450a  and  a46447a );
 a46452a <=( a46451a  and  a46444a );
 a46456a <=( (not A168)  and  (not A169) );
 a46457a <=( (not A170)  and  a46456a );
 a46460a <=( A201  and  A199 );
 a46463a <=( (not A233)  and  (not A232) );
 a46464a <=( a46463a  and  a46460a );
 a46465a <=( a46464a  and  a46457a );
 a46469a <=( (not A268)  and  (not A267) );
 a46470a <=( (not A235)  and  a46469a );
 a46473a <=( (not A298)  and  (not A269) );
 a46476a <=( A302  and  A299 );
 a46477a <=( a46476a  and  a46473a );
 a46478a <=( a46477a  and  a46470a );
 a46482a <=( (not A168)  and  (not A169) );
 a46483a <=( (not A170)  and  a46482a );
 a46486a <=( A201  and  A199 );
 a46489a <=( (not A233)  and  (not A232) );
 a46490a <=( a46489a  and  a46486a );
 a46491a <=( a46490a  and  a46483a );
 a46495a <=( A266  and  A265 );
 a46496a <=( (not A235)  and  a46495a );
 a46499a <=( (not A268)  and  (not A267) );
 a46502a <=( A300  and  A299 );
 a46503a <=( a46502a  and  a46499a );
 a46504a <=( a46503a  and  a46496a );
 a46508a <=( (not A168)  and  (not A169) );
 a46509a <=( (not A170)  and  a46508a );
 a46512a <=( A201  and  A199 );
 a46515a <=( (not A233)  and  (not A232) );
 a46516a <=( a46515a  and  a46512a );
 a46517a <=( a46516a  and  a46509a );
 a46521a <=( A266  and  A265 );
 a46522a <=( (not A235)  and  a46521a );
 a46525a <=( (not A268)  and  (not A267) );
 a46528a <=( A300  and  A298 );
 a46529a <=( a46528a  and  a46525a );
 a46530a <=( a46529a  and  a46522a );
 a46534a <=( (not A168)  and  (not A169) );
 a46535a <=( (not A170)  and  a46534a );
 a46538a <=( A201  and  A199 );
 a46541a <=( (not A233)  and  (not A232) );
 a46542a <=( a46541a  and  a46538a );
 a46543a <=( a46542a  and  a46535a );
 a46547a <=( (not A266)  and  (not A265) );
 a46548a <=( (not A235)  and  a46547a );
 a46551a <=( A298  and  (not A268) );
 a46554a <=( A302  and  (not A299) );
 a46555a <=( a46554a  and  a46551a );
 a46556a <=( a46555a  and  a46548a );
 a46560a <=( (not A168)  and  (not A169) );
 a46561a <=( (not A170)  and  a46560a );
 a46564a <=( A201  and  A199 );
 a46567a <=( (not A233)  and  (not A232) );
 a46568a <=( a46567a  and  a46564a );
 a46569a <=( a46568a  and  a46561a );
 a46573a <=( (not A266)  and  (not A265) );
 a46574a <=( (not A235)  and  a46573a );
 a46577a <=( (not A298)  and  (not A268) );
 a46580a <=( A302  and  A299 );
 a46581a <=( a46580a  and  a46577a );
 a46582a <=( a46581a  and  a46574a );
 a46586a <=( (not A168)  and  (not A169) );
 a46587a <=( (not A170)  and  a46586a );
 a46590a <=( A201  and  A200 );
 a46593a <=( (not A235)  and  (not A234) );
 a46594a <=( a46593a  and  a46590a );
 a46595a <=( a46594a  and  a46587a );
 a46599a <=( (not A268)  and  (not A267) );
 a46600a <=( (not A236)  and  a46599a );
 a46603a <=( A298  and  (not A269) );
 a46606a <=( A302  and  (not A299) );
 a46607a <=( a46606a  and  a46603a );
 a46608a <=( a46607a  and  a46600a );
 a46612a <=( (not A168)  and  (not A169) );
 a46613a <=( (not A170)  and  a46612a );
 a46616a <=( A201  and  A200 );
 a46619a <=( (not A235)  and  (not A234) );
 a46620a <=( a46619a  and  a46616a );
 a46621a <=( a46620a  and  a46613a );
 a46625a <=( (not A268)  and  (not A267) );
 a46626a <=( (not A236)  and  a46625a );
 a46629a <=( (not A298)  and  (not A269) );
 a46632a <=( A302  and  A299 );
 a46633a <=( a46632a  and  a46629a );
 a46634a <=( a46633a  and  a46626a );
 a46638a <=( (not A168)  and  (not A169) );
 a46639a <=( (not A170)  and  a46638a );
 a46642a <=( A201  and  A200 );
 a46645a <=( (not A235)  and  (not A234) );
 a46646a <=( a46645a  and  a46642a );
 a46647a <=( a46646a  and  a46639a );
 a46651a <=( A266  and  A265 );
 a46652a <=( (not A236)  and  a46651a );
 a46655a <=( (not A268)  and  (not A267) );
 a46658a <=( A300  and  A299 );
 a46659a <=( a46658a  and  a46655a );
 a46660a <=( a46659a  and  a46652a );
 a46664a <=( (not A168)  and  (not A169) );
 a46665a <=( (not A170)  and  a46664a );
 a46668a <=( A201  and  A200 );
 a46671a <=( (not A235)  and  (not A234) );
 a46672a <=( a46671a  and  a46668a );
 a46673a <=( a46672a  and  a46665a );
 a46677a <=( A266  and  A265 );
 a46678a <=( (not A236)  and  a46677a );
 a46681a <=( (not A268)  and  (not A267) );
 a46684a <=( A300  and  A298 );
 a46685a <=( a46684a  and  a46681a );
 a46686a <=( a46685a  and  a46678a );
 a46690a <=( (not A168)  and  (not A169) );
 a46691a <=( (not A170)  and  a46690a );
 a46694a <=( A201  and  A200 );
 a46697a <=( (not A235)  and  (not A234) );
 a46698a <=( a46697a  and  a46694a );
 a46699a <=( a46698a  and  a46691a );
 a46703a <=( (not A266)  and  (not A265) );
 a46704a <=( (not A236)  and  a46703a );
 a46707a <=( A298  and  (not A268) );
 a46710a <=( A302  and  (not A299) );
 a46711a <=( a46710a  and  a46707a );
 a46712a <=( a46711a  and  a46704a );
 a46716a <=( (not A168)  and  (not A169) );
 a46717a <=( (not A170)  and  a46716a );
 a46720a <=( A201  and  A200 );
 a46723a <=( (not A235)  and  (not A234) );
 a46724a <=( a46723a  and  a46720a );
 a46725a <=( a46724a  and  a46717a );
 a46729a <=( (not A266)  and  (not A265) );
 a46730a <=( (not A236)  and  a46729a );
 a46733a <=( (not A298)  and  (not A268) );
 a46736a <=( A302  and  A299 );
 a46737a <=( a46736a  and  a46733a );
 a46738a <=( a46737a  and  a46730a );
 a46742a <=( (not A168)  and  (not A169) );
 a46743a <=( (not A170)  and  a46742a );
 a46746a <=( A201  and  A200 );
 a46749a <=( A233  and  A232 );
 a46750a <=( a46749a  and  a46746a );
 a46751a <=( a46750a  and  a46743a );
 a46755a <=( (not A267)  and  (not A235) );
 a46756a <=( (not A234)  and  a46755a );
 a46759a <=( (not A269)  and  (not A268) );
 a46762a <=( A300  and  A299 );
 a46763a <=( a46762a  and  a46759a );
 a46764a <=( a46763a  and  a46756a );
 a46768a <=( (not A168)  and  (not A169) );
 a46769a <=( (not A170)  and  a46768a );
 a46772a <=( A201  and  A200 );
 a46775a <=( A233  and  A232 );
 a46776a <=( a46775a  and  a46772a );
 a46777a <=( a46776a  and  a46769a );
 a46781a <=( (not A267)  and  (not A235) );
 a46782a <=( (not A234)  and  a46781a );
 a46785a <=( (not A269)  and  (not A268) );
 a46788a <=( A300  and  A298 );
 a46789a <=( a46788a  and  a46785a );
 a46790a <=( a46789a  and  a46782a );
 a46794a <=( (not A168)  and  (not A169) );
 a46795a <=( (not A170)  and  a46794a );
 a46798a <=( A201  and  A200 );
 a46801a <=( A233  and  A232 );
 a46802a <=( a46801a  and  a46798a );
 a46803a <=( a46802a  and  a46795a );
 a46807a <=( A265  and  (not A235) );
 a46808a <=( (not A234)  and  a46807a );
 a46811a <=( (not A267)  and  A266 );
 a46814a <=( A301  and  (not A268) );
 a46815a <=( a46814a  and  a46811a );
 a46816a <=( a46815a  and  a46808a );
 a46820a <=( (not A168)  and  (not A169) );
 a46821a <=( (not A170)  and  a46820a );
 a46824a <=( A201  and  A200 );
 a46827a <=( A233  and  A232 );
 a46828a <=( a46827a  and  a46824a );
 a46829a <=( a46828a  and  a46821a );
 a46833a <=( (not A265)  and  (not A235) );
 a46834a <=( (not A234)  and  a46833a );
 a46837a <=( (not A268)  and  (not A266) );
 a46840a <=( A300  and  A299 );
 a46841a <=( a46840a  and  a46837a );
 a46842a <=( a46841a  and  a46834a );
 a46846a <=( (not A168)  and  (not A169) );
 a46847a <=( (not A170)  and  a46846a );
 a46850a <=( A201  and  A200 );
 a46853a <=( A233  and  A232 );
 a46854a <=( a46853a  and  a46850a );
 a46855a <=( a46854a  and  a46847a );
 a46859a <=( (not A265)  and  (not A235) );
 a46860a <=( (not A234)  and  a46859a );
 a46863a <=( (not A268)  and  (not A266) );
 a46866a <=( A300  and  A298 );
 a46867a <=( a46866a  and  a46863a );
 a46868a <=( a46867a  and  a46860a );
 a46872a <=( (not A168)  and  (not A169) );
 a46873a <=( (not A170)  and  a46872a );
 a46876a <=( A201  and  A200 );
 a46879a <=( (not A233)  and  (not A232) );
 a46880a <=( a46879a  and  a46876a );
 a46881a <=( a46880a  and  a46873a );
 a46885a <=( (not A268)  and  (not A267) );
 a46886a <=( (not A235)  and  a46885a );
 a46889a <=( A298  and  (not A269) );
 a46892a <=( A302  and  (not A299) );
 a46893a <=( a46892a  and  a46889a );
 a46894a <=( a46893a  and  a46886a );
 a46898a <=( (not A168)  and  (not A169) );
 a46899a <=( (not A170)  and  a46898a );
 a46902a <=( A201  and  A200 );
 a46905a <=( (not A233)  and  (not A232) );
 a46906a <=( a46905a  and  a46902a );
 a46907a <=( a46906a  and  a46899a );
 a46911a <=( (not A268)  and  (not A267) );
 a46912a <=( (not A235)  and  a46911a );
 a46915a <=( (not A298)  and  (not A269) );
 a46918a <=( A302  and  A299 );
 a46919a <=( a46918a  and  a46915a );
 a46920a <=( a46919a  and  a46912a );
 a46924a <=( (not A168)  and  (not A169) );
 a46925a <=( (not A170)  and  a46924a );
 a46928a <=( A201  and  A200 );
 a46931a <=( (not A233)  and  (not A232) );
 a46932a <=( a46931a  and  a46928a );
 a46933a <=( a46932a  and  a46925a );
 a46937a <=( A266  and  A265 );
 a46938a <=( (not A235)  and  a46937a );
 a46941a <=( (not A268)  and  (not A267) );
 a46944a <=( A300  and  A299 );
 a46945a <=( a46944a  and  a46941a );
 a46946a <=( a46945a  and  a46938a );
 a46950a <=( (not A168)  and  (not A169) );
 a46951a <=( (not A170)  and  a46950a );
 a46954a <=( A201  and  A200 );
 a46957a <=( (not A233)  and  (not A232) );
 a46958a <=( a46957a  and  a46954a );
 a46959a <=( a46958a  and  a46951a );
 a46963a <=( A266  and  A265 );
 a46964a <=( (not A235)  and  a46963a );
 a46967a <=( (not A268)  and  (not A267) );
 a46970a <=( A300  and  A298 );
 a46971a <=( a46970a  and  a46967a );
 a46972a <=( a46971a  and  a46964a );
 a46976a <=( (not A168)  and  (not A169) );
 a46977a <=( (not A170)  and  a46976a );
 a46980a <=( A201  and  A200 );
 a46983a <=( (not A233)  and  (not A232) );
 a46984a <=( a46983a  and  a46980a );
 a46985a <=( a46984a  and  a46977a );
 a46989a <=( (not A266)  and  (not A265) );
 a46990a <=( (not A235)  and  a46989a );
 a46993a <=( A298  and  (not A268) );
 a46996a <=( A302  and  (not A299) );
 a46997a <=( a46996a  and  a46993a );
 a46998a <=( a46997a  and  a46990a );
 a47002a <=( (not A168)  and  (not A169) );
 a47003a <=( (not A170)  and  a47002a );
 a47006a <=( A201  and  A200 );
 a47009a <=( (not A233)  and  (not A232) );
 a47010a <=( a47009a  and  a47006a );
 a47011a <=( a47010a  and  a47003a );
 a47015a <=( (not A266)  and  (not A265) );
 a47016a <=( (not A235)  and  a47015a );
 a47019a <=( (not A298)  and  (not A268) );
 a47022a <=( A302  and  A299 );
 a47023a <=( a47022a  and  a47019a );
 a47024a <=( a47023a  and  a47016a );
 a47028a <=( (not A168)  and  (not A169) );
 a47029a <=( (not A170)  and  a47028a );
 a47032a <=( A200  and  (not A199) );
 a47035a <=( (not A234)  and  A203 );
 a47036a <=( a47035a  and  a47032a );
 a47037a <=( a47036a  and  a47029a );
 a47041a <=( (not A267)  and  (not A236) );
 a47042a <=( (not A235)  and  a47041a );
 a47045a <=( (not A269)  and  (not A268) );
 a47048a <=( A300  and  A299 );
 a47049a <=( a47048a  and  a47045a );
 a47050a <=( a47049a  and  a47042a );
 a47054a <=( (not A168)  and  (not A169) );
 a47055a <=( (not A170)  and  a47054a );
 a47058a <=( A200  and  (not A199) );
 a47061a <=( (not A234)  and  A203 );
 a47062a <=( a47061a  and  a47058a );
 a47063a <=( a47062a  and  a47055a );
 a47067a <=( (not A267)  and  (not A236) );
 a47068a <=( (not A235)  and  a47067a );
 a47071a <=( (not A269)  and  (not A268) );
 a47074a <=( A300  and  A298 );
 a47075a <=( a47074a  and  a47071a );
 a47076a <=( a47075a  and  a47068a );
 a47080a <=( (not A168)  and  (not A169) );
 a47081a <=( (not A170)  and  a47080a );
 a47084a <=( A200  and  (not A199) );
 a47087a <=( (not A234)  and  A203 );
 a47088a <=( a47087a  and  a47084a );
 a47089a <=( a47088a  and  a47081a );
 a47093a <=( A265  and  (not A236) );
 a47094a <=( (not A235)  and  a47093a );
 a47097a <=( (not A267)  and  A266 );
 a47100a <=( A301  and  (not A268) );
 a47101a <=( a47100a  and  a47097a );
 a47102a <=( a47101a  and  a47094a );
 a47106a <=( (not A168)  and  (not A169) );
 a47107a <=( (not A170)  and  a47106a );
 a47110a <=( A200  and  (not A199) );
 a47113a <=( (not A234)  and  A203 );
 a47114a <=( a47113a  and  a47110a );
 a47115a <=( a47114a  and  a47107a );
 a47119a <=( (not A265)  and  (not A236) );
 a47120a <=( (not A235)  and  a47119a );
 a47123a <=( (not A268)  and  (not A266) );
 a47126a <=( A300  and  A299 );
 a47127a <=( a47126a  and  a47123a );
 a47128a <=( a47127a  and  a47120a );
 a47132a <=( (not A168)  and  (not A169) );
 a47133a <=( (not A170)  and  a47132a );
 a47136a <=( A200  and  (not A199) );
 a47139a <=( (not A234)  and  A203 );
 a47140a <=( a47139a  and  a47136a );
 a47141a <=( a47140a  and  a47133a );
 a47145a <=( (not A265)  and  (not A236) );
 a47146a <=( (not A235)  and  a47145a );
 a47149a <=( (not A268)  and  (not A266) );
 a47152a <=( A300  and  A298 );
 a47153a <=( a47152a  and  a47149a );
 a47154a <=( a47153a  and  a47146a );
 a47158a <=( (not A168)  and  (not A169) );
 a47159a <=( (not A170)  and  a47158a );
 a47162a <=( A200  and  (not A199) );
 a47165a <=( A232  and  A203 );
 a47166a <=( a47165a  and  a47162a );
 a47167a <=( a47166a  and  a47159a );
 a47171a <=( (not A235)  and  (not A234) );
 a47172a <=( A233  and  a47171a );
 a47175a <=( (not A268)  and  (not A267) );
 a47178a <=( A301  and  (not A269) );
 a47179a <=( a47178a  and  a47175a );
 a47180a <=( a47179a  and  a47172a );
 a47184a <=( (not A168)  and  (not A169) );
 a47185a <=( (not A170)  and  a47184a );
 a47188a <=( A200  and  (not A199) );
 a47191a <=( A232  and  A203 );
 a47192a <=( a47191a  and  a47188a );
 a47193a <=( a47192a  and  a47185a );
 a47197a <=( (not A235)  and  (not A234) );
 a47198a <=( A233  and  a47197a );
 a47201a <=( (not A266)  and  (not A265) );
 a47204a <=( A301  and  (not A268) );
 a47205a <=( a47204a  and  a47201a );
 a47206a <=( a47205a  and  a47198a );
 a47210a <=( (not A168)  and  (not A169) );
 a47211a <=( (not A170)  and  a47210a );
 a47214a <=( A200  and  (not A199) );
 a47217a <=( (not A232)  and  A203 );
 a47218a <=( a47217a  and  a47214a );
 a47219a <=( a47218a  and  a47211a );
 a47223a <=( (not A267)  and  (not A235) );
 a47224a <=( (not A233)  and  a47223a );
 a47227a <=( (not A269)  and  (not A268) );
 a47230a <=( A300  and  A299 );
 a47231a <=( a47230a  and  a47227a );
 a47232a <=( a47231a  and  a47224a );
 a47236a <=( (not A168)  and  (not A169) );
 a47237a <=( (not A170)  and  a47236a );
 a47240a <=( A200  and  (not A199) );
 a47243a <=( (not A232)  and  A203 );
 a47244a <=( a47243a  and  a47240a );
 a47245a <=( a47244a  and  a47237a );
 a47249a <=( (not A267)  and  (not A235) );
 a47250a <=( (not A233)  and  a47249a );
 a47253a <=( (not A269)  and  (not A268) );
 a47256a <=( A300  and  A298 );
 a47257a <=( a47256a  and  a47253a );
 a47258a <=( a47257a  and  a47250a );
 a47262a <=( (not A168)  and  (not A169) );
 a47263a <=( (not A170)  and  a47262a );
 a47266a <=( A200  and  (not A199) );
 a47269a <=( (not A232)  and  A203 );
 a47270a <=( a47269a  and  a47266a );
 a47271a <=( a47270a  and  a47263a );
 a47275a <=( A265  and  (not A235) );
 a47276a <=( (not A233)  and  a47275a );
 a47279a <=( (not A267)  and  A266 );
 a47282a <=( A301  and  (not A268) );
 a47283a <=( a47282a  and  a47279a );
 a47284a <=( a47283a  and  a47276a );
 a47288a <=( (not A168)  and  (not A169) );
 a47289a <=( (not A170)  and  a47288a );
 a47292a <=( A200  and  (not A199) );
 a47295a <=( (not A232)  and  A203 );
 a47296a <=( a47295a  and  a47292a );
 a47297a <=( a47296a  and  a47289a );
 a47301a <=( (not A265)  and  (not A235) );
 a47302a <=( (not A233)  and  a47301a );
 a47305a <=( (not A268)  and  (not A266) );
 a47308a <=( A300  and  A299 );
 a47309a <=( a47308a  and  a47305a );
 a47310a <=( a47309a  and  a47302a );
 a47314a <=( (not A168)  and  (not A169) );
 a47315a <=( (not A170)  and  a47314a );
 a47318a <=( A200  and  (not A199) );
 a47321a <=( (not A232)  and  A203 );
 a47322a <=( a47321a  and  a47318a );
 a47323a <=( a47322a  and  a47315a );
 a47327a <=( (not A265)  and  (not A235) );
 a47328a <=( (not A233)  and  a47327a );
 a47331a <=( (not A268)  and  (not A266) );
 a47334a <=( A300  and  A298 );
 a47335a <=( a47334a  and  a47331a );
 a47336a <=( a47335a  and  a47328a );
 a47340a <=( (not A168)  and  (not A169) );
 a47341a <=( (not A170)  and  a47340a );
 a47344a <=( (not A200)  and  A199 );
 a47347a <=( (not A234)  and  A203 );
 a47348a <=( a47347a  and  a47344a );
 a47349a <=( a47348a  and  a47341a );
 a47353a <=( (not A267)  and  (not A236) );
 a47354a <=( (not A235)  and  a47353a );
 a47357a <=( (not A269)  and  (not A268) );
 a47360a <=( A300  and  A299 );
 a47361a <=( a47360a  and  a47357a );
 a47362a <=( a47361a  and  a47354a );
 a47366a <=( (not A168)  and  (not A169) );
 a47367a <=( (not A170)  and  a47366a );
 a47370a <=( (not A200)  and  A199 );
 a47373a <=( (not A234)  and  A203 );
 a47374a <=( a47373a  and  a47370a );
 a47375a <=( a47374a  and  a47367a );
 a47379a <=( (not A267)  and  (not A236) );
 a47380a <=( (not A235)  and  a47379a );
 a47383a <=( (not A269)  and  (not A268) );
 a47386a <=( A300  and  A298 );
 a47387a <=( a47386a  and  a47383a );
 a47388a <=( a47387a  and  a47380a );
 a47392a <=( (not A168)  and  (not A169) );
 a47393a <=( (not A170)  and  a47392a );
 a47396a <=( (not A200)  and  A199 );
 a47399a <=( (not A234)  and  A203 );
 a47400a <=( a47399a  and  a47396a );
 a47401a <=( a47400a  and  a47393a );
 a47405a <=( A265  and  (not A236) );
 a47406a <=( (not A235)  and  a47405a );
 a47409a <=( (not A267)  and  A266 );
 a47412a <=( A301  and  (not A268) );
 a47413a <=( a47412a  and  a47409a );
 a47414a <=( a47413a  and  a47406a );
 a47418a <=( (not A168)  and  (not A169) );
 a47419a <=( (not A170)  and  a47418a );
 a47422a <=( (not A200)  and  A199 );
 a47425a <=( (not A234)  and  A203 );
 a47426a <=( a47425a  and  a47422a );
 a47427a <=( a47426a  and  a47419a );
 a47431a <=( (not A265)  and  (not A236) );
 a47432a <=( (not A235)  and  a47431a );
 a47435a <=( (not A268)  and  (not A266) );
 a47438a <=( A300  and  A299 );
 a47439a <=( a47438a  and  a47435a );
 a47440a <=( a47439a  and  a47432a );
 a47444a <=( (not A168)  and  (not A169) );
 a47445a <=( (not A170)  and  a47444a );
 a47448a <=( (not A200)  and  A199 );
 a47451a <=( (not A234)  and  A203 );
 a47452a <=( a47451a  and  a47448a );
 a47453a <=( a47452a  and  a47445a );
 a47457a <=( (not A265)  and  (not A236) );
 a47458a <=( (not A235)  and  a47457a );
 a47461a <=( (not A268)  and  (not A266) );
 a47464a <=( A300  and  A298 );
 a47465a <=( a47464a  and  a47461a );
 a47466a <=( a47465a  and  a47458a );
 a47470a <=( (not A168)  and  (not A169) );
 a47471a <=( (not A170)  and  a47470a );
 a47474a <=( (not A200)  and  A199 );
 a47477a <=( A232  and  A203 );
 a47478a <=( a47477a  and  a47474a );
 a47479a <=( a47478a  and  a47471a );
 a47483a <=( (not A235)  and  (not A234) );
 a47484a <=( A233  and  a47483a );
 a47487a <=( (not A268)  and  (not A267) );
 a47490a <=( A301  and  (not A269) );
 a47491a <=( a47490a  and  a47487a );
 a47492a <=( a47491a  and  a47484a );
 a47496a <=( (not A168)  and  (not A169) );
 a47497a <=( (not A170)  and  a47496a );
 a47500a <=( (not A200)  and  A199 );
 a47503a <=( A232  and  A203 );
 a47504a <=( a47503a  and  a47500a );
 a47505a <=( a47504a  and  a47497a );
 a47509a <=( (not A235)  and  (not A234) );
 a47510a <=( A233  and  a47509a );
 a47513a <=( (not A266)  and  (not A265) );
 a47516a <=( A301  and  (not A268) );
 a47517a <=( a47516a  and  a47513a );
 a47518a <=( a47517a  and  a47510a );
 a47522a <=( (not A168)  and  (not A169) );
 a47523a <=( (not A170)  and  a47522a );
 a47526a <=( (not A200)  and  A199 );
 a47529a <=( (not A232)  and  A203 );
 a47530a <=( a47529a  and  a47526a );
 a47531a <=( a47530a  and  a47523a );
 a47535a <=( (not A267)  and  (not A235) );
 a47536a <=( (not A233)  and  a47535a );
 a47539a <=( (not A269)  and  (not A268) );
 a47542a <=( A300  and  A299 );
 a47543a <=( a47542a  and  a47539a );
 a47544a <=( a47543a  and  a47536a );
 a47548a <=( (not A168)  and  (not A169) );
 a47549a <=( (not A170)  and  a47548a );
 a47552a <=( (not A200)  and  A199 );
 a47555a <=( (not A232)  and  A203 );
 a47556a <=( a47555a  and  a47552a );
 a47557a <=( a47556a  and  a47549a );
 a47561a <=( (not A267)  and  (not A235) );
 a47562a <=( (not A233)  and  a47561a );
 a47565a <=( (not A269)  and  (not A268) );
 a47568a <=( A300  and  A298 );
 a47569a <=( a47568a  and  a47565a );
 a47570a <=( a47569a  and  a47562a );
 a47574a <=( (not A168)  and  (not A169) );
 a47575a <=( (not A170)  and  a47574a );
 a47578a <=( (not A200)  and  A199 );
 a47581a <=( (not A232)  and  A203 );
 a47582a <=( a47581a  and  a47578a );
 a47583a <=( a47582a  and  a47575a );
 a47587a <=( A265  and  (not A235) );
 a47588a <=( (not A233)  and  a47587a );
 a47591a <=( (not A267)  and  A266 );
 a47594a <=( A301  and  (not A268) );
 a47595a <=( a47594a  and  a47591a );
 a47596a <=( a47595a  and  a47588a );
 a47600a <=( (not A168)  and  (not A169) );
 a47601a <=( (not A170)  and  a47600a );
 a47604a <=( (not A200)  and  A199 );
 a47607a <=( (not A232)  and  A203 );
 a47608a <=( a47607a  and  a47604a );
 a47609a <=( a47608a  and  a47601a );
 a47613a <=( (not A265)  and  (not A235) );
 a47614a <=( (not A233)  and  a47613a );
 a47617a <=( (not A268)  and  (not A266) );
 a47620a <=( A300  and  A299 );
 a47621a <=( a47620a  and  a47617a );
 a47622a <=( a47621a  and  a47614a );
 a47626a <=( (not A168)  and  (not A169) );
 a47627a <=( (not A170)  and  a47626a );
 a47630a <=( (not A200)  and  A199 );
 a47633a <=( (not A232)  and  A203 );
 a47634a <=( a47633a  and  a47630a );
 a47635a <=( a47634a  and  a47627a );
 a47639a <=( (not A265)  and  (not A235) );
 a47640a <=( (not A233)  and  a47639a );
 a47643a <=( (not A268)  and  (not A266) );
 a47646a <=( A300  and  A298 );
 a47647a <=( a47646a  and  a47643a );
 a47648a <=( a47647a  and  a47640a );
 a47652a <=( (not A201)  and  A166 );
 a47653a <=( A168  and  a47652a );
 a47656a <=( (not A203)  and  (not A202) );
 a47659a <=( (not A235)  and  (not A234) );
 a47660a <=( a47659a  and  a47656a );
 a47661a <=( a47660a  and  a47653a );
 a47664a <=( A265  and  (not A236) );
 a47667a <=( (not A267)  and  A266 );
 a47668a <=( a47667a  and  a47664a );
 a47671a <=( A298  and  (not A268) );
 a47674a <=( A302  and  (not A299) );
 a47675a <=( a47674a  and  a47671a );
 a47676a <=( a47675a  and  a47668a );
 a47680a <=( (not A201)  and  A166 );
 a47681a <=( A168  and  a47680a );
 a47684a <=( (not A203)  and  (not A202) );
 a47687a <=( (not A235)  and  (not A234) );
 a47688a <=( a47687a  and  a47684a );
 a47689a <=( a47688a  and  a47681a );
 a47692a <=( A265  and  (not A236) );
 a47695a <=( (not A267)  and  A266 );
 a47696a <=( a47695a  and  a47692a );
 a47699a <=( (not A298)  and  (not A268) );
 a47702a <=( A302  and  A299 );
 a47703a <=( a47702a  and  a47699a );
 a47704a <=( a47703a  and  a47696a );
 a47708a <=( (not A201)  and  A166 );
 a47709a <=( A168  and  a47708a );
 a47712a <=( (not A203)  and  (not A202) );
 a47715a <=( A233  and  A232 );
 a47716a <=( a47715a  and  a47712a );
 a47717a <=( a47716a  and  a47709a );
 a47720a <=( (not A235)  and  (not A234) );
 a47723a <=( (not A268)  and  (not A267) );
 a47724a <=( a47723a  and  a47720a );
 a47727a <=( A298  and  (not A269) );
 a47730a <=( A302  and  (not A299) );
 a47731a <=( a47730a  and  a47727a );
 a47732a <=( a47731a  and  a47724a );
 a47736a <=( (not A201)  and  A166 );
 a47737a <=( A168  and  a47736a );
 a47740a <=( (not A203)  and  (not A202) );
 a47743a <=( A233  and  A232 );
 a47744a <=( a47743a  and  a47740a );
 a47745a <=( a47744a  and  a47737a );
 a47748a <=( (not A235)  and  (not A234) );
 a47751a <=( (not A268)  and  (not A267) );
 a47752a <=( a47751a  and  a47748a );
 a47755a <=( (not A298)  and  (not A269) );
 a47758a <=( A302  and  A299 );
 a47759a <=( a47758a  and  a47755a );
 a47760a <=( a47759a  and  a47752a );
 a47764a <=( (not A201)  and  A166 );
 a47765a <=( A168  and  a47764a );
 a47768a <=( (not A203)  and  (not A202) );
 a47771a <=( A233  and  A232 );
 a47772a <=( a47771a  and  a47768a );
 a47773a <=( a47772a  and  a47765a );
 a47776a <=( (not A235)  and  (not A234) );
 a47779a <=( A266  and  A265 );
 a47780a <=( a47779a  and  a47776a );
 a47783a <=( (not A268)  and  (not A267) );
 a47786a <=( A300  and  A299 );
 a47787a <=( a47786a  and  a47783a );
 a47788a <=( a47787a  and  a47780a );
 a47792a <=( (not A201)  and  A166 );
 a47793a <=( A168  and  a47792a );
 a47796a <=( (not A203)  and  (not A202) );
 a47799a <=( A233  and  A232 );
 a47800a <=( a47799a  and  a47796a );
 a47801a <=( a47800a  and  a47793a );
 a47804a <=( (not A235)  and  (not A234) );
 a47807a <=( A266  and  A265 );
 a47808a <=( a47807a  and  a47804a );
 a47811a <=( (not A268)  and  (not A267) );
 a47814a <=( A300  and  A298 );
 a47815a <=( a47814a  and  a47811a );
 a47816a <=( a47815a  and  a47808a );
 a47820a <=( (not A201)  and  A166 );
 a47821a <=( A168  and  a47820a );
 a47824a <=( (not A203)  and  (not A202) );
 a47827a <=( A233  and  A232 );
 a47828a <=( a47827a  and  a47824a );
 a47829a <=( a47828a  and  a47821a );
 a47832a <=( (not A235)  and  (not A234) );
 a47835a <=( (not A266)  and  (not A265) );
 a47836a <=( a47835a  and  a47832a );
 a47839a <=( A298  and  (not A268) );
 a47842a <=( A302  and  (not A299) );
 a47843a <=( a47842a  and  a47839a );
 a47844a <=( a47843a  and  a47836a );
 a47848a <=( (not A201)  and  A166 );
 a47849a <=( A168  and  a47848a );
 a47852a <=( (not A203)  and  (not A202) );
 a47855a <=( A233  and  A232 );
 a47856a <=( a47855a  and  a47852a );
 a47857a <=( a47856a  and  a47849a );
 a47860a <=( (not A235)  and  (not A234) );
 a47863a <=( (not A266)  and  (not A265) );
 a47864a <=( a47863a  and  a47860a );
 a47867a <=( (not A298)  and  (not A268) );
 a47870a <=( A302  and  A299 );
 a47871a <=( a47870a  and  a47867a );
 a47872a <=( a47871a  and  a47864a );
 a47876a <=( (not A201)  and  A166 );
 a47877a <=( A168  and  a47876a );
 a47880a <=( (not A203)  and  (not A202) );
 a47883a <=( (not A233)  and  (not A232) );
 a47884a <=( a47883a  and  a47880a );
 a47885a <=( a47884a  and  a47877a );
 a47888a <=( A265  and  (not A235) );
 a47891a <=( (not A267)  and  A266 );
 a47892a <=( a47891a  and  a47888a );
 a47895a <=( A298  and  (not A268) );
 a47898a <=( A302  and  (not A299) );
 a47899a <=( a47898a  and  a47895a );
 a47900a <=( a47899a  and  a47892a );
 a47904a <=( (not A201)  and  A166 );
 a47905a <=( A168  and  a47904a );
 a47908a <=( (not A203)  and  (not A202) );
 a47911a <=( (not A233)  and  (not A232) );
 a47912a <=( a47911a  and  a47908a );
 a47913a <=( a47912a  and  a47905a );
 a47916a <=( A265  and  (not A235) );
 a47919a <=( (not A267)  and  A266 );
 a47920a <=( a47919a  and  a47916a );
 a47923a <=( (not A298)  and  (not A268) );
 a47926a <=( A302  and  A299 );
 a47927a <=( a47926a  and  a47923a );
 a47928a <=( a47927a  and  a47920a );
 a47932a <=( A199  and  A166 );
 a47933a <=( A168  and  a47932a );
 a47936a <=( (not A201)  and  A200 );
 a47939a <=( (not A234)  and  (not A202) );
 a47940a <=( a47939a  and  a47936a );
 a47941a <=( a47940a  and  a47933a );
 a47944a <=( (not A236)  and  (not A235) );
 a47947a <=( (not A268)  and  (not A267) );
 a47948a <=( a47947a  and  a47944a );
 a47951a <=( A298  and  (not A269) );
 a47954a <=( A302  and  (not A299) );
 a47955a <=( a47954a  and  a47951a );
 a47956a <=( a47955a  and  a47948a );
 a47960a <=( A199  and  A166 );
 a47961a <=( A168  and  a47960a );
 a47964a <=( (not A201)  and  A200 );
 a47967a <=( (not A234)  and  (not A202) );
 a47968a <=( a47967a  and  a47964a );
 a47969a <=( a47968a  and  a47961a );
 a47972a <=( (not A236)  and  (not A235) );
 a47975a <=( (not A268)  and  (not A267) );
 a47976a <=( a47975a  and  a47972a );
 a47979a <=( (not A298)  and  (not A269) );
 a47982a <=( A302  and  A299 );
 a47983a <=( a47982a  and  a47979a );
 a47984a <=( a47983a  and  a47976a );
 a47988a <=( A199  and  A166 );
 a47989a <=( A168  and  a47988a );
 a47992a <=( (not A201)  and  A200 );
 a47995a <=( (not A234)  and  (not A202) );
 a47996a <=( a47995a  and  a47992a );
 a47997a <=( a47996a  and  a47989a );
 a48000a <=( (not A236)  and  (not A235) );
 a48003a <=( A266  and  A265 );
 a48004a <=( a48003a  and  a48000a );
 a48007a <=( (not A268)  and  (not A267) );
 a48010a <=( A300  and  A299 );
 a48011a <=( a48010a  and  a48007a );
 a48012a <=( a48011a  and  a48004a );
 a48016a <=( A199  and  A166 );
 a48017a <=( A168  and  a48016a );
 a48020a <=( (not A201)  and  A200 );
 a48023a <=( (not A234)  and  (not A202) );
 a48024a <=( a48023a  and  a48020a );
 a48025a <=( a48024a  and  a48017a );
 a48028a <=( (not A236)  and  (not A235) );
 a48031a <=( A266  and  A265 );
 a48032a <=( a48031a  and  a48028a );
 a48035a <=( (not A268)  and  (not A267) );
 a48038a <=( A300  and  A298 );
 a48039a <=( a48038a  and  a48035a );
 a48040a <=( a48039a  and  a48032a );
 a48044a <=( A199  and  A166 );
 a48045a <=( A168  and  a48044a );
 a48048a <=( (not A201)  and  A200 );
 a48051a <=( (not A234)  and  (not A202) );
 a48052a <=( a48051a  and  a48048a );
 a48053a <=( a48052a  and  a48045a );
 a48056a <=( (not A236)  and  (not A235) );
 a48059a <=( (not A266)  and  (not A265) );
 a48060a <=( a48059a  and  a48056a );
 a48063a <=( A298  and  (not A268) );
 a48066a <=( A302  and  (not A299) );
 a48067a <=( a48066a  and  a48063a );
 a48068a <=( a48067a  and  a48060a );
 a48072a <=( A199  and  A166 );
 a48073a <=( A168  and  a48072a );
 a48076a <=( (not A201)  and  A200 );
 a48079a <=( (not A234)  and  (not A202) );
 a48080a <=( a48079a  and  a48076a );
 a48081a <=( a48080a  and  a48073a );
 a48084a <=( (not A236)  and  (not A235) );
 a48087a <=( (not A266)  and  (not A265) );
 a48088a <=( a48087a  and  a48084a );
 a48091a <=( (not A298)  and  (not A268) );
 a48094a <=( A302  and  A299 );
 a48095a <=( a48094a  and  a48091a );
 a48096a <=( a48095a  and  a48088a );
 a48100a <=( A199  and  A166 );
 a48101a <=( A168  and  a48100a );
 a48104a <=( (not A201)  and  A200 );
 a48107a <=( A232  and  (not A202) );
 a48108a <=( a48107a  and  a48104a );
 a48109a <=( a48108a  and  a48101a );
 a48112a <=( (not A234)  and  A233 );
 a48115a <=( (not A267)  and  (not A235) );
 a48116a <=( a48115a  and  a48112a );
 a48119a <=( (not A269)  and  (not A268) );
 a48122a <=( A300  and  A299 );
 a48123a <=( a48122a  and  a48119a );
 a48124a <=( a48123a  and  a48116a );
 a48128a <=( A199  and  A166 );
 a48129a <=( A168  and  a48128a );
 a48132a <=( (not A201)  and  A200 );
 a48135a <=( A232  and  (not A202) );
 a48136a <=( a48135a  and  a48132a );
 a48137a <=( a48136a  and  a48129a );
 a48140a <=( (not A234)  and  A233 );
 a48143a <=( (not A267)  and  (not A235) );
 a48144a <=( a48143a  and  a48140a );
 a48147a <=( (not A269)  and  (not A268) );
 a48150a <=( A300  and  A298 );
 a48151a <=( a48150a  and  a48147a );
 a48152a <=( a48151a  and  a48144a );
 a48156a <=( A199  and  A166 );
 a48157a <=( A168  and  a48156a );
 a48160a <=( (not A201)  and  A200 );
 a48163a <=( A232  and  (not A202) );
 a48164a <=( a48163a  and  a48160a );
 a48165a <=( a48164a  and  a48157a );
 a48168a <=( (not A234)  and  A233 );
 a48171a <=( A265  and  (not A235) );
 a48172a <=( a48171a  and  a48168a );
 a48175a <=( (not A267)  and  A266 );
 a48178a <=( A301  and  (not A268) );
 a48179a <=( a48178a  and  a48175a );
 a48180a <=( a48179a  and  a48172a );
 a48184a <=( A199  and  A166 );
 a48185a <=( A168  and  a48184a );
 a48188a <=( (not A201)  and  A200 );
 a48191a <=( A232  and  (not A202) );
 a48192a <=( a48191a  and  a48188a );
 a48193a <=( a48192a  and  a48185a );
 a48196a <=( (not A234)  and  A233 );
 a48199a <=( (not A265)  and  (not A235) );
 a48200a <=( a48199a  and  a48196a );
 a48203a <=( (not A268)  and  (not A266) );
 a48206a <=( A300  and  A299 );
 a48207a <=( a48206a  and  a48203a );
 a48208a <=( a48207a  and  a48200a );
 a48212a <=( A199  and  A166 );
 a48213a <=( A168  and  a48212a );
 a48216a <=( (not A201)  and  A200 );
 a48219a <=( A232  and  (not A202) );
 a48220a <=( a48219a  and  a48216a );
 a48221a <=( a48220a  and  a48213a );
 a48224a <=( (not A234)  and  A233 );
 a48227a <=( (not A265)  and  (not A235) );
 a48228a <=( a48227a  and  a48224a );
 a48231a <=( (not A268)  and  (not A266) );
 a48234a <=( A300  and  A298 );
 a48235a <=( a48234a  and  a48231a );
 a48236a <=( a48235a  and  a48228a );
 a48240a <=( A199  and  A166 );
 a48241a <=( A168  and  a48240a );
 a48244a <=( (not A201)  and  A200 );
 a48247a <=( (not A232)  and  (not A202) );
 a48248a <=( a48247a  and  a48244a );
 a48249a <=( a48248a  and  a48241a );
 a48252a <=( (not A235)  and  (not A233) );
 a48255a <=( (not A268)  and  (not A267) );
 a48256a <=( a48255a  and  a48252a );
 a48259a <=( A298  and  (not A269) );
 a48262a <=( A302  and  (not A299) );
 a48263a <=( a48262a  and  a48259a );
 a48264a <=( a48263a  and  a48256a );
 a48268a <=( A199  and  A166 );
 a48269a <=( A168  and  a48268a );
 a48272a <=( (not A201)  and  A200 );
 a48275a <=( (not A232)  and  (not A202) );
 a48276a <=( a48275a  and  a48272a );
 a48277a <=( a48276a  and  a48269a );
 a48280a <=( (not A235)  and  (not A233) );
 a48283a <=( (not A268)  and  (not A267) );
 a48284a <=( a48283a  and  a48280a );
 a48287a <=( (not A298)  and  (not A269) );
 a48290a <=( A302  and  A299 );
 a48291a <=( a48290a  and  a48287a );
 a48292a <=( a48291a  and  a48284a );
 a48296a <=( A199  and  A166 );
 a48297a <=( A168  and  a48296a );
 a48300a <=( (not A201)  and  A200 );
 a48303a <=( (not A232)  and  (not A202) );
 a48304a <=( a48303a  and  a48300a );
 a48305a <=( a48304a  and  a48297a );
 a48308a <=( (not A235)  and  (not A233) );
 a48311a <=( A266  and  A265 );
 a48312a <=( a48311a  and  a48308a );
 a48315a <=( (not A268)  and  (not A267) );
 a48318a <=( A300  and  A299 );
 a48319a <=( a48318a  and  a48315a );
 a48320a <=( a48319a  and  a48312a );
 a48324a <=( A199  and  A166 );
 a48325a <=( A168  and  a48324a );
 a48328a <=( (not A201)  and  A200 );
 a48331a <=( (not A232)  and  (not A202) );
 a48332a <=( a48331a  and  a48328a );
 a48333a <=( a48332a  and  a48325a );
 a48336a <=( (not A235)  and  (not A233) );
 a48339a <=( A266  and  A265 );
 a48340a <=( a48339a  and  a48336a );
 a48343a <=( (not A268)  and  (not A267) );
 a48346a <=( A300  and  A298 );
 a48347a <=( a48346a  and  a48343a );
 a48348a <=( a48347a  and  a48340a );
 a48352a <=( A199  and  A166 );
 a48353a <=( A168  and  a48352a );
 a48356a <=( (not A201)  and  A200 );
 a48359a <=( (not A232)  and  (not A202) );
 a48360a <=( a48359a  and  a48356a );
 a48361a <=( a48360a  and  a48353a );
 a48364a <=( (not A235)  and  (not A233) );
 a48367a <=( (not A266)  and  (not A265) );
 a48368a <=( a48367a  and  a48364a );
 a48371a <=( A298  and  (not A268) );
 a48374a <=( A302  and  (not A299) );
 a48375a <=( a48374a  and  a48371a );
 a48376a <=( a48375a  and  a48368a );
 a48380a <=( A199  and  A166 );
 a48381a <=( A168  and  a48380a );
 a48384a <=( (not A201)  and  A200 );
 a48387a <=( (not A232)  and  (not A202) );
 a48388a <=( a48387a  and  a48384a );
 a48389a <=( a48388a  and  a48381a );
 a48392a <=( (not A235)  and  (not A233) );
 a48395a <=( (not A266)  and  (not A265) );
 a48396a <=( a48395a  and  a48392a );
 a48399a <=( (not A298)  and  (not A268) );
 a48402a <=( A302  and  A299 );
 a48403a <=( a48402a  and  a48399a );
 a48404a <=( a48403a  and  a48396a );
 a48408a <=( (not A199)  and  A166 );
 a48409a <=( A168  and  a48408a );
 a48412a <=( (not A202)  and  (not A200) );
 a48415a <=( (not A235)  and  (not A234) );
 a48416a <=( a48415a  and  a48412a );
 a48417a <=( a48416a  and  a48409a );
 a48420a <=( A265  and  (not A236) );
 a48423a <=( (not A267)  and  A266 );
 a48424a <=( a48423a  and  a48420a );
 a48427a <=( A298  and  (not A268) );
 a48430a <=( A302  and  (not A299) );
 a48431a <=( a48430a  and  a48427a );
 a48432a <=( a48431a  and  a48424a );
 a48436a <=( (not A199)  and  A166 );
 a48437a <=( A168  and  a48436a );
 a48440a <=( (not A202)  and  (not A200) );
 a48443a <=( (not A235)  and  (not A234) );
 a48444a <=( a48443a  and  a48440a );
 a48445a <=( a48444a  and  a48437a );
 a48448a <=( A265  and  (not A236) );
 a48451a <=( (not A267)  and  A266 );
 a48452a <=( a48451a  and  a48448a );
 a48455a <=( (not A298)  and  (not A268) );
 a48458a <=( A302  and  A299 );
 a48459a <=( a48458a  and  a48455a );
 a48460a <=( a48459a  and  a48452a );
 a48464a <=( (not A199)  and  A166 );
 a48465a <=( A168  and  a48464a );
 a48468a <=( (not A202)  and  (not A200) );
 a48471a <=( A233  and  A232 );
 a48472a <=( a48471a  and  a48468a );
 a48473a <=( a48472a  and  a48465a );
 a48476a <=( (not A235)  and  (not A234) );
 a48479a <=( (not A268)  and  (not A267) );
 a48480a <=( a48479a  and  a48476a );
 a48483a <=( A298  and  (not A269) );
 a48486a <=( A302  and  (not A299) );
 a48487a <=( a48486a  and  a48483a );
 a48488a <=( a48487a  and  a48480a );
 a48492a <=( (not A199)  and  A166 );
 a48493a <=( A168  and  a48492a );
 a48496a <=( (not A202)  and  (not A200) );
 a48499a <=( A233  and  A232 );
 a48500a <=( a48499a  and  a48496a );
 a48501a <=( a48500a  and  a48493a );
 a48504a <=( (not A235)  and  (not A234) );
 a48507a <=( (not A268)  and  (not A267) );
 a48508a <=( a48507a  and  a48504a );
 a48511a <=( (not A298)  and  (not A269) );
 a48514a <=( A302  and  A299 );
 a48515a <=( a48514a  and  a48511a );
 a48516a <=( a48515a  and  a48508a );
 a48520a <=( (not A199)  and  A166 );
 a48521a <=( A168  and  a48520a );
 a48524a <=( (not A202)  and  (not A200) );
 a48527a <=( A233  and  A232 );
 a48528a <=( a48527a  and  a48524a );
 a48529a <=( a48528a  and  a48521a );
 a48532a <=( (not A235)  and  (not A234) );
 a48535a <=( A266  and  A265 );
 a48536a <=( a48535a  and  a48532a );
 a48539a <=( (not A268)  and  (not A267) );
 a48542a <=( A300  and  A299 );
 a48543a <=( a48542a  and  a48539a );
 a48544a <=( a48543a  and  a48536a );
 a48548a <=( (not A199)  and  A166 );
 a48549a <=( A168  and  a48548a );
 a48552a <=( (not A202)  and  (not A200) );
 a48555a <=( A233  and  A232 );
 a48556a <=( a48555a  and  a48552a );
 a48557a <=( a48556a  and  a48549a );
 a48560a <=( (not A235)  and  (not A234) );
 a48563a <=( A266  and  A265 );
 a48564a <=( a48563a  and  a48560a );
 a48567a <=( (not A268)  and  (not A267) );
 a48570a <=( A300  and  A298 );
 a48571a <=( a48570a  and  a48567a );
 a48572a <=( a48571a  and  a48564a );
 a48576a <=( (not A199)  and  A166 );
 a48577a <=( A168  and  a48576a );
 a48580a <=( (not A202)  and  (not A200) );
 a48583a <=( A233  and  A232 );
 a48584a <=( a48583a  and  a48580a );
 a48585a <=( a48584a  and  a48577a );
 a48588a <=( (not A235)  and  (not A234) );
 a48591a <=( (not A266)  and  (not A265) );
 a48592a <=( a48591a  and  a48588a );
 a48595a <=( A298  and  (not A268) );
 a48598a <=( A302  and  (not A299) );
 a48599a <=( a48598a  and  a48595a );
 a48600a <=( a48599a  and  a48592a );
 a48604a <=( (not A199)  and  A166 );
 a48605a <=( A168  and  a48604a );
 a48608a <=( (not A202)  and  (not A200) );
 a48611a <=( A233  and  A232 );
 a48612a <=( a48611a  and  a48608a );
 a48613a <=( a48612a  and  a48605a );
 a48616a <=( (not A235)  and  (not A234) );
 a48619a <=( (not A266)  and  (not A265) );
 a48620a <=( a48619a  and  a48616a );
 a48623a <=( (not A298)  and  (not A268) );
 a48626a <=( A302  and  A299 );
 a48627a <=( a48626a  and  a48623a );
 a48628a <=( a48627a  and  a48620a );
 a48632a <=( (not A199)  and  A166 );
 a48633a <=( A168  and  a48632a );
 a48636a <=( (not A202)  and  (not A200) );
 a48639a <=( (not A233)  and  (not A232) );
 a48640a <=( a48639a  and  a48636a );
 a48641a <=( a48640a  and  a48633a );
 a48644a <=( A265  and  (not A235) );
 a48647a <=( (not A267)  and  A266 );
 a48648a <=( a48647a  and  a48644a );
 a48651a <=( A298  and  (not A268) );
 a48654a <=( A302  and  (not A299) );
 a48655a <=( a48654a  and  a48651a );
 a48656a <=( a48655a  and  a48648a );
 a48660a <=( (not A199)  and  A166 );
 a48661a <=( A168  and  a48660a );
 a48664a <=( (not A202)  and  (not A200) );
 a48667a <=( (not A233)  and  (not A232) );
 a48668a <=( a48667a  and  a48664a );
 a48669a <=( a48668a  and  a48661a );
 a48672a <=( A265  and  (not A235) );
 a48675a <=( (not A267)  and  A266 );
 a48676a <=( a48675a  and  a48672a );
 a48679a <=( (not A298)  and  (not A268) );
 a48682a <=( A302  and  A299 );
 a48683a <=( a48682a  and  a48679a );
 a48684a <=( a48683a  and  a48676a );
 a48688a <=( (not A201)  and  A167 );
 a48689a <=( A168  and  a48688a );
 a48692a <=( (not A203)  and  (not A202) );
 a48695a <=( (not A235)  and  (not A234) );
 a48696a <=( a48695a  and  a48692a );
 a48697a <=( a48696a  and  a48689a );
 a48700a <=( A265  and  (not A236) );
 a48703a <=( (not A267)  and  A266 );
 a48704a <=( a48703a  and  a48700a );
 a48707a <=( A298  and  (not A268) );
 a48710a <=( A302  and  (not A299) );
 a48711a <=( a48710a  and  a48707a );
 a48712a <=( a48711a  and  a48704a );
 a48716a <=( (not A201)  and  A167 );
 a48717a <=( A168  and  a48716a );
 a48720a <=( (not A203)  and  (not A202) );
 a48723a <=( (not A235)  and  (not A234) );
 a48724a <=( a48723a  and  a48720a );
 a48725a <=( a48724a  and  a48717a );
 a48728a <=( A265  and  (not A236) );
 a48731a <=( (not A267)  and  A266 );
 a48732a <=( a48731a  and  a48728a );
 a48735a <=( (not A298)  and  (not A268) );
 a48738a <=( A302  and  A299 );
 a48739a <=( a48738a  and  a48735a );
 a48740a <=( a48739a  and  a48732a );
 a48744a <=( (not A201)  and  A167 );
 a48745a <=( A168  and  a48744a );
 a48748a <=( (not A203)  and  (not A202) );
 a48751a <=( A233  and  A232 );
 a48752a <=( a48751a  and  a48748a );
 a48753a <=( a48752a  and  a48745a );
 a48756a <=( (not A235)  and  (not A234) );
 a48759a <=( (not A268)  and  (not A267) );
 a48760a <=( a48759a  and  a48756a );
 a48763a <=( A298  and  (not A269) );
 a48766a <=( A302  and  (not A299) );
 a48767a <=( a48766a  and  a48763a );
 a48768a <=( a48767a  and  a48760a );
 a48772a <=( (not A201)  and  A167 );
 a48773a <=( A168  and  a48772a );
 a48776a <=( (not A203)  and  (not A202) );
 a48779a <=( A233  and  A232 );
 a48780a <=( a48779a  and  a48776a );
 a48781a <=( a48780a  and  a48773a );
 a48784a <=( (not A235)  and  (not A234) );
 a48787a <=( (not A268)  and  (not A267) );
 a48788a <=( a48787a  and  a48784a );
 a48791a <=( (not A298)  and  (not A269) );
 a48794a <=( A302  and  A299 );
 a48795a <=( a48794a  and  a48791a );
 a48796a <=( a48795a  and  a48788a );
 a48800a <=( (not A201)  and  A167 );
 a48801a <=( A168  and  a48800a );
 a48804a <=( (not A203)  and  (not A202) );
 a48807a <=( A233  and  A232 );
 a48808a <=( a48807a  and  a48804a );
 a48809a <=( a48808a  and  a48801a );
 a48812a <=( (not A235)  and  (not A234) );
 a48815a <=( A266  and  A265 );
 a48816a <=( a48815a  and  a48812a );
 a48819a <=( (not A268)  and  (not A267) );
 a48822a <=( A300  and  A299 );
 a48823a <=( a48822a  and  a48819a );
 a48824a <=( a48823a  and  a48816a );
 a48828a <=( (not A201)  and  A167 );
 a48829a <=( A168  and  a48828a );
 a48832a <=( (not A203)  and  (not A202) );
 a48835a <=( A233  and  A232 );
 a48836a <=( a48835a  and  a48832a );
 a48837a <=( a48836a  and  a48829a );
 a48840a <=( (not A235)  and  (not A234) );
 a48843a <=( A266  and  A265 );
 a48844a <=( a48843a  and  a48840a );
 a48847a <=( (not A268)  and  (not A267) );
 a48850a <=( A300  and  A298 );
 a48851a <=( a48850a  and  a48847a );
 a48852a <=( a48851a  and  a48844a );
 a48856a <=( (not A201)  and  A167 );
 a48857a <=( A168  and  a48856a );
 a48860a <=( (not A203)  and  (not A202) );
 a48863a <=( A233  and  A232 );
 a48864a <=( a48863a  and  a48860a );
 a48865a <=( a48864a  and  a48857a );
 a48868a <=( (not A235)  and  (not A234) );
 a48871a <=( (not A266)  and  (not A265) );
 a48872a <=( a48871a  and  a48868a );
 a48875a <=( A298  and  (not A268) );
 a48878a <=( A302  and  (not A299) );
 a48879a <=( a48878a  and  a48875a );
 a48880a <=( a48879a  and  a48872a );
 a48884a <=( (not A201)  and  A167 );
 a48885a <=( A168  and  a48884a );
 a48888a <=( (not A203)  and  (not A202) );
 a48891a <=( A233  and  A232 );
 a48892a <=( a48891a  and  a48888a );
 a48893a <=( a48892a  and  a48885a );
 a48896a <=( (not A235)  and  (not A234) );
 a48899a <=( (not A266)  and  (not A265) );
 a48900a <=( a48899a  and  a48896a );
 a48903a <=( (not A298)  and  (not A268) );
 a48906a <=( A302  and  A299 );
 a48907a <=( a48906a  and  a48903a );
 a48908a <=( a48907a  and  a48900a );
 a48912a <=( (not A201)  and  A167 );
 a48913a <=( A168  and  a48912a );
 a48916a <=( (not A203)  and  (not A202) );
 a48919a <=( (not A233)  and  (not A232) );
 a48920a <=( a48919a  and  a48916a );
 a48921a <=( a48920a  and  a48913a );
 a48924a <=( A265  and  (not A235) );
 a48927a <=( (not A267)  and  A266 );
 a48928a <=( a48927a  and  a48924a );
 a48931a <=( A298  and  (not A268) );
 a48934a <=( A302  and  (not A299) );
 a48935a <=( a48934a  and  a48931a );
 a48936a <=( a48935a  and  a48928a );
 a48940a <=( (not A201)  and  A167 );
 a48941a <=( A168  and  a48940a );
 a48944a <=( (not A203)  and  (not A202) );
 a48947a <=( (not A233)  and  (not A232) );
 a48948a <=( a48947a  and  a48944a );
 a48949a <=( a48948a  and  a48941a );
 a48952a <=( A265  and  (not A235) );
 a48955a <=( (not A267)  and  A266 );
 a48956a <=( a48955a  and  a48952a );
 a48959a <=( (not A298)  and  (not A268) );
 a48962a <=( A302  and  A299 );
 a48963a <=( a48962a  and  a48959a );
 a48964a <=( a48963a  and  a48956a );
 a48968a <=( A199  and  A167 );
 a48969a <=( A168  and  a48968a );
 a48972a <=( (not A201)  and  A200 );
 a48975a <=( (not A234)  and  (not A202) );
 a48976a <=( a48975a  and  a48972a );
 a48977a <=( a48976a  and  a48969a );
 a48980a <=( (not A236)  and  (not A235) );
 a48983a <=( (not A268)  and  (not A267) );
 a48984a <=( a48983a  and  a48980a );
 a48987a <=( A298  and  (not A269) );
 a48990a <=( A302  and  (not A299) );
 a48991a <=( a48990a  and  a48987a );
 a48992a <=( a48991a  and  a48984a );
 a48996a <=( A199  and  A167 );
 a48997a <=( A168  and  a48996a );
 a49000a <=( (not A201)  and  A200 );
 a49003a <=( (not A234)  and  (not A202) );
 a49004a <=( a49003a  and  a49000a );
 a49005a <=( a49004a  and  a48997a );
 a49008a <=( (not A236)  and  (not A235) );
 a49011a <=( (not A268)  and  (not A267) );
 a49012a <=( a49011a  and  a49008a );
 a49015a <=( (not A298)  and  (not A269) );
 a49018a <=( A302  and  A299 );
 a49019a <=( a49018a  and  a49015a );
 a49020a <=( a49019a  and  a49012a );
 a49024a <=( A199  and  A167 );
 a49025a <=( A168  and  a49024a );
 a49028a <=( (not A201)  and  A200 );
 a49031a <=( (not A234)  and  (not A202) );
 a49032a <=( a49031a  and  a49028a );
 a49033a <=( a49032a  and  a49025a );
 a49036a <=( (not A236)  and  (not A235) );
 a49039a <=( A266  and  A265 );
 a49040a <=( a49039a  and  a49036a );
 a49043a <=( (not A268)  and  (not A267) );
 a49046a <=( A300  and  A299 );
 a49047a <=( a49046a  and  a49043a );
 a49048a <=( a49047a  and  a49040a );
 a49052a <=( A199  and  A167 );
 a49053a <=( A168  and  a49052a );
 a49056a <=( (not A201)  and  A200 );
 a49059a <=( (not A234)  and  (not A202) );
 a49060a <=( a49059a  and  a49056a );
 a49061a <=( a49060a  and  a49053a );
 a49064a <=( (not A236)  and  (not A235) );
 a49067a <=( A266  and  A265 );
 a49068a <=( a49067a  and  a49064a );
 a49071a <=( (not A268)  and  (not A267) );
 a49074a <=( A300  and  A298 );
 a49075a <=( a49074a  and  a49071a );
 a49076a <=( a49075a  and  a49068a );
 a49080a <=( A199  and  A167 );
 a49081a <=( A168  and  a49080a );
 a49084a <=( (not A201)  and  A200 );
 a49087a <=( (not A234)  and  (not A202) );
 a49088a <=( a49087a  and  a49084a );
 a49089a <=( a49088a  and  a49081a );
 a49092a <=( (not A236)  and  (not A235) );
 a49095a <=( (not A266)  and  (not A265) );
 a49096a <=( a49095a  and  a49092a );
 a49099a <=( A298  and  (not A268) );
 a49102a <=( A302  and  (not A299) );
 a49103a <=( a49102a  and  a49099a );
 a49104a <=( a49103a  and  a49096a );
 a49108a <=( A199  and  A167 );
 a49109a <=( A168  and  a49108a );
 a49112a <=( (not A201)  and  A200 );
 a49115a <=( (not A234)  and  (not A202) );
 a49116a <=( a49115a  and  a49112a );
 a49117a <=( a49116a  and  a49109a );
 a49120a <=( (not A236)  and  (not A235) );
 a49123a <=( (not A266)  and  (not A265) );
 a49124a <=( a49123a  and  a49120a );
 a49127a <=( (not A298)  and  (not A268) );
 a49130a <=( A302  and  A299 );
 a49131a <=( a49130a  and  a49127a );
 a49132a <=( a49131a  and  a49124a );
 a49136a <=( A199  and  A167 );
 a49137a <=( A168  and  a49136a );
 a49140a <=( (not A201)  and  A200 );
 a49143a <=( A232  and  (not A202) );
 a49144a <=( a49143a  and  a49140a );
 a49145a <=( a49144a  and  a49137a );
 a49148a <=( (not A234)  and  A233 );
 a49151a <=( (not A267)  and  (not A235) );
 a49152a <=( a49151a  and  a49148a );
 a49155a <=( (not A269)  and  (not A268) );
 a49158a <=( A300  and  A299 );
 a49159a <=( a49158a  and  a49155a );
 a49160a <=( a49159a  and  a49152a );
 a49164a <=( A199  and  A167 );
 a49165a <=( A168  and  a49164a );
 a49168a <=( (not A201)  and  A200 );
 a49171a <=( A232  and  (not A202) );
 a49172a <=( a49171a  and  a49168a );
 a49173a <=( a49172a  and  a49165a );
 a49176a <=( (not A234)  and  A233 );
 a49179a <=( (not A267)  and  (not A235) );
 a49180a <=( a49179a  and  a49176a );
 a49183a <=( (not A269)  and  (not A268) );
 a49186a <=( A300  and  A298 );
 a49187a <=( a49186a  and  a49183a );
 a49188a <=( a49187a  and  a49180a );
 a49192a <=( A199  and  A167 );
 a49193a <=( A168  and  a49192a );
 a49196a <=( (not A201)  and  A200 );
 a49199a <=( A232  and  (not A202) );
 a49200a <=( a49199a  and  a49196a );
 a49201a <=( a49200a  and  a49193a );
 a49204a <=( (not A234)  and  A233 );
 a49207a <=( A265  and  (not A235) );
 a49208a <=( a49207a  and  a49204a );
 a49211a <=( (not A267)  and  A266 );
 a49214a <=( A301  and  (not A268) );
 a49215a <=( a49214a  and  a49211a );
 a49216a <=( a49215a  and  a49208a );
 a49220a <=( A199  and  A167 );
 a49221a <=( A168  and  a49220a );
 a49224a <=( (not A201)  and  A200 );
 a49227a <=( A232  and  (not A202) );
 a49228a <=( a49227a  and  a49224a );
 a49229a <=( a49228a  and  a49221a );
 a49232a <=( (not A234)  and  A233 );
 a49235a <=( (not A265)  and  (not A235) );
 a49236a <=( a49235a  and  a49232a );
 a49239a <=( (not A268)  and  (not A266) );
 a49242a <=( A300  and  A299 );
 a49243a <=( a49242a  and  a49239a );
 a49244a <=( a49243a  and  a49236a );
 a49248a <=( A199  and  A167 );
 a49249a <=( A168  and  a49248a );
 a49252a <=( (not A201)  and  A200 );
 a49255a <=( A232  and  (not A202) );
 a49256a <=( a49255a  and  a49252a );
 a49257a <=( a49256a  and  a49249a );
 a49260a <=( (not A234)  and  A233 );
 a49263a <=( (not A265)  and  (not A235) );
 a49264a <=( a49263a  and  a49260a );
 a49267a <=( (not A268)  and  (not A266) );
 a49270a <=( A300  and  A298 );
 a49271a <=( a49270a  and  a49267a );
 a49272a <=( a49271a  and  a49264a );
 a49276a <=( A199  and  A167 );
 a49277a <=( A168  and  a49276a );
 a49280a <=( (not A201)  and  A200 );
 a49283a <=( (not A232)  and  (not A202) );
 a49284a <=( a49283a  and  a49280a );
 a49285a <=( a49284a  and  a49277a );
 a49288a <=( (not A235)  and  (not A233) );
 a49291a <=( (not A268)  and  (not A267) );
 a49292a <=( a49291a  and  a49288a );
 a49295a <=( A298  and  (not A269) );
 a49298a <=( A302  and  (not A299) );
 a49299a <=( a49298a  and  a49295a );
 a49300a <=( a49299a  and  a49292a );
 a49304a <=( A199  and  A167 );
 a49305a <=( A168  and  a49304a );
 a49308a <=( (not A201)  and  A200 );
 a49311a <=( (not A232)  and  (not A202) );
 a49312a <=( a49311a  and  a49308a );
 a49313a <=( a49312a  and  a49305a );
 a49316a <=( (not A235)  and  (not A233) );
 a49319a <=( (not A268)  and  (not A267) );
 a49320a <=( a49319a  and  a49316a );
 a49323a <=( (not A298)  and  (not A269) );
 a49326a <=( A302  and  A299 );
 a49327a <=( a49326a  and  a49323a );
 a49328a <=( a49327a  and  a49320a );
 a49332a <=( A199  and  A167 );
 a49333a <=( A168  and  a49332a );
 a49336a <=( (not A201)  and  A200 );
 a49339a <=( (not A232)  and  (not A202) );
 a49340a <=( a49339a  and  a49336a );
 a49341a <=( a49340a  and  a49333a );
 a49344a <=( (not A235)  and  (not A233) );
 a49347a <=( A266  and  A265 );
 a49348a <=( a49347a  and  a49344a );
 a49351a <=( (not A268)  and  (not A267) );
 a49354a <=( A300  and  A299 );
 a49355a <=( a49354a  and  a49351a );
 a49356a <=( a49355a  and  a49348a );
 a49360a <=( A199  and  A167 );
 a49361a <=( A168  and  a49360a );
 a49364a <=( (not A201)  and  A200 );
 a49367a <=( (not A232)  and  (not A202) );
 a49368a <=( a49367a  and  a49364a );
 a49369a <=( a49368a  and  a49361a );
 a49372a <=( (not A235)  and  (not A233) );
 a49375a <=( A266  and  A265 );
 a49376a <=( a49375a  and  a49372a );
 a49379a <=( (not A268)  and  (not A267) );
 a49382a <=( A300  and  A298 );
 a49383a <=( a49382a  and  a49379a );
 a49384a <=( a49383a  and  a49376a );
 a49388a <=( A199  and  A167 );
 a49389a <=( A168  and  a49388a );
 a49392a <=( (not A201)  and  A200 );
 a49395a <=( (not A232)  and  (not A202) );
 a49396a <=( a49395a  and  a49392a );
 a49397a <=( a49396a  and  a49389a );
 a49400a <=( (not A235)  and  (not A233) );
 a49403a <=( (not A266)  and  (not A265) );
 a49404a <=( a49403a  and  a49400a );
 a49407a <=( A298  and  (not A268) );
 a49410a <=( A302  and  (not A299) );
 a49411a <=( a49410a  and  a49407a );
 a49412a <=( a49411a  and  a49404a );
 a49416a <=( A199  and  A167 );
 a49417a <=( A168  and  a49416a );
 a49420a <=( (not A201)  and  A200 );
 a49423a <=( (not A232)  and  (not A202) );
 a49424a <=( a49423a  and  a49420a );
 a49425a <=( a49424a  and  a49417a );
 a49428a <=( (not A235)  and  (not A233) );
 a49431a <=( (not A266)  and  (not A265) );
 a49432a <=( a49431a  and  a49428a );
 a49435a <=( (not A298)  and  (not A268) );
 a49438a <=( A302  and  A299 );
 a49439a <=( a49438a  and  a49435a );
 a49440a <=( a49439a  and  a49432a );
 a49444a <=( (not A199)  and  A167 );
 a49445a <=( A168  and  a49444a );
 a49448a <=( (not A202)  and  (not A200) );
 a49451a <=( (not A235)  and  (not A234) );
 a49452a <=( a49451a  and  a49448a );
 a49453a <=( a49452a  and  a49445a );
 a49456a <=( A265  and  (not A236) );
 a49459a <=( (not A267)  and  A266 );
 a49460a <=( a49459a  and  a49456a );
 a49463a <=( A298  and  (not A268) );
 a49466a <=( A302  and  (not A299) );
 a49467a <=( a49466a  and  a49463a );
 a49468a <=( a49467a  and  a49460a );
 a49472a <=( (not A199)  and  A167 );
 a49473a <=( A168  and  a49472a );
 a49476a <=( (not A202)  and  (not A200) );
 a49479a <=( (not A235)  and  (not A234) );
 a49480a <=( a49479a  and  a49476a );
 a49481a <=( a49480a  and  a49473a );
 a49484a <=( A265  and  (not A236) );
 a49487a <=( (not A267)  and  A266 );
 a49488a <=( a49487a  and  a49484a );
 a49491a <=( (not A298)  and  (not A268) );
 a49494a <=( A302  and  A299 );
 a49495a <=( a49494a  and  a49491a );
 a49496a <=( a49495a  and  a49488a );
 a49500a <=( (not A199)  and  A167 );
 a49501a <=( A168  and  a49500a );
 a49504a <=( (not A202)  and  (not A200) );
 a49507a <=( A233  and  A232 );
 a49508a <=( a49507a  and  a49504a );
 a49509a <=( a49508a  and  a49501a );
 a49512a <=( (not A235)  and  (not A234) );
 a49515a <=( (not A268)  and  (not A267) );
 a49516a <=( a49515a  and  a49512a );
 a49519a <=( A298  and  (not A269) );
 a49522a <=( A302  and  (not A299) );
 a49523a <=( a49522a  and  a49519a );
 a49524a <=( a49523a  and  a49516a );
 a49528a <=( (not A199)  and  A167 );
 a49529a <=( A168  and  a49528a );
 a49532a <=( (not A202)  and  (not A200) );
 a49535a <=( A233  and  A232 );
 a49536a <=( a49535a  and  a49532a );
 a49537a <=( a49536a  and  a49529a );
 a49540a <=( (not A235)  and  (not A234) );
 a49543a <=( (not A268)  and  (not A267) );
 a49544a <=( a49543a  and  a49540a );
 a49547a <=( (not A298)  and  (not A269) );
 a49550a <=( A302  and  A299 );
 a49551a <=( a49550a  and  a49547a );
 a49552a <=( a49551a  and  a49544a );
 a49556a <=( (not A199)  and  A167 );
 a49557a <=( A168  and  a49556a );
 a49560a <=( (not A202)  and  (not A200) );
 a49563a <=( A233  and  A232 );
 a49564a <=( a49563a  and  a49560a );
 a49565a <=( a49564a  and  a49557a );
 a49568a <=( (not A235)  and  (not A234) );
 a49571a <=( A266  and  A265 );
 a49572a <=( a49571a  and  a49568a );
 a49575a <=( (not A268)  and  (not A267) );
 a49578a <=( A300  and  A299 );
 a49579a <=( a49578a  and  a49575a );
 a49580a <=( a49579a  and  a49572a );
 a49584a <=( (not A199)  and  A167 );
 a49585a <=( A168  and  a49584a );
 a49588a <=( (not A202)  and  (not A200) );
 a49591a <=( A233  and  A232 );
 a49592a <=( a49591a  and  a49588a );
 a49593a <=( a49592a  and  a49585a );
 a49596a <=( (not A235)  and  (not A234) );
 a49599a <=( A266  and  A265 );
 a49600a <=( a49599a  and  a49596a );
 a49603a <=( (not A268)  and  (not A267) );
 a49606a <=( A300  and  A298 );
 a49607a <=( a49606a  and  a49603a );
 a49608a <=( a49607a  and  a49600a );
 a49612a <=( (not A199)  and  A167 );
 a49613a <=( A168  and  a49612a );
 a49616a <=( (not A202)  and  (not A200) );
 a49619a <=( A233  and  A232 );
 a49620a <=( a49619a  and  a49616a );
 a49621a <=( a49620a  and  a49613a );
 a49624a <=( (not A235)  and  (not A234) );
 a49627a <=( (not A266)  and  (not A265) );
 a49628a <=( a49627a  and  a49624a );
 a49631a <=( A298  and  (not A268) );
 a49634a <=( A302  and  (not A299) );
 a49635a <=( a49634a  and  a49631a );
 a49636a <=( a49635a  and  a49628a );
 a49640a <=( (not A199)  and  A167 );
 a49641a <=( A168  and  a49640a );
 a49644a <=( (not A202)  and  (not A200) );
 a49647a <=( A233  and  A232 );
 a49648a <=( a49647a  and  a49644a );
 a49649a <=( a49648a  and  a49641a );
 a49652a <=( (not A235)  and  (not A234) );
 a49655a <=( (not A266)  and  (not A265) );
 a49656a <=( a49655a  and  a49652a );
 a49659a <=( (not A298)  and  (not A268) );
 a49662a <=( A302  and  A299 );
 a49663a <=( a49662a  and  a49659a );
 a49664a <=( a49663a  and  a49656a );
 a49668a <=( (not A199)  and  A167 );
 a49669a <=( A168  and  a49668a );
 a49672a <=( (not A202)  and  (not A200) );
 a49675a <=( (not A233)  and  (not A232) );
 a49676a <=( a49675a  and  a49672a );
 a49677a <=( a49676a  and  a49669a );
 a49680a <=( A265  and  (not A235) );
 a49683a <=( (not A267)  and  A266 );
 a49684a <=( a49683a  and  a49680a );
 a49687a <=( A298  and  (not A268) );
 a49690a <=( A302  and  (not A299) );
 a49691a <=( a49690a  and  a49687a );
 a49692a <=( a49691a  and  a49684a );
 a49696a <=( (not A199)  and  A167 );
 a49697a <=( A168  and  a49696a );
 a49700a <=( (not A202)  and  (not A200) );
 a49703a <=( (not A233)  and  (not A232) );
 a49704a <=( a49703a  and  a49700a );
 a49705a <=( a49704a  and  a49697a );
 a49708a <=( A265  and  (not A235) );
 a49711a <=( (not A267)  and  A266 );
 a49712a <=( a49711a  and  a49708a );
 a49715a <=( (not A298)  and  (not A268) );
 a49718a <=( A302  and  A299 );
 a49719a <=( a49718a  and  a49715a );
 a49720a <=( a49719a  and  a49712a );
 a49724a <=( (not A166)  and  A167 );
 a49725a <=( A170  and  a49724a );
 a49728a <=( (not A202)  and  (not A201) );
 a49731a <=( (not A234)  and  (not A203) );
 a49732a <=( a49731a  and  a49728a );
 a49733a <=( a49732a  and  a49725a );
 a49736a <=( (not A236)  and  (not A235) );
 a49739a <=( (not A268)  and  (not A267) );
 a49740a <=( a49739a  and  a49736a );
 a49743a <=( A298  and  (not A269) );
 a49746a <=( A302  and  (not A299) );
 a49747a <=( a49746a  and  a49743a );
 a49748a <=( a49747a  and  a49740a );
 a49752a <=( (not A166)  and  A167 );
 a49753a <=( A170  and  a49752a );
 a49756a <=( (not A202)  and  (not A201) );
 a49759a <=( (not A234)  and  (not A203) );
 a49760a <=( a49759a  and  a49756a );
 a49761a <=( a49760a  and  a49753a );
 a49764a <=( (not A236)  and  (not A235) );
 a49767a <=( (not A268)  and  (not A267) );
 a49768a <=( a49767a  and  a49764a );
 a49771a <=( (not A298)  and  (not A269) );
 a49774a <=( A302  and  A299 );
 a49775a <=( a49774a  and  a49771a );
 a49776a <=( a49775a  and  a49768a );
 a49780a <=( (not A166)  and  A167 );
 a49781a <=( A170  and  a49780a );
 a49784a <=( (not A202)  and  (not A201) );
 a49787a <=( (not A234)  and  (not A203) );
 a49788a <=( a49787a  and  a49784a );
 a49789a <=( a49788a  and  a49781a );
 a49792a <=( (not A236)  and  (not A235) );
 a49795a <=( A266  and  A265 );
 a49796a <=( a49795a  and  a49792a );
 a49799a <=( (not A268)  and  (not A267) );
 a49802a <=( A300  and  A299 );
 a49803a <=( a49802a  and  a49799a );
 a49804a <=( a49803a  and  a49796a );
 a49808a <=( (not A166)  and  A167 );
 a49809a <=( A170  and  a49808a );
 a49812a <=( (not A202)  and  (not A201) );
 a49815a <=( (not A234)  and  (not A203) );
 a49816a <=( a49815a  and  a49812a );
 a49817a <=( a49816a  and  a49809a );
 a49820a <=( (not A236)  and  (not A235) );
 a49823a <=( A266  and  A265 );
 a49824a <=( a49823a  and  a49820a );
 a49827a <=( (not A268)  and  (not A267) );
 a49830a <=( A300  and  A298 );
 a49831a <=( a49830a  and  a49827a );
 a49832a <=( a49831a  and  a49824a );
 a49836a <=( (not A166)  and  A167 );
 a49837a <=( A170  and  a49836a );
 a49840a <=( (not A202)  and  (not A201) );
 a49843a <=( (not A234)  and  (not A203) );
 a49844a <=( a49843a  and  a49840a );
 a49845a <=( a49844a  and  a49837a );
 a49848a <=( (not A236)  and  (not A235) );
 a49851a <=( (not A266)  and  (not A265) );
 a49852a <=( a49851a  and  a49848a );
 a49855a <=( A298  and  (not A268) );
 a49858a <=( A302  and  (not A299) );
 a49859a <=( a49858a  and  a49855a );
 a49860a <=( a49859a  and  a49852a );
 a49864a <=( (not A166)  and  A167 );
 a49865a <=( A170  and  a49864a );
 a49868a <=( (not A202)  and  (not A201) );
 a49871a <=( (not A234)  and  (not A203) );
 a49872a <=( a49871a  and  a49868a );
 a49873a <=( a49872a  and  a49865a );
 a49876a <=( (not A236)  and  (not A235) );
 a49879a <=( (not A266)  and  (not A265) );
 a49880a <=( a49879a  and  a49876a );
 a49883a <=( (not A298)  and  (not A268) );
 a49886a <=( A302  and  A299 );
 a49887a <=( a49886a  and  a49883a );
 a49888a <=( a49887a  and  a49880a );
 a49892a <=( (not A166)  and  A167 );
 a49893a <=( A170  and  a49892a );
 a49896a <=( (not A202)  and  (not A201) );
 a49899a <=( A232  and  (not A203) );
 a49900a <=( a49899a  and  a49896a );
 a49901a <=( a49900a  and  a49893a );
 a49904a <=( (not A234)  and  A233 );
 a49907a <=( (not A267)  and  (not A235) );
 a49908a <=( a49907a  and  a49904a );
 a49911a <=( (not A269)  and  (not A268) );
 a49914a <=( A300  and  A299 );
 a49915a <=( a49914a  and  a49911a );
 a49916a <=( a49915a  and  a49908a );
 a49920a <=( (not A166)  and  A167 );
 a49921a <=( A170  and  a49920a );
 a49924a <=( (not A202)  and  (not A201) );
 a49927a <=( A232  and  (not A203) );
 a49928a <=( a49927a  and  a49924a );
 a49929a <=( a49928a  and  a49921a );
 a49932a <=( (not A234)  and  A233 );
 a49935a <=( (not A267)  and  (not A235) );
 a49936a <=( a49935a  and  a49932a );
 a49939a <=( (not A269)  and  (not A268) );
 a49942a <=( A300  and  A298 );
 a49943a <=( a49942a  and  a49939a );
 a49944a <=( a49943a  and  a49936a );
 a49948a <=( (not A166)  and  A167 );
 a49949a <=( A170  and  a49948a );
 a49952a <=( (not A202)  and  (not A201) );
 a49955a <=( A232  and  (not A203) );
 a49956a <=( a49955a  and  a49952a );
 a49957a <=( a49956a  and  a49949a );
 a49960a <=( (not A234)  and  A233 );
 a49963a <=( A265  and  (not A235) );
 a49964a <=( a49963a  and  a49960a );
 a49967a <=( (not A267)  and  A266 );
 a49970a <=( A301  and  (not A268) );
 a49971a <=( a49970a  and  a49967a );
 a49972a <=( a49971a  and  a49964a );
 a49976a <=( (not A166)  and  A167 );
 a49977a <=( A170  and  a49976a );
 a49980a <=( (not A202)  and  (not A201) );
 a49983a <=( A232  and  (not A203) );
 a49984a <=( a49983a  and  a49980a );
 a49985a <=( a49984a  and  a49977a );
 a49988a <=( (not A234)  and  A233 );
 a49991a <=( (not A265)  and  (not A235) );
 a49992a <=( a49991a  and  a49988a );
 a49995a <=( (not A268)  and  (not A266) );
 a49998a <=( A300  and  A299 );
 a49999a <=( a49998a  and  a49995a );
 a50000a <=( a49999a  and  a49992a );
 a50004a <=( (not A166)  and  A167 );
 a50005a <=( A170  and  a50004a );
 a50008a <=( (not A202)  and  (not A201) );
 a50011a <=( A232  and  (not A203) );
 a50012a <=( a50011a  and  a50008a );
 a50013a <=( a50012a  and  a50005a );
 a50016a <=( (not A234)  and  A233 );
 a50019a <=( (not A265)  and  (not A235) );
 a50020a <=( a50019a  and  a50016a );
 a50023a <=( (not A268)  and  (not A266) );
 a50026a <=( A300  and  A298 );
 a50027a <=( a50026a  and  a50023a );
 a50028a <=( a50027a  and  a50020a );
 a50032a <=( (not A166)  and  A167 );
 a50033a <=( A170  and  a50032a );
 a50036a <=( (not A202)  and  (not A201) );
 a50039a <=( (not A232)  and  (not A203) );
 a50040a <=( a50039a  and  a50036a );
 a50041a <=( a50040a  and  a50033a );
 a50044a <=( (not A235)  and  (not A233) );
 a50047a <=( (not A268)  and  (not A267) );
 a50048a <=( a50047a  and  a50044a );
 a50051a <=( A298  and  (not A269) );
 a50054a <=( A302  and  (not A299) );
 a50055a <=( a50054a  and  a50051a );
 a50056a <=( a50055a  and  a50048a );
 a50060a <=( (not A166)  and  A167 );
 a50061a <=( A170  and  a50060a );
 a50064a <=( (not A202)  and  (not A201) );
 a50067a <=( (not A232)  and  (not A203) );
 a50068a <=( a50067a  and  a50064a );
 a50069a <=( a50068a  and  a50061a );
 a50072a <=( (not A235)  and  (not A233) );
 a50075a <=( (not A268)  and  (not A267) );
 a50076a <=( a50075a  and  a50072a );
 a50079a <=( (not A298)  and  (not A269) );
 a50082a <=( A302  and  A299 );
 a50083a <=( a50082a  and  a50079a );
 a50084a <=( a50083a  and  a50076a );
 a50088a <=( (not A166)  and  A167 );
 a50089a <=( A170  and  a50088a );
 a50092a <=( (not A202)  and  (not A201) );
 a50095a <=( (not A232)  and  (not A203) );
 a50096a <=( a50095a  and  a50092a );
 a50097a <=( a50096a  and  a50089a );
 a50100a <=( (not A235)  and  (not A233) );
 a50103a <=( A266  and  A265 );
 a50104a <=( a50103a  and  a50100a );
 a50107a <=( (not A268)  and  (not A267) );
 a50110a <=( A300  and  A299 );
 a50111a <=( a50110a  and  a50107a );
 a50112a <=( a50111a  and  a50104a );
 a50116a <=( (not A166)  and  A167 );
 a50117a <=( A170  and  a50116a );
 a50120a <=( (not A202)  and  (not A201) );
 a50123a <=( (not A232)  and  (not A203) );
 a50124a <=( a50123a  and  a50120a );
 a50125a <=( a50124a  and  a50117a );
 a50128a <=( (not A235)  and  (not A233) );
 a50131a <=( A266  and  A265 );
 a50132a <=( a50131a  and  a50128a );
 a50135a <=( (not A268)  and  (not A267) );
 a50138a <=( A300  and  A298 );
 a50139a <=( a50138a  and  a50135a );
 a50140a <=( a50139a  and  a50132a );
 a50144a <=( (not A166)  and  A167 );
 a50145a <=( A170  and  a50144a );
 a50148a <=( (not A202)  and  (not A201) );
 a50151a <=( (not A232)  and  (not A203) );
 a50152a <=( a50151a  and  a50148a );
 a50153a <=( a50152a  and  a50145a );
 a50156a <=( (not A235)  and  (not A233) );
 a50159a <=( (not A266)  and  (not A265) );
 a50160a <=( a50159a  and  a50156a );
 a50163a <=( A298  and  (not A268) );
 a50166a <=( A302  and  (not A299) );
 a50167a <=( a50166a  and  a50163a );
 a50168a <=( a50167a  and  a50160a );
 a50172a <=( (not A166)  and  A167 );
 a50173a <=( A170  and  a50172a );
 a50176a <=( (not A202)  and  (not A201) );
 a50179a <=( (not A232)  and  (not A203) );
 a50180a <=( a50179a  and  a50176a );
 a50181a <=( a50180a  and  a50173a );
 a50184a <=( (not A235)  and  (not A233) );
 a50187a <=( (not A266)  and  (not A265) );
 a50188a <=( a50187a  and  a50184a );
 a50191a <=( (not A298)  and  (not A268) );
 a50194a <=( A302  and  A299 );
 a50195a <=( a50194a  and  a50191a );
 a50196a <=( a50195a  and  a50188a );
 a50200a <=( (not A166)  and  A167 );
 a50201a <=( A170  and  a50200a );
 a50204a <=( A200  and  A199 );
 a50207a <=( (not A202)  and  (not A201) );
 a50208a <=( a50207a  and  a50204a );
 a50209a <=( a50208a  and  a50201a );
 a50212a <=( (not A235)  and  (not A234) );
 a50215a <=( (not A267)  and  (not A236) );
 a50216a <=( a50215a  and  a50212a );
 a50219a <=( (not A269)  and  (not A268) );
 a50222a <=( A300  and  A299 );
 a50223a <=( a50222a  and  a50219a );
 a50224a <=( a50223a  and  a50216a );
 a50228a <=( (not A166)  and  A167 );
 a50229a <=( A170  and  a50228a );
 a50232a <=( A200  and  A199 );
 a50235a <=( (not A202)  and  (not A201) );
 a50236a <=( a50235a  and  a50232a );
 a50237a <=( a50236a  and  a50229a );
 a50240a <=( (not A235)  and  (not A234) );
 a50243a <=( (not A267)  and  (not A236) );
 a50244a <=( a50243a  and  a50240a );
 a50247a <=( (not A269)  and  (not A268) );
 a50250a <=( A300  and  A298 );
 a50251a <=( a50250a  and  a50247a );
 a50252a <=( a50251a  and  a50244a );
 a50256a <=( (not A166)  and  A167 );
 a50257a <=( A170  and  a50256a );
 a50260a <=( A200  and  A199 );
 a50263a <=( (not A202)  and  (not A201) );
 a50264a <=( a50263a  and  a50260a );
 a50265a <=( a50264a  and  a50257a );
 a50268a <=( (not A235)  and  (not A234) );
 a50271a <=( A265  and  (not A236) );
 a50272a <=( a50271a  and  a50268a );
 a50275a <=( (not A267)  and  A266 );
 a50278a <=( A301  and  (not A268) );
 a50279a <=( a50278a  and  a50275a );
 a50280a <=( a50279a  and  a50272a );
 a50284a <=( (not A166)  and  A167 );
 a50285a <=( A170  and  a50284a );
 a50288a <=( A200  and  A199 );
 a50291a <=( (not A202)  and  (not A201) );
 a50292a <=( a50291a  and  a50288a );
 a50293a <=( a50292a  and  a50285a );
 a50296a <=( (not A235)  and  (not A234) );
 a50299a <=( (not A265)  and  (not A236) );
 a50300a <=( a50299a  and  a50296a );
 a50303a <=( (not A268)  and  (not A266) );
 a50306a <=( A300  and  A299 );
 a50307a <=( a50306a  and  a50303a );
 a50308a <=( a50307a  and  a50300a );
 a50312a <=( (not A166)  and  A167 );
 a50313a <=( A170  and  a50312a );
 a50316a <=( A200  and  A199 );
 a50319a <=( (not A202)  and  (not A201) );
 a50320a <=( a50319a  and  a50316a );
 a50321a <=( a50320a  and  a50313a );
 a50324a <=( (not A235)  and  (not A234) );
 a50327a <=( (not A265)  and  (not A236) );
 a50328a <=( a50327a  and  a50324a );
 a50331a <=( (not A268)  and  (not A266) );
 a50334a <=( A300  and  A298 );
 a50335a <=( a50334a  and  a50331a );
 a50336a <=( a50335a  and  a50328a );
 a50340a <=( (not A166)  and  A167 );
 a50341a <=( A170  and  a50340a );
 a50344a <=( A200  and  A199 );
 a50347a <=( (not A202)  and  (not A201) );
 a50348a <=( a50347a  and  a50344a );
 a50349a <=( a50348a  and  a50341a );
 a50352a <=( A233  and  A232 );
 a50355a <=( (not A235)  and  (not A234) );
 a50356a <=( a50355a  and  a50352a );
 a50359a <=( (not A268)  and  (not A267) );
 a50362a <=( A301  and  (not A269) );
 a50363a <=( a50362a  and  a50359a );
 a50364a <=( a50363a  and  a50356a );
 a50368a <=( (not A166)  and  A167 );
 a50369a <=( A170  and  a50368a );
 a50372a <=( A200  and  A199 );
 a50375a <=( (not A202)  and  (not A201) );
 a50376a <=( a50375a  and  a50372a );
 a50377a <=( a50376a  and  a50369a );
 a50380a <=( A233  and  A232 );
 a50383a <=( (not A235)  and  (not A234) );
 a50384a <=( a50383a  and  a50380a );
 a50387a <=( (not A266)  and  (not A265) );
 a50390a <=( A301  and  (not A268) );
 a50391a <=( a50390a  and  a50387a );
 a50392a <=( a50391a  and  a50384a );
 a50396a <=( (not A166)  and  A167 );
 a50397a <=( A170  and  a50396a );
 a50400a <=( A200  and  A199 );
 a50403a <=( (not A202)  and  (not A201) );
 a50404a <=( a50403a  and  a50400a );
 a50405a <=( a50404a  and  a50397a );
 a50408a <=( (not A233)  and  (not A232) );
 a50411a <=( (not A267)  and  (not A235) );
 a50412a <=( a50411a  and  a50408a );
 a50415a <=( (not A269)  and  (not A268) );
 a50418a <=( A300  and  A299 );
 a50419a <=( a50418a  and  a50415a );
 a50420a <=( a50419a  and  a50412a );
 a50424a <=( (not A166)  and  A167 );
 a50425a <=( A170  and  a50424a );
 a50428a <=( A200  and  A199 );
 a50431a <=( (not A202)  and  (not A201) );
 a50432a <=( a50431a  and  a50428a );
 a50433a <=( a50432a  and  a50425a );
 a50436a <=( (not A233)  and  (not A232) );
 a50439a <=( (not A267)  and  (not A235) );
 a50440a <=( a50439a  and  a50436a );
 a50443a <=( (not A269)  and  (not A268) );
 a50446a <=( A300  and  A298 );
 a50447a <=( a50446a  and  a50443a );
 a50448a <=( a50447a  and  a50440a );
 a50452a <=( (not A166)  and  A167 );
 a50453a <=( A170  and  a50452a );
 a50456a <=( A200  and  A199 );
 a50459a <=( (not A202)  and  (not A201) );
 a50460a <=( a50459a  and  a50456a );
 a50461a <=( a50460a  and  a50453a );
 a50464a <=( (not A233)  and  (not A232) );
 a50467a <=( A265  and  (not A235) );
 a50468a <=( a50467a  and  a50464a );
 a50471a <=( (not A267)  and  A266 );
 a50474a <=( A301  and  (not A268) );
 a50475a <=( a50474a  and  a50471a );
 a50476a <=( a50475a  and  a50468a );
 a50480a <=( (not A166)  and  A167 );
 a50481a <=( A170  and  a50480a );
 a50484a <=( A200  and  A199 );
 a50487a <=( (not A202)  and  (not A201) );
 a50488a <=( a50487a  and  a50484a );
 a50489a <=( a50488a  and  a50481a );
 a50492a <=( (not A233)  and  (not A232) );
 a50495a <=( (not A265)  and  (not A235) );
 a50496a <=( a50495a  and  a50492a );
 a50499a <=( (not A268)  and  (not A266) );
 a50502a <=( A300  and  A299 );
 a50503a <=( a50502a  and  a50499a );
 a50504a <=( a50503a  and  a50496a );
 a50508a <=( (not A166)  and  A167 );
 a50509a <=( A170  and  a50508a );
 a50512a <=( A200  and  A199 );
 a50515a <=( (not A202)  and  (not A201) );
 a50516a <=( a50515a  and  a50512a );
 a50517a <=( a50516a  and  a50509a );
 a50520a <=( (not A233)  and  (not A232) );
 a50523a <=( (not A265)  and  (not A235) );
 a50524a <=( a50523a  and  a50520a );
 a50527a <=( (not A268)  and  (not A266) );
 a50530a <=( A300  and  A298 );
 a50531a <=( a50530a  and  a50527a );
 a50532a <=( a50531a  and  a50524a );
 a50536a <=( (not A166)  and  A167 );
 a50537a <=( A170  and  a50536a );
 a50540a <=( (not A200)  and  (not A199) );
 a50543a <=( (not A234)  and  (not A202) );
 a50544a <=( a50543a  and  a50540a );
 a50545a <=( a50544a  and  a50537a );
 a50548a <=( (not A236)  and  (not A235) );
 a50551a <=( (not A268)  and  (not A267) );
 a50552a <=( a50551a  and  a50548a );
 a50555a <=( A298  and  (not A269) );
 a50558a <=( A302  and  (not A299) );
 a50559a <=( a50558a  and  a50555a );
 a50560a <=( a50559a  and  a50552a );
 a50564a <=( (not A166)  and  A167 );
 a50565a <=( A170  and  a50564a );
 a50568a <=( (not A200)  and  (not A199) );
 a50571a <=( (not A234)  and  (not A202) );
 a50572a <=( a50571a  and  a50568a );
 a50573a <=( a50572a  and  a50565a );
 a50576a <=( (not A236)  and  (not A235) );
 a50579a <=( (not A268)  and  (not A267) );
 a50580a <=( a50579a  and  a50576a );
 a50583a <=( (not A298)  and  (not A269) );
 a50586a <=( A302  and  A299 );
 a50587a <=( a50586a  and  a50583a );
 a50588a <=( a50587a  and  a50580a );
 a50592a <=( (not A166)  and  A167 );
 a50593a <=( A170  and  a50592a );
 a50596a <=( (not A200)  and  (not A199) );
 a50599a <=( (not A234)  and  (not A202) );
 a50600a <=( a50599a  and  a50596a );
 a50601a <=( a50600a  and  a50593a );
 a50604a <=( (not A236)  and  (not A235) );
 a50607a <=( A266  and  A265 );
 a50608a <=( a50607a  and  a50604a );
 a50611a <=( (not A268)  and  (not A267) );
 a50614a <=( A300  and  A299 );
 a50615a <=( a50614a  and  a50611a );
 a50616a <=( a50615a  and  a50608a );
 a50620a <=( (not A166)  and  A167 );
 a50621a <=( A170  and  a50620a );
 a50624a <=( (not A200)  and  (not A199) );
 a50627a <=( (not A234)  and  (not A202) );
 a50628a <=( a50627a  and  a50624a );
 a50629a <=( a50628a  and  a50621a );
 a50632a <=( (not A236)  and  (not A235) );
 a50635a <=( A266  and  A265 );
 a50636a <=( a50635a  and  a50632a );
 a50639a <=( (not A268)  and  (not A267) );
 a50642a <=( A300  and  A298 );
 a50643a <=( a50642a  and  a50639a );
 a50644a <=( a50643a  and  a50636a );
 a50648a <=( (not A166)  and  A167 );
 a50649a <=( A170  and  a50648a );
 a50652a <=( (not A200)  and  (not A199) );
 a50655a <=( (not A234)  and  (not A202) );
 a50656a <=( a50655a  and  a50652a );
 a50657a <=( a50656a  and  a50649a );
 a50660a <=( (not A236)  and  (not A235) );
 a50663a <=( (not A266)  and  (not A265) );
 a50664a <=( a50663a  and  a50660a );
 a50667a <=( A298  and  (not A268) );
 a50670a <=( A302  and  (not A299) );
 a50671a <=( a50670a  and  a50667a );
 a50672a <=( a50671a  and  a50664a );
 a50676a <=( (not A166)  and  A167 );
 a50677a <=( A170  and  a50676a );
 a50680a <=( (not A200)  and  (not A199) );
 a50683a <=( (not A234)  and  (not A202) );
 a50684a <=( a50683a  and  a50680a );
 a50685a <=( a50684a  and  a50677a );
 a50688a <=( (not A236)  and  (not A235) );
 a50691a <=( (not A266)  and  (not A265) );
 a50692a <=( a50691a  and  a50688a );
 a50695a <=( (not A298)  and  (not A268) );
 a50698a <=( A302  and  A299 );
 a50699a <=( a50698a  and  a50695a );
 a50700a <=( a50699a  and  a50692a );
 a50704a <=( (not A166)  and  A167 );
 a50705a <=( A170  and  a50704a );
 a50708a <=( (not A200)  and  (not A199) );
 a50711a <=( A232  and  (not A202) );
 a50712a <=( a50711a  and  a50708a );
 a50713a <=( a50712a  and  a50705a );
 a50716a <=( (not A234)  and  A233 );
 a50719a <=( (not A267)  and  (not A235) );
 a50720a <=( a50719a  and  a50716a );
 a50723a <=( (not A269)  and  (not A268) );
 a50726a <=( A300  and  A299 );
 a50727a <=( a50726a  and  a50723a );
 a50728a <=( a50727a  and  a50720a );
 a50732a <=( (not A166)  and  A167 );
 a50733a <=( A170  and  a50732a );
 a50736a <=( (not A200)  and  (not A199) );
 a50739a <=( A232  and  (not A202) );
 a50740a <=( a50739a  and  a50736a );
 a50741a <=( a50740a  and  a50733a );
 a50744a <=( (not A234)  and  A233 );
 a50747a <=( (not A267)  and  (not A235) );
 a50748a <=( a50747a  and  a50744a );
 a50751a <=( (not A269)  and  (not A268) );
 a50754a <=( A300  and  A298 );
 a50755a <=( a50754a  and  a50751a );
 a50756a <=( a50755a  and  a50748a );
 a50760a <=( (not A166)  and  A167 );
 a50761a <=( A170  and  a50760a );
 a50764a <=( (not A200)  and  (not A199) );
 a50767a <=( A232  and  (not A202) );
 a50768a <=( a50767a  and  a50764a );
 a50769a <=( a50768a  and  a50761a );
 a50772a <=( (not A234)  and  A233 );
 a50775a <=( A265  and  (not A235) );
 a50776a <=( a50775a  and  a50772a );
 a50779a <=( (not A267)  and  A266 );
 a50782a <=( A301  and  (not A268) );
 a50783a <=( a50782a  and  a50779a );
 a50784a <=( a50783a  and  a50776a );
 a50788a <=( (not A166)  and  A167 );
 a50789a <=( A170  and  a50788a );
 a50792a <=( (not A200)  and  (not A199) );
 a50795a <=( A232  and  (not A202) );
 a50796a <=( a50795a  and  a50792a );
 a50797a <=( a50796a  and  a50789a );
 a50800a <=( (not A234)  and  A233 );
 a50803a <=( (not A265)  and  (not A235) );
 a50804a <=( a50803a  and  a50800a );
 a50807a <=( (not A268)  and  (not A266) );
 a50810a <=( A300  and  A299 );
 a50811a <=( a50810a  and  a50807a );
 a50812a <=( a50811a  and  a50804a );
 a50816a <=( (not A166)  and  A167 );
 a50817a <=( A170  and  a50816a );
 a50820a <=( (not A200)  and  (not A199) );
 a50823a <=( A232  and  (not A202) );
 a50824a <=( a50823a  and  a50820a );
 a50825a <=( a50824a  and  a50817a );
 a50828a <=( (not A234)  and  A233 );
 a50831a <=( (not A265)  and  (not A235) );
 a50832a <=( a50831a  and  a50828a );
 a50835a <=( (not A268)  and  (not A266) );
 a50838a <=( A300  and  A298 );
 a50839a <=( a50838a  and  a50835a );
 a50840a <=( a50839a  and  a50832a );
 a50844a <=( (not A166)  and  A167 );
 a50845a <=( A170  and  a50844a );
 a50848a <=( (not A200)  and  (not A199) );
 a50851a <=( (not A232)  and  (not A202) );
 a50852a <=( a50851a  and  a50848a );
 a50853a <=( a50852a  and  a50845a );
 a50856a <=( (not A235)  and  (not A233) );
 a50859a <=( (not A268)  and  (not A267) );
 a50860a <=( a50859a  and  a50856a );
 a50863a <=( A298  and  (not A269) );
 a50866a <=( A302  and  (not A299) );
 a50867a <=( a50866a  and  a50863a );
 a50868a <=( a50867a  and  a50860a );
 a50872a <=( (not A166)  and  A167 );
 a50873a <=( A170  and  a50872a );
 a50876a <=( (not A200)  and  (not A199) );
 a50879a <=( (not A232)  and  (not A202) );
 a50880a <=( a50879a  and  a50876a );
 a50881a <=( a50880a  and  a50873a );
 a50884a <=( (not A235)  and  (not A233) );
 a50887a <=( (not A268)  and  (not A267) );
 a50888a <=( a50887a  and  a50884a );
 a50891a <=( (not A298)  and  (not A269) );
 a50894a <=( A302  and  A299 );
 a50895a <=( a50894a  and  a50891a );
 a50896a <=( a50895a  and  a50888a );
 a50900a <=( (not A166)  and  A167 );
 a50901a <=( A170  and  a50900a );
 a50904a <=( (not A200)  and  (not A199) );
 a50907a <=( (not A232)  and  (not A202) );
 a50908a <=( a50907a  and  a50904a );
 a50909a <=( a50908a  and  a50901a );
 a50912a <=( (not A235)  and  (not A233) );
 a50915a <=( A266  and  A265 );
 a50916a <=( a50915a  and  a50912a );
 a50919a <=( (not A268)  and  (not A267) );
 a50922a <=( A300  and  A299 );
 a50923a <=( a50922a  and  a50919a );
 a50924a <=( a50923a  and  a50916a );
 a50928a <=( (not A166)  and  A167 );
 a50929a <=( A170  and  a50928a );
 a50932a <=( (not A200)  and  (not A199) );
 a50935a <=( (not A232)  and  (not A202) );
 a50936a <=( a50935a  and  a50932a );
 a50937a <=( a50936a  and  a50929a );
 a50940a <=( (not A235)  and  (not A233) );
 a50943a <=( A266  and  A265 );
 a50944a <=( a50943a  and  a50940a );
 a50947a <=( (not A268)  and  (not A267) );
 a50950a <=( A300  and  A298 );
 a50951a <=( a50950a  and  a50947a );
 a50952a <=( a50951a  and  a50944a );
 a50956a <=( (not A166)  and  A167 );
 a50957a <=( A170  and  a50956a );
 a50960a <=( (not A200)  and  (not A199) );
 a50963a <=( (not A232)  and  (not A202) );
 a50964a <=( a50963a  and  a50960a );
 a50965a <=( a50964a  and  a50957a );
 a50968a <=( (not A235)  and  (not A233) );
 a50971a <=( (not A266)  and  (not A265) );
 a50972a <=( a50971a  and  a50968a );
 a50975a <=( A298  and  (not A268) );
 a50978a <=( A302  and  (not A299) );
 a50979a <=( a50978a  and  a50975a );
 a50980a <=( a50979a  and  a50972a );
 a50984a <=( (not A166)  and  A167 );
 a50985a <=( A170  and  a50984a );
 a50988a <=( (not A200)  and  (not A199) );
 a50991a <=( (not A232)  and  (not A202) );
 a50992a <=( a50991a  and  a50988a );
 a50993a <=( a50992a  and  a50985a );
 a50996a <=( (not A235)  and  (not A233) );
 a50999a <=( (not A266)  and  (not A265) );
 a51000a <=( a50999a  and  a50996a );
 a51003a <=( (not A298)  and  (not A268) );
 a51006a <=( A302  and  A299 );
 a51007a <=( a51006a  and  a51003a );
 a51008a <=( a51007a  and  a51000a );
 a51012a <=( A166  and  (not A167) );
 a51013a <=( A170  and  a51012a );
 a51016a <=( (not A202)  and  (not A201) );
 a51019a <=( (not A234)  and  (not A203) );
 a51020a <=( a51019a  and  a51016a );
 a51021a <=( a51020a  and  a51013a );
 a51024a <=( (not A236)  and  (not A235) );
 a51027a <=( (not A268)  and  (not A267) );
 a51028a <=( a51027a  and  a51024a );
 a51031a <=( A298  and  (not A269) );
 a51034a <=( A302  and  (not A299) );
 a51035a <=( a51034a  and  a51031a );
 a51036a <=( a51035a  and  a51028a );
 a51040a <=( A166  and  (not A167) );
 a51041a <=( A170  and  a51040a );
 a51044a <=( (not A202)  and  (not A201) );
 a51047a <=( (not A234)  and  (not A203) );
 a51048a <=( a51047a  and  a51044a );
 a51049a <=( a51048a  and  a51041a );
 a51052a <=( (not A236)  and  (not A235) );
 a51055a <=( (not A268)  and  (not A267) );
 a51056a <=( a51055a  and  a51052a );
 a51059a <=( (not A298)  and  (not A269) );
 a51062a <=( A302  and  A299 );
 a51063a <=( a51062a  and  a51059a );
 a51064a <=( a51063a  and  a51056a );
 a51068a <=( A166  and  (not A167) );
 a51069a <=( A170  and  a51068a );
 a51072a <=( (not A202)  and  (not A201) );
 a51075a <=( (not A234)  and  (not A203) );
 a51076a <=( a51075a  and  a51072a );
 a51077a <=( a51076a  and  a51069a );
 a51080a <=( (not A236)  and  (not A235) );
 a51083a <=( A266  and  A265 );
 a51084a <=( a51083a  and  a51080a );
 a51087a <=( (not A268)  and  (not A267) );
 a51090a <=( A300  and  A299 );
 a51091a <=( a51090a  and  a51087a );
 a51092a <=( a51091a  and  a51084a );
 a51096a <=( A166  and  (not A167) );
 a51097a <=( A170  and  a51096a );
 a51100a <=( (not A202)  and  (not A201) );
 a51103a <=( (not A234)  and  (not A203) );
 a51104a <=( a51103a  and  a51100a );
 a51105a <=( a51104a  and  a51097a );
 a51108a <=( (not A236)  and  (not A235) );
 a51111a <=( A266  and  A265 );
 a51112a <=( a51111a  and  a51108a );
 a51115a <=( (not A268)  and  (not A267) );
 a51118a <=( A300  and  A298 );
 a51119a <=( a51118a  and  a51115a );
 a51120a <=( a51119a  and  a51112a );
 a51124a <=( A166  and  (not A167) );
 a51125a <=( A170  and  a51124a );
 a51128a <=( (not A202)  and  (not A201) );
 a51131a <=( (not A234)  and  (not A203) );
 a51132a <=( a51131a  and  a51128a );
 a51133a <=( a51132a  and  a51125a );
 a51136a <=( (not A236)  and  (not A235) );
 a51139a <=( (not A266)  and  (not A265) );
 a51140a <=( a51139a  and  a51136a );
 a51143a <=( A298  and  (not A268) );
 a51146a <=( A302  and  (not A299) );
 a51147a <=( a51146a  and  a51143a );
 a51148a <=( a51147a  and  a51140a );
 a51152a <=( A166  and  (not A167) );
 a51153a <=( A170  and  a51152a );
 a51156a <=( (not A202)  and  (not A201) );
 a51159a <=( (not A234)  and  (not A203) );
 a51160a <=( a51159a  and  a51156a );
 a51161a <=( a51160a  and  a51153a );
 a51164a <=( (not A236)  and  (not A235) );
 a51167a <=( (not A266)  and  (not A265) );
 a51168a <=( a51167a  and  a51164a );
 a51171a <=( (not A298)  and  (not A268) );
 a51174a <=( A302  and  A299 );
 a51175a <=( a51174a  and  a51171a );
 a51176a <=( a51175a  and  a51168a );
 a51180a <=( A166  and  (not A167) );
 a51181a <=( A170  and  a51180a );
 a51184a <=( (not A202)  and  (not A201) );
 a51187a <=( A232  and  (not A203) );
 a51188a <=( a51187a  and  a51184a );
 a51189a <=( a51188a  and  a51181a );
 a51192a <=( (not A234)  and  A233 );
 a51195a <=( (not A267)  and  (not A235) );
 a51196a <=( a51195a  and  a51192a );
 a51199a <=( (not A269)  and  (not A268) );
 a51202a <=( A300  and  A299 );
 a51203a <=( a51202a  and  a51199a );
 a51204a <=( a51203a  and  a51196a );
 a51208a <=( A166  and  (not A167) );
 a51209a <=( A170  and  a51208a );
 a51212a <=( (not A202)  and  (not A201) );
 a51215a <=( A232  and  (not A203) );
 a51216a <=( a51215a  and  a51212a );
 a51217a <=( a51216a  and  a51209a );
 a51220a <=( (not A234)  and  A233 );
 a51223a <=( (not A267)  and  (not A235) );
 a51224a <=( a51223a  and  a51220a );
 a51227a <=( (not A269)  and  (not A268) );
 a51230a <=( A300  and  A298 );
 a51231a <=( a51230a  and  a51227a );
 a51232a <=( a51231a  and  a51224a );
 a51236a <=( A166  and  (not A167) );
 a51237a <=( A170  and  a51236a );
 a51240a <=( (not A202)  and  (not A201) );
 a51243a <=( A232  and  (not A203) );
 a51244a <=( a51243a  and  a51240a );
 a51245a <=( a51244a  and  a51237a );
 a51248a <=( (not A234)  and  A233 );
 a51251a <=( A265  and  (not A235) );
 a51252a <=( a51251a  and  a51248a );
 a51255a <=( (not A267)  and  A266 );
 a51258a <=( A301  and  (not A268) );
 a51259a <=( a51258a  and  a51255a );
 a51260a <=( a51259a  and  a51252a );
 a51264a <=( A166  and  (not A167) );
 a51265a <=( A170  and  a51264a );
 a51268a <=( (not A202)  and  (not A201) );
 a51271a <=( A232  and  (not A203) );
 a51272a <=( a51271a  and  a51268a );
 a51273a <=( a51272a  and  a51265a );
 a51276a <=( (not A234)  and  A233 );
 a51279a <=( (not A265)  and  (not A235) );
 a51280a <=( a51279a  and  a51276a );
 a51283a <=( (not A268)  and  (not A266) );
 a51286a <=( A300  and  A299 );
 a51287a <=( a51286a  and  a51283a );
 a51288a <=( a51287a  and  a51280a );
 a51292a <=( A166  and  (not A167) );
 a51293a <=( A170  and  a51292a );
 a51296a <=( (not A202)  and  (not A201) );
 a51299a <=( A232  and  (not A203) );
 a51300a <=( a51299a  and  a51296a );
 a51301a <=( a51300a  and  a51293a );
 a51304a <=( (not A234)  and  A233 );
 a51307a <=( (not A265)  and  (not A235) );
 a51308a <=( a51307a  and  a51304a );
 a51311a <=( (not A268)  and  (not A266) );
 a51314a <=( A300  and  A298 );
 a51315a <=( a51314a  and  a51311a );
 a51316a <=( a51315a  and  a51308a );
 a51320a <=( A166  and  (not A167) );
 a51321a <=( A170  and  a51320a );
 a51324a <=( (not A202)  and  (not A201) );
 a51327a <=( (not A232)  and  (not A203) );
 a51328a <=( a51327a  and  a51324a );
 a51329a <=( a51328a  and  a51321a );
 a51332a <=( (not A235)  and  (not A233) );
 a51335a <=( (not A268)  and  (not A267) );
 a51336a <=( a51335a  and  a51332a );
 a51339a <=( A298  and  (not A269) );
 a51342a <=( A302  and  (not A299) );
 a51343a <=( a51342a  and  a51339a );
 a51344a <=( a51343a  and  a51336a );
 a51348a <=( A166  and  (not A167) );
 a51349a <=( A170  and  a51348a );
 a51352a <=( (not A202)  and  (not A201) );
 a51355a <=( (not A232)  and  (not A203) );
 a51356a <=( a51355a  and  a51352a );
 a51357a <=( a51356a  and  a51349a );
 a51360a <=( (not A235)  and  (not A233) );
 a51363a <=( (not A268)  and  (not A267) );
 a51364a <=( a51363a  and  a51360a );
 a51367a <=( (not A298)  and  (not A269) );
 a51370a <=( A302  and  A299 );
 a51371a <=( a51370a  and  a51367a );
 a51372a <=( a51371a  and  a51364a );
 a51376a <=( A166  and  (not A167) );
 a51377a <=( A170  and  a51376a );
 a51380a <=( (not A202)  and  (not A201) );
 a51383a <=( (not A232)  and  (not A203) );
 a51384a <=( a51383a  and  a51380a );
 a51385a <=( a51384a  and  a51377a );
 a51388a <=( (not A235)  and  (not A233) );
 a51391a <=( A266  and  A265 );
 a51392a <=( a51391a  and  a51388a );
 a51395a <=( (not A268)  and  (not A267) );
 a51398a <=( A300  and  A299 );
 a51399a <=( a51398a  and  a51395a );
 a51400a <=( a51399a  and  a51392a );
 a51404a <=( A166  and  (not A167) );
 a51405a <=( A170  and  a51404a );
 a51408a <=( (not A202)  and  (not A201) );
 a51411a <=( (not A232)  and  (not A203) );
 a51412a <=( a51411a  and  a51408a );
 a51413a <=( a51412a  and  a51405a );
 a51416a <=( (not A235)  and  (not A233) );
 a51419a <=( A266  and  A265 );
 a51420a <=( a51419a  and  a51416a );
 a51423a <=( (not A268)  and  (not A267) );
 a51426a <=( A300  and  A298 );
 a51427a <=( a51426a  and  a51423a );
 a51428a <=( a51427a  and  a51420a );
 a51432a <=( A166  and  (not A167) );
 a51433a <=( A170  and  a51432a );
 a51436a <=( (not A202)  and  (not A201) );
 a51439a <=( (not A232)  and  (not A203) );
 a51440a <=( a51439a  and  a51436a );
 a51441a <=( a51440a  and  a51433a );
 a51444a <=( (not A235)  and  (not A233) );
 a51447a <=( (not A266)  and  (not A265) );
 a51448a <=( a51447a  and  a51444a );
 a51451a <=( A298  and  (not A268) );
 a51454a <=( A302  and  (not A299) );
 a51455a <=( a51454a  and  a51451a );
 a51456a <=( a51455a  and  a51448a );
 a51460a <=( A166  and  (not A167) );
 a51461a <=( A170  and  a51460a );
 a51464a <=( (not A202)  and  (not A201) );
 a51467a <=( (not A232)  and  (not A203) );
 a51468a <=( a51467a  and  a51464a );
 a51469a <=( a51468a  and  a51461a );
 a51472a <=( (not A235)  and  (not A233) );
 a51475a <=( (not A266)  and  (not A265) );
 a51476a <=( a51475a  and  a51472a );
 a51479a <=( (not A298)  and  (not A268) );
 a51482a <=( A302  and  A299 );
 a51483a <=( a51482a  and  a51479a );
 a51484a <=( a51483a  and  a51476a );
 a51488a <=( A166  and  (not A167) );
 a51489a <=( A170  and  a51488a );
 a51492a <=( A200  and  A199 );
 a51495a <=( (not A202)  and  (not A201) );
 a51496a <=( a51495a  and  a51492a );
 a51497a <=( a51496a  and  a51489a );
 a51500a <=( (not A235)  and  (not A234) );
 a51503a <=( (not A267)  and  (not A236) );
 a51504a <=( a51503a  and  a51500a );
 a51507a <=( (not A269)  and  (not A268) );
 a51510a <=( A300  and  A299 );
 a51511a <=( a51510a  and  a51507a );
 a51512a <=( a51511a  and  a51504a );
 a51516a <=( A166  and  (not A167) );
 a51517a <=( A170  and  a51516a );
 a51520a <=( A200  and  A199 );
 a51523a <=( (not A202)  and  (not A201) );
 a51524a <=( a51523a  and  a51520a );
 a51525a <=( a51524a  and  a51517a );
 a51528a <=( (not A235)  and  (not A234) );
 a51531a <=( (not A267)  and  (not A236) );
 a51532a <=( a51531a  and  a51528a );
 a51535a <=( (not A269)  and  (not A268) );
 a51538a <=( A300  and  A298 );
 a51539a <=( a51538a  and  a51535a );
 a51540a <=( a51539a  and  a51532a );
 a51544a <=( A166  and  (not A167) );
 a51545a <=( A170  and  a51544a );
 a51548a <=( A200  and  A199 );
 a51551a <=( (not A202)  and  (not A201) );
 a51552a <=( a51551a  and  a51548a );
 a51553a <=( a51552a  and  a51545a );
 a51556a <=( (not A235)  and  (not A234) );
 a51559a <=( A265  and  (not A236) );
 a51560a <=( a51559a  and  a51556a );
 a51563a <=( (not A267)  and  A266 );
 a51566a <=( A301  and  (not A268) );
 a51567a <=( a51566a  and  a51563a );
 a51568a <=( a51567a  and  a51560a );
 a51572a <=( A166  and  (not A167) );
 a51573a <=( A170  and  a51572a );
 a51576a <=( A200  and  A199 );
 a51579a <=( (not A202)  and  (not A201) );
 a51580a <=( a51579a  and  a51576a );
 a51581a <=( a51580a  and  a51573a );
 a51584a <=( (not A235)  and  (not A234) );
 a51587a <=( (not A265)  and  (not A236) );
 a51588a <=( a51587a  and  a51584a );
 a51591a <=( (not A268)  and  (not A266) );
 a51594a <=( A300  and  A299 );
 a51595a <=( a51594a  and  a51591a );
 a51596a <=( a51595a  and  a51588a );
 a51600a <=( A166  and  (not A167) );
 a51601a <=( A170  and  a51600a );
 a51604a <=( A200  and  A199 );
 a51607a <=( (not A202)  and  (not A201) );
 a51608a <=( a51607a  and  a51604a );
 a51609a <=( a51608a  and  a51601a );
 a51612a <=( (not A235)  and  (not A234) );
 a51615a <=( (not A265)  and  (not A236) );
 a51616a <=( a51615a  and  a51612a );
 a51619a <=( (not A268)  and  (not A266) );
 a51622a <=( A300  and  A298 );
 a51623a <=( a51622a  and  a51619a );
 a51624a <=( a51623a  and  a51616a );
 a51628a <=( A166  and  (not A167) );
 a51629a <=( A170  and  a51628a );
 a51632a <=( A200  and  A199 );
 a51635a <=( (not A202)  and  (not A201) );
 a51636a <=( a51635a  and  a51632a );
 a51637a <=( a51636a  and  a51629a );
 a51640a <=( A233  and  A232 );
 a51643a <=( (not A235)  and  (not A234) );
 a51644a <=( a51643a  and  a51640a );
 a51647a <=( (not A268)  and  (not A267) );
 a51650a <=( A301  and  (not A269) );
 a51651a <=( a51650a  and  a51647a );
 a51652a <=( a51651a  and  a51644a );
 a51656a <=( A166  and  (not A167) );
 a51657a <=( A170  and  a51656a );
 a51660a <=( A200  and  A199 );
 a51663a <=( (not A202)  and  (not A201) );
 a51664a <=( a51663a  and  a51660a );
 a51665a <=( a51664a  and  a51657a );
 a51668a <=( A233  and  A232 );
 a51671a <=( (not A235)  and  (not A234) );
 a51672a <=( a51671a  and  a51668a );
 a51675a <=( (not A266)  and  (not A265) );
 a51678a <=( A301  and  (not A268) );
 a51679a <=( a51678a  and  a51675a );
 a51680a <=( a51679a  and  a51672a );
 a51684a <=( A166  and  (not A167) );
 a51685a <=( A170  and  a51684a );
 a51688a <=( A200  and  A199 );
 a51691a <=( (not A202)  and  (not A201) );
 a51692a <=( a51691a  and  a51688a );
 a51693a <=( a51692a  and  a51685a );
 a51696a <=( (not A233)  and  (not A232) );
 a51699a <=( (not A267)  and  (not A235) );
 a51700a <=( a51699a  and  a51696a );
 a51703a <=( (not A269)  and  (not A268) );
 a51706a <=( A300  and  A299 );
 a51707a <=( a51706a  and  a51703a );
 a51708a <=( a51707a  and  a51700a );
 a51712a <=( A166  and  (not A167) );
 a51713a <=( A170  and  a51712a );
 a51716a <=( A200  and  A199 );
 a51719a <=( (not A202)  and  (not A201) );
 a51720a <=( a51719a  and  a51716a );
 a51721a <=( a51720a  and  a51713a );
 a51724a <=( (not A233)  and  (not A232) );
 a51727a <=( (not A267)  and  (not A235) );
 a51728a <=( a51727a  and  a51724a );
 a51731a <=( (not A269)  and  (not A268) );
 a51734a <=( A300  and  A298 );
 a51735a <=( a51734a  and  a51731a );
 a51736a <=( a51735a  and  a51728a );
 a51740a <=( A166  and  (not A167) );
 a51741a <=( A170  and  a51740a );
 a51744a <=( A200  and  A199 );
 a51747a <=( (not A202)  and  (not A201) );
 a51748a <=( a51747a  and  a51744a );
 a51749a <=( a51748a  and  a51741a );
 a51752a <=( (not A233)  and  (not A232) );
 a51755a <=( A265  and  (not A235) );
 a51756a <=( a51755a  and  a51752a );
 a51759a <=( (not A267)  and  A266 );
 a51762a <=( A301  and  (not A268) );
 a51763a <=( a51762a  and  a51759a );
 a51764a <=( a51763a  and  a51756a );
 a51768a <=( A166  and  (not A167) );
 a51769a <=( A170  and  a51768a );
 a51772a <=( A200  and  A199 );
 a51775a <=( (not A202)  and  (not A201) );
 a51776a <=( a51775a  and  a51772a );
 a51777a <=( a51776a  and  a51769a );
 a51780a <=( (not A233)  and  (not A232) );
 a51783a <=( (not A265)  and  (not A235) );
 a51784a <=( a51783a  and  a51780a );
 a51787a <=( (not A268)  and  (not A266) );
 a51790a <=( A300  and  A299 );
 a51791a <=( a51790a  and  a51787a );
 a51792a <=( a51791a  and  a51784a );
 a51796a <=( A166  and  (not A167) );
 a51797a <=( A170  and  a51796a );
 a51800a <=( A200  and  A199 );
 a51803a <=( (not A202)  and  (not A201) );
 a51804a <=( a51803a  and  a51800a );
 a51805a <=( a51804a  and  a51797a );
 a51808a <=( (not A233)  and  (not A232) );
 a51811a <=( (not A265)  and  (not A235) );
 a51812a <=( a51811a  and  a51808a );
 a51815a <=( (not A268)  and  (not A266) );
 a51818a <=( A300  and  A298 );
 a51819a <=( a51818a  and  a51815a );
 a51820a <=( a51819a  and  a51812a );
 a51824a <=( A166  and  (not A167) );
 a51825a <=( A170  and  a51824a );
 a51828a <=( (not A200)  and  (not A199) );
 a51831a <=( (not A234)  and  (not A202) );
 a51832a <=( a51831a  and  a51828a );
 a51833a <=( a51832a  and  a51825a );
 a51836a <=( (not A236)  and  (not A235) );
 a51839a <=( (not A268)  and  (not A267) );
 a51840a <=( a51839a  and  a51836a );
 a51843a <=( A298  and  (not A269) );
 a51846a <=( A302  and  (not A299) );
 a51847a <=( a51846a  and  a51843a );
 a51848a <=( a51847a  and  a51840a );
 a51852a <=( A166  and  (not A167) );
 a51853a <=( A170  and  a51852a );
 a51856a <=( (not A200)  and  (not A199) );
 a51859a <=( (not A234)  and  (not A202) );
 a51860a <=( a51859a  and  a51856a );
 a51861a <=( a51860a  and  a51853a );
 a51864a <=( (not A236)  and  (not A235) );
 a51867a <=( (not A268)  and  (not A267) );
 a51868a <=( a51867a  and  a51864a );
 a51871a <=( (not A298)  and  (not A269) );
 a51874a <=( A302  and  A299 );
 a51875a <=( a51874a  and  a51871a );
 a51876a <=( a51875a  and  a51868a );
 a51880a <=( A166  and  (not A167) );
 a51881a <=( A170  and  a51880a );
 a51884a <=( (not A200)  and  (not A199) );
 a51887a <=( (not A234)  and  (not A202) );
 a51888a <=( a51887a  and  a51884a );
 a51889a <=( a51888a  and  a51881a );
 a51892a <=( (not A236)  and  (not A235) );
 a51895a <=( A266  and  A265 );
 a51896a <=( a51895a  and  a51892a );
 a51899a <=( (not A268)  and  (not A267) );
 a51902a <=( A300  and  A299 );
 a51903a <=( a51902a  and  a51899a );
 a51904a <=( a51903a  and  a51896a );
 a51908a <=( A166  and  (not A167) );
 a51909a <=( A170  and  a51908a );
 a51912a <=( (not A200)  and  (not A199) );
 a51915a <=( (not A234)  and  (not A202) );
 a51916a <=( a51915a  and  a51912a );
 a51917a <=( a51916a  and  a51909a );
 a51920a <=( (not A236)  and  (not A235) );
 a51923a <=( A266  and  A265 );
 a51924a <=( a51923a  and  a51920a );
 a51927a <=( (not A268)  and  (not A267) );
 a51930a <=( A300  and  A298 );
 a51931a <=( a51930a  and  a51927a );
 a51932a <=( a51931a  and  a51924a );
 a51936a <=( A166  and  (not A167) );
 a51937a <=( A170  and  a51936a );
 a51940a <=( (not A200)  and  (not A199) );
 a51943a <=( (not A234)  and  (not A202) );
 a51944a <=( a51943a  and  a51940a );
 a51945a <=( a51944a  and  a51937a );
 a51948a <=( (not A236)  and  (not A235) );
 a51951a <=( (not A266)  and  (not A265) );
 a51952a <=( a51951a  and  a51948a );
 a51955a <=( A298  and  (not A268) );
 a51958a <=( A302  and  (not A299) );
 a51959a <=( a51958a  and  a51955a );
 a51960a <=( a51959a  and  a51952a );
 a51964a <=( A166  and  (not A167) );
 a51965a <=( A170  and  a51964a );
 a51968a <=( (not A200)  and  (not A199) );
 a51971a <=( (not A234)  and  (not A202) );
 a51972a <=( a51971a  and  a51968a );
 a51973a <=( a51972a  and  a51965a );
 a51976a <=( (not A236)  and  (not A235) );
 a51979a <=( (not A266)  and  (not A265) );
 a51980a <=( a51979a  and  a51976a );
 a51983a <=( (not A298)  and  (not A268) );
 a51986a <=( A302  and  A299 );
 a51987a <=( a51986a  and  a51983a );
 a51988a <=( a51987a  and  a51980a );
 a51992a <=( A166  and  (not A167) );
 a51993a <=( A170  and  a51992a );
 a51996a <=( (not A200)  and  (not A199) );
 a51999a <=( A232  and  (not A202) );
 a52000a <=( a51999a  and  a51996a );
 a52001a <=( a52000a  and  a51993a );
 a52004a <=( (not A234)  and  A233 );
 a52007a <=( (not A267)  and  (not A235) );
 a52008a <=( a52007a  and  a52004a );
 a52011a <=( (not A269)  and  (not A268) );
 a52014a <=( A300  and  A299 );
 a52015a <=( a52014a  and  a52011a );
 a52016a <=( a52015a  and  a52008a );
 a52020a <=( A166  and  (not A167) );
 a52021a <=( A170  and  a52020a );
 a52024a <=( (not A200)  and  (not A199) );
 a52027a <=( A232  and  (not A202) );
 a52028a <=( a52027a  and  a52024a );
 a52029a <=( a52028a  and  a52021a );
 a52032a <=( (not A234)  and  A233 );
 a52035a <=( (not A267)  and  (not A235) );
 a52036a <=( a52035a  and  a52032a );
 a52039a <=( (not A269)  and  (not A268) );
 a52042a <=( A300  and  A298 );
 a52043a <=( a52042a  and  a52039a );
 a52044a <=( a52043a  and  a52036a );
 a52048a <=( A166  and  (not A167) );
 a52049a <=( A170  and  a52048a );
 a52052a <=( (not A200)  and  (not A199) );
 a52055a <=( A232  and  (not A202) );
 a52056a <=( a52055a  and  a52052a );
 a52057a <=( a52056a  and  a52049a );
 a52060a <=( (not A234)  and  A233 );
 a52063a <=( A265  and  (not A235) );
 a52064a <=( a52063a  and  a52060a );
 a52067a <=( (not A267)  and  A266 );
 a52070a <=( A301  and  (not A268) );
 a52071a <=( a52070a  and  a52067a );
 a52072a <=( a52071a  and  a52064a );
 a52076a <=( A166  and  (not A167) );
 a52077a <=( A170  and  a52076a );
 a52080a <=( (not A200)  and  (not A199) );
 a52083a <=( A232  and  (not A202) );
 a52084a <=( a52083a  and  a52080a );
 a52085a <=( a52084a  and  a52077a );
 a52088a <=( (not A234)  and  A233 );
 a52091a <=( (not A265)  and  (not A235) );
 a52092a <=( a52091a  and  a52088a );
 a52095a <=( (not A268)  and  (not A266) );
 a52098a <=( A300  and  A299 );
 a52099a <=( a52098a  and  a52095a );
 a52100a <=( a52099a  and  a52092a );
 a52104a <=( A166  and  (not A167) );
 a52105a <=( A170  and  a52104a );
 a52108a <=( (not A200)  and  (not A199) );
 a52111a <=( A232  and  (not A202) );
 a52112a <=( a52111a  and  a52108a );
 a52113a <=( a52112a  and  a52105a );
 a52116a <=( (not A234)  and  A233 );
 a52119a <=( (not A265)  and  (not A235) );
 a52120a <=( a52119a  and  a52116a );
 a52123a <=( (not A268)  and  (not A266) );
 a52126a <=( A300  and  A298 );
 a52127a <=( a52126a  and  a52123a );
 a52128a <=( a52127a  and  a52120a );
 a52132a <=( A166  and  (not A167) );
 a52133a <=( A170  and  a52132a );
 a52136a <=( (not A200)  and  (not A199) );
 a52139a <=( (not A232)  and  (not A202) );
 a52140a <=( a52139a  and  a52136a );
 a52141a <=( a52140a  and  a52133a );
 a52144a <=( (not A235)  and  (not A233) );
 a52147a <=( (not A268)  and  (not A267) );
 a52148a <=( a52147a  and  a52144a );
 a52151a <=( A298  and  (not A269) );
 a52154a <=( A302  and  (not A299) );
 a52155a <=( a52154a  and  a52151a );
 a52156a <=( a52155a  and  a52148a );
 a52160a <=( A166  and  (not A167) );
 a52161a <=( A170  and  a52160a );
 a52164a <=( (not A200)  and  (not A199) );
 a52167a <=( (not A232)  and  (not A202) );
 a52168a <=( a52167a  and  a52164a );
 a52169a <=( a52168a  and  a52161a );
 a52172a <=( (not A235)  and  (not A233) );
 a52175a <=( (not A268)  and  (not A267) );
 a52176a <=( a52175a  and  a52172a );
 a52179a <=( (not A298)  and  (not A269) );
 a52182a <=( A302  and  A299 );
 a52183a <=( a52182a  and  a52179a );
 a52184a <=( a52183a  and  a52176a );
 a52188a <=( A166  and  (not A167) );
 a52189a <=( A170  and  a52188a );
 a52192a <=( (not A200)  and  (not A199) );
 a52195a <=( (not A232)  and  (not A202) );
 a52196a <=( a52195a  and  a52192a );
 a52197a <=( a52196a  and  a52189a );
 a52200a <=( (not A235)  and  (not A233) );
 a52203a <=( A266  and  A265 );
 a52204a <=( a52203a  and  a52200a );
 a52207a <=( (not A268)  and  (not A267) );
 a52210a <=( A300  and  A299 );
 a52211a <=( a52210a  and  a52207a );
 a52212a <=( a52211a  and  a52204a );
 a52216a <=( A166  and  (not A167) );
 a52217a <=( A170  and  a52216a );
 a52220a <=( (not A200)  and  (not A199) );
 a52223a <=( (not A232)  and  (not A202) );
 a52224a <=( a52223a  and  a52220a );
 a52225a <=( a52224a  and  a52217a );
 a52228a <=( (not A235)  and  (not A233) );
 a52231a <=( A266  and  A265 );
 a52232a <=( a52231a  and  a52228a );
 a52235a <=( (not A268)  and  (not A267) );
 a52238a <=( A300  and  A298 );
 a52239a <=( a52238a  and  a52235a );
 a52240a <=( a52239a  and  a52232a );
 a52244a <=( A166  and  (not A167) );
 a52245a <=( A170  and  a52244a );
 a52248a <=( (not A200)  and  (not A199) );
 a52251a <=( (not A232)  and  (not A202) );
 a52252a <=( a52251a  and  a52248a );
 a52253a <=( a52252a  and  a52245a );
 a52256a <=( (not A235)  and  (not A233) );
 a52259a <=( (not A266)  and  (not A265) );
 a52260a <=( a52259a  and  a52256a );
 a52263a <=( A298  and  (not A268) );
 a52266a <=( A302  and  (not A299) );
 a52267a <=( a52266a  and  a52263a );
 a52268a <=( a52267a  and  a52260a );
 a52272a <=( A166  and  (not A167) );
 a52273a <=( A170  and  a52272a );
 a52276a <=( (not A200)  and  (not A199) );
 a52279a <=( (not A232)  and  (not A202) );
 a52280a <=( a52279a  and  a52276a );
 a52281a <=( a52280a  and  a52273a );
 a52284a <=( (not A235)  and  (not A233) );
 a52287a <=( (not A266)  and  (not A265) );
 a52288a <=( a52287a  and  a52284a );
 a52291a <=( (not A298)  and  (not A268) );
 a52294a <=( A302  and  A299 );
 a52295a <=( a52294a  and  a52291a );
 a52296a <=( a52295a  and  a52288a );
 a52300a <=( (not A202)  and  (not A201) );
 a52301a <=( A169  and  a52300a );
 a52304a <=( A232  and  (not A203) );
 a52307a <=( (not A234)  and  A233 );
 a52308a <=( a52307a  and  a52304a );
 a52309a <=( a52308a  and  a52301a );
 a52312a <=( A265  and  (not A235) );
 a52315a <=( (not A267)  and  A266 );
 a52316a <=( a52315a  and  a52312a );
 a52319a <=( A298  and  (not A268) );
 a52322a <=( A302  and  (not A299) );
 a52323a <=( a52322a  and  a52319a );
 a52324a <=( a52323a  and  a52316a );
 a52328a <=( (not A202)  and  (not A201) );
 a52329a <=( A169  and  a52328a );
 a52332a <=( A232  and  (not A203) );
 a52335a <=( (not A234)  and  A233 );
 a52336a <=( a52335a  and  a52332a );
 a52337a <=( a52336a  and  a52329a );
 a52340a <=( A265  and  (not A235) );
 a52343a <=( (not A267)  and  A266 );
 a52344a <=( a52343a  and  a52340a );
 a52347a <=( (not A298)  and  (not A268) );
 a52350a <=( A302  and  A299 );
 a52351a <=( a52350a  and  a52347a );
 a52352a <=( a52351a  and  a52344a );
 a52356a <=( A200  and  A199 );
 a52357a <=( A169  and  a52356a );
 a52360a <=( (not A202)  and  (not A201) );
 a52363a <=( (not A235)  and  (not A234) );
 a52364a <=( a52363a  and  a52360a );
 a52365a <=( a52364a  and  a52357a );
 a52368a <=( A265  and  (not A236) );
 a52371a <=( (not A267)  and  A266 );
 a52372a <=( a52371a  and  a52368a );
 a52375a <=( A298  and  (not A268) );
 a52378a <=( A302  and  (not A299) );
 a52379a <=( a52378a  and  a52375a );
 a52380a <=( a52379a  and  a52372a );
 a52384a <=( A200  and  A199 );
 a52385a <=( A169  and  a52384a );
 a52388a <=( (not A202)  and  (not A201) );
 a52391a <=( (not A235)  and  (not A234) );
 a52392a <=( a52391a  and  a52388a );
 a52393a <=( a52392a  and  a52385a );
 a52396a <=( A265  and  (not A236) );
 a52399a <=( (not A267)  and  A266 );
 a52400a <=( a52399a  and  a52396a );
 a52403a <=( (not A298)  and  (not A268) );
 a52406a <=( A302  and  A299 );
 a52407a <=( a52406a  and  a52403a );
 a52408a <=( a52407a  and  a52400a );
 a52412a <=( A200  and  A199 );
 a52413a <=( A169  and  a52412a );
 a52416a <=( (not A202)  and  (not A201) );
 a52419a <=( A233  and  A232 );
 a52420a <=( a52419a  and  a52416a );
 a52421a <=( a52420a  and  a52413a );
 a52424a <=( (not A235)  and  (not A234) );
 a52427a <=( (not A268)  and  (not A267) );
 a52428a <=( a52427a  and  a52424a );
 a52431a <=( A298  and  (not A269) );
 a52434a <=( A302  and  (not A299) );
 a52435a <=( a52434a  and  a52431a );
 a52436a <=( a52435a  and  a52428a );
 a52440a <=( A200  and  A199 );
 a52441a <=( A169  and  a52440a );
 a52444a <=( (not A202)  and  (not A201) );
 a52447a <=( A233  and  A232 );
 a52448a <=( a52447a  and  a52444a );
 a52449a <=( a52448a  and  a52441a );
 a52452a <=( (not A235)  and  (not A234) );
 a52455a <=( (not A268)  and  (not A267) );
 a52456a <=( a52455a  and  a52452a );
 a52459a <=( (not A298)  and  (not A269) );
 a52462a <=( A302  and  A299 );
 a52463a <=( a52462a  and  a52459a );
 a52464a <=( a52463a  and  a52456a );
 a52468a <=( A200  and  A199 );
 a52469a <=( A169  and  a52468a );
 a52472a <=( (not A202)  and  (not A201) );
 a52475a <=( A233  and  A232 );
 a52476a <=( a52475a  and  a52472a );
 a52477a <=( a52476a  and  a52469a );
 a52480a <=( (not A235)  and  (not A234) );
 a52483a <=( A266  and  A265 );
 a52484a <=( a52483a  and  a52480a );
 a52487a <=( (not A268)  and  (not A267) );
 a52490a <=( A300  and  A299 );
 a52491a <=( a52490a  and  a52487a );
 a52492a <=( a52491a  and  a52484a );
 a52496a <=( A200  and  A199 );
 a52497a <=( A169  and  a52496a );
 a52500a <=( (not A202)  and  (not A201) );
 a52503a <=( A233  and  A232 );
 a52504a <=( a52503a  and  a52500a );
 a52505a <=( a52504a  and  a52497a );
 a52508a <=( (not A235)  and  (not A234) );
 a52511a <=( A266  and  A265 );
 a52512a <=( a52511a  and  a52508a );
 a52515a <=( (not A268)  and  (not A267) );
 a52518a <=( A300  and  A298 );
 a52519a <=( a52518a  and  a52515a );
 a52520a <=( a52519a  and  a52512a );
 a52524a <=( A200  and  A199 );
 a52525a <=( A169  and  a52524a );
 a52528a <=( (not A202)  and  (not A201) );
 a52531a <=( A233  and  A232 );
 a52532a <=( a52531a  and  a52528a );
 a52533a <=( a52532a  and  a52525a );
 a52536a <=( (not A235)  and  (not A234) );
 a52539a <=( (not A266)  and  (not A265) );
 a52540a <=( a52539a  and  a52536a );
 a52543a <=( A298  and  (not A268) );
 a52546a <=( A302  and  (not A299) );
 a52547a <=( a52546a  and  a52543a );
 a52548a <=( a52547a  and  a52540a );
 a52552a <=( A200  and  A199 );
 a52553a <=( A169  and  a52552a );
 a52556a <=( (not A202)  and  (not A201) );
 a52559a <=( A233  and  A232 );
 a52560a <=( a52559a  and  a52556a );
 a52561a <=( a52560a  and  a52553a );
 a52564a <=( (not A235)  and  (not A234) );
 a52567a <=( (not A266)  and  (not A265) );
 a52568a <=( a52567a  and  a52564a );
 a52571a <=( (not A298)  and  (not A268) );
 a52574a <=( A302  and  A299 );
 a52575a <=( a52574a  and  a52571a );
 a52576a <=( a52575a  and  a52568a );
 a52580a <=( A200  and  A199 );
 a52581a <=( A169  and  a52580a );
 a52584a <=( (not A202)  and  (not A201) );
 a52587a <=( (not A233)  and  (not A232) );
 a52588a <=( a52587a  and  a52584a );
 a52589a <=( a52588a  and  a52581a );
 a52592a <=( A265  and  (not A235) );
 a52595a <=( (not A267)  and  A266 );
 a52596a <=( a52595a  and  a52592a );
 a52599a <=( A298  and  (not A268) );
 a52602a <=( A302  and  (not A299) );
 a52603a <=( a52602a  and  a52599a );
 a52604a <=( a52603a  and  a52596a );
 a52608a <=( A200  and  A199 );
 a52609a <=( A169  and  a52608a );
 a52612a <=( (not A202)  and  (not A201) );
 a52615a <=( (not A233)  and  (not A232) );
 a52616a <=( a52615a  and  a52612a );
 a52617a <=( a52616a  and  a52609a );
 a52620a <=( A265  and  (not A235) );
 a52623a <=( (not A267)  and  A266 );
 a52624a <=( a52623a  and  a52620a );
 a52627a <=( (not A298)  and  (not A268) );
 a52630a <=( A302  and  A299 );
 a52631a <=( a52630a  and  a52627a );
 a52632a <=( a52631a  and  a52624a );
 a52636a <=( (not A200)  and  (not A199) );
 a52637a <=( A169  and  a52636a );
 a52640a <=( A232  and  (not A202) );
 a52643a <=( (not A234)  and  A233 );
 a52644a <=( a52643a  and  a52640a );
 a52645a <=( a52644a  and  a52637a );
 a52648a <=( A265  and  (not A235) );
 a52651a <=( (not A267)  and  A266 );
 a52652a <=( a52651a  and  a52648a );
 a52655a <=( A298  and  (not A268) );
 a52658a <=( A302  and  (not A299) );
 a52659a <=( a52658a  and  a52655a );
 a52660a <=( a52659a  and  a52652a );
 a52664a <=( (not A200)  and  (not A199) );
 a52665a <=( A169  and  a52664a );
 a52668a <=( A232  and  (not A202) );
 a52671a <=( (not A234)  and  A233 );
 a52672a <=( a52671a  and  a52668a );
 a52673a <=( a52672a  and  a52665a );
 a52676a <=( A265  and  (not A235) );
 a52679a <=( (not A267)  and  A266 );
 a52680a <=( a52679a  and  a52676a );
 a52683a <=( (not A298)  and  (not A268) );
 a52686a <=( A302  and  A299 );
 a52687a <=( a52686a  and  a52683a );
 a52688a <=( a52687a  and  a52680a );
 a52692a <=( (not A166)  and  (not A167) );
 a52693a <=( (not A169)  and  a52692a );
 a52696a <=( A232  and  A202 );
 a52699a <=( (not A234)  and  A233 );
 a52700a <=( a52699a  and  a52696a );
 a52701a <=( a52700a  and  a52693a );
 a52704a <=( A265  and  (not A235) );
 a52707a <=( (not A267)  and  A266 );
 a52708a <=( a52707a  and  a52704a );
 a52711a <=( A298  and  (not A268) );
 a52714a <=( A302  and  (not A299) );
 a52715a <=( a52714a  and  a52711a );
 a52716a <=( a52715a  and  a52708a );
 a52720a <=( (not A166)  and  (not A167) );
 a52721a <=( (not A169)  and  a52720a );
 a52724a <=( A232  and  A202 );
 a52727a <=( (not A234)  and  A233 );
 a52728a <=( a52727a  and  a52724a );
 a52729a <=( a52728a  and  a52721a );
 a52732a <=( A265  and  (not A235) );
 a52735a <=( (not A267)  and  A266 );
 a52736a <=( a52735a  and  a52732a );
 a52739a <=( (not A298)  and  (not A268) );
 a52742a <=( A302  and  A299 );
 a52743a <=( a52742a  and  a52739a );
 a52744a <=( a52743a  and  a52736a );
 a52748a <=( (not A166)  and  (not A167) );
 a52749a <=( (not A169)  and  a52748a );
 a52752a <=( A201  and  A199 );
 a52755a <=( (not A235)  and  (not A234) );
 a52756a <=( a52755a  and  a52752a );
 a52757a <=( a52756a  and  a52749a );
 a52760a <=( A265  and  (not A236) );
 a52763a <=( (not A267)  and  A266 );
 a52764a <=( a52763a  and  a52760a );
 a52767a <=( A298  and  (not A268) );
 a52770a <=( A302  and  (not A299) );
 a52771a <=( a52770a  and  a52767a );
 a52772a <=( a52771a  and  a52764a );
 a52776a <=( (not A166)  and  (not A167) );
 a52777a <=( (not A169)  and  a52776a );
 a52780a <=( A201  and  A199 );
 a52783a <=( (not A235)  and  (not A234) );
 a52784a <=( a52783a  and  a52780a );
 a52785a <=( a52784a  and  a52777a );
 a52788a <=( A265  and  (not A236) );
 a52791a <=( (not A267)  and  A266 );
 a52792a <=( a52791a  and  a52788a );
 a52795a <=( (not A298)  and  (not A268) );
 a52798a <=( A302  and  A299 );
 a52799a <=( a52798a  and  a52795a );
 a52800a <=( a52799a  and  a52792a );
 a52804a <=( (not A166)  and  (not A167) );
 a52805a <=( (not A169)  and  a52804a );
 a52808a <=( A201  and  A199 );
 a52811a <=( A233  and  A232 );
 a52812a <=( a52811a  and  a52808a );
 a52813a <=( a52812a  and  a52805a );
 a52816a <=( (not A235)  and  (not A234) );
 a52819a <=( (not A268)  and  (not A267) );
 a52820a <=( a52819a  and  a52816a );
 a52823a <=( A298  and  (not A269) );
 a52826a <=( A302  and  (not A299) );
 a52827a <=( a52826a  and  a52823a );
 a52828a <=( a52827a  and  a52820a );
 a52832a <=( (not A166)  and  (not A167) );
 a52833a <=( (not A169)  and  a52832a );
 a52836a <=( A201  and  A199 );
 a52839a <=( A233  and  A232 );
 a52840a <=( a52839a  and  a52836a );
 a52841a <=( a52840a  and  a52833a );
 a52844a <=( (not A235)  and  (not A234) );
 a52847a <=( (not A268)  and  (not A267) );
 a52848a <=( a52847a  and  a52844a );
 a52851a <=( (not A298)  and  (not A269) );
 a52854a <=( A302  and  A299 );
 a52855a <=( a52854a  and  a52851a );
 a52856a <=( a52855a  and  a52848a );
 a52860a <=( (not A166)  and  (not A167) );
 a52861a <=( (not A169)  and  a52860a );
 a52864a <=( A201  and  A199 );
 a52867a <=( A233  and  A232 );
 a52868a <=( a52867a  and  a52864a );
 a52869a <=( a52868a  and  a52861a );
 a52872a <=( (not A235)  and  (not A234) );
 a52875a <=( A266  and  A265 );
 a52876a <=( a52875a  and  a52872a );
 a52879a <=( (not A268)  and  (not A267) );
 a52882a <=( A300  and  A299 );
 a52883a <=( a52882a  and  a52879a );
 a52884a <=( a52883a  and  a52876a );
 a52888a <=( (not A166)  and  (not A167) );
 a52889a <=( (not A169)  and  a52888a );
 a52892a <=( A201  and  A199 );
 a52895a <=( A233  and  A232 );
 a52896a <=( a52895a  and  a52892a );
 a52897a <=( a52896a  and  a52889a );
 a52900a <=( (not A235)  and  (not A234) );
 a52903a <=( A266  and  A265 );
 a52904a <=( a52903a  and  a52900a );
 a52907a <=( (not A268)  and  (not A267) );
 a52910a <=( A300  and  A298 );
 a52911a <=( a52910a  and  a52907a );
 a52912a <=( a52911a  and  a52904a );
 a52916a <=( (not A166)  and  (not A167) );
 a52917a <=( (not A169)  and  a52916a );
 a52920a <=( A201  and  A199 );
 a52923a <=( A233  and  A232 );
 a52924a <=( a52923a  and  a52920a );
 a52925a <=( a52924a  and  a52917a );
 a52928a <=( (not A235)  and  (not A234) );
 a52931a <=( (not A266)  and  (not A265) );
 a52932a <=( a52931a  and  a52928a );
 a52935a <=( A298  and  (not A268) );
 a52938a <=( A302  and  (not A299) );
 a52939a <=( a52938a  and  a52935a );
 a52940a <=( a52939a  and  a52932a );
 a52944a <=( (not A166)  and  (not A167) );
 a52945a <=( (not A169)  and  a52944a );
 a52948a <=( A201  and  A199 );
 a52951a <=( A233  and  A232 );
 a52952a <=( a52951a  and  a52948a );
 a52953a <=( a52952a  and  a52945a );
 a52956a <=( (not A235)  and  (not A234) );
 a52959a <=( (not A266)  and  (not A265) );
 a52960a <=( a52959a  and  a52956a );
 a52963a <=( (not A298)  and  (not A268) );
 a52966a <=( A302  and  A299 );
 a52967a <=( a52966a  and  a52963a );
 a52968a <=( a52967a  and  a52960a );
 a52972a <=( (not A166)  and  (not A167) );
 a52973a <=( (not A169)  and  a52972a );
 a52976a <=( A201  and  A199 );
 a52979a <=( (not A233)  and  (not A232) );
 a52980a <=( a52979a  and  a52976a );
 a52981a <=( a52980a  and  a52973a );
 a52984a <=( A265  and  (not A235) );
 a52987a <=( (not A267)  and  A266 );
 a52988a <=( a52987a  and  a52984a );
 a52991a <=( A298  and  (not A268) );
 a52994a <=( A302  and  (not A299) );
 a52995a <=( a52994a  and  a52991a );
 a52996a <=( a52995a  and  a52988a );
 a53000a <=( (not A166)  and  (not A167) );
 a53001a <=( (not A169)  and  a53000a );
 a53004a <=( A201  and  A199 );
 a53007a <=( (not A233)  and  (not A232) );
 a53008a <=( a53007a  and  a53004a );
 a53009a <=( a53008a  and  a53001a );
 a53012a <=( A265  and  (not A235) );
 a53015a <=( (not A267)  and  A266 );
 a53016a <=( a53015a  and  a53012a );
 a53019a <=( (not A298)  and  (not A268) );
 a53022a <=( A302  and  A299 );
 a53023a <=( a53022a  and  a53019a );
 a53024a <=( a53023a  and  a53016a );
 a53028a <=( (not A166)  and  (not A167) );
 a53029a <=( (not A169)  and  a53028a );
 a53032a <=( A201  and  A200 );
 a53035a <=( (not A235)  and  (not A234) );
 a53036a <=( a53035a  and  a53032a );
 a53037a <=( a53036a  and  a53029a );
 a53040a <=( A265  and  (not A236) );
 a53043a <=( (not A267)  and  A266 );
 a53044a <=( a53043a  and  a53040a );
 a53047a <=( A298  and  (not A268) );
 a53050a <=( A302  and  (not A299) );
 a53051a <=( a53050a  and  a53047a );
 a53052a <=( a53051a  and  a53044a );
 a53056a <=( (not A166)  and  (not A167) );
 a53057a <=( (not A169)  and  a53056a );
 a53060a <=( A201  and  A200 );
 a53063a <=( (not A235)  and  (not A234) );
 a53064a <=( a53063a  and  a53060a );
 a53065a <=( a53064a  and  a53057a );
 a53068a <=( A265  and  (not A236) );
 a53071a <=( (not A267)  and  A266 );
 a53072a <=( a53071a  and  a53068a );
 a53075a <=( (not A298)  and  (not A268) );
 a53078a <=( A302  and  A299 );
 a53079a <=( a53078a  and  a53075a );
 a53080a <=( a53079a  and  a53072a );
 a53084a <=( (not A166)  and  (not A167) );
 a53085a <=( (not A169)  and  a53084a );
 a53088a <=( A201  and  A200 );
 a53091a <=( A233  and  A232 );
 a53092a <=( a53091a  and  a53088a );
 a53093a <=( a53092a  and  a53085a );
 a53096a <=( (not A235)  and  (not A234) );
 a53099a <=( (not A268)  and  (not A267) );
 a53100a <=( a53099a  and  a53096a );
 a53103a <=( A298  and  (not A269) );
 a53106a <=( A302  and  (not A299) );
 a53107a <=( a53106a  and  a53103a );
 a53108a <=( a53107a  and  a53100a );
 a53112a <=( (not A166)  and  (not A167) );
 a53113a <=( (not A169)  and  a53112a );
 a53116a <=( A201  and  A200 );
 a53119a <=( A233  and  A232 );
 a53120a <=( a53119a  and  a53116a );
 a53121a <=( a53120a  and  a53113a );
 a53124a <=( (not A235)  and  (not A234) );
 a53127a <=( (not A268)  and  (not A267) );
 a53128a <=( a53127a  and  a53124a );
 a53131a <=( (not A298)  and  (not A269) );
 a53134a <=( A302  and  A299 );
 a53135a <=( a53134a  and  a53131a );
 a53136a <=( a53135a  and  a53128a );
 a53140a <=( (not A166)  and  (not A167) );
 a53141a <=( (not A169)  and  a53140a );
 a53144a <=( A201  and  A200 );
 a53147a <=( A233  and  A232 );
 a53148a <=( a53147a  and  a53144a );
 a53149a <=( a53148a  and  a53141a );
 a53152a <=( (not A235)  and  (not A234) );
 a53155a <=( A266  and  A265 );
 a53156a <=( a53155a  and  a53152a );
 a53159a <=( (not A268)  and  (not A267) );
 a53162a <=( A300  and  A299 );
 a53163a <=( a53162a  and  a53159a );
 a53164a <=( a53163a  and  a53156a );
 a53168a <=( (not A166)  and  (not A167) );
 a53169a <=( (not A169)  and  a53168a );
 a53172a <=( A201  and  A200 );
 a53175a <=( A233  and  A232 );
 a53176a <=( a53175a  and  a53172a );
 a53177a <=( a53176a  and  a53169a );
 a53180a <=( (not A235)  and  (not A234) );
 a53183a <=( A266  and  A265 );
 a53184a <=( a53183a  and  a53180a );
 a53187a <=( (not A268)  and  (not A267) );
 a53190a <=( A300  and  A298 );
 a53191a <=( a53190a  and  a53187a );
 a53192a <=( a53191a  and  a53184a );
 a53196a <=( (not A166)  and  (not A167) );
 a53197a <=( (not A169)  and  a53196a );
 a53200a <=( A201  and  A200 );
 a53203a <=( A233  and  A232 );
 a53204a <=( a53203a  and  a53200a );
 a53205a <=( a53204a  and  a53197a );
 a53208a <=( (not A235)  and  (not A234) );
 a53211a <=( (not A266)  and  (not A265) );
 a53212a <=( a53211a  and  a53208a );
 a53215a <=( A298  and  (not A268) );
 a53218a <=( A302  and  (not A299) );
 a53219a <=( a53218a  and  a53215a );
 a53220a <=( a53219a  and  a53212a );
 a53224a <=( (not A166)  and  (not A167) );
 a53225a <=( (not A169)  and  a53224a );
 a53228a <=( A201  and  A200 );
 a53231a <=( A233  and  A232 );
 a53232a <=( a53231a  and  a53228a );
 a53233a <=( a53232a  and  a53225a );
 a53236a <=( (not A235)  and  (not A234) );
 a53239a <=( (not A266)  and  (not A265) );
 a53240a <=( a53239a  and  a53236a );
 a53243a <=( (not A298)  and  (not A268) );
 a53246a <=( A302  and  A299 );
 a53247a <=( a53246a  and  a53243a );
 a53248a <=( a53247a  and  a53240a );
 a53252a <=( (not A166)  and  (not A167) );
 a53253a <=( (not A169)  and  a53252a );
 a53256a <=( A201  and  A200 );
 a53259a <=( (not A233)  and  (not A232) );
 a53260a <=( a53259a  and  a53256a );
 a53261a <=( a53260a  and  a53253a );
 a53264a <=( A265  and  (not A235) );
 a53267a <=( (not A267)  and  A266 );
 a53268a <=( a53267a  and  a53264a );
 a53271a <=( A298  and  (not A268) );
 a53274a <=( A302  and  (not A299) );
 a53275a <=( a53274a  and  a53271a );
 a53276a <=( a53275a  and  a53268a );
 a53280a <=( (not A166)  and  (not A167) );
 a53281a <=( (not A169)  and  a53280a );
 a53284a <=( A201  and  A200 );
 a53287a <=( (not A233)  and  (not A232) );
 a53288a <=( a53287a  and  a53284a );
 a53289a <=( a53288a  and  a53281a );
 a53292a <=( A265  and  (not A235) );
 a53295a <=( (not A267)  and  A266 );
 a53296a <=( a53295a  and  a53292a );
 a53299a <=( (not A298)  and  (not A268) );
 a53302a <=( A302  and  A299 );
 a53303a <=( a53302a  and  a53299a );
 a53304a <=( a53303a  and  a53296a );
 a53308a <=( (not A166)  and  (not A167) );
 a53309a <=( (not A169)  and  a53308a );
 a53312a <=( A200  and  (not A199) );
 a53315a <=( (not A234)  and  A203 );
 a53316a <=( a53315a  and  a53312a );
 a53317a <=( a53316a  and  a53309a );
 a53320a <=( (not A236)  and  (not A235) );
 a53323a <=( (not A268)  and  (not A267) );
 a53324a <=( a53323a  and  a53320a );
 a53327a <=( A298  and  (not A269) );
 a53330a <=( A302  and  (not A299) );
 a53331a <=( a53330a  and  a53327a );
 a53332a <=( a53331a  and  a53324a );
 a53336a <=( (not A166)  and  (not A167) );
 a53337a <=( (not A169)  and  a53336a );
 a53340a <=( A200  and  (not A199) );
 a53343a <=( (not A234)  and  A203 );
 a53344a <=( a53343a  and  a53340a );
 a53345a <=( a53344a  and  a53337a );
 a53348a <=( (not A236)  and  (not A235) );
 a53351a <=( (not A268)  and  (not A267) );
 a53352a <=( a53351a  and  a53348a );
 a53355a <=( (not A298)  and  (not A269) );
 a53358a <=( A302  and  A299 );
 a53359a <=( a53358a  and  a53355a );
 a53360a <=( a53359a  and  a53352a );
 a53364a <=( (not A166)  and  (not A167) );
 a53365a <=( (not A169)  and  a53364a );
 a53368a <=( A200  and  (not A199) );
 a53371a <=( (not A234)  and  A203 );
 a53372a <=( a53371a  and  a53368a );
 a53373a <=( a53372a  and  a53365a );
 a53376a <=( (not A236)  and  (not A235) );
 a53379a <=( A266  and  A265 );
 a53380a <=( a53379a  and  a53376a );
 a53383a <=( (not A268)  and  (not A267) );
 a53386a <=( A300  and  A299 );
 a53387a <=( a53386a  and  a53383a );
 a53388a <=( a53387a  and  a53380a );
 a53392a <=( (not A166)  and  (not A167) );
 a53393a <=( (not A169)  and  a53392a );
 a53396a <=( A200  and  (not A199) );
 a53399a <=( (not A234)  and  A203 );
 a53400a <=( a53399a  and  a53396a );
 a53401a <=( a53400a  and  a53393a );
 a53404a <=( (not A236)  and  (not A235) );
 a53407a <=( A266  and  A265 );
 a53408a <=( a53407a  and  a53404a );
 a53411a <=( (not A268)  and  (not A267) );
 a53414a <=( A300  and  A298 );
 a53415a <=( a53414a  and  a53411a );
 a53416a <=( a53415a  and  a53408a );
 a53420a <=( (not A166)  and  (not A167) );
 a53421a <=( (not A169)  and  a53420a );
 a53424a <=( A200  and  (not A199) );
 a53427a <=( (not A234)  and  A203 );
 a53428a <=( a53427a  and  a53424a );
 a53429a <=( a53428a  and  a53421a );
 a53432a <=( (not A236)  and  (not A235) );
 a53435a <=( (not A266)  and  (not A265) );
 a53436a <=( a53435a  and  a53432a );
 a53439a <=( A298  and  (not A268) );
 a53442a <=( A302  and  (not A299) );
 a53443a <=( a53442a  and  a53439a );
 a53444a <=( a53443a  and  a53436a );
 a53448a <=( (not A166)  and  (not A167) );
 a53449a <=( (not A169)  and  a53448a );
 a53452a <=( A200  and  (not A199) );
 a53455a <=( (not A234)  and  A203 );
 a53456a <=( a53455a  and  a53452a );
 a53457a <=( a53456a  and  a53449a );
 a53460a <=( (not A236)  and  (not A235) );
 a53463a <=( (not A266)  and  (not A265) );
 a53464a <=( a53463a  and  a53460a );
 a53467a <=( (not A298)  and  (not A268) );
 a53470a <=( A302  and  A299 );
 a53471a <=( a53470a  and  a53467a );
 a53472a <=( a53471a  and  a53464a );
 a53476a <=( (not A166)  and  (not A167) );
 a53477a <=( (not A169)  and  a53476a );
 a53480a <=( A200  and  (not A199) );
 a53483a <=( A232  and  A203 );
 a53484a <=( a53483a  and  a53480a );
 a53485a <=( a53484a  and  a53477a );
 a53488a <=( (not A234)  and  A233 );
 a53491a <=( (not A267)  and  (not A235) );
 a53492a <=( a53491a  and  a53488a );
 a53495a <=( (not A269)  and  (not A268) );
 a53498a <=( A300  and  A299 );
 a53499a <=( a53498a  and  a53495a );
 a53500a <=( a53499a  and  a53492a );
 a53504a <=( (not A166)  and  (not A167) );
 a53505a <=( (not A169)  and  a53504a );
 a53508a <=( A200  and  (not A199) );
 a53511a <=( A232  and  A203 );
 a53512a <=( a53511a  and  a53508a );
 a53513a <=( a53512a  and  a53505a );
 a53516a <=( (not A234)  and  A233 );
 a53519a <=( (not A267)  and  (not A235) );
 a53520a <=( a53519a  and  a53516a );
 a53523a <=( (not A269)  and  (not A268) );
 a53526a <=( A300  and  A298 );
 a53527a <=( a53526a  and  a53523a );
 a53528a <=( a53527a  and  a53520a );
 a53532a <=( (not A166)  and  (not A167) );
 a53533a <=( (not A169)  and  a53532a );
 a53536a <=( A200  and  (not A199) );
 a53539a <=( A232  and  A203 );
 a53540a <=( a53539a  and  a53536a );
 a53541a <=( a53540a  and  a53533a );
 a53544a <=( (not A234)  and  A233 );
 a53547a <=( A265  and  (not A235) );
 a53548a <=( a53547a  and  a53544a );
 a53551a <=( (not A267)  and  A266 );
 a53554a <=( A301  and  (not A268) );
 a53555a <=( a53554a  and  a53551a );
 a53556a <=( a53555a  and  a53548a );
 a53560a <=( (not A166)  and  (not A167) );
 a53561a <=( (not A169)  and  a53560a );
 a53564a <=( A200  and  (not A199) );
 a53567a <=( A232  and  A203 );
 a53568a <=( a53567a  and  a53564a );
 a53569a <=( a53568a  and  a53561a );
 a53572a <=( (not A234)  and  A233 );
 a53575a <=( (not A265)  and  (not A235) );
 a53576a <=( a53575a  and  a53572a );
 a53579a <=( (not A268)  and  (not A266) );
 a53582a <=( A300  and  A299 );
 a53583a <=( a53582a  and  a53579a );
 a53584a <=( a53583a  and  a53576a );
 a53588a <=( (not A166)  and  (not A167) );
 a53589a <=( (not A169)  and  a53588a );
 a53592a <=( A200  and  (not A199) );
 a53595a <=( A232  and  A203 );
 a53596a <=( a53595a  and  a53592a );
 a53597a <=( a53596a  and  a53589a );
 a53600a <=( (not A234)  and  A233 );
 a53603a <=( (not A265)  and  (not A235) );
 a53604a <=( a53603a  and  a53600a );
 a53607a <=( (not A268)  and  (not A266) );
 a53610a <=( A300  and  A298 );
 a53611a <=( a53610a  and  a53607a );
 a53612a <=( a53611a  and  a53604a );
 a53616a <=( (not A166)  and  (not A167) );
 a53617a <=( (not A169)  and  a53616a );
 a53620a <=( A200  and  (not A199) );
 a53623a <=( (not A232)  and  A203 );
 a53624a <=( a53623a  and  a53620a );
 a53625a <=( a53624a  and  a53617a );
 a53628a <=( (not A235)  and  (not A233) );
 a53631a <=( (not A268)  and  (not A267) );
 a53632a <=( a53631a  and  a53628a );
 a53635a <=( A298  and  (not A269) );
 a53638a <=( A302  and  (not A299) );
 a53639a <=( a53638a  and  a53635a );
 a53640a <=( a53639a  and  a53632a );
 a53644a <=( (not A166)  and  (not A167) );
 a53645a <=( (not A169)  and  a53644a );
 a53648a <=( A200  and  (not A199) );
 a53651a <=( (not A232)  and  A203 );
 a53652a <=( a53651a  and  a53648a );
 a53653a <=( a53652a  and  a53645a );
 a53656a <=( (not A235)  and  (not A233) );
 a53659a <=( (not A268)  and  (not A267) );
 a53660a <=( a53659a  and  a53656a );
 a53663a <=( (not A298)  and  (not A269) );
 a53666a <=( A302  and  A299 );
 a53667a <=( a53666a  and  a53663a );
 a53668a <=( a53667a  and  a53660a );
 a53672a <=( (not A166)  and  (not A167) );
 a53673a <=( (not A169)  and  a53672a );
 a53676a <=( A200  and  (not A199) );
 a53679a <=( (not A232)  and  A203 );
 a53680a <=( a53679a  and  a53676a );
 a53681a <=( a53680a  and  a53673a );
 a53684a <=( (not A235)  and  (not A233) );
 a53687a <=( A266  and  A265 );
 a53688a <=( a53687a  and  a53684a );
 a53691a <=( (not A268)  and  (not A267) );
 a53694a <=( A300  and  A299 );
 a53695a <=( a53694a  and  a53691a );
 a53696a <=( a53695a  and  a53688a );
 a53700a <=( (not A166)  and  (not A167) );
 a53701a <=( (not A169)  and  a53700a );
 a53704a <=( A200  and  (not A199) );
 a53707a <=( (not A232)  and  A203 );
 a53708a <=( a53707a  and  a53704a );
 a53709a <=( a53708a  and  a53701a );
 a53712a <=( (not A235)  and  (not A233) );
 a53715a <=( A266  and  A265 );
 a53716a <=( a53715a  and  a53712a );
 a53719a <=( (not A268)  and  (not A267) );
 a53722a <=( A300  and  A298 );
 a53723a <=( a53722a  and  a53719a );
 a53724a <=( a53723a  and  a53716a );
 a53728a <=( (not A166)  and  (not A167) );
 a53729a <=( (not A169)  and  a53728a );
 a53732a <=( A200  and  (not A199) );
 a53735a <=( (not A232)  and  A203 );
 a53736a <=( a53735a  and  a53732a );
 a53737a <=( a53736a  and  a53729a );
 a53740a <=( (not A235)  and  (not A233) );
 a53743a <=( (not A266)  and  (not A265) );
 a53744a <=( a53743a  and  a53740a );
 a53747a <=( A298  and  (not A268) );
 a53750a <=( A302  and  (not A299) );
 a53751a <=( a53750a  and  a53747a );
 a53752a <=( a53751a  and  a53744a );
 a53756a <=( (not A166)  and  (not A167) );
 a53757a <=( (not A169)  and  a53756a );
 a53760a <=( A200  and  (not A199) );
 a53763a <=( (not A232)  and  A203 );
 a53764a <=( a53763a  and  a53760a );
 a53765a <=( a53764a  and  a53757a );
 a53768a <=( (not A235)  and  (not A233) );
 a53771a <=( (not A266)  and  (not A265) );
 a53772a <=( a53771a  and  a53768a );
 a53775a <=( (not A298)  and  (not A268) );
 a53778a <=( A302  and  A299 );
 a53779a <=( a53778a  and  a53775a );
 a53780a <=( a53779a  and  a53772a );
 a53784a <=( (not A166)  and  (not A167) );
 a53785a <=( (not A169)  and  a53784a );
 a53788a <=( (not A200)  and  A199 );
 a53791a <=( (not A234)  and  A203 );
 a53792a <=( a53791a  and  a53788a );
 a53793a <=( a53792a  and  a53785a );
 a53796a <=( (not A236)  and  (not A235) );
 a53799a <=( (not A268)  and  (not A267) );
 a53800a <=( a53799a  and  a53796a );
 a53803a <=( A298  and  (not A269) );
 a53806a <=( A302  and  (not A299) );
 a53807a <=( a53806a  and  a53803a );
 a53808a <=( a53807a  and  a53800a );
 a53812a <=( (not A166)  and  (not A167) );
 a53813a <=( (not A169)  and  a53812a );
 a53816a <=( (not A200)  and  A199 );
 a53819a <=( (not A234)  and  A203 );
 a53820a <=( a53819a  and  a53816a );
 a53821a <=( a53820a  and  a53813a );
 a53824a <=( (not A236)  and  (not A235) );
 a53827a <=( (not A268)  and  (not A267) );
 a53828a <=( a53827a  and  a53824a );
 a53831a <=( (not A298)  and  (not A269) );
 a53834a <=( A302  and  A299 );
 a53835a <=( a53834a  and  a53831a );
 a53836a <=( a53835a  and  a53828a );
 a53840a <=( (not A166)  and  (not A167) );
 a53841a <=( (not A169)  and  a53840a );
 a53844a <=( (not A200)  and  A199 );
 a53847a <=( (not A234)  and  A203 );
 a53848a <=( a53847a  and  a53844a );
 a53849a <=( a53848a  and  a53841a );
 a53852a <=( (not A236)  and  (not A235) );
 a53855a <=( A266  and  A265 );
 a53856a <=( a53855a  and  a53852a );
 a53859a <=( (not A268)  and  (not A267) );
 a53862a <=( A300  and  A299 );
 a53863a <=( a53862a  and  a53859a );
 a53864a <=( a53863a  and  a53856a );
 a53868a <=( (not A166)  and  (not A167) );
 a53869a <=( (not A169)  and  a53868a );
 a53872a <=( (not A200)  and  A199 );
 a53875a <=( (not A234)  and  A203 );
 a53876a <=( a53875a  and  a53872a );
 a53877a <=( a53876a  and  a53869a );
 a53880a <=( (not A236)  and  (not A235) );
 a53883a <=( A266  and  A265 );
 a53884a <=( a53883a  and  a53880a );
 a53887a <=( (not A268)  and  (not A267) );
 a53890a <=( A300  and  A298 );
 a53891a <=( a53890a  and  a53887a );
 a53892a <=( a53891a  and  a53884a );
 a53896a <=( (not A166)  and  (not A167) );
 a53897a <=( (not A169)  and  a53896a );
 a53900a <=( (not A200)  and  A199 );
 a53903a <=( (not A234)  and  A203 );
 a53904a <=( a53903a  and  a53900a );
 a53905a <=( a53904a  and  a53897a );
 a53908a <=( (not A236)  and  (not A235) );
 a53911a <=( (not A266)  and  (not A265) );
 a53912a <=( a53911a  and  a53908a );
 a53915a <=( A298  and  (not A268) );
 a53918a <=( A302  and  (not A299) );
 a53919a <=( a53918a  and  a53915a );
 a53920a <=( a53919a  and  a53912a );
 a53924a <=( (not A166)  and  (not A167) );
 a53925a <=( (not A169)  and  a53924a );
 a53928a <=( (not A200)  and  A199 );
 a53931a <=( (not A234)  and  A203 );
 a53932a <=( a53931a  and  a53928a );
 a53933a <=( a53932a  and  a53925a );
 a53936a <=( (not A236)  and  (not A235) );
 a53939a <=( (not A266)  and  (not A265) );
 a53940a <=( a53939a  and  a53936a );
 a53943a <=( (not A298)  and  (not A268) );
 a53946a <=( A302  and  A299 );
 a53947a <=( a53946a  and  a53943a );
 a53948a <=( a53947a  and  a53940a );
 a53952a <=( (not A166)  and  (not A167) );
 a53953a <=( (not A169)  and  a53952a );
 a53956a <=( (not A200)  and  A199 );
 a53959a <=( A232  and  A203 );
 a53960a <=( a53959a  and  a53956a );
 a53961a <=( a53960a  and  a53953a );
 a53964a <=( (not A234)  and  A233 );
 a53967a <=( (not A267)  and  (not A235) );
 a53968a <=( a53967a  and  a53964a );
 a53971a <=( (not A269)  and  (not A268) );
 a53974a <=( A300  and  A299 );
 a53975a <=( a53974a  and  a53971a );
 a53976a <=( a53975a  and  a53968a );
 a53980a <=( (not A166)  and  (not A167) );
 a53981a <=( (not A169)  and  a53980a );
 a53984a <=( (not A200)  and  A199 );
 a53987a <=( A232  and  A203 );
 a53988a <=( a53987a  and  a53984a );
 a53989a <=( a53988a  and  a53981a );
 a53992a <=( (not A234)  and  A233 );
 a53995a <=( (not A267)  and  (not A235) );
 a53996a <=( a53995a  and  a53992a );
 a53999a <=( (not A269)  and  (not A268) );
 a54002a <=( A300  and  A298 );
 a54003a <=( a54002a  and  a53999a );
 a54004a <=( a54003a  and  a53996a );
 a54008a <=( (not A166)  and  (not A167) );
 a54009a <=( (not A169)  and  a54008a );
 a54012a <=( (not A200)  and  A199 );
 a54015a <=( A232  and  A203 );
 a54016a <=( a54015a  and  a54012a );
 a54017a <=( a54016a  and  a54009a );
 a54020a <=( (not A234)  and  A233 );
 a54023a <=( A265  and  (not A235) );
 a54024a <=( a54023a  and  a54020a );
 a54027a <=( (not A267)  and  A266 );
 a54030a <=( A301  and  (not A268) );
 a54031a <=( a54030a  and  a54027a );
 a54032a <=( a54031a  and  a54024a );
 a54036a <=( (not A166)  and  (not A167) );
 a54037a <=( (not A169)  and  a54036a );
 a54040a <=( (not A200)  and  A199 );
 a54043a <=( A232  and  A203 );
 a54044a <=( a54043a  and  a54040a );
 a54045a <=( a54044a  and  a54037a );
 a54048a <=( (not A234)  and  A233 );
 a54051a <=( (not A265)  and  (not A235) );
 a54052a <=( a54051a  and  a54048a );
 a54055a <=( (not A268)  and  (not A266) );
 a54058a <=( A300  and  A299 );
 a54059a <=( a54058a  and  a54055a );
 a54060a <=( a54059a  and  a54052a );
 a54064a <=( (not A166)  and  (not A167) );
 a54065a <=( (not A169)  and  a54064a );
 a54068a <=( (not A200)  and  A199 );
 a54071a <=( A232  and  A203 );
 a54072a <=( a54071a  and  a54068a );
 a54073a <=( a54072a  and  a54065a );
 a54076a <=( (not A234)  and  A233 );
 a54079a <=( (not A265)  and  (not A235) );
 a54080a <=( a54079a  and  a54076a );
 a54083a <=( (not A268)  and  (not A266) );
 a54086a <=( A300  and  A298 );
 a54087a <=( a54086a  and  a54083a );
 a54088a <=( a54087a  and  a54080a );
 a54092a <=( (not A166)  and  (not A167) );
 a54093a <=( (not A169)  and  a54092a );
 a54096a <=( (not A200)  and  A199 );
 a54099a <=( (not A232)  and  A203 );
 a54100a <=( a54099a  and  a54096a );
 a54101a <=( a54100a  and  a54093a );
 a54104a <=( (not A235)  and  (not A233) );
 a54107a <=( (not A268)  and  (not A267) );
 a54108a <=( a54107a  and  a54104a );
 a54111a <=( A298  and  (not A269) );
 a54114a <=( A302  and  (not A299) );
 a54115a <=( a54114a  and  a54111a );
 a54116a <=( a54115a  and  a54108a );
 a54120a <=( (not A166)  and  (not A167) );
 a54121a <=( (not A169)  and  a54120a );
 a54124a <=( (not A200)  and  A199 );
 a54127a <=( (not A232)  and  A203 );
 a54128a <=( a54127a  and  a54124a );
 a54129a <=( a54128a  and  a54121a );
 a54132a <=( (not A235)  and  (not A233) );
 a54135a <=( (not A268)  and  (not A267) );
 a54136a <=( a54135a  and  a54132a );
 a54139a <=( (not A298)  and  (not A269) );
 a54142a <=( A302  and  A299 );
 a54143a <=( a54142a  and  a54139a );
 a54144a <=( a54143a  and  a54136a );
 a54148a <=( (not A166)  and  (not A167) );
 a54149a <=( (not A169)  and  a54148a );
 a54152a <=( (not A200)  and  A199 );
 a54155a <=( (not A232)  and  A203 );
 a54156a <=( a54155a  and  a54152a );
 a54157a <=( a54156a  and  a54149a );
 a54160a <=( (not A235)  and  (not A233) );
 a54163a <=( A266  and  A265 );
 a54164a <=( a54163a  and  a54160a );
 a54167a <=( (not A268)  and  (not A267) );
 a54170a <=( A300  and  A299 );
 a54171a <=( a54170a  and  a54167a );
 a54172a <=( a54171a  and  a54164a );
 a54176a <=( (not A166)  and  (not A167) );
 a54177a <=( (not A169)  and  a54176a );
 a54180a <=( (not A200)  and  A199 );
 a54183a <=( (not A232)  and  A203 );
 a54184a <=( a54183a  and  a54180a );
 a54185a <=( a54184a  and  a54177a );
 a54188a <=( (not A235)  and  (not A233) );
 a54191a <=( A266  and  A265 );
 a54192a <=( a54191a  and  a54188a );
 a54195a <=( (not A268)  and  (not A267) );
 a54198a <=( A300  and  A298 );
 a54199a <=( a54198a  and  a54195a );
 a54200a <=( a54199a  and  a54192a );
 a54204a <=( (not A166)  and  (not A167) );
 a54205a <=( (not A169)  and  a54204a );
 a54208a <=( (not A200)  and  A199 );
 a54211a <=( (not A232)  and  A203 );
 a54212a <=( a54211a  and  a54208a );
 a54213a <=( a54212a  and  a54205a );
 a54216a <=( (not A235)  and  (not A233) );
 a54219a <=( (not A266)  and  (not A265) );
 a54220a <=( a54219a  and  a54216a );
 a54223a <=( A298  and  (not A268) );
 a54226a <=( A302  and  (not A299) );
 a54227a <=( a54226a  and  a54223a );
 a54228a <=( a54227a  and  a54220a );
 a54232a <=( (not A166)  and  (not A167) );
 a54233a <=( (not A169)  and  a54232a );
 a54236a <=( (not A200)  and  A199 );
 a54239a <=( (not A232)  and  A203 );
 a54240a <=( a54239a  and  a54236a );
 a54241a <=( a54240a  and  a54233a );
 a54244a <=( (not A235)  and  (not A233) );
 a54247a <=( (not A266)  and  (not A265) );
 a54248a <=( a54247a  and  a54244a );
 a54251a <=( (not A298)  and  (not A268) );
 a54254a <=( A302  and  A299 );
 a54255a <=( a54254a  and  a54251a );
 a54256a <=( a54255a  and  a54248a );
 a54260a <=( A167  and  (not A168) );
 a54261a <=( (not A169)  and  a54260a );
 a54264a <=( A202  and  A166 );
 a54267a <=( (not A235)  and  (not A234) );
 a54268a <=( a54267a  and  a54264a );
 a54269a <=( a54268a  and  a54261a );
 a54272a <=( A265  and  (not A236) );
 a54275a <=( (not A267)  and  A266 );
 a54276a <=( a54275a  and  a54272a );
 a54279a <=( A298  and  (not A268) );
 a54282a <=( A302  and  (not A299) );
 a54283a <=( a54282a  and  a54279a );
 a54284a <=( a54283a  and  a54276a );
 a54288a <=( A167  and  (not A168) );
 a54289a <=( (not A169)  and  a54288a );
 a54292a <=( A202  and  A166 );
 a54295a <=( (not A235)  and  (not A234) );
 a54296a <=( a54295a  and  a54292a );
 a54297a <=( a54296a  and  a54289a );
 a54300a <=( A265  and  (not A236) );
 a54303a <=( (not A267)  and  A266 );
 a54304a <=( a54303a  and  a54300a );
 a54307a <=( (not A298)  and  (not A268) );
 a54310a <=( A302  and  A299 );
 a54311a <=( a54310a  and  a54307a );
 a54312a <=( a54311a  and  a54304a );
 a54316a <=( A167  and  (not A168) );
 a54317a <=( (not A169)  and  a54316a );
 a54320a <=( A202  and  A166 );
 a54323a <=( A233  and  A232 );
 a54324a <=( a54323a  and  a54320a );
 a54325a <=( a54324a  and  a54317a );
 a54328a <=( (not A235)  and  (not A234) );
 a54331a <=( (not A268)  and  (not A267) );
 a54332a <=( a54331a  and  a54328a );
 a54335a <=( A298  and  (not A269) );
 a54338a <=( A302  and  (not A299) );
 a54339a <=( a54338a  and  a54335a );
 a54340a <=( a54339a  and  a54332a );
 a54344a <=( A167  and  (not A168) );
 a54345a <=( (not A169)  and  a54344a );
 a54348a <=( A202  and  A166 );
 a54351a <=( A233  and  A232 );
 a54352a <=( a54351a  and  a54348a );
 a54353a <=( a54352a  and  a54345a );
 a54356a <=( (not A235)  and  (not A234) );
 a54359a <=( (not A268)  and  (not A267) );
 a54360a <=( a54359a  and  a54356a );
 a54363a <=( (not A298)  and  (not A269) );
 a54366a <=( A302  and  A299 );
 a54367a <=( a54366a  and  a54363a );
 a54368a <=( a54367a  and  a54360a );
 a54372a <=( A167  and  (not A168) );
 a54373a <=( (not A169)  and  a54372a );
 a54376a <=( A202  and  A166 );
 a54379a <=( A233  and  A232 );
 a54380a <=( a54379a  and  a54376a );
 a54381a <=( a54380a  and  a54373a );
 a54384a <=( (not A235)  and  (not A234) );
 a54387a <=( A266  and  A265 );
 a54388a <=( a54387a  and  a54384a );
 a54391a <=( (not A268)  and  (not A267) );
 a54394a <=( A300  and  A299 );
 a54395a <=( a54394a  and  a54391a );
 a54396a <=( a54395a  and  a54388a );
 a54400a <=( A167  and  (not A168) );
 a54401a <=( (not A169)  and  a54400a );
 a54404a <=( A202  and  A166 );
 a54407a <=( A233  and  A232 );
 a54408a <=( a54407a  and  a54404a );
 a54409a <=( a54408a  and  a54401a );
 a54412a <=( (not A235)  and  (not A234) );
 a54415a <=( A266  and  A265 );
 a54416a <=( a54415a  and  a54412a );
 a54419a <=( (not A268)  and  (not A267) );
 a54422a <=( A300  and  A298 );
 a54423a <=( a54422a  and  a54419a );
 a54424a <=( a54423a  and  a54416a );
 a54428a <=( A167  and  (not A168) );
 a54429a <=( (not A169)  and  a54428a );
 a54432a <=( A202  and  A166 );
 a54435a <=( A233  and  A232 );
 a54436a <=( a54435a  and  a54432a );
 a54437a <=( a54436a  and  a54429a );
 a54440a <=( (not A235)  and  (not A234) );
 a54443a <=( (not A266)  and  (not A265) );
 a54444a <=( a54443a  and  a54440a );
 a54447a <=( A298  and  (not A268) );
 a54450a <=( A302  and  (not A299) );
 a54451a <=( a54450a  and  a54447a );
 a54452a <=( a54451a  and  a54444a );
 a54456a <=( A167  and  (not A168) );
 a54457a <=( (not A169)  and  a54456a );
 a54460a <=( A202  and  A166 );
 a54463a <=( A233  and  A232 );
 a54464a <=( a54463a  and  a54460a );
 a54465a <=( a54464a  and  a54457a );
 a54468a <=( (not A235)  and  (not A234) );
 a54471a <=( (not A266)  and  (not A265) );
 a54472a <=( a54471a  and  a54468a );
 a54475a <=( (not A298)  and  (not A268) );
 a54478a <=( A302  and  A299 );
 a54479a <=( a54478a  and  a54475a );
 a54480a <=( a54479a  and  a54472a );
 a54484a <=( A167  and  (not A168) );
 a54485a <=( (not A169)  and  a54484a );
 a54488a <=( A202  and  A166 );
 a54491a <=( (not A233)  and  (not A232) );
 a54492a <=( a54491a  and  a54488a );
 a54493a <=( a54492a  and  a54485a );
 a54496a <=( A265  and  (not A235) );
 a54499a <=( (not A267)  and  A266 );
 a54500a <=( a54499a  and  a54496a );
 a54503a <=( A298  and  (not A268) );
 a54506a <=( A302  and  (not A299) );
 a54507a <=( a54506a  and  a54503a );
 a54508a <=( a54507a  and  a54500a );
 a54512a <=( A167  and  (not A168) );
 a54513a <=( (not A169)  and  a54512a );
 a54516a <=( A202  and  A166 );
 a54519a <=( (not A233)  and  (not A232) );
 a54520a <=( a54519a  and  a54516a );
 a54521a <=( a54520a  and  a54513a );
 a54524a <=( A265  and  (not A235) );
 a54527a <=( (not A267)  and  A266 );
 a54528a <=( a54527a  and  a54524a );
 a54531a <=( (not A298)  and  (not A268) );
 a54534a <=( A302  and  A299 );
 a54535a <=( a54534a  and  a54531a );
 a54536a <=( a54535a  and  a54528a );
 a54540a <=( A167  and  (not A168) );
 a54541a <=( (not A169)  and  a54540a );
 a54544a <=( A199  and  A166 );
 a54547a <=( (not A234)  and  A201 );
 a54548a <=( a54547a  and  a54544a );
 a54549a <=( a54548a  and  a54541a );
 a54552a <=( (not A236)  and  (not A235) );
 a54555a <=( (not A268)  and  (not A267) );
 a54556a <=( a54555a  and  a54552a );
 a54559a <=( A298  and  (not A269) );
 a54562a <=( A302  and  (not A299) );
 a54563a <=( a54562a  and  a54559a );
 a54564a <=( a54563a  and  a54556a );
 a54568a <=( A167  and  (not A168) );
 a54569a <=( (not A169)  and  a54568a );
 a54572a <=( A199  and  A166 );
 a54575a <=( (not A234)  and  A201 );
 a54576a <=( a54575a  and  a54572a );
 a54577a <=( a54576a  and  a54569a );
 a54580a <=( (not A236)  and  (not A235) );
 a54583a <=( (not A268)  and  (not A267) );
 a54584a <=( a54583a  and  a54580a );
 a54587a <=( (not A298)  and  (not A269) );
 a54590a <=( A302  and  A299 );
 a54591a <=( a54590a  and  a54587a );
 a54592a <=( a54591a  and  a54584a );
 a54596a <=( A167  and  (not A168) );
 a54597a <=( (not A169)  and  a54596a );
 a54600a <=( A199  and  A166 );
 a54603a <=( (not A234)  and  A201 );
 a54604a <=( a54603a  and  a54600a );
 a54605a <=( a54604a  and  a54597a );
 a54608a <=( (not A236)  and  (not A235) );
 a54611a <=( A266  and  A265 );
 a54612a <=( a54611a  and  a54608a );
 a54615a <=( (not A268)  and  (not A267) );
 a54618a <=( A300  and  A299 );
 a54619a <=( a54618a  and  a54615a );
 a54620a <=( a54619a  and  a54612a );
 a54624a <=( A167  and  (not A168) );
 a54625a <=( (not A169)  and  a54624a );
 a54628a <=( A199  and  A166 );
 a54631a <=( (not A234)  and  A201 );
 a54632a <=( a54631a  and  a54628a );
 a54633a <=( a54632a  and  a54625a );
 a54636a <=( (not A236)  and  (not A235) );
 a54639a <=( A266  and  A265 );
 a54640a <=( a54639a  and  a54636a );
 a54643a <=( (not A268)  and  (not A267) );
 a54646a <=( A300  and  A298 );
 a54647a <=( a54646a  and  a54643a );
 a54648a <=( a54647a  and  a54640a );
 a54652a <=( A167  and  (not A168) );
 a54653a <=( (not A169)  and  a54652a );
 a54656a <=( A199  and  A166 );
 a54659a <=( (not A234)  and  A201 );
 a54660a <=( a54659a  and  a54656a );
 a54661a <=( a54660a  and  a54653a );
 a54664a <=( (not A236)  and  (not A235) );
 a54667a <=( (not A266)  and  (not A265) );
 a54668a <=( a54667a  and  a54664a );
 a54671a <=( A298  and  (not A268) );
 a54674a <=( A302  and  (not A299) );
 a54675a <=( a54674a  and  a54671a );
 a54676a <=( a54675a  and  a54668a );
 a54680a <=( A167  and  (not A168) );
 a54681a <=( (not A169)  and  a54680a );
 a54684a <=( A199  and  A166 );
 a54687a <=( (not A234)  and  A201 );
 a54688a <=( a54687a  and  a54684a );
 a54689a <=( a54688a  and  a54681a );
 a54692a <=( (not A236)  and  (not A235) );
 a54695a <=( (not A266)  and  (not A265) );
 a54696a <=( a54695a  and  a54692a );
 a54699a <=( (not A298)  and  (not A268) );
 a54702a <=( A302  and  A299 );
 a54703a <=( a54702a  and  a54699a );
 a54704a <=( a54703a  and  a54696a );
 a54708a <=( A167  and  (not A168) );
 a54709a <=( (not A169)  and  a54708a );
 a54712a <=( A199  and  A166 );
 a54715a <=( A232  and  A201 );
 a54716a <=( a54715a  and  a54712a );
 a54717a <=( a54716a  and  a54709a );
 a54720a <=( (not A234)  and  A233 );
 a54723a <=( (not A267)  and  (not A235) );
 a54724a <=( a54723a  and  a54720a );
 a54727a <=( (not A269)  and  (not A268) );
 a54730a <=( A300  and  A299 );
 a54731a <=( a54730a  and  a54727a );
 a54732a <=( a54731a  and  a54724a );
 a54736a <=( A167  and  (not A168) );
 a54737a <=( (not A169)  and  a54736a );
 a54740a <=( A199  and  A166 );
 a54743a <=( A232  and  A201 );
 a54744a <=( a54743a  and  a54740a );
 a54745a <=( a54744a  and  a54737a );
 a54748a <=( (not A234)  and  A233 );
 a54751a <=( (not A267)  and  (not A235) );
 a54752a <=( a54751a  and  a54748a );
 a54755a <=( (not A269)  and  (not A268) );
 a54758a <=( A300  and  A298 );
 a54759a <=( a54758a  and  a54755a );
 a54760a <=( a54759a  and  a54752a );
 a54764a <=( A167  and  (not A168) );
 a54765a <=( (not A169)  and  a54764a );
 a54768a <=( A199  and  A166 );
 a54771a <=( A232  and  A201 );
 a54772a <=( a54771a  and  a54768a );
 a54773a <=( a54772a  and  a54765a );
 a54776a <=( (not A234)  and  A233 );
 a54779a <=( A265  and  (not A235) );
 a54780a <=( a54779a  and  a54776a );
 a54783a <=( (not A267)  and  A266 );
 a54786a <=( A301  and  (not A268) );
 a54787a <=( a54786a  and  a54783a );
 a54788a <=( a54787a  and  a54780a );
 a54792a <=( A167  and  (not A168) );
 a54793a <=( (not A169)  and  a54792a );
 a54796a <=( A199  and  A166 );
 a54799a <=( A232  and  A201 );
 a54800a <=( a54799a  and  a54796a );
 a54801a <=( a54800a  and  a54793a );
 a54804a <=( (not A234)  and  A233 );
 a54807a <=( (not A265)  and  (not A235) );
 a54808a <=( a54807a  and  a54804a );
 a54811a <=( (not A268)  and  (not A266) );
 a54814a <=( A300  and  A299 );
 a54815a <=( a54814a  and  a54811a );
 a54816a <=( a54815a  and  a54808a );
 a54820a <=( A167  and  (not A168) );
 a54821a <=( (not A169)  and  a54820a );
 a54824a <=( A199  and  A166 );
 a54827a <=( A232  and  A201 );
 a54828a <=( a54827a  and  a54824a );
 a54829a <=( a54828a  and  a54821a );
 a54832a <=( (not A234)  and  A233 );
 a54835a <=( (not A265)  and  (not A235) );
 a54836a <=( a54835a  and  a54832a );
 a54839a <=( (not A268)  and  (not A266) );
 a54842a <=( A300  and  A298 );
 a54843a <=( a54842a  and  a54839a );
 a54844a <=( a54843a  and  a54836a );
 a54848a <=( A167  and  (not A168) );
 a54849a <=( (not A169)  and  a54848a );
 a54852a <=( A199  and  A166 );
 a54855a <=( (not A232)  and  A201 );
 a54856a <=( a54855a  and  a54852a );
 a54857a <=( a54856a  and  a54849a );
 a54860a <=( (not A235)  and  (not A233) );
 a54863a <=( (not A268)  and  (not A267) );
 a54864a <=( a54863a  and  a54860a );
 a54867a <=( A298  and  (not A269) );
 a54870a <=( A302  and  (not A299) );
 a54871a <=( a54870a  and  a54867a );
 a54872a <=( a54871a  and  a54864a );
 a54876a <=( A167  and  (not A168) );
 a54877a <=( (not A169)  and  a54876a );
 a54880a <=( A199  and  A166 );
 a54883a <=( (not A232)  and  A201 );
 a54884a <=( a54883a  and  a54880a );
 a54885a <=( a54884a  and  a54877a );
 a54888a <=( (not A235)  and  (not A233) );
 a54891a <=( (not A268)  and  (not A267) );
 a54892a <=( a54891a  and  a54888a );
 a54895a <=( (not A298)  and  (not A269) );
 a54898a <=( A302  and  A299 );
 a54899a <=( a54898a  and  a54895a );
 a54900a <=( a54899a  and  a54892a );
 a54904a <=( A167  and  (not A168) );
 a54905a <=( (not A169)  and  a54904a );
 a54908a <=( A199  and  A166 );
 a54911a <=( (not A232)  and  A201 );
 a54912a <=( a54911a  and  a54908a );
 a54913a <=( a54912a  and  a54905a );
 a54916a <=( (not A235)  and  (not A233) );
 a54919a <=( A266  and  A265 );
 a54920a <=( a54919a  and  a54916a );
 a54923a <=( (not A268)  and  (not A267) );
 a54926a <=( A300  and  A299 );
 a54927a <=( a54926a  and  a54923a );
 a54928a <=( a54927a  and  a54920a );
 a54932a <=( A167  and  (not A168) );
 a54933a <=( (not A169)  and  a54932a );
 a54936a <=( A199  and  A166 );
 a54939a <=( (not A232)  and  A201 );
 a54940a <=( a54939a  and  a54936a );
 a54941a <=( a54940a  and  a54933a );
 a54944a <=( (not A235)  and  (not A233) );
 a54947a <=( A266  and  A265 );
 a54948a <=( a54947a  and  a54944a );
 a54951a <=( (not A268)  and  (not A267) );
 a54954a <=( A300  and  A298 );
 a54955a <=( a54954a  and  a54951a );
 a54956a <=( a54955a  and  a54948a );
 a54960a <=( A167  and  (not A168) );
 a54961a <=( (not A169)  and  a54960a );
 a54964a <=( A199  and  A166 );
 a54967a <=( (not A232)  and  A201 );
 a54968a <=( a54967a  and  a54964a );
 a54969a <=( a54968a  and  a54961a );
 a54972a <=( (not A235)  and  (not A233) );
 a54975a <=( (not A266)  and  (not A265) );
 a54976a <=( a54975a  and  a54972a );
 a54979a <=( A298  and  (not A268) );
 a54982a <=( A302  and  (not A299) );
 a54983a <=( a54982a  and  a54979a );
 a54984a <=( a54983a  and  a54976a );
 a54988a <=( A167  and  (not A168) );
 a54989a <=( (not A169)  and  a54988a );
 a54992a <=( A199  and  A166 );
 a54995a <=( (not A232)  and  A201 );
 a54996a <=( a54995a  and  a54992a );
 a54997a <=( a54996a  and  a54989a );
 a55000a <=( (not A235)  and  (not A233) );
 a55003a <=( (not A266)  and  (not A265) );
 a55004a <=( a55003a  and  a55000a );
 a55007a <=( (not A298)  and  (not A268) );
 a55010a <=( A302  and  A299 );
 a55011a <=( a55010a  and  a55007a );
 a55012a <=( a55011a  and  a55004a );
 a55016a <=( A167  and  (not A168) );
 a55017a <=( (not A169)  and  a55016a );
 a55020a <=( A200  and  A166 );
 a55023a <=( (not A234)  and  A201 );
 a55024a <=( a55023a  and  a55020a );
 a55025a <=( a55024a  and  a55017a );
 a55028a <=( (not A236)  and  (not A235) );
 a55031a <=( (not A268)  and  (not A267) );
 a55032a <=( a55031a  and  a55028a );
 a55035a <=( A298  and  (not A269) );
 a55038a <=( A302  and  (not A299) );
 a55039a <=( a55038a  and  a55035a );
 a55040a <=( a55039a  and  a55032a );
 a55044a <=( A167  and  (not A168) );
 a55045a <=( (not A169)  and  a55044a );
 a55048a <=( A200  and  A166 );
 a55051a <=( (not A234)  and  A201 );
 a55052a <=( a55051a  and  a55048a );
 a55053a <=( a55052a  and  a55045a );
 a55056a <=( (not A236)  and  (not A235) );
 a55059a <=( (not A268)  and  (not A267) );
 a55060a <=( a55059a  and  a55056a );
 a55063a <=( (not A298)  and  (not A269) );
 a55066a <=( A302  and  A299 );
 a55067a <=( a55066a  and  a55063a );
 a55068a <=( a55067a  and  a55060a );
 a55072a <=( A167  and  (not A168) );
 a55073a <=( (not A169)  and  a55072a );
 a55076a <=( A200  and  A166 );
 a55079a <=( (not A234)  and  A201 );
 a55080a <=( a55079a  and  a55076a );
 a55081a <=( a55080a  and  a55073a );
 a55084a <=( (not A236)  and  (not A235) );
 a55087a <=( A266  and  A265 );
 a55088a <=( a55087a  and  a55084a );
 a55091a <=( (not A268)  and  (not A267) );
 a55094a <=( A300  and  A299 );
 a55095a <=( a55094a  and  a55091a );
 a55096a <=( a55095a  and  a55088a );
 a55100a <=( A167  and  (not A168) );
 a55101a <=( (not A169)  and  a55100a );
 a55104a <=( A200  and  A166 );
 a55107a <=( (not A234)  and  A201 );
 a55108a <=( a55107a  and  a55104a );
 a55109a <=( a55108a  and  a55101a );
 a55112a <=( (not A236)  and  (not A235) );
 a55115a <=( A266  and  A265 );
 a55116a <=( a55115a  and  a55112a );
 a55119a <=( (not A268)  and  (not A267) );
 a55122a <=( A300  and  A298 );
 a55123a <=( a55122a  and  a55119a );
 a55124a <=( a55123a  and  a55116a );
 a55128a <=( A167  and  (not A168) );
 a55129a <=( (not A169)  and  a55128a );
 a55132a <=( A200  and  A166 );
 a55135a <=( (not A234)  and  A201 );
 a55136a <=( a55135a  and  a55132a );
 a55137a <=( a55136a  and  a55129a );
 a55140a <=( (not A236)  and  (not A235) );
 a55143a <=( (not A266)  and  (not A265) );
 a55144a <=( a55143a  and  a55140a );
 a55147a <=( A298  and  (not A268) );
 a55150a <=( A302  and  (not A299) );
 a55151a <=( a55150a  and  a55147a );
 a55152a <=( a55151a  and  a55144a );
 a55156a <=( A167  and  (not A168) );
 a55157a <=( (not A169)  and  a55156a );
 a55160a <=( A200  and  A166 );
 a55163a <=( (not A234)  and  A201 );
 a55164a <=( a55163a  and  a55160a );
 a55165a <=( a55164a  and  a55157a );
 a55168a <=( (not A236)  and  (not A235) );
 a55171a <=( (not A266)  and  (not A265) );
 a55172a <=( a55171a  and  a55168a );
 a55175a <=( (not A298)  and  (not A268) );
 a55178a <=( A302  and  A299 );
 a55179a <=( a55178a  and  a55175a );
 a55180a <=( a55179a  and  a55172a );
 a55184a <=( A167  and  (not A168) );
 a55185a <=( (not A169)  and  a55184a );
 a55188a <=( A200  and  A166 );
 a55191a <=( A232  and  A201 );
 a55192a <=( a55191a  and  a55188a );
 a55193a <=( a55192a  and  a55185a );
 a55196a <=( (not A234)  and  A233 );
 a55199a <=( (not A267)  and  (not A235) );
 a55200a <=( a55199a  and  a55196a );
 a55203a <=( (not A269)  and  (not A268) );
 a55206a <=( A300  and  A299 );
 a55207a <=( a55206a  and  a55203a );
 a55208a <=( a55207a  and  a55200a );
 a55212a <=( A167  and  (not A168) );
 a55213a <=( (not A169)  and  a55212a );
 a55216a <=( A200  and  A166 );
 a55219a <=( A232  and  A201 );
 a55220a <=( a55219a  and  a55216a );
 a55221a <=( a55220a  and  a55213a );
 a55224a <=( (not A234)  and  A233 );
 a55227a <=( (not A267)  and  (not A235) );
 a55228a <=( a55227a  and  a55224a );
 a55231a <=( (not A269)  and  (not A268) );
 a55234a <=( A300  and  A298 );
 a55235a <=( a55234a  and  a55231a );
 a55236a <=( a55235a  and  a55228a );
 a55240a <=( A167  and  (not A168) );
 a55241a <=( (not A169)  and  a55240a );
 a55244a <=( A200  and  A166 );
 a55247a <=( A232  and  A201 );
 a55248a <=( a55247a  and  a55244a );
 a55249a <=( a55248a  and  a55241a );
 a55252a <=( (not A234)  and  A233 );
 a55255a <=( A265  and  (not A235) );
 a55256a <=( a55255a  and  a55252a );
 a55259a <=( (not A267)  and  A266 );
 a55262a <=( A301  and  (not A268) );
 a55263a <=( a55262a  and  a55259a );
 a55264a <=( a55263a  and  a55256a );
 a55268a <=( A167  and  (not A168) );
 a55269a <=( (not A169)  and  a55268a );
 a55272a <=( A200  and  A166 );
 a55275a <=( A232  and  A201 );
 a55276a <=( a55275a  and  a55272a );
 a55277a <=( a55276a  and  a55269a );
 a55280a <=( (not A234)  and  A233 );
 a55283a <=( (not A265)  and  (not A235) );
 a55284a <=( a55283a  and  a55280a );
 a55287a <=( (not A268)  and  (not A266) );
 a55290a <=( A300  and  A299 );
 a55291a <=( a55290a  and  a55287a );
 a55292a <=( a55291a  and  a55284a );
 a55296a <=( A167  and  (not A168) );
 a55297a <=( (not A169)  and  a55296a );
 a55300a <=( A200  and  A166 );
 a55303a <=( A232  and  A201 );
 a55304a <=( a55303a  and  a55300a );
 a55305a <=( a55304a  and  a55297a );
 a55308a <=( (not A234)  and  A233 );
 a55311a <=( (not A265)  and  (not A235) );
 a55312a <=( a55311a  and  a55308a );
 a55315a <=( (not A268)  and  (not A266) );
 a55318a <=( A300  and  A298 );
 a55319a <=( a55318a  and  a55315a );
 a55320a <=( a55319a  and  a55312a );
 a55324a <=( A167  and  (not A168) );
 a55325a <=( (not A169)  and  a55324a );
 a55328a <=( A200  and  A166 );
 a55331a <=( (not A232)  and  A201 );
 a55332a <=( a55331a  and  a55328a );
 a55333a <=( a55332a  and  a55325a );
 a55336a <=( (not A235)  and  (not A233) );
 a55339a <=( (not A268)  and  (not A267) );
 a55340a <=( a55339a  and  a55336a );
 a55343a <=( A298  and  (not A269) );
 a55346a <=( A302  and  (not A299) );
 a55347a <=( a55346a  and  a55343a );
 a55348a <=( a55347a  and  a55340a );
 a55352a <=( A167  and  (not A168) );
 a55353a <=( (not A169)  and  a55352a );
 a55356a <=( A200  and  A166 );
 a55359a <=( (not A232)  and  A201 );
 a55360a <=( a55359a  and  a55356a );
 a55361a <=( a55360a  and  a55353a );
 a55364a <=( (not A235)  and  (not A233) );
 a55367a <=( (not A268)  and  (not A267) );
 a55368a <=( a55367a  and  a55364a );
 a55371a <=( (not A298)  and  (not A269) );
 a55374a <=( A302  and  A299 );
 a55375a <=( a55374a  and  a55371a );
 a55376a <=( a55375a  and  a55368a );
 a55380a <=( A167  and  (not A168) );
 a55381a <=( (not A169)  and  a55380a );
 a55384a <=( A200  and  A166 );
 a55387a <=( (not A232)  and  A201 );
 a55388a <=( a55387a  and  a55384a );
 a55389a <=( a55388a  and  a55381a );
 a55392a <=( (not A235)  and  (not A233) );
 a55395a <=( A266  and  A265 );
 a55396a <=( a55395a  and  a55392a );
 a55399a <=( (not A268)  and  (not A267) );
 a55402a <=( A300  and  A299 );
 a55403a <=( a55402a  and  a55399a );
 a55404a <=( a55403a  and  a55396a );
 a55408a <=( A167  and  (not A168) );
 a55409a <=( (not A169)  and  a55408a );
 a55412a <=( A200  and  A166 );
 a55415a <=( (not A232)  and  A201 );
 a55416a <=( a55415a  and  a55412a );
 a55417a <=( a55416a  and  a55409a );
 a55420a <=( (not A235)  and  (not A233) );
 a55423a <=( A266  and  A265 );
 a55424a <=( a55423a  and  a55420a );
 a55427a <=( (not A268)  and  (not A267) );
 a55430a <=( A300  and  A298 );
 a55431a <=( a55430a  and  a55427a );
 a55432a <=( a55431a  and  a55424a );
 a55436a <=( A167  and  (not A168) );
 a55437a <=( (not A169)  and  a55436a );
 a55440a <=( A200  and  A166 );
 a55443a <=( (not A232)  and  A201 );
 a55444a <=( a55443a  and  a55440a );
 a55445a <=( a55444a  and  a55437a );
 a55448a <=( (not A235)  and  (not A233) );
 a55451a <=( (not A266)  and  (not A265) );
 a55452a <=( a55451a  and  a55448a );
 a55455a <=( A298  and  (not A268) );
 a55458a <=( A302  and  (not A299) );
 a55459a <=( a55458a  and  a55455a );
 a55460a <=( a55459a  and  a55452a );
 a55464a <=( A167  and  (not A168) );
 a55465a <=( (not A169)  and  a55464a );
 a55468a <=( A200  and  A166 );
 a55471a <=( (not A232)  and  A201 );
 a55472a <=( a55471a  and  a55468a );
 a55473a <=( a55472a  and  a55465a );
 a55476a <=( (not A235)  and  (not A233) );
 a55479a <=( (not A266)  and  (not A265) );
 a55480a <=( a55479a  and  a55476a );
 a55483a <=( (not A298)  and  (not A268) );
 a55486a <=( A302  and  A299 );
 a55487a <=( a55486a  and  a55483a );
 a55488a <=( a55487a  and  a55480a );
 a55492a <=( A167  and  (not A168) );
 a55493a <=( (not A169)  and  a55492a );
 a55496a <=( (not A199)  and  A166 );
 a55499a <=( A203  and  A200 );
 a55500a <=( a55499a  and  a55496a );
 a55501a <=( a55500a  and  a55493a );
 a55504a <=( (not A235)  and  (not A234) );
 a55507a <=( (not A267)  and  (not A236) );
 a55508a <=( a55507a  and  a55504a );
 a55511a <=( (not A269)  and  (not A268) );
 a55514a <=( A300  and  A299 );
 a55515a <=( a55514a  and  a55511a );
 a55516a <=( a55515a  and  a55508a );
 a55520a <=( A167  and  (not A168) );
 a55521a <=( (not A169)  and  a55520a );
 a55524a <=( (not A199)  and  A166 );
 a55527a <=( A203  and  A200 );
 a55528a <=( a55527a  and  a55524a );
 a55529a <=( a55528a  and  a55521a );
 a55532a <=( (not A235)  and  (not A234) );
 a55535a <=( (not A267)  and  (not A236) );
 a55536a <=( a55535a  and  a55532a );
 a55539a <=( (not A269)  and  (not A268) );
 a55542a <=( A300  and  A298 );
 a55543a <=( a55542a  and  a55539a );
 a55544a <=( a55543a  and  a55536a );
 a55548a <=( A167  and  (not A168) );
 a55549a <=( (not A169)  and  a55548a );
 a55552a <=( (not A199)  and  A166 );
 a55555a <=( A203  and  A200 );
 a55556a <=( a55555a  and  a55552a );
 a55557a <=( a55556a  and  a55549a );
 a55560a <=( (not A235)  and  (not A234) );
 a55563a <=( A265  and  (not A236) );
 a55564a <=( a55563a  and  a55560a );
 a55567a <=( (not A267)  and  A266 );
 a55570a <=( A301  and  (not A268) );
 a55571a <=( a55570a  and  a55567a );
 a55572a <=( a55571a  and  a55564a );
 a55576a <=( A167  and  (not A168) );
 a55577a <=( (not A169)  and  a55576a );
 a55580a <=( (not A199)  and  A166 );
 a55583a <=( A203  and  A200 );
 a55584a <=( a55583a  and  a55580a );
 a55585a <=( a55584a  and  a55577a );
 a55588a <=( (not A235)  and  (not A234) );
 a55591a <=( (not A265)  and  (not A236) );
 a55592a <=( a55591a  and  a55588a );
 a55595a <=( (not A268)  and  (not A266) );
 a55598a <=( A300  and  A299 );
 a55599a <=( a55598a  and  a55595a );
 a55600a <=( a55599a  and  a55592a );
 a55604a <=( A167  and  (not A168) );
 a55605a <=( (not A169)  and  a55604a );
 a55608a <=( (not A199)  and  A166 );
 a55611a <=( A203  and  A200 );
 a55612a <=( a55611a  and  a55608a );
 a55613a <=( a55612a  and  a55605a );
 a55616a <=( (not A235)  and  (not A234) );
 a55619a <=( (not A265)  and  (not A236) );
 a55620a <=( a55619a  and  a55616a );
 a55623a <=( (not A268)  and  (not A266) );
 a55626a <=( A300  and  A298 );
 a55627a <=( a55626a  and  a55623a );
 a55628a <=( a55627a  and  a55620a );
 a55632a <=( A167  and  (not A168) );
 a55633a <=( (not A169)  and  a55632a );
 a55636a <=( (not A199)  and  A166 );
 a55639a <=( A203  and  A200 );
 a55640a <=( a55639a  and  a55636a );
 a55641a <=( a55640a  and  a55633a );
 a55644a <=( A233  and  A232 );
 a55647a <=( (not A235)  and  (not A234) );
 a55648a <=( a55647a  and  a55644a );
 a55651a <=( (not A268)  and  (not A267) );
 a55654a <=( A301  and  (not A269) );
 a55655a <=( a55654a  and  a55651a );
 a55656a <=( a55655a  and  a55648a );
 a55660a <=( A167  and  (not A168) );
 a55661a <=( (not A169)  and  a55660a );
 a55664a <=( (not A199)  and  A166 );
 a55667a <=( A203  and  A200 );
 a55668a <=( a55667a  and  a55664a );
 a55669a <=( a55668a  and  a55661a );
 a55672a <=( A233  and  A232 );
 a55675a <=( (not A235)  and  (not A234) );
 a55676a <=( a55675a  and  a55672a );
 a55679a <=( (not A266)  and  (not A265) );
 a55682a <=( A301  and  (not A268) );
 a55683a <=( a55682a  and  a55679a );
 a55684a <=( a55683a  and  a55676a );
 a55688a <=( A167  and  (not A168) );
 a55689a <=( (not A169)  and  a55688a );
 a55692a <=( (not A199)  and  A166 );
 a55695a <=( A203  and  A200 );
 a55696a <=( a55695a  and  a55692a );
 a55697a <=( a55696a  and  a55689a );
 a55700a <=( (not A233)  and  (not A232) );
 a55703a <=( (not A267)  and  (not A235) );
 a55704a <=( a55703a  and  a55700a );
 a55707a <=( (not A269)  and  (not A268) );
 a55710a <=( A300  and  A299 );
 a55711a <=( a55710a  and  a55707a );
 a55712a <=( a55711a  and  a55704a );
 a55716a <=( A167  and  (not A168) );
 a55717a <=( (not A169)  and  a55716a );
 a55720a <=( (not A199)  and  A166 );
 a55723a <=( A203  and  A200 );
 a55724a <=( a55723a  and  a55720a );
 a55725a <=( a55724a  and  a55717a );
 a55728a <=( (not A233)  and  (not A232) );
 a55731a <=( (not A267)  and  (not A235) );
 a55732a <=( a55731a  and  a55728a );
 a55735a <=( (not A269)  and  (not A268) );
 a55738a <=( A300  and  A298 );
 a55739a <=( a55738a  and  a55735a );
 a55740a <=( a55739a  and  a55732a );
 a55744a <=( A167  and  (not A168) );
 a55745a <=( (not A169)  and  a55744a );
 a55748a <=( (not A199)  and  A166 );
 a55751a <=( A203  and  A200 );
 a55752a <=( a55751a  and  a55748a );
 a55753a <=( a55752a  and  a55745a );
 a55756a <=( (not A233)  and  (not A232) );
 a55759a <=( A265  and  (not A235) );
 a55760a <=( a55759a  and  a55756a );
 a55763a <=( (not A267)  and  A266 );
 a55766a <=( A301  and  (not A268) );
 a55767a <=( a55766a  and  a55763a );
 a55768a <=( a55767a  and  a55760a );
 a55772a <=( A167  and  (not A168) );
 a55773a <=( (not A169)  and  a55772a );
 a55776a <=( (not A199)  and  A166 );
 a55779a <=( A203  and  A200 );
 a55780a <=( a55779a  and  a55776a );
 a55781a <=( a55780a  and  a55773a );
 a55784a <=( (not A233)  and  (not A232) );
 a55787a <=( (not A265)  and  (not A235) );
 a55788a <=( a55787a  and  a55784a );
 a55791a <=( (not A268)  and  (not A266) );
 a55794a <=( A300  and  A299 );
 a55795a <=( a55794a  and  a55791a );
 a55796a <=( a55795a  and  a55788a );
 a55800a <=( A167  and  (not A168) );
 a55801a <=( (not A169)  and  a55800a );
 a55804a <=( (not A199)  and  A166 );
 a55807a <=( A203  and  A200 );
 a55808a <=( a55807a  and  a55804a );
 a55809a <=( a55808a  and  a55801a );
 a55812a <=( (not A233)  and  (not A232) );
 a55815a <=( (not A265)  and  (not A235) );
 a55816a <=( a55815a  and  a55812a );
 a55819a <=( (not A268)  and  (not A266) );
 a55822a <=( A300  and  A298 );
 a55823a <=( a55822a  and  a55819a );
 a55824a <=( a55823a  and  a55816a );
 a55828a <=( A167  and  (not A168) );
 a55829a <=( (not A169)  and  a55828a );
 a55832a <=( A199  and  A166 );
 a55835a <=( A203  and  (not A200) );
 a55836a <=( a55835a  and  a55832a );
 a55837a <=( a55836a  and  a55829a );
 a55840a <=( (not A235)  and  (not A234) );
 a55843a <=( (not A267)  and  (not A236) );
 a55844a <=( a55843a  and  a55840a );
 a55847a <=( (not A269)  and  (not A268) );
 a55850a <=( A300  and  A299 );
 a55851a <=( a55850a  and  a55847a );
 a55852a <=( a55851a  and  a55844a );
 a55856a <=( A167  and  (not A168) );
 a55857a <=( (not A169)  and  a55856a );
 a55860a <=( A199  and  A166 );
 a55863a <=( A203  and  (not A200) );
 a55864a <=( a55863a  and  a55860a );
 a55865a <=( a55864a  and  a55857a );
 a55868a <=( (not A235)  and  (not A234) );
 a55871a <=( (not A267)  and  (not A236) );
 a55872a <=( a55871a  and  a55868a );
 a55875a <=( (not A269)  and  (not A268) );
 a55878a <=( A300  and  A298 );
 a55879a <=( a55878a  and  a55875a );
 a55880a <=( a55879a  and  a55872a );
 a55884a <=( A167  and  (not A168) );
 a55885a <=( (not A169)  and  a55884a );
 a55888a <=( A199  and  A166 );
 a55891a <=( A203  and  (not A200) );
 a55892a <=( a55891a  and  a55888a );
 a55893a <=( a55892a  and  a55885a );
 a55896a <=( (not A235)  and  (not A234) );
 a55899a <=( A265  and  (not A236) );
 a55900a <=( a55899a  and  a55896a );
 a55903a <=( (not A267)  and  A266 );
 a55906a <=( A301  and  (not A268) );
 a55907a <=( a55906a  and  a55903a );
 a55908a <=( a55907a  and  a55900a );
 a55912a <=( A167  and  (not A168) );
 a55913a <=( (not A169)  and  a55912a );
 a55916a <=( A199  and  A166 );
 a55919a <=( A203  and  (not A200) );
 a55920a <=( a55919a  and  a55916a );
 a55921a <=( a55920a  and  a55913a );
 a55924a <=( (not A235)  and  (not A234) );
 a55927a <=( (not A265)  and  (not A236) );
 a55928a <=( a55927a  and  a55924a );
 a55931a <=( (not A268)  and  (not A266) );
 a55934a <=( A300  and  A299 );
 a55935a <=( a55934a  and  a55931a );
 a55936a <=( a55935a  and  a55928a );
 a55940a <=( A167  and  (not A168) );
 a55941a <=( (not A169)  and  a55940a );
 a55944a <=( A199  and  A166 );
 a55947a <=( A203  and  (not A200) );
 a55948a <=( a55947a  and  a55944a );
 a55949a <=( a55948a  and  a55941a );
 a55952a <=( (not A235)  and  (not A234) );
 a55955a <=( (not A265)  and  (not A236) );
 a55956a <=( a55955a  and  a55952a );
 a55959a <=( (not A268)  and  (not A266) );
 a55962a <=( A300  and  A298 );
 a55963a <=( a55962a  and  a55959a );
 a55964a <=( a55963a  and  a55956a );
 a55968a <=( A167  and  (not A168) );
 a55969a <=( (not A169)  and  a55968a );
 a55972a <=( A199  and  A166 );
 a55975a <=( A203  and  (not A200) );
 a55976a <=( a55975a  and  a55972a );
 a55977a <=( a55976a  and  a55969a );
 a55980a <=( A233  and  A232 );
 a55983a <=( (not A235)  and  (not A234) );
 a55984a <=( a55983a  and  a55980a );
 a55987a <=( (not A268)  and  (not A267) );
 a55990a <=( A301  and  (not A269) );
 a55991a <=( a55990a  and  a55987a );
 a55992a <=( a55991a  and  a55984a );
 a55996a <=( A167  and  (not A168) );
 a55997a <=( (not A169)  and  a55996a );
 a56000a <=( A199  and  A166 );
 a56003a <=( A203  and  (not A200) );
 a56004a <=( a56003a  and  a56000a );
 a56005a <=( a56004a  and  a55997a );
 a56008a <=( A233  and  A232 );
 a56011a <=( (not A235)  and  (not A234) );
 a56012a <=( a56011a  and  a56008a );
 a56015a <=( (not A266)  and  (not A265) );
 a56018a <=( A301  and  (not A268) );
 a56019a <=( a56018a  and  a56015a );
 a56020a <=( a56019a  and  a56012a );
 a56024a <=( A167  and  (not A168) );
 a56025a <=( (not A169)  and  a56024a );
 a56028a <=( A199  and  A166 );
 a56031a <=( A203  and  (not A200) );
 a56032a <=( a56031a  and  a56028a );
 a56033a <=( a56032a  and  a56025a );
 a56036a <=( (not A233)  and  (not A232) );
 a56039a <=( (not A267)  and  (not A235) );
 a56040a <=( a56039a  and  a56036a );
 a56043a <=( (not A269)  and  (not A268) );
 a56046a <=( A300  and  A299 );
 a56047a <=( a56046a  and  a56043a );
 a56048a <=( a56047a  and  a56040a );
 a56052a <=( A167  and  (not A168) );
 a56053a <=( (not A169)  and  a56052a );
 a56056a <=( A199  and  A166 );
 a56059a <=( A203  and  (not A200) );
 a56060a <=( a56059a  and  a56056a );
 a56061a <=( a56060a  and  a56053a );
 a56064a <=( (not A233)  and  (not A232) );
 a56067a <=( (not A267)  and  (not A235) );
 a56068a <=( a56067a  and  a56064a );
 a56071a <=( (not A269)  and  (not A268) );
 a56074a <=( A300  and  A298 );
 a56075a <=( a56074a  and  a56071a );
 a56076a <=( a56075a  and  a56068a );
 a56080a <=( A167  and  (not A168) );
 a56081a <=( (not A169)  and  a56080a );
 a56084a <=( A199  and  A166 );
 a56087a <=( A203  and  (not A200) );
 a56088a <=( a56087a  and  a56084a );
 a56089a <=( a56088a  and  a56081a );
 a56092a <=( (not A233)  and  (not A232) );
 a56095a <=( A265  and  (not A235) );
 a56096a <=( a56095a  and  a56092a );
 a56099a <=( (not A267)  and  A266 );
 a56102a <=( A301  and  (not A268) );
 a56103a <=( a56102a  and  a56099a );
 a56104a <=( a56103a  and  a56096a );
 a56108a <=( A167  and  (not A168) );
 a56109a <=( (not A169)  and  a56108a );
 a56112a <=( A199  and  A166 );
 a56115a <=( A203  and  (not A200) );
 a56116a <=( a56115a  and  a56112a );
 a56117a <=( a56116a  and  a56109a );
 a56120a <=( (not A233)  and  (not A232) );
 a56123a <=( (not A265)  and  (not A235) );
 a56124a <=( a56123a  and  a56120a );
 a56127a <=( (not A268)  and  (not A266) );
 a56130a <=( A300  and  A299 );
 a56131a <=( a56130a  and  a56127a );
 a56132a <=( a56131a  and  a56124a );
 a56136a <=( A167  and  (not A168) );
 a56137a <=( (not A169)  and  a56136a );
 a56140a <=( A199  and  A166 );
 a56143a <=( A203  and  (not A200) );
 a56144a <=( a56143a  and  a56140a );
 a56145a <=( a56144a  and  a56137a );
 a56148a <=( (not A233)  and  (not A232) );
 a56151a <=( (not A265)  and  (not A235) );
 a56152a <=( a56151a  and  a56148a );
 a56155a <=( (not A268)  and  (not A266) );
 a56158a <=( A300  and  A298 );
 a56159a <=( a56158a  and  a56155a );
 a56160a <=( a56159a  and  a56152a );
 a56164a <=( (not A168)  and  (not A169) );
 a56165a <=( (not A170)  and  a56164a );
 a56168a <=( A232  and  A202 );
 a56171a <=( (not A234)  and  A233 );
 a56172a <=( a56171a  and  a56168a );
 a56173a <=( a56172a  and  a56165a );
 a56176a <=( A265  and  (not A235) );
 a56179a <=( (not A267)  and  A266 );
 a56180a <=( a56179a  and  a56176a );
 a56183a <=( A298  and  (not A268) );
 a56186a <=( A302  and  (not A299) );
 a56187a <=( a56186a  and  a56183a );
 a56188a <=( a56187a  and  a56180a );
 a56192a <=( (not A168)  and  (not A169) );
 a56193a <=( (not A170)  and  a56192a );
 a56196a <=( A232  and  A202 );
 a56199a <=( (not A234)  and  A233 );
 a56200a <=( a56199a  and  a56196a );
 a56201a <=( a56200a  and  a56193a );
 a56204a <=( A265  and  (not A235) );
 a56207a <=( (not A267)  and  A266 );
 a56208a <=( a56207a  and  a56204a );
 a56211a <=( (not A298)  and  (not A268) );
 a56214a <=( A302  and  A299 );
 a56215a <=( a56214a  and  a56211a );
 a56216a <=( a56215a  and  a56208a );
 a56220a <=( (not A168)  and  (not A169) );
 a56221a <=( (not A170)  and  a56220a );
 a56224a <=( A201  and  A199 );
 a56227a <=( (not A235)  and  (not A234) );
 a56228a <=( a56227a  and  a56224a );
 a56229a <=( a56228a  and  a56221a );
 a56232a <=( A265  and  (not A236) );
 a56235a <=( (not A267)  and  A266 );
 a56236a <=( a56235a  and  a56232a );
 a56239a <=( A298  and  (not A268) );
 a56242a <=( A302  and  (not A299) );
 a56243a <=( a56242a  and  a56239a );
 a56244a <=( a56243a  and  a56236a );
 a56248a <=( (not A168)  and  (not A169) );
 a56249a <=( (not A170)  and  a56248a );
 a56252a <=( A201  and  A199 );
 a56255a <=( (not A235)  and  (not A234) );
 a56256a <=( a56255a  and  a56252a );
 a56257a <=( a56256a  and  a56249a );
 a56260a <=( A265  and  (not A236) );
 a56263a <=( (not A267)  and  A266 );
 a56264a <=( a56263a  and  a56260a );
 a56267a <=( (not A298)  and  (not A268) );
 a56270a <=( A302  and  A299 );
 a56271a <=( a56270a  and  a56267a );
 a56272a <=( a56271a  and  a56264a );
 a56276a <=( (not A168)  and  (not A169) );
 a56277a <=( (not A170)  and  a56276a );
 a56280a <=( A201  and  A199 );
 a56283a <=( A233  and  A232 );
 a56284a <=( a56283a  and  a56280a );
 a56285a <=( a56284a  and  a56277a );
 a56288a <=( (not A235)  and  (not A234) );
 a56291a <=( (not A268)  and  (not A267) );
 a56292a <=( a56291a  and  a56288a );
 a56295a <=( A298  and  (not A269) );
 a56298a <=( A302  and  (not A299) );
 a56299a <=( a56298a  and  a56295a );
 a56300a <=( a56299a  and  a56292a );
 a56304a <=( (not A168)  and  (not A169) );
 a56305a <=( (not A170)  and  a56304a );
 a56308a <=( A201  and  A199 );
 a56311a <=( A233  and  A232 );
 a56312a <=( a56311a  and  a56308a );
 a56313a <=( a56312a  and  a56305a );
 a56316a <=( (not A235)  and  (not A234) );
 a56319a <=( (not A268)  and  (not A267) );
 a56320a <=( a56319a  and  a56316a );
 a56323a <=( (not A298)  and  (not A269) );
 a56326a <=( A302  and  A299 );
 a56327a <=( a56326a  and  a56323a );
 a56328a <=( a56327a  and  a56320a );
 a56332a <=( (not A168)  and  (not A169) );
 a56333a <=( (not A170)  and  a56332a );
 a56336a <=( A201  and  A199 );
 a56339a <=( A233  and  A232 );
 a56340a <=( a56339a  and  a56336a );
 a56341a <=( a56340a  and  a56333a );
 a56344a <=( (not A235)  and  (not A234) );
 a56347a <=( A266  and  A265 );
 a56348a <=( a56347a  and  a56344a );
 a56351a <=( (not A268)  and  (not A267) );
 a56354a <=( A300  and  A299 );
 a56355a <=( a56354a  and  a56351a );
 a56356a <=( a56355a  and  a56348a );
 a56360a <=( (not A168)  and  (not A169) );
 a56361a <=( (not A170)  and  a56360a );
 a56364a <=( A201  and  A199 );
 a56367a <=( A233  and  A232 );
 a56368a <=( a56367a  and  a56364a );
 a56369a <=( a56368a  and  a56361a );
 a56372a <=( (not A235)  and  (not A234) );
 a56375a <=( A266  and  A265 );
 a56376a <=( a56375a  and  a56372a );
 a56379a <=( (not A268)  and  (not A267) );
 a56382a <=( A300  and  A298 );
 a56383a <=( a56382a  and  a56379a );
 a56384a <=( a56383a  and  a56376a );
 a56388a <=( (not A168)  and  (not A169) );
 a56389a <=( (not A170)  and  a56388a );
 a56392a <=( A201  and  A199 );
 a56395a <=( A233  and  A232 );
 a56396a <=( a56395a  and  a56392a );
 a56397a <=( a56396a  and  a56389a );
 a56400a <=( (not A235)  and  (not A234) );
 a56403a <=( (not A266)  and  (not A265) );
 a56404a <=( a56403a  and  a56400a );
 a56407a <=( A298  and  (not A268) );
 a56410a <=( A302  and  (not A299) );
 a56411a <=( a56410a  and  a56407a );
 a56412a <=( a56411a  and  a56404a );
 a56416a <=( (not A168)  and  (not A169) );
 a56417a <=( (not A170)  and  a56416a );
 a56420a <=( A201  and  A199 );
 a56423a <=( A233  and  A232 );
 a56424a <=( a56423a  and  a56420a );
 a56425a <=( a56424a  and  a56417a );
 a56428a <=( (not A235)  and  (not A234) );
 a56431a <=( (not A266)  and  (not A265) );
 a56432a <=( a56431a  and  a56428a );
 a56435a <=( (not A298)  and  (not A268) );
 a56438a <=( A302  and  A299 );
 a56439a <=( a56438a  and  a56435a );
 a56440a <=( a56439a  and  a56432a );
 a56444a <=( (not A168)  and  (not A169) );
 a56445a <=( (not A170)  and  a56444a );
 a56448a <=( A201  and  A199 );
 a56451a <=( (not A233)  and  (not A232) );
 a56452a <=( a56451a  and  a56448a );
 a56453a <=( a56452a  and  a56445a );
 a56456a <=( A265  and  (not A235) );
 a56459a <=( (not A267)  and  A266 );
 a56460a <=( a56459a  and  a56456a );
 a56463a <=( A298  and  (not A268) );
 a56466a <=( A302  and  (not A299) );
 a56467a <=( a56466a  and  a56463a );
 a56468a <=( a56467a  and  a56460a );
 a56472a <=( (not A168)  and  (not A169) );
 a56473a <=( (not A170)  and  a56472a );
 a56476a <=( A201  and  A199 );
 a56479a <=( (not A233)  and  (not A232) );
 a56480a <=( a56479a  and  a56476a );
 a56481a <=( a56480a  and  a56473a );
 a56484a <=( A265  and  (not A235) );
 a56487a <=( (not A267)  and  A266 );
 a56488a <=( a56487a  and  a56484a );
 a56491a <=( (not A298)  and  (not A268) );
 a56494a <=( A302  and  A299 );
 a56495a <=( a56494a  and  a56491a );
 a56496a <=( a56495a  and  a56488a );
 a56500a <=( (not A168)  and  (not A169) );
 a56501a <=( (not A170)  and  a56500a );
 a56504a <=( A201  and  A200 );
 a56507a <=( (not A235)  and  (not A234) );
 a56508a <=( a56507a  and  a56504a );
 a56509a <=( a56508a  and  a56501a );
 a56512a <=( A265  and  (not A236) );
 a56515a <=( (not A267)  and  A266 );
 a56516a <=( a56515a  and  a56512a );
 a56519a <=( A298  and  (not A268) );
 a56522a <=( A302  and  (not A299) );
 a56523a <=( a56522a  and  a56519a );
 a56524a <=( a56523a  and  a56516a );
 a56528a <=( (not A168)  and  (not A169) );
 a56529a <=( (not A170)  and  a56528a );
 a56532a <=( A201  and  A200 );
 a56535a <=( (not A235)  and  (not A234) );
 a56536a <=( a56535a  and  a56532a );
 a56537a <=( a56536a  and  a56529a );
 a56540a <=( A265  and  (not A236) );
 a56543a <=( (not A267)  and  A266 );
 a56544a <=( a56543a  and  a56540a );
 a56547a <=( (not A298)  and  (not A268) );
 a56550a <=( A302  and  A299 );
 a56551a <=( a56550a  and  a56547a );
 a56552a <=( a56551a  and  a56544a );
 a56556a <=( (not A168)  and  (not A169) );
 a56557a <=( (not A170)  and  a56556a );
 a56560a <=( A201  and  A200 );
 a56563a <=( A233  and  A232 );
 a56564a <=( a56563a  and  a56560a );
 a56565a <=( a56564a  and  a56557a );
 a56568a <=( (not A235)  and  (not A234) );
 a56571a <=( (not A268)  and  (not A267) );
 a56572a <=( a56571a  and  a56568a );
 a56575a <=( A298  and  (not A269) );
 a56578a <=( A302  and  (not A299) );
 a56579a <=( a56578a  and  a56575a );
 a56580a <=( a56579a  and  a56572a );
 a56584a <=( (not A168)  and  (not A169) );
 a56585a <=( (not A170)  and  a56584a );
 a56588a <=( A201  and  A200 );
 a56591a <=( A233  and  A232 );
 a56592a <=( a56591a  and  a56588a );
 a56593a <=( a56592a  and  a56585a );
 a56596a <=( (not A235)  and  (not A234) );
 a56599a <=( (not A268)  and  (not A267) );
 a56600a <=( a56599a  and  a56596a );
 a56603a <=( (not A298)  and  (not A269) );
 a56606a <=( A302  and  A299 );
 a56607a <=( a56606a  and  a56603a );
 a56608a <=( a56607a  and  a56600a );
 a56612a <=( (not A168)  and  (not A169) );
 a56613a <=( (not A170)  and  a56612a );
 a56616a <=( A201  and  A200 );
 a56619a <=( A233  and  A232 );
 a56620a <=( a56619a  and  a56616a );
 a56621a <=( a56620a  and  a56613a );
 a56624a <=( (not A235)  and  (not A234) );
 a56627a <=( A266  and  A265 );
 a56628a <=( a56627a  and  a56624a );
 a56631a <=( (not A268)  and  (not A267) );
 a56634a <=( A300  and  A299 );
 a56635a <=( a56634a  and  a56631a );
 a56636a <=( a56635a  and  a56628a );
 a56640a <=( (not A168)  and  (not A169) );
 a56641a <=( (not A170)  and  a56640a );
 a56644a <=( A201  and  A200 );
 a56647a <=( A233  and  A232 );
 a56648a <=( a56647a  and  a56644a );
 a56649a <=( a56648a  and  a56641a );
 a56652a <=( (not A235)  and  (not A234) );
 a56655a <=( A266  and  A265 );
 a56656a <=( a56655a  and  a56652a );
 a56659a <=( (not A268)  and  (not A267) );
 a56662a <=( A300  and  A298 );
 a56663a <=( a56662a  and  a56659a );
 a56664a <=( a56663a  and  a56656a );
 a56668a <=( (not A168)  and  (not A169) );
 a56669a <=( (not A170)  and  a56668a );
 a56672a <=( A201  and  A200 );
 a56675a <=( A233  and  A232 );
 a56676a <=( a56675a  and  a56672a );
 a56677a <=( a56676a  and  a56669a );
 a56680a <=( (not A235)  and  (not A234) );
 a56683a <=( (not A266)  and  (not A265) );
 a56684a <=( a56683a  and  a56680a );
 a56687a <=( A298  and  (not A268) );
 a56690a <=( A302  and  (not A299) );
 a56691a <=( a56690a  and  a56687a );
 a56692a <=( a56691a  and  a56684a );
 a56696a <=( (not A168)  and  (not A169) );
 a56697a <=( (not A170)  and  a56696a );
 a56700a <=( A201  and  A200 );
 a56703a <=( A233  and  A232 );
 a56704a <=( a56703a  and  a56700a );
 a56705a <=( a56704a  and  a56697a );
 a56708a <=( (not A235)  and  (not A234) );
 a56711a <=( (not A266)  and  (not A265) );
 a56712a <=( a56711a  and  a56708a );
 a56715a <=( (not A298)  and  (not A268) );
 a56718a <=( A302  and  A299 );
 a56719a <=( a56718a  and  a56715a );
 a56720a <=( a56719a  and  a56712a );
 a56724a <=( (not A168)  and  (not A169) );
 a56725a <=( (not A170)  and  a56724a );
 a56728a <=( A201  and  A200 );
 a56731a <=( (not A233)  and  (not A232) );
 a56732a <=( a56731a  and  a56728a );
 a56733a <=( a56732a  and  a56725a );
 a56736a <=( A265  and  (not A235) );
 a56739a <=( (not A267)  and  A266 );
 a56740a <=( a56739a  and  a56736a );
 a56743a <=( A298  and  (not A268) );
 a56746a <=( A302  and  (not A299) );
 a56747a <=( a56746a  and  a56743a );
 a56748a <=( a56747a  and  a56740a );
 a56752a <=( (not A168)  and  (not A169) );
 a56753a <=( (not A170)  and  a56752a );
 a56756a <=( A201  and  A200 );
 a56759a <=( (not A233)  and  (not A232) );
 a56760a <=( a56759a  and  a56756a );
 a56761a <=( a56760a  and  a56753a );
 a56764a <=( A265  and  (not A235) );
 a56767a <=( (not A267)  and  A266 );
 a56768a <=( a56767a  and  a56764a );
 a56771a <=( (not A298)  and  (not A268) );
 a56774a <=( A302  and  A299 );
 a56775a <=( a56774a  and  a56771a );
 a56776a <=( a56775a  and  a56768a );
 a56780a <=( (not A168)  and  (not A169) );
 a56781a <=( (not A170)  and  a56780a );
 a56784a <=( A200  and  (not A199) );
 a56787a <=( (not A234)  and  A203 );
 a56788a <=( a56787a  and  a56784a );
 a56789a <=( a56788a  and  a56781a );
 a56792a <=( (not A236)  and  (not A235) );
 a56795a <=( (not A268)  and  (not A267) );
 a56796a <=( a56795a  and  a56792a );
 a56799a <=( A298  and  (not A269) );
 a56802a <=( A302  and  (not A299) );
 a56803a <=( a56802a  and  a56799a );
 a56804a <=( a56803a  and  a56796a );
 a56808a <=( (not A168)  and  (not A169) );
 a56809a <=( (not A170)  and  a56808a );
 a56812a <=( A200  and  (not A199) );
 a56815a <=( (not A234)  and  A203 );
 a56816a <=( a56815a  and  a56812a );
 a56817a <=( a56816a  and  a56809a );
 a56820a <=( (not A236)  and  (not A235) );
 a56823a <=( (not A268)  and  (not A267) );
 a56824a <=( a56823a  and  a56820a );
 a56827a <=( (not A298)  and  (not A269) );
 a56830a <=( A302  and  A299 );
 a56831a <=( a56830a  and  a56827a );
 a56832a <=( a56831a  and  a56824a );
 a56836a <=( (not A168)  and  (not A169) );
 a56837a <=( (not A170)  and  a56836a );
 a56840a <=( A200  and  (not A199) );
 a56843a <=( (not A234)  and  A203 );
 a56844a <=( a56843a  and  a56840a );
 a56845a <=( a56844a  and  a56837a );
 a56848a <=( (not A236)  and  (not A235) );
 a56851a <=( A266  and  A265 );
 a56852a <=( a56851a  and  a56848a );
 a56855a <=( (not A268)  and  (not A267) );
 a56858a <=( A300  and  A299 );
 a56859a <=( a56858a  and  a56855a );
 a56860a <=( a56859a  and  a56852a );
 a56864a <=( (not A168)  and  (not A169) );
 a56865a <=( (not A170)  and  a56864a );
 a56868a <=( A200  and  (not A199) );
 a56871a <=( (not A234)  and  A203 );
 a56872a <=( a56871a  and  a56868a );
 a56873a <=( a56872a  and  a56865a );
 a56876a <=( (not A236)  and  (not A235) );
 a56879a <=( A266  and  A265 );
 a56880a <=( a56879a  and  a56876a );
 a56883a <=( (not A268)  and  (not A267) );
 a56886a <=( A300  and  A298 );
 a56887a <=( a56886a  and  a56883a );
 a56888a <=( a56887a  and  a56880a );
 a56892a <=( (not A168)  and  (not A169) );
 a56893a <=( (not A170)  and  a56892a );
 a56896a <=( A200  and  (not A199) );
 a56899a <=( (not A234)  and  A203 );
 a56900a <=( a56899a  and  a56896a );
 a56901a <=( a56900a  and  a56893a );
 a56904a <=( (not A236)  and  (not A235) );
 a56907a <=( (not A266)  and  (not A265) );
 a56908a <=( a56907a  and  a56904a );
 a56911a <=( A298  and  (not A268) );
 a56914a <=( A302  and  (not A299) );
 a56915a <=( a56914a  and  a56911a );
 a56916a <=( a56915a  and  a56908a );
 a56920a <=( (not A168)  and  (not A169) );
 a56921a <=( (not A170)  and  a56920a );
 a56924a <=( A200  and  (not A199) );
 a56927a <=( (not A234)  and  A203 );
 a56928a <=( a56927a  and  a56924a );
 a56929a <=( a56928a  and  a56921a );
 a56932a <=( (not A236)  and  (not A235) );
 a56935a <=( (not A266)  and  (not A265) );
 a56936a <=( a56935a  and  a56932a );
 a56939a <=( (not A298)  and  (not A268) );
 a56942a <=( A302  and  A299 );
 a56943a <=( a56942a  and  a56939a );
 a56944a <=( a56943a  and  a56936a );
 a56948a <=( (not A168)  and  (not A169) );
 a56949a <=( (not A170)  and  a56948a );
 a56952a <=( A200  and  (not A199) );
 a56955a <=( A232  and  A203 );
 a56956a <=( a56955a  and  a56952a );
 a56957a <=( a56956a  and  a56949a );
 a56960a <=( (not A234)  and  A233 );
 a56963a <=( (not A267)  and  (not A235) );
 a56964a <=( a56963a  and  a56960a );
 a56967a <=( (not A269)  and  (not A268) );
 a56970a <=( A300  and  A299 );
 a56971a <=( a56970a  and  a56967a );
 a56972a <=( a56971a  and  a56964a );
 a56976a <=( (not A168)  and  (not A169) );
 a56977a <=( (not A170)  and  a56976a );
 a56980a <=( A200  and  (not A199) );
 a56983a <=( A232  and  A203 );
 a56984a <=( a56983a  and  a56980a );
 a56985a <=( a56984a  and  a56977a );
 a56988a <=( (not A234)  and  A233 );
 a56991a <=( (not A267)  and  (not A235) );
 a56992a <=( a56991a  and  a56988a );
 a56995a <=( (not A269)  and  (not A268) );
 a56998a <=( A300  and  A298 );
 a56999a <=( a56998a  and  a56995a );
 a57000a <=( a56999a  and  a56992a );
 a57004a <=( (not A168)  and  (not A169) );
 a57005a <=( (not A170)  and  a57004a );
 a57008a <=( A200  and  (not A199) );
 a57011a <=( A232  and  A203 );
 a57012a <=( a57011a  and  a57008a );
 a57013a <=( a57012a  and  a57005a );
 a57016a <=( (not A234)  and  A233 );
 a57019a <=( A265  and  (not A235) );
 a57020a <=( a57019a  and  a57016a );
 a57023a <=( (not A267)  and  A266 );
 a57026a <=( A301  and  (not A268) );
 a57027a <=( a57026a  and  a57023a );
 a57028a <=( a57027a  and  a57020a );
 a57032a <=( (not A168)  and  (not A169) );
 a57033a <=( (not A170)  and  a57032a );
 a57036a <=( A200  and  (not A199) );
 a57039a <=( A232  and  A203 );
 a57040a <=( a57039a  and  a57036a );
 a57041a <=( a57040a  and  a57033a );
 a57044a <=( (not A234)  and  A233 );
 a57047a <=( (not A265)  and  (not A235) );
 a57048a <=( a57047a  and  a57044a );
 a57051a <=( (not A268)  and  (not A266) );
 a57054a <=( A300  and  A299 );
 a57055a <=( a57054a  and  a57051a );
 a57056a <=( a57055a  and  a57048a );
 a57060a <=( (not A168)  and  (not A169) );
 a57061a <=( (not A170)  and  a57060a );
 a57064a <=( A200  and  (not A199) );
 a57067a <=( A232  and  A203 );
 a57068a <=( a57067a  and  a57064a );
 a57069a <=( a57068a  and  a57061a );
 a57072a <=( (not A234)  and  A233 );
 a57075a <=( (not A265)  and  (not A235) );
 a57076a <=( a57075a  and  a57072a );
 a57079a <=( (not A268)  and  (not A266) );
 a57082a <=( A300  and  A298 );
 a57083a <=( a57082a  and  a57079a );
 a57084a <=( a57083a  and  a57076a );
 a57088a <=( (not A168)  and  (not A169) );
 a57089a <=( (not A170)  and  a57088a );
 a57092a <=( A200  and  (not A199) );
 a57095a <=( (not A232)  and  A203 );
 a57096a <=( a57095a  and  a57092a );
 a57097a <=( a57096a  and  a57089a );
 a57100a <=( (not A235)  and  (not A233) );
 a57103a <=( (not A268)  and  (not A267) );
 a57104a <=( a57103a  and  a57100a );
 a57107a <=( A298  and  (not A269) );
 a57110a <=( A302  and  (not A299) );
 a57111a <=( a57110a  and  a57107a );
 a57112a <=( a57111a  and  a57104a );
 a57116a <=( (not A168)  and  (not A169) );
 a57117a <=( (not A170)  and  a57116a );
 a57120a <=( A200  and  (not A199) );
 a57123a <=( (not A232)  and  A203 );
 a57124a <=( a57123a  and  a57120a );
 a57125a <=( a57124a  and  a57117a );
 a57128a <=( (not A235)  and  (not A233) );
 a57131a <=( (not A268)  and  (not A267) );
 a57132a <=( a57131a  and  a57128a );
 a57135a <=( (not A298)  and  (not A269) );
 a57138a <=( A302  and  A299 );
 a57139a <=( a57138a  and  a57135a );
 a57140a <=( a57139a  and  a57132a );
 a57144a <=( (not A168)  and  (not A169) );
 a57145a <=( (not A170)  and  a57144a );
 a57148a <=( A200  and  (not A199) );
 a57151a <=( (not A232)  and  A203 );
 a57152a <=( a57151a  and  a57148a );
 a57153a <=( a57152a  and  a57145a );
 a57156a <=( (not A235)  and  (not A233) );
 a57159a <=( A266  and  A265 );
 a57160a <=( a57159a  and  a57156a );
 a57163a <=( (not A268)  and  (not A267) );
 a57166a <=( A300  and  A299 );
 a57167a <=( a57166a  and  a57163a );
 a57168a <=( a57167a  and  a57160a );
 a57172a <=( (not A168)  and  (not A169) );
 a57173a <=( (not A170)  and  a57172a );
 a57176a <=( A200  and  (not A199) );
 a57179a <=( (not A232)  and  A203 );
 a57180a <=( a57179a  and  a57176a );
 a57181a <=( a57180a  and  a57173a );
 a57184a <=( (not A235)  and  (not A233) );
 a57187a <=( A266  and  A265 );
 a57188a <=( a57187a  and  a57184a );
 a57191a <=( (not A268)  and  (not A267) );
 a57194a <=( A300  and  A298 );
 a57195a <=( a57194a  and  a57191a );
 a57196a <=( a57195a  and  a57188a );
 a57200a <=( (not A168)  and  (not A169) );
 a57201a <=( (not A170)  and  a57200a );
 a57204a <=( A200  and  (not A199) );
 a57207a <=( (not A232)  and  A203 );
 a57208a <=( a57207a  and  a57204a );
 a57209a <=( a57208a  and  a57201a );
 a57212a <=( (not A235)  and  (not A233) );
 a57215a <=( (not A266)  and  (not A265) );
 a57216a <=( a57215a  and  a57212a );
 a57219a <=( A298  and  (not A268) );
 a57222a <=( A302  and  (not A299) );
 a57223a <=( a57222a  and  a57219a );
 a57224a <=( a57223a  and  a57216a );
 a57228a <=( (not A168)  and  (not A169) );
 a57229a <=( (not A170)  and  a57228a );
 a57232a <=( A200  and  (not A199) );
 a57235a <=( (not A232)  and  A203 );
 a57236a <=( a57235a  and  a57232a );
 a57237a <=( a57236a  and  a57229a );
 a57240a <=( (not A235)  and  (not A233) );
 a57243a <=( (not A266)  and  (not A265) );
 a57244a <=( a57243a  and  a57240a );
 a57247a <=( (not A298)  and  (not A268) );
 a57250a <=( A302  and  A299 );
 a57251a <=( a57250a  and  a57247a );
 a57252a <=( a57251a  and  a57244a );
 a57256a <=( (not A168)  and  (not A169) );
 a57257a <=( (not A170)  and  a57256a );
 a57260a <=( (not A200)  and  A199 );
 a57263a <=( (not A234)  and  A203 );
 a57264a <=( a57263a  and  a57260a );
 a57265a <=( a57264a  and  a57257a );
 a57268a <=( (not A236)  and  (not A235) );
 a57271a <=( (not A268)  and  (not A267) );
 a57272a <=( a57271a  and  a57268a );
 a57275a <=( A298  and  (not A269) );
 a57278a <=( A302  and  (not A299) );
 a57279a <=( a57278a  and  a57275a );
 a57280a <=( a57279a  and  a57272a );
 a57284a <=( (not A168)  and  (not A169) );
 a57285a <=( (not A170)  and  a57284a );
 a57288a <=( (not A200)  and  A199 );
 a57291a <=( (not A234)  and  A203 );
 a57292a <=( a57291a  and  a57288a );
 a57293a <=( a57292a  and  a57285a );
 a57296a <=( (not A236)  and  (not A235) );
 a57299a <=( (not A268)  and  (not A267) );
 a57300a <=( a57299a  and  a57296a );
 a57303a <=( (not A298)  and  (not A269) );
 a57306a <=( A302  and  A299 );
 a57307a <=( a57306a  and  a57303a );
 a57308a <=( a57307a  and  a57300a );
 a57312a <=( (not A168)  and  (not A169) );
 a57313a <=( (not A170)  and  a57312a );
 a57316a <=( (not A200)  and  A199 );
 a57319a <=( (not A234)  and  A203 );
 a57320a <=( a57319a  and  a57316a );
 a57321a <=( a57320a  and  a57313a );
 a57324a <=( (not A236)  and  (not A235) );
 a57327a <=( A266  and  A265 );
 a57328a <=( a57327a  and  a57324a );
 a57331a <=( (not A268)  and  (not A267) );
 a57334a <=( A300  and  A299 );
 a57335a <=( a57334a  and  a57331a );
 a57336a <=( a57335a  and  a57328a );
 a57340a <=( (not A168)  and  (not A169) );
 a57341a <=( (not A170)  and  a57340a );
 a57344a <=( (not A200)  and  A199 );
 a57347a <=( (not A234)  and  A203 );
 a57348a <=( a57347a  and  a57344a );
 a57349a <=( a57348a  and  a57341a );
 a57352a <=( (not A236)  and  (not A235) );
 a57355a <=( A266  and  A265 );
 a57356a <=( a57355a  and  a57352a );
 a57359a <=( (not A268)  and  (not A267) );
 a57362a <=( A300  and  A298 );
 a57363a <=( a57362a  and  a57359a );
 a57364a <=( a57363a  and  a57356a );
 a57368a <=( (not A168)  and  (not A169) );
 a57369a <=( (not A170)  and  a57368a );
 a57372a <=( (not A200)  and  A199 );
 a57375a <=( (not A234)  and  A203 );
 a57376a <=( a57375a  and  a57372a );
 a57377a <=( a57376a  and  a57369a );
 a57380a <=( (not A236)  and  (not A235) );
 a57383a <=( (not A266)  and  (not A265) );
 a57384a <=( a57383a  and  a57380a );
 a57387a <=( A298  and  (not A268) );
 a57390a <=( A302  and  (not A299) );
 a57391a <=( a57390a  and  a57387a );
 a57392a <=( a57391a  and  a57384a );
 a57396a <=( (not A168)  and  (not A169) );
 a57397a <=( (not A170)  and  a57396a );
 a57400a <=( (not A200)  and  A199 );
 a57403a <=( (not A234)  and  A203 );
 a57404a <=( a57403a  and  a57400a );
 a57405a <=( a57404a  and  a57397a );
 a57408a <=( (not A236)  and  (not A235) );
 a57411a <=( (not A266)  and  (not A265) );
 a57412a <=( a57411a  and  a57408a );
 a57415a <=( (not A298)  and  (not A268) );
 a57418a <=( A302  and  A299 );
 a57419a <=( a57418a  and  a57415a );
 a57420a <=( a57419a  and  a57412a );
 a57424a <=( (not A168)  and  (not A169) );
 a57425a <=( (not A170)  and  a57424a );
 a57428a <=( (not A200)  and  A199 );
 a57431a <=( A232  and  A203 );
 a57432a <=( a57431a  and  a57428a );
 a57433a <=( a57432a  and  a57425a );
 a57436a <=( (not A234)  and  A233 );
 a57439a <=( (not A267)  and  (not A235) );
 a57440a <=( a57439a  and  a57436a );
 a57443a <=( (not A269)  and  (not A268) );
 a57446a <=( A300  and  A299 );
 a57447a <=( a57446a  and  a57443a );
 a57448a <=( a57447a  and  a57440a );
 a57452a <=( (not A168)  and  (not A169) );
 a57453a <=( (not A170)  and  a57452a );
 a57456a <=( (not A200)  and  A199 );
 a57459a <=( A232  and  A203 );
 a57460a <=( a57459a  and  a57456a );
 a57461a <=( a57460a  and  a57453a );
 a57464a <=( (not A234)  and  A233 );
 a57467a <=( (not A267)  and  (not A235) );
 a57468a <=( a57467a  and  a57464a );
 a57471a <=( (not A269)  and  (not A268) );
 a57474a <=( A300  and  A298 );
 a57475a <=( a57474a  and  a57471a );
 a57476a <=( a57475a  and  a57468a );
 a57480a <=( (not A168)  and  (not A169) );
 a57481a <=( (not A170)  and  a57480a );
 a57484a <=( (not A200)  and  A199 );
 a57487a <=( A232  and  A203 );
 a57488a <=( a57487a  and  a57484a );
 a57489a <=( a57488a  and  a57481a );
 a57492a <=( (not A234)  and  A233 );
 a57495a <=( A265  and  (not A235) );
 a57496a <=( a57495a  and  a57492a );
 a57499a <=( (not A267)  and  A266 );
 a57502a <=( A301  and  (not A268) );
 a57503a <=( a57502a  and  a57499a );
 a57504a <=( a57503a  and  a57496a );
 a57508a <=( (not A168)  and  (not A169) );
 a57509a <=( (not A170)  and  a57508a );
 a57512a <=( (not A200)  and  A199 );
 a57515a <=( A232  and  A203 );
 a57516a <=( a57515a  and  a57512a );
 a57517a <=( a57516a  and  a57509a );
 a57520a <=( (not A234)  and  A233 );
 a57523a <=( (not A265)  and  (not A235) );
 a57524a <=( a57523a  and  a57520a );
 a57527a <=( (not A268)  and  (not A266) );
 a57530a <=( A300  and  A299 );
 a57531a <=( a57530a  and  a57527a );
 a57532a <=( a57531a  and  a57524a );
 a57536a <=( (not A168)  and  (not A169) );
 a57537a <=( (not A170)  and  a57536a );
 a57540a <=( (not A200)  and  A199 );
 a57543a <=( A232  and  A203 );
 a57544a <=( a57543a  and  a57540a );
 a57545a <=( a57544a  and  a57537a );
 a57548a <=( (not A234)  and  A233 );
 a57551a <=( (not A265)  and  (not A235) );
 a57552a <=( a57551a  and  a57548a );
 a57555a <=( (not A268)  and  (not A266) );
 a57558a <=( A300  and  A298 );
 a57559a <=( a57558a  and  a57555a );
 a57560a <=( a57559a  and  a57552a );
 a57564a <=( (not A168)  and  (not A169) );
 a57565a <=( (not A170)  and  a57564a );
 a57568a <=( (not A200)  and  A199 );
 a57571a <=( (not A232)  and  A203 );
 a57572a <=( a57571a  and  a57568a );
 a57573a <=( a57572a  and  a57565a );
 a57576a <=( (not A235)  and  (not A233) );
 a57579a <=( (not A268)  and  (not A267) );
 a57580a <=( a57579a  and  a57576a );
 a57583a <=( A298  and  (not A269) );
 a57586a <=( A302  and  (not A299) );
 a57587a <=( a57586a  and  a57583a );
 a57588a <=( a57587a  and  a57580a );
 a57592a <=( (not A168)  and  (not A169) );
 a57593a <=( (not A170)  and  a57592a );
 a57596a <=( (not A200)  and  A199 );
 a57599a <=( (not A232)  and  A203 );
 a57600a <=( a57599a  and  a57596a );
 a57601a <=( a57600a  and  a57593a );
 a57604a <=( (not A235)  and  (not A233) );
 a57607a <=( (not A268)  and  (not A267) );
 a57608a <=( a57607a  and  a57604a );
 a57611a <=( (not A298)  and  (not A269) );
 a57614a <=( A302  and  A299 );
 a57615a <=( a57614a  and  a57611a );
 a57616a <=( a57615a  and  a57608a );
 a57620a <=( (not A168)  and  (not A169) );
 a57621a <=( (not A170)  and  a57620a );
 a57624a <=( (not A200)  and  A199 );
 a57627a <=( (not A232)  and  A203 );
 a57628a <=( a57627a  and  a57624a );
 a57629a <=( a57628a  and  a57621a );
 a57632a <=( (not A235)  and  (not A233) );
 a57635a <=( A266  and  A265 );
 a57636a <=( a57635a  and  a57632a );
 a57639a <=( (not A268)  and  (not A267) );
 a57642a <=( A300  and  A299 );
 a57643a <=( a57642a  and  a57639a );
 a57644a <=( a57643a  and  a57636a );
 a57648a <=( (not A168)  and  (not A169) );
 a57649a <=( (not A170)  and  a57648a );
 a57652a <=( (not A200)  and  A199 );
 a57655a <=( (not A232)  and  A203 );
 a57656a <=( a57655a  and  a57652a );
 a57657a <=( a57656a  and  a57649a );
 a57660a <=( (not A235)  and  (not A233) );
 a57663a <=( A266  and  A265 );
 a57664a <=( a57663a  and  a57660a );
 a57667a <=( (not A268)  and  (not A267) );
 a57670a <=( A300  and  A298 );
 a57671a <=( a57670a  and  a57667a );
 a57672a <=( a57671a  and  a57664a );
 a57676a <=( (not A168)  and  (not A169) );
 a57677a <=( (not A170)  and  a57676a );
 a57680a <=( (not A200)  and  A199 );
 a57683a <=( (not A232)  and  A203 );
 a57684a <=( a57683a  and  a57680a );
 a57685a <=( a57684a  and  a57677a );
 a57688a <=( (not A235)  and  (not A233) );
 a57691a <=( (not A266)  and  (not A265) );
 a57692a <=( a57691a  and  a57688a );
 a57695a <=( A298  and  (not A268) );
 a57698a <=( A302  and  (not A299) );
 a57699a <=( a57698a  and  a57695a );
 a57700a <=( a57699a  and  a57692a );
 a57704a <=( (not A168)  and  (not A169) );
 a57705a <=( (not A170)  and  a57704a );
 a57708a <=( (not A200)  and  A199 );
 a57711a <=( (not A232)  and  A203 );
 a57712a <=( a57711a  and  a57708a );
 a57713a <=( a57712a  and  a57705a );
 a57716a <=( (not A235)  and  (not A233) );
 a57719a <=( (not A266)  and  (not A265) );
 a57720a <=( a57719a  and  a57716a );
 a57723a <=( (not A298)  and  (not A268) );
 a57726a <=( A302  and  A299 );
 a57727a <=( a57726a  and  a57723a );
 a57728a <=( a57727a  and  a57720a );
 a57731a <=( A166  and  A168 );
 a57734a <=( (not A202)  and  (not A201) );
 a57735a <=( a57734a  and  a57731a );
 a57738a <=( A232  and  (not A203) );
 a57741a <=( (not A234)  and  A233 );
 a57742a <=( a57741a  and  a57738a );
 a57743a <=( a57742a  and  a57735a );
 a57746a <=( A265  and  (not A235) );
 a57749a <=( (not A267)  and  A266 );
 a57750a <=( a57749a  and  a57746a );
 a57753a <=( A298  and  (not A268) );
 a57756a <=( A302  and  (not A299) );
 a57757a <=( a57756a  and  a57753a );
 a57758a <=( a57757a  and  a57750a );
 a57761a <=( A166  and  A168 );
 a57764a <=( (not A202)  and  (not A201) );
 a57765a <=( a57764a  and  a57761a );
 a57768a <=( A232  and  (not A203) );
 a57771a <=( (not A234)  and  A233 );
 a57772a <=( a57771a  and  a57768a );
 a57773a <=( a57772a  and  a57765a );
 a57776a <=( A265  and  (not A235) );
 a57779a <=( (not A267)  and  A266 );
 a57780a <=( a57779a  and  a57776a );
 a57783a <=( (not A298)  and  (not A268) );
 a57786a <=( A302  and  A299 );
 a57787a <=( a57786a  and  a57783a );
 a57788a <=( a57787a  and  a57780a );
 a57791a <=( A166  and  A168 );
 a57794a <=( A200  and  A199 );
 a57795a <=( a57794a  and  a57791a );
 a57798a <=( (not A202)  and  (not A201) );
 a57801a <=( (not A235)  and  (not A234) );
 a57802a <=( a57801a  and  a57798a );
 a57803a <=( a57802a  and  a57795a );
 a57806a <=( A265  and  (not A236) );
 a57809a <=( (not A267)  and  A266 );
 a57810a <=( a57809a  and  a57806a );
 a57813a <=( A298  and  (not A268) );
 a57816a <=( A302  and  (not A299) );
 a57817a <=( a57816a  and  a57813a );
 a57818a <=( a57817a  and  a57810a );
 a57821a <=( A166  and  A168 );
 a57824a <=( A200  and  A199 );
 a57825a <=( a57824a  and  a57821a );
 a57828a <=( (not A202)  and  (not A201) );
 a57831a <=( (not A235)  and  (not A234) );
 a57832a <=( a57831a  and  a57828a );
 a57833a <=( a57832a  and  a57825a );
 a57836a <=( A265  and  (not A236) );
 a57839a <=( (not A267)  and  A266 );
 a57840a <=( a57839a  and  a57836a );
 a57843a <=( (not A298)  and  (not A268) );
 a57846a <=( A302  and  A299 );
 a57847a <=( a57846a  and  a57843a );
 a57848a <=( a57847a  and  a57840a );
 a57851a <=( A166  and  A168 );
 a57854a <=( A200  and  A199 );
 a57855a <=( a57854a  and  a57851a );
 a57858a <=( (not A202)  and  (not A201) );
 a57861a <=( A233  and  A232 );
 a57862a <=( a57861a  and  a57858a );
 a57863a <=( a57862a  and  a57855a );
 a57866a <=( (not A235)  and  (not A234) );
 a57869a <=( (not A268)  and  (not A267) );
 a57870a <=( a57869a  and  a57866a );
 a57873a <=( A298  and  (not A269) );
 a57876a <=( A302  and  (not A299) );
 a57877a <=( a57876a  and  a57873a );
 a57878a <=( a57877a  and  a57870a );
 a57881a <=( A166  and  A168 );
 a57884a <=( A200  and  A199 );
 a57885a <=( a57884a  and  a57881a );
 a57888a <=( (not A202)  and  (not A201) );
 a57891a <=( A233  and  A232 );
 a57892a <=( a57891a  and  a57888a );
 a57893a <=( a57892a  and  a57885a );
 a57896a <=( (not A235)  and  (not A234) );
 a57899a <=( (not A268)  and  (not A267) );
 a57900a <=( a57899a  and  a57896a );
 a57903a <=( (not A298)  and  (not A269) );
 a57906a <=( A302  and  A299 );
 a57907a <=( a57906a  and  a57903a );
 a57908a <=( a57907a  and  a57900a );
 a57911a <=( A166  and  A168 );
 a57914a <=( A200  and  A199 );
 a57915a <=( a57914a  and  a57911a );
 a57918a <=( (not A202)  and  (not A201) );
 a57921a <=( A233  and  A232 );
 a57922a <=( a57921a  and  a57918a );
 a57923a <=( a57922a  and  a57915a );
 a57926a <=( (not A235)  and  (not A234) );
 a57929a <=( A266  and  A265 );
 a57930a <=( a57929a  and  a57926a );
 a57933a <=( (not A268)  and  (not A267) );
 a57936a <=( A300  and  A299 );
 a57937a <=( a57936a  and  a57933a );
 a57938a <=( a57937a  and  a57930a );
 a57941a <=( A166  and  A168 );
 a57944a <=( A200  and  A199 );
 a57945a <=( a57944a  and  a57941a );
 a57948a <=( (not A202)  and  (not A201) );
 a57951a <=( A233  and  A232 );
 a57952a <=( a57951a  and  a57948a );
 a57953a <=( a57952a  and  a57945a );
 a57956a <=( (not A235)  and  (not A234) );
 a57959a <=( A266  and  A265 );
 a57960a <=( a57959a  and  a57956a );
 a57963a <=( (not A268)  and  (not A267) );
 a57966a <=( A300  and  A298 );
 a57967a <=( a57966a  and  a57963a );
 a57968a <=( a57967a  and  a57960a );
 a57971a <=( A166  and  A168 );
 a57974a <=( A200  and  A199 );
 a57975a <=( a57974a  and  a57971a );
 a57978a <=( (not A202)  and  (not A201) );
 a57981a <=( A233  and  A232 );
 a57982a <=( a57981a  and  a57978a );
 a57983a <=( a57982a  and  a57975a );
 a57986a <=( (not A235)  and  (not A234) );
 a57989a <=( (not A266)  and  (not A265) );
 a57990a <=( a57989a  and  a57986a );
 a57993a <=( A298  and  (not A268) );
 a57996a <=( A302  and  (not A299) );
 a57997a <=( a57996a  and  a57993a );
 a57998a <=( a57997a  and  a57990a );
 a58001a <=( A166  and  A168 );
 a58004a <=( A200  and  A199 );
 a58005a <=( a58004a  and  a58001a );
 a58008a <=( (not A202)  and  (not A201) );
 a58011a <=( A233  and  A232 );
 a58012a <=( a58011a  and  a58008a );
 a58013a <=( a58012a  and  a58005a );
 a58016a <=( (not A235)  and  (not A234) );
 a58019a <=( (not A266)  and  (not A265) );
 a58020a <=( a58019a  and  a58016a );
 a58023a <=( (not A298)  and  (not A268) );
 a58026a <=( A302  and  A299 );
 a58027a <=( a58026a  and  a58023a );
 a58028a <=( a58027a  and  a58020a );
 a58031a <=( A166  and  A168 );
 a58034a <=( A200  and  A199 );
 a58035a <=( a58034a  and  a58031a );
 a58038a <=( (not A202)  and  (not A201) );
 a58041a <=( (not A233)  and  (not A232) );
 a58042a <=( a58041a  and  a58038a );
 a58043a <=( a58042a  and  a58035a );
 a58046a <=( A265  and  (not A235) );
 a58049a <=( (not A267)  and  A266 );
 a58050a <=( a58049a  and  a58046a );
 a58053a <=( A298  and  (not A268) );
 a58056a <=( A302  and  (not A299) );
 a58057a <=( a58056a  and  a58053a );
 a58058a <=( a58057a  and  a58050a );
 a58061a <=( A166  and  A168 );
 a58064a <=( A200  and  A199 );
 a58065a <=( a58064a  and  a58061a );
 a58068a <=( (not A202)  and  (not A201) );
 a58071a <=( (not A233)  and  (not A232) );
 a58072a <=( a58071a  and  a58068a );
 a58073a <=( a58072a  and  a58065a );
 a58076a <=( A265  and  (not A235) );
 a58079a <=( (not A267)  and  A266 );
 a58080a <=( a58079a  and  a58076a );
 a58083a <=( (not A298)  and  (not A268) );
 a58086a <=( A302  and  A299 );
 a58087a <=( a58086a  and  a58083a );
 a58088a <=( a58087a  and  a58080a );
 a58091a <=( A166  and  A168 );
 a58094a <=( (not A200)  and  (not A199) );
 a58095a <=( a58094a  and  a58091a );
 a58098a <=( A232  and  (not A202) );
 a58101a <=( (not A234)  and  A233 );
 a58102a <=( a58101a  and  a58098a );
 a58103a <=( a58102a  and  a58095a );
 a58106a <=( A265  and  (not A235) );
 a58109a <=( (not A267)  and  A266 );
 a58110a <=( a58109a  and  a58106a );
 a58113a <=( A298  and  (not A268) );
 a58116a <=( A302  and  (not A299) );
 a58117a <=( a58116a  and  a58113a );
 a58118a <=( a58117a  and  a58110a );
 a58121a <=( A166  and  A168 );
 a58124a <=( (not A200)  and  (not A199) );
 a58125a <=( a58124a  and  a58121a );
 a58128a <=( A232  and  (not A202) );
 a58131a <=( (not A234)  and  A233 );
 a58132a <=( a58131a  and  a58128a );
 a58133a <=( a58132a  and  a58125a );
 a58136a <=( A265  and  (not A235) );
 a58139a <=( (not A267)  and  A266 );
 a58140a <=( a58139a  and  a58136a );
 a58143a <=( (not A298)  and  (not A268) );
 a58146a <=( A302  and  A299 );
 a58147a <=( a58146a  and  a58143a );
 a58148a <=( a58147a  and  a58140a );
 a58151a <=( A167  and  A168 );
 a58154a <=( (not A202)  and  (not A201) );
 a58155a <=( a58154a  and  a58151a );
 a58158a <=( A232  and  (not A203) );
 a58161a <=( (not A234)  and  A233 );
 a58162a <=( a58161a  and  a58158a );
 a58163a <=( a58162a  and  a58155a );
 a58166a <=( A265  and  (not A235) );
 a58169a <=( (not A267)  and  A266 );
 a58170a <=( a58169a  and  a58166a );
 a58173a <=( A298  and  (not A268) );
 a58176a <=( A302  and  (not A299) );
 a58177a <=( a58176a  and  a58173a );
 a58178a <=( a58177a  and  a58170a );
 a58181a <=( A167  and  A168 );
 a58184a <=( (not A202)  and  (not A201) );
 a58185a <=( a58184a  and  a58181a );
 a58188a <=( A232  and  (not A203) );
 a58191a <=( (not A234)  and  A233 );
 a58192a <=( a58191a  and  a58188a );
 a58193a <=( a58192a  and  a58185a );
 a58196a <=( A265  and  (not A235) );
 a58199a <=( (not A267)  and  A266 );
 a58200a <=( a58199a  and  a58196a );
 a58203a <=( (not A298)  and  (not A268) );
 a58206a <=( A302  and  A299 );
 a58207a <=( a58206a  and  a58203a );
 a58208a <=( a58207a  and  a58200a );
 a58211a <=( A167  and  A168 );
 a58214a <=( A200  and  A199 );
 a58215a <=( a58214a  and  a58211a );
 a58218a <=( (not A202)  and  (not A201) );
 a58221a <=( (not A235)  and  (not A234) );
 a58222a <=( a58221a  and  a58218a );
 a58223a <=( a58222a  and  a58215a );
 a58226a <=( A265  and  (not A236) );
 a58229a <=( (not A267)  and  A266 );
 a58230a <=( a58229a  and  a58226a );
 a58233a <=( A298  and  (not A268) );
 a58236a <=( A302  and  (not A299) );
 a58237a <=( a58236a  and  a58233a );
 a58238a <=( a58237a  and  a58230a );
 a58241a <=( A167  and  A168 );
 a58244a <=( A200  and  A199 );
 a58245a <=( a58244a  and  a58241a );
 a58248a <=( (not A202)  and  (not A201) );
 a58251a <=( (not A235)  and  (not A234) );
 a58252a <=( a58251a  and  a58248a );
 a58253a <=( a58252a  and  a58245a );
 a58256a <=( A265  and  (not A236) );
 a58259a <=( (not A267)  and  A266 );
 a58260a <=( a58259a  and  a58256a );
 a58263a <=( (not A298)  and  (not A268) );
 a58266a <=( A302  and  A299 );
 a58267a <=( a58266a  and  a58263a );
 a58268a <=( a58267a  and  a58260a );
 a58271a <=( A167  and  A168 );
 a58274a <=( A200  and  A199 );
 a58275a <=( a58274a  and  a58271a );
 a58278a <=( (not A202)  and  (not A201) );
 a58281a <=( A233  and  A232 );
 a58282a <=( a58281a  and  a58278a );
 a58283a <=( a58282a  and  a58275a );
 a58286a <=( (not A235)  and  (not A234) );
 a58289a <=( (not A268)  and  (not A267) );
 a58290a <=( a58289a  and  a58286a );
 a58293a <=( A298  and  (not A269) );
 a58296a <=( A302  and  (not A299) );
 a58297a <=( a58296a  and  a58293a );
 a58298a <=( a58297a  and  a58290a );
 a58301a <=( A167  and  A168 );
 a58304a <=( A200  and  A199 );
 a58305a <=( a58304a  and  a58301a );
 a58308a <=( (not A202)  and  (not A201) );
 a58311a <=( A233  and  A232 );
 a58312a <=( a58311a  and  a58308a );
 a58313a <=( a58312a  and  a58305a );
 a58316a <=( (not A235)  and  (not A234) );
 a58319a <=( (not A268)  and  (not A267) );
 a58320a <=( a58319a  and  a58316a );
 a58323a <=( (not A298)  and  (not A269) );
 a58326a <=( A302  and  A299 );
 a58327a <=( a58326a  and  a58323a );
 a58328a <=( a58327a  and  a58320a );
 a58331a <=( A167  and  A168 );
 a58334a <=( A200  and  A199 );
 a58335a <=( a58334a  and  a58331a );
 a58338a <=( (not A202)  and  (not A201) );
 a58341a <=( A233  and  A232 );
 a58342a <=( a58341a  and  a58338a );
 a58343a <=( a58342a  and  a58335a );
 a58346a <=( (not A235)  and  (not A234) );
 a58349a <=( A266  and  A265 );
 a58350a <=( a58349a  and  a58346a );
 a58353a <=( (not A268)  and  (not A267) );
 a58356a <=( A300  and  A299 );
 a58357a <=( a58356a  and  a58353a );
 a58358a <=( a58357a  and  a58350a );
 a58361a <=( A167  and  A168 );
 a58364a <=( A200  and  A199 );
 a58365a <=( a58364a  and  a58361a );
 a58368a <=( (not A202)  and  (not A201) );
 a58371a <=( A233  and  A232 );
 a58372a <=( a58371a  and  a58368a );
 a58373a <=( a58372a  and  a58365a );
 a58376a <=( (not A235)  and  (not A234) );
 a58379a <=( A266  and  A265 );
 a58380a <=( a58379a  and  a58376a );
 a58383a <=( (not A268)  and  (not A267) );
 a58386a <=( A300  and  A298 );
 a58387a <=( a58386a  and  a58383a );
 a58388a <=( a58387a  and  a58380a );
 a58391a <=( A167  and  A168 );
 a58394a <=( A200  and  A199 );
 a58395a <=( a58394a  and  a58391a );
 a58398a <=( (not A202)  and  (not A201) );
 a58401a <=( A233  and  A232 );
 a58402a <=( a58401a  and  a58398a );
 a58403a <=( a58402a  and  a58395a );
 a58406a <=( (not A235)  and  (not A234) );
 a58409a <=( (not A266)  and  (not A265) );
 a58410a <=( a58409a  and  a58406a );
 a58413a <=( A298  and  (not A268) );
 a58416a <=( A302  and  (not A299) );
 a58417a <=( a58416a  and  a58413a );
 a58418a <=( a58417a  and  a58410a );
 a58421a <=( A167  and  A168 );
 a58424a <=( A200  and  A199 );
 a58425a <=( a58424a  and  a58421a );
 a58428a <=( (not A202)  and  (not A201) );
 a58431a <=( A233  and  A232 );
 a58432a <=( a58431a  and  a58428a );
 a58433a <=( a58432a  and  a58425a );
 a58436a <=( (not A235)  and  (not A234) );
 a58439a <=( (not A266)  and  (not A265) );
 a58440a <=( a58439a  and  a58436a );
 a58443a <=( (not A298)  and  (not A268) );
 a58446a <=( A302  and  A299 );
 a58447a <=( a58446a  and  a58443a );
 a58448a <=( a58447a  and  a58440a );
 a58451a <=( A167  and  A168 );
 a58454a <=( A200  and  A199 );
 a58455a <=( a58454a  and  a58451a );
 a58458a <=( (not A202)  and  (not A201) );
 a58461a <=( (not A233)  and  (not A232) );
 a58462a <=( a58461a  and  a58458a );
 a58463a <=( a58462a  and  a58455a );
 a58466a <=( A265  and  (not A235) );
 a58469a <=( (not A267)  and  A266 );
 a58470a <=( a58469a  and  a58466a );
 a58473a <=( A298  and  (not A268) );
 a58476a <=( A302  and  (not A299) );
 a58477a <=( a58476a  and  a58473a );
 a58478a <=( a58477a  and  a58470a );
 a58481a <=( A167  and  A168 );
 a58484a <=( A200  and  A199 );
 a58485a <=( a58484a  and  a58481a );
 a58488a <=( (not A202)  and  (not A201) );
 a58491a <=( (not A233)  and  (not A232) );
 a58492a <=( a58491a  and  a58488a );
 a58493a <=( a58492a  and  a58485a );
 a58496a <=( A265  and  (not A235) );
 a58499a <=( (not A267)  and  A266 );
 a58500a <=( a58499a  and  a58496a );
 a58503a <=( (not A298)  and  (not A268) );
 a58506a <=( A302  and  A299 );
 a58507a <=( a58506a  and  a58503a );
 a58508a <=( a58507a  and  a58500a );
 a58511a <=( A167  and  A168 );
 a58514a <=( (not A200)  and  (not A199) );
 a58515a <=( a58514a  and  a58511a );
 a58518a <=( A232  and  (not A202) );
 a58521a <=( (not A234)  and  A233 );
 a58522a <=( a58521a  and  a58518a );
 a58523a <=( a58522a  and  a58515a );
 a58526a <=( A265  and  (not A235) );
 a58529a <=( (not A267)  and  A266 );
 a58530a <=( a58529a  and  a58526a );
 a58533a <=( A298  and  (not A268) );
 a58536a <=( A302  and  (not A299) );
 a58537a <=( a58536a  and  a58533a );
 a58538a <=( a58537a  and  a58530a );
 a58541a <=( A167  and  A168 );
 a58544a <=( (not A200)  and  (not A199) );
 a58545a <=( a58544a  and  a58541a );
 a58548a <=( A232  and  (not A202) );
 a58551a <=( (not A234)  and  A233 );
 a58552a <=( a58551a  and  a58548a );
 a58553a <=( a58552a  and  a58545a );
 a58556a <=( A265  and  (not A235) );
 a58559a <=( (not A267)  and  A266 );
 a58560a <=( a58559a  and  a58556a );
 a58563a <=( (not A298)  and  (not A268) );
 a58566a <=( A302  and  A299 );
 a58567a <=( a58566a  and  a58563a );
 a58568a <=( a58567a  and  a58560a );
 a58571a <=( A167  and  A170 );
 a58574a <=( (not A201)  and  (not A166) );
 a58575a <=( a58574a  and  a58571a );
 a58578a <=( (not A203)  and  (not A202) );
 a58581a <=( (not A235)  and  (not A234) );
 a58582a <=( a58581a  and  a58578a );
 a58583a <=( a58582a  and  a58575a );
 a58586a <=( A265  and  (not A236) );
 a58589a <=( (not A267)  and  A266 );
 a58590a <=( a58589a  and  a58586a );
 a58593a <=( A298  and  (not A268) );
 a58596a <=( A302  and  (not A299) );
 a58597a <=( a58596a  and  a58593a );
 a58598a <=( a58597a  and  a58590a );
 a58601a <=( A167  and  A170 );
 a58604a <=( (not A201)  and  (not A166) );
 a58605a <=( a58604a  and  a58601a );
 a58608a <=( (not A203)  and  (not A202) );
 a58611a <=( (not A235)  and  (not A234) );
 a58612a <=( a58611a  and  a58608a );
 a58613a <=( a58612a  and  a58605a );
 a58616a <=( A265  and  (not A236) );
 a58619a <=( (not A267)  and  A266 );
 a58620a <=( a58619a  and  a58616a );
 a58623a <=( (not A298)  and  (not A268) );
 a58626a <=( A302  and  A299 );
 a58627a <=( a58626a  and  a58623a );
 a58628a <=( a58627a  and  a58620a );
 a58631a <=( A167  and  A170 );
 a58634a <=( (not A201)  and  (not A166) );
 a58635a <=( a58634a  and  a58631a );
 a58638a <=( (not A203)  and  (not A202) );
 a58641a <=( A233  and  A232 );
 a58642a <=( a58641a  and  a58638a );
 a58643a <=( a58642a  and  a58635a );
 a58646a <=( (not A235)  and  (not A234) );
 a58649a <=( (not A268)  and  (not A267) );
 a58650a <=( a58649a  and  a58646a );
 a58653a <=( A298  and  (not A269) );
 a58656a <=( A302  and  (not A299) );
 a58657a <=( a58656a  and  a58653a );
 a58658a <=( a58657a  and  a58650a );
 a58661a <=( A167  and  A170 );
 a58664a <=( (not A201)  and  (not A166) );
 a58665a <=( a58664a  and  a58661a );
 a58668a <=( (not A203)  and  (not A202) );
 a58671a <=( A233  and  A232 );
 a58672a <=( a58671a  and  a58668a );
 a58673a <=( a58672a  and  a58665a );
 a58676a <=( (not A235)  and  (not A234) );
 a58679a <=( (not A268)  and  (not A267) );
 a58680a <=( a58679a  and  a58676a );
 a58683a <=( (not A298)  and  (not A269) );
 a58686a <=( A302  and  A299 );
 a58687a <=( a58686a  and  a58683a );
 a58688a <=( a58687a  and  a58680a );
 a58691a <=( A167  and  A170 );
 a58694a <=( (not A201)  and  (not A166) );
 a58695a <=( a58694a  and  a58691a );
 a58698a <=( (not A203)  and  (not A202) );
 a58701a <=( A233  and  A232 );
 a58702a <=( a58701a  and  a58698a );
 a58703a <=( a58702a  and  a58695a );
 a58706a <=( (not A235)  and  (not A234) );
 a58709a <=( A266  and  A265 );
 a58710a <=( a58709a  and  a58706a );
 a58713a <=( (not A268)  and  (not A267) );
 a58716a <=( A300  and  A299 );
 a58717a <=( a58716a  and  a58713a );
 a58718a <=( a58717a  and  a58710a );
 a58721a <=( A167  and  A170 );
 a58724a <=( (not A201)  and  (not A166) );
 a58725a <=( a58724a  and  a58721a );
 a58728a <=( (not A203)  and  (not A202) );
 a58731a <=( A233  and  A232 );
 a58732a <=( a58731a  and  a58728a );
 a58733a <=( a58732a  and  a58725a );
 a58736a <=( (not A235)  and  (not A234) );
 a58739a <=( A266  and  A265 );
 a58740a <=( a58739a  and  a58736a );
 a58743a <=( (not A268)  and  (not A267) );
 a58746a <=( A300  and  A298 );
 a58747a <=( a58746a  and  a58743a );
 a58748a <=( a58747a  and  a58740a );
 a58751a <=( A167  and  A170 );
 a58754a <=( (not A201)  and  (not A166) );
 a58755a <=( a58754a  and  a58751a );
 a58758a <=( (not A203)  and  (not A202) );
 a58761a <=( A233  and  A232 );
 a58762a <=( a58761a  and  a58758a );
 a58763a <=( a58762a  and  a58755a );
 a58766a <=( (not A235)  and  (not A234) );
 a58769a <=( (not A266)  and  (not A265) );
 a58770a <=( a58769a  and  a58766a );
 a58773a <=( A298  and  (not A268) );
 a58776a <=( A302  and  (not A299) );
 a58777a <=( a58776a  and  a58773a );
 a58778a <=( a58777a  and  a58770a );
 a58781a <=( A167  and  A170 );
 a58784a <=( (not A201)  and  (not A166) );
 a58785a <=( a58784a  and  a58781a );
 a58788a <=( (not A203)  and  (not A202) );
 a58791a <=( A233  and  A232 );
 a58792a <=( a58791a  and  a58788a );
 a58793a <=( a58792a  and  a58785a );
 a58796a <=( (not A235)  and  (not A234) );
 a58799a <=( (not A266)  and  (not A265) );
 a58800a <=( a58799a  and  a58796a );
 a58803a <=( (not A298)  and  (not A268) );
 a58806a <=( A302  and  A299 );
 a58807a <=( a58806a  and  a58803a );
 a58808a <=( a58807a  and  a58800a );
 a58811a <=( A167  and  A170 );
 a58814a <=( (not A201)  and  (not A166) );
 a58815a <=( a58814a  and  a58811a );
 a58818a <=( (not A203)  and  (not A202) );
 a58821a <=( (not A233)  and  (not A232) );
 a58822a <=( a58821a  and  a58818a );
 a58823a <=( a58822a  and  a58815a );
 a58826a <=( A265  and  (not A235) );
 a58829a <=( (not A267)  and  A266 );
 a58830a <=( a58829a  and  a58826a );
 a58833a <=( A298  and  (not A268) );
 a58836a <=( A302  and  (not A299) );
 a58837a <=( a58836a  and  a58833a );
 a58838a <=( a58837a  and  a58830a );
 a58841a <=( A167  and  A170 );
 a58844a <=( (not A201)  and  (not A166) );
 a58845a <=( a58844a  and  a58841a );
 a58848a <=( (not A203)  and  (not A202) );
 a58851a <=( (not A233)  and  (not A232) );
 a58852a <=( a58851a  and  a58848a );
 a58853a <=( a58852a  and  a58845a );
 a58856a <=( A265  and  (not A235) );
 a58859a <=( (not A267)  and  A266 );
 a58860a <=( a58859a  and  a58856a );
 a58863a <=( (not A298)  and  (not A268) );
 a58866a <=( A302  and  A299 );
 a58867a <=( a58866a  and  a58863a );
 a58868a <=( a58867a  and  a58860a );
 a58871a <=( A167  and  A170 );
 a58874a <=( A199  and  (not A166) );
 a58875a <=( a58874a  and  a58871a );
 a58878a <=( (not A201)  and  A200 );
 a58881a <=( (not A234)  and  (not A202) );
 a58882a <=( a58881a  and  a58878a );
 a58883a <=( a58882a  and  a58875a );
 a58886a <=( (not A236)  and  (not A235) );
 a58889a <=( (not A268)  and  (not A267) );
 a58890a <=( a58889a  and  a58886a );
 a58893a <=( A298  and  (not A269) );
 a58896a <=( A302  and  (not A299) );
 a58897a <=( a58896a  and  a58893a );
 a58898a <=( a58897a  and  a58890a );
 a58901a <=( A167  and  A170 );
 a58904a <=( A199  and  (not A166) );
 a58905a <=( a58904a  and  a58901a );
 a58908a <=( (not A201)  and  A200 );
 a58911a <=( (not A234)  and  (not A202) );
 a58912a <=( a58911a  and  a58908a );
 a58913a <=( a58912a  and  a58905a );
 a58916a <=( (not A236)  and  (not A235) );
 a58919a <=( (not A268)  and  (not A267) );
 a58920a <=( a58919a  and  a58916a );
 a58923a <=( (not A298)  and  (not A269) );
 a58926a <=( A302  and  A299 );
 a58927a <=( a58926a  and  a58923a );
 a58928a <=( a58927a  and  a58920a );
 a58931a <=( A167  and  A170 );
 a58934a <=( A199  and  (not A166) );
 a58935a <=( a58934a  and  a58931a );
 a58938a <=( (not A201)  and  A200 );
 a58941a <=( (not A234)  and  (not A202) );
 a58942a <=( a58941a  and  a58938a );
 a58943a <=( a58942a  and  a58935a );
 a58946a <=( (not A236)  and  (not A235) );
 a58949a <=( A266  and  A265 );
 a58950a <=( a58949a  and  a58946a );
 a58953a <=( (not A268)  and  (not A267) );
 a58956a <=( A300  and  A299 );
 a58957a <=( a58956a  and  a58953a );
 a58958a <=( a58957a  and  a58950a );
 a58961a <=( A167  and  A170 );
 a58964a <=( A199  and  (not A166) );
 a58965a <=( a58964a  and  a58961a );
 a58968a <=( (not A201)  and  A200 );
 a58971a <=( (not A234)  and  (not A202) );
 a58972a <=( a58971a  and  a58968a );
 a58973a <=( a58972a  and  a58965a );
 a58976a <=( (not A236)  and  (not A235) );
 a58979a <=( A266  and  A265 );
 a58980a <=( a58979a  and  a58976a );
 a58983a <=( (not A268)  and  (not A267) );
 a58986a <=( A300  and  A298 );
 a58987a <=( a58986a  and  a58983a );
 a58988a <=( a58987a  and  a58980a );
 a58991a <=( A167  and  A170 );
 a58994a <=( A199  and  (not A166) );
 a58995a <=( a58994a  and  a58991a );
 a58998a <=( (not A201)  and  A200 );
 a59001a <=( (not A234)  and  (not A202) );
 a59002a <=( a59001a  and  a58998a );
 a59003a <=( a59002a  and  a58995a );
 a59006a <=( (not A236)  and  (not A235) );
 a59009a <=( (not A266)  and  (not A265) );
 a59010a <=( a59009a  and  a59006a );
 a59013a <=( A298  and  (not A268) );
 a59016a <=( A302  and  (not A299) );
 a59017a <=( a59016a  and  a59013a );
 a59018a <=( a59017a  and  a59010a );
 a59021a <=( A167  and  A170 );
 a59024a <=( A199  and  (not A166) );
 a59025a <=( a59024a  and  a59021a );
 a59028a <=( (not A201)  and  A200 );
 a59031a <=( (not A234)  and  (not A202) );
 a59032a <=( a59031a  and  a59028a );
 a59033a <=( a59032a  and  a59025a );
 a59036a <=( (not A236)  and  (not A235) );
 a59039a <=( (not A266)  and  (not A265) );
 a59040a <=( a59039a  and  a59036a );
 a59043a <=( (not A298)  and  (not A268) );
 a59046a <=( A302  and  A299 );
 a59047a <=( a59046a  and  a59043a );
 a59048a <=( a59047a  and  a59040a );
 a59051a <=( A167  and  A170 );
 a59054a <=( A199  and  (not A166) );
 a59055a <=( a59054a  and  a59051a );
 a59058a <=( (not A201)  and  A200 );
 a59061a <=( A232  and  (not A202) );
 a59062a <=( a59061a  and  a59058a );
 a59063a <=( a59062a  and  a59055a );
 a59066a <=( (not A234)  and  A233 );
 a59069a <=( (not A267)  and  (not A235) );
 a59070a <=( a59069a  and  a59066a );
 a59073a <=( (not A269)  and  (not A268) );
 a59076a <=( A300  and  A299 );
 a59077a <=( a59076a  and  a59073a );
 a59078a <=( a59077a  and  a59070a );
 a59081a <=( A167  and  A170 );
 a59084a <=( A199  and  (not A166) );
 a59085a <=( a59084a  and  a59081a );
 a59088a <=( (not A201)  and  A200 );
 a59091a <=( A232  and  (not A202) );
 a59092a <=( a59091a  and  a59088a );
 a59093a <=( a59092a  and  a59085a );
 a59096a <=( (not A234)  and  A233 );
 a59099a <=( (not A267)  and  (not A235) );
 a59100a <=( a59099a  and  a59096a );
 a59103a <=( (not A269)  and  (not A268) );
 a59106a <=( A300  and  A298 );
 a59107a <=( a59106a  and  a59103a );
 a59108a <=( a59107a  and  a59100a );
 a59111a <=( A167  and  A170 );
 a59114a <=( A199  and  (not A166) );
 a59115a <=( a59114a  and  a59111a );
 a59118a <=( (not A201)  and  A200 );
 a59121a <=( A232  and  (not A202) );
 a59122a <=( a59121a  and  a59118a );
 a59123a <=( a59122a  and  a59115a );
 a59126a <=( (not A234)  and  A233 );
 a59129a <=( A265  and  (not A235) );
 a59130a <=( a59129a  and  a59126a );
 a59133a <=( (not A267)  and  A266 );
 a59136a <=( A301  and  (not A268) );
 a59137a <=( a59136a  and  a59133a );
 a59138a <=( a59137a  and  a59130a );
 a59141a <=( A167  and  A170 );
 a59144a <=( A199  and  (not A166) );
 a59145a <=( a59144a  and  a59141a );
 a59148a <=( (not A201)  and  A200 );
 a59151a <=( A232  and  (not A202) );
 a59152a <=( a59151a  and  a59148a );
 a59153a <=( a59152a  and  a59145a );
 a59156a <=( (not A234)  and  A233 );
 a59159a <=( (not A265)  and  (not A235) );
 a59160a <=( a59159a  and  a59156a );
 a59163a <=( (not A268)  and  (not A266) );
 a59166a <=( A300  and  A299 );
 a59167a <=( a59166a  and  a59163a );
 a59168a <=( a59167a  and  a59160a );
 a59171a <=( A167  and  A170 );
 a59174a <=( A199  and  (not A166) );
 a59175a <=( a59174a  and  a59171a );
 a59178a <=( (not A201)  and  A200 );
 a59181a <=( A232  and  (not A202) );
 a59182a <=( a59181a  and  a59178a );
 a59183a <=( a59182a  and  a59175a );
 a59186a <=( (not A234)  and  A233 );
 a59189a <=( (not A265)  and  (not A235) );
 a59190a <=( a59189a  and  a59186a );
 a59193a <=( (not A268)  and  (not A266) );
 a59196a <=( A300  and  A298 );
 a59197a <=( a59196a  and  a59193a );
 a59198a <=( a59197a  and  a59190a );
 a59201a <=( A167  and  A170 );
 a59204a <=( A199  and  (not A166) );
 a59205a <=( a59204a  and  a59201a );
 a59208a <=( (not A201)  and  A200 );
 a59211a <=( (not A232)  and  (not A202) );
 a59212a <=( a59211a  and  a59208a );
 a59213a <=( a59212a  and  a59205a );
 a59216a <=( (not A235)  and  (not A233) );
 a59219a <=( (not A268)  and  (not A267) );
 a59220a <=( a59219a  and  a59216a );
 a59223a <=( A298  and  (not A269) );
 a59226a <=( A302  and  (not A299) );
 a59227a <=( a59226a  and  a59223a );
 a59228a <=( a59227a  and  a59220a );
 a59231a <=( A167  and  A170 );
 a59234a <=( A199  and  (not A166) );
 a59235a <=( a59234a  and  a59231a );
 a59238a <=( (not A201)  and  A200 );
 a59241a <=( (not A232)  and  (not A202) );
 a59242a <=( a59241a  and  a59238a );
 a59243a <=( a59242a  and  a59235a );
 a59246a <=( (not A235)  and  (not A233) );
 a59249a <=( (not A268)  and  (not A267) );
 a59250a <=( a59249a  and  a59246a );
 a59253a <=( (not A298)  and  (not A269) );
 a59256a <=( A302  and  A299 );
 a59257a <=( a59256a  and  a59253a );
 a59258a <=( a59257a  and  a59250a );
 a59261a <=( A167  and  A170 );
 a59264a <=( A199  and  (not A166) );
 a59265a <=( a59264a  and  a59261a );
 a59268a <=( (not A201)  and  A200 );
 a59271a <=( (not A232)  and  (not A202) );
 a59272a <=( a59271a  and  a59268a );
 a59273a <=( a59272a  and  a59265a );
 a59276a <=( (not A235)  and  (not A233) );
 a59279a <=( A266  and  A265 );
 a59280a <=( a59279a  and  a59276a );
 a59283a <=( (not A268)  and  (not A267) );
 a59286a <=( A300  and  A299 );
 a59287a <=( a59286a  and  a59283a );
 a59288a <=( a59287a  and  a59280a );
 a59291a <=( A167  and  A170 );
 a59294a <=( A199  and  (not A166) );
 a59295a <=( a59294a  and  a59291a );
 a59298a <=( (not A201)  and  A200 );
 a59301a <=( (not A232)  and  (not A202) );
 a59302a <=( a59301a  and  a59298a );
 a59303a <=( a59302a  and  a59295a );
 a59306a <=( (not A235)  and  (not A233) );
 a59309a <=( A266  and  A265 );
 a59310a <=( a59309a  and  a59306a );
 a59313a <=( (not A268)  and  (not A267) );
 a59316a <=( A300  and  A298 );
 a59317a <=( a59316a  and  a59313a );
 a59318a <=( a59317a  and  a59310a );
 a59321a <=( A167  and  A170 );
 a59324a <=( A199  and  (not A166) );
 a59325a <=( a59324a  and  a59321a );
 a59328a <=( (not A201)  and  A200 );
 a59331a <=( (not A232)  and  (not A202) );
 a59332a <=( a59331a  and  a59328a );
 a59333a <=( a59332a  and  a59325a );
 a59336a <=( (not A235)  and  (not A233) );
 a59339a <=( (not A266)  and  (not A265) );
 a59340a <=( a59339a  and  a59336a );
 a59343a <=( A298  and  (not A268) );
 a59346a <=( A302  and  (not A299) );
 a59347a <=( a59346a  and  a59343a );
 a59348a <=( a59347a  and  a59340a );
 a59351a <=( A167  and  A170 );
 a59354a <=( A199  and  (not A166) );
 a59355a <=( a59354a  and  a59351a );
 a59358a <=( (not A201)  and  A200 );
 a59361a <=( (not A232)  and  (not A202) );
 a59362a <=( a59361a  and  a59358a );
 a59363a <=( a59362a  and  a59355a );
 a59366a <=( (not A235)  and  (not A233) );
 a59369a <=( (not A266)  and  (not A265) );
 a59370a <=( a59369a  and  a59366a );
 a59373a <=( (not A298)  and  (not A268) );
 a59376a <=( A302  and  A299 );
 a59377a <=( a59376a  and  a59373a );
 a59378a <=( a59377a  and  a59370a );
 a59381a <=( A167  and  A170 );
 a59384a <=( (not A199)  and  (not A166) );
 a59385a <=( a59384a  and  a59381a );
 a59388a <=( (not A202)  and  (not A200) );
 a59391a <=( (not A235)  and  (not A234) );
 a59392a <=( a59391a  and  a59388a );
 a59393a <=( a59392a  and  a59385a );
 a59396a <=( A265  and  (not A236) );
 a59399a <=( (not A267)  and  A266 );
 a59400a <=( a59399a  and  a59396a );
 a59403a <=( A298  and  (not A268) );
 a59406a <=( A302  and  (not A299) );
 a59407a <=( a59406a  and  a59403a );
 a59408a <=( a59407a  and  a59400a );
 a59411a <=( A167  and  A170 );
 a59414a <=( (not A199)  and  (not A166) );
 a59415a <=( a59414a  and  a59411a );
 a59418a <=( (not A202)  and  (not A200) );
 a59421a <=( (not A235)  and  (not A234) );
 a59422a <=( a59421a  and  a59418a );
 a59423a <=( a59422a  and  a59415a );
 a59426a <=( A265  and  (not A236) );
 a59429a <=( (not A267)  and  A266 );
 a59430a <=( a59429a  and  a59426a );
 a59433a <=( (not A298)  and  (not A268) );
 a59436a <=( A302  and  A299 );
 a59437a <=( a59436a  and  a59433a );
 a59438a <=( a59437a  and  a59430a );
 a59441a <=( A167  and  A170 );
 a59444a <=( (not A199)  and  (not A166) );
 a59445a <=( a59444a  and  a59441a );
 a59448a <=( (not A202)  and  (not A200) );
 a59451a <=( A233  and  A232 );
 a59452a <=( a59451a  and  a59448a );
 a59453a <=( a59452a  and  a59445a );
 a59456a <=( (not A235)  and  (not A234) );
 a59459a <=( (not A268)  and  (not A267) );
 a59460a <=( a59459a  and  a59456a );
 a59463a <=( A298  and  (not A269) );
 a59466a <=( A302  and  (not A299) );
 a59467a <=( a59466a  and  a59463a );
 a59468a <=( a59467a  and  a59460a );
 a59471a <=( A167  and  A170 );
 a59474a <=( (not A199)  and  (not A166) );
 a59475a <=( a59474a  and  a59471a );
 a59478a <=( (not A202)  and  (not A200) );
 a59481a <=( A233  and  A232 );
 a59482a <=( a59481a  and  a59478a );
 a59483a <=( a59482a  and  a59475a );
 a59486a <=( (not A235)  and  (not A234) );
 a59489a <=( (not A268)  and  (not A267) );
 a59490a <=( a59489a  and  a59486a );
 a59493a <=( (not A298)  and  (not A269) );
 a59496a <=( A302  and  A299 );
 a59497a <=( a59496a  and  a59493a );
 a59498a <=( a59497a  and  a59490a );
 a59501a <=( A167  and  A170 );
 a59504a <=( (not A199)  and  (not A166) );
 a59505a <=( a59504a  and  a59501a );
 a59508a <=( (not A202)  and  (not A200) );
 a59511a <=( A233  and  A232 );
 a59512a <=( a59511a  and  a59508a );
 a59513a <=( a59512a  and  a59505a );
 a59516a <=( (not A235)  and  (not A234) );
 a59519a <=( A266  and  A265 );
 a59520a <=( a59519a  and  a59516a );
 a59523a <=( (not A268)  and  (not A267) );
 a59526a <=( A300  and  A299 );
 a59527a <=( a59526a  and  a59523a );
 a59528a <=( a59527a  and  a59520a );
 a59531a <=( A167  and  A170 );
 a59534a <=( (not A199)  and  (not A166) );
 a59535a <=( a59534a  and  a59531a );
 a59538a <=( (not A202)  and  (not A200) );
 a59541a <=( A233  and  A232 );
 a59542a <=( a59541a  and  a59538a );
 a59543a <=( a59542a  and  a59535a );
 a59546a <=( (not A235)  and  (not A234) );
 a59549a <=( A266  and  A265 );
 a59550a <=( a59549a  and  a59546a );
 a59553a <=( (not A268)  and  (not A267) );
 a59556a <=( A300  and  A298 );
 a59557a <=( a59556a  and  a59553a );
 a59558a <=( a59557a  and  a59550a );
 a59561a <=( A167  and  A170 );
 a59564a <=( (not A199)  and  (not A166) );
 a59565a <=( a59564a  and  a59561a );
 a59568a <=( (not A202)  and  (not A200) );
 a59571a <=( A233  and  A232 );
 a59572a <=( a59571a  and  a59568a );
 a59573a <=( a59572a  and  a59565a );
 a59576a <=( (not A235)  and  (not A234) );
 a59579a <=( (not A266)  and  (not A265) );
 a59580a <=( a59579a  and  a59576a );
 a59583a <=( A298  and  (not A268) );
 a59586a <=( A302  and  (not A299) );
 a59587a <=( a59586a  and  a59583a );
 a59588a <=( a59587a  and  a59580a );
 a59591a <=( A167  and  A170 );
 a59594a <=( (not A199)  and  (not A166) );
 a59595a <=( a59594a  and  a59591a );
 a59598a <=( (not A202)  and  (not A200) );
 a59601a <=( A233  and  A232 );
 a59602a <=( a59601a  and  a59598a );
 a59603a <=( a59602a  and  a59595a );
 a59606a <=( (not A235)  and  (not A234) );
 a59609a <=( (not A266)  and  (not A265) );
 a59610a <=( a59609a  and  a59606a );
 a59613a <=( (not A298)  and  (not A268) );
 a59616a <=( A302  and  A299 );
 a59617a <=( a59616a  and  a59613a );
 a59618a <=( a59617a  and  a59610a );
 a59621a <=( A167  and  A170 );
 a59624a <=( (not A199)  and  (not A166) );
 a59625a <=( a59624a  and  a59621a );
 a59628a <=( (not A202)  and  (not A200) );
 a59631a <=( (not A233)  and  (not A232) );
 a59632a <=( a59631a  and  a59628a );
 a59633a <=( a59632a  and  a59625a );
 a59636a <=( A265  and  (not A235) );
 a59639a <=( (not A267)  and  A266 );
 a59640a <=( a59639a  and  a59636a );
 a59643a <=( A298  and  (not A268) );
 a59646a <=( A302  and  (not A299) );
 a59647a <=( a59646a  and  a59643a );
 a59648a <=( a59647a  and  a59640a );
 a59651a <=( A167  and  A170 );
 a59654a <=( (not A199)  and  (not A166) );
 a59655a <=( a59654a  and  a59651a );
 a59658a <=( (not A202)  and  (not A200) );
 a59661a <=( (not A233)  and  (not A232) );
 a59662a <=( a59661a  and  a59658a );
 a59663a <=( a59662a  and  a59655a );
 a59666a <=( A265  and  (not A235) );
 a59669a <=( (not A267)  and  A266 );
 a59670a <=( a59669a  and  a59666a );
 a59673a <=( (not A298)  and  (not A268) );
 a59676a <=( A302  and  A299 );
 a59677a <=( a59676a  and  a59673a );
 a59678a <=( a59677a  and  a59670a );
 a59681a <=( (not A167)  and  A170 );
 a59684a <=( (not A201)  and  A166 );
 a59685a <=( a59684a  and  a59681a );
 a59688a <=( (not A203)  and  (not A202) );
 a59691a <=( (not A235)  and  (not A234) );
 a59692a <=( a59691a  and  a59688a );
 a59693a <=( a59692a  and  a59685a );
 a59696a <=( A265  and  (not A236) );
 a59699a <=( (not A267)  and  A266 );
 a59700a <=( a59699a  and  a59696a );
 a59703a <=( A298  and  (not A268) );
 a59706a <=( A302  and  (not A299) );
 a59707a <=( a59706a  and  a59703a );
 a59708a <=( a59707a  and  a59700a );
 a59711a <=( (not A167)  and  A170 );
 a59714a <=( (not A201)  and  A166 );
 a59715a <=( a59714a  and  a59711a );
 a59718a <=( (not A203)  and  (not A202) );
 a59721a <=( (not A235)  and  (not A234) );
 a59722a <=( a59721a  and  a59718a );
 a59723a <=( a59722a  and  a59715a );
 a59726a <=( A265  and  (not A236) );
 a59729a <=( (not A267)  and  A266 );
 a59730a <=( a59729a  and  a59726a );
 a59733a <=( (not A298)  and  (not A268) );
 a59736a <=( A302  and  A299 );
 a59737a <=( a59736a  and  a59733a );
 a59738a <=( a59737a  and  a59730a );
 a59741a <=( (not A167)  and  A170 );
 a59744a <=( (not A201)  and  A166 );
 a59745a <=( a59744a  and  a59741a );
 a59748a <=( (not A203)  and  (not A202) );
 a59751a <=( A233  and  A232 );
 a59752a <=( a59751a  and  a59748a );
 a59753a <=( a59752a  and  a59745a );
 a59756a <=( (not A235)  and  (not A234) );
 a59759a <=( (not A268)  and  (not A267) );
 a59760a <=( a59759a  and  a59756a );
 a59763a <=( A298  and  (not A269) );
 a59766a <=( A302  and  (not A299) );
 a59767a <=( a59766a  and  a59763a );
 a59768a <=( a59767a  and  a59760a );
 a59771a <=( (not A167)  and  A170 );
 a59774a <=( (not A201)  and  A166 );
 a59775a <=( a59774a  and  a59771a );
 a59778a <=( (not A203)  and  (not A202) );
 a59781a <=( A233  and  A232 );
 a59782a <=( a59781a  and  a59778a );
 a59783a <=( a59782a  and  a59775a );
 a59786a <=( (not A235)  and  (not A234) );
 a59789a <=( (not A268)  and  (not A267) );
 a59790a <=( a59789a  and  a59786a );
 a59793a <=( (not A298)  and  (not A269) );
 a59796a <=( A302  and  A299 );
 a59797a <=( a59796a  and  a59793a );
 a59798a <=( a59797a  and  a59790a );
 a59801a <=( (not A167)  and  A170 );
 a59804a <=( (not A201)  and  A166 );
 a59805a <=( a59804a  and  a59801a );
 a59808a <=( (not A203)  and  (not A202) );
 a59811a <=( A233  and  A232 );
 a59812a <=( a59811a  and  a59808a );
 a59813a <=( a59812a  and  a59805a );
 a59816a <=( (not A235)  and  (not A234) );
 a59819a <=( A266  and  A265 );
 a59820a <=( a59819a  and  a59816a );
 a59823a <=( (not A268)  and  (not A267) );
 a59826a <=( A300  and  A299 );
 a59827a <=( a59826a  and  a59823a );
 a59828a <=( a59827a  and  a59820a );
 a59831a <=( (not A167)  and  A170 );
 a59834a <=( (not A201)  and  A166 );
 a59835a <=( a59834a  and  a59831a );
 a59838a <=( (not A203)  and  (not A202) );
 a59841a <=( A233  and  A232 );
 a59842a <=( a59841a  and  a59838a );
 a59843a <=( a59842a  and  a59835a );
 a59846a <=( (not A235)  and  (not A234) );
 a59849a <=( A266  and  A265 );
 a59850a <=( a59849a  and  a59846a );
 a59853a <=( (not A268)  and  (not A267) );
 a59856a <=( A300  and  A298 );
 a59857a <=( a59856a  and  a59853a );
 a59858a <=( a59857a  and  a59850a );
 a59861a <=( (not A167)  and  A170 );
 a59864a <=( (not A201)  and  A166 );
 a59865a <=( a59864a  and  a59861a );
 a59868a <=( (not A203)  and  (not A202) );
 a59871a <=( A233  and  A232 );
 a59872a <=( a59871a  and  a59868a );
 a59873a <=( a59872a  and  a59865a );
 a59876a <=( (not A235)  and  (not A234) );
 a59879a <=( (not A266)  and  (not A265) );
 a59880a <=( a59879a  and  a59876a );
 a59883a <=( A298  and  (not A268) );
 a59886a <=( A302  and  (not A299) );
 a59887a <=( a59886a  and  a59883a );
 a59888a <=( a59887a  and  a59880a );
 a59891a <=( (not A167)  and  A170 );
 a59894a <=( (not A201)  and  A166 );
 a59895a <=( a59894a  and  a59891a );
 a59898a <=( (not A203)  and  (not A202) );
 a59901a <=( A233  and  A232 );
 a59902a <=( a59901a  and  a59898a );
 a59903a <=( a59902a  and  a59895a );
 a59906a <=( (not A235)  and  (not A234) );
 a59909a <=( (not A266)  and  (not A265) );
 a59910a <=( a59909a  and  a59906a );
 a59913a <=( (not A298)  and  (not A268) );
 a59916a <=( A302  and  A299 );
 a59917a <=( a59916a  and  a59913a );
 a59918a <=( a59917a  and  a59910a );
 a59921a <=( (not A167)  and  A170 );
 a59924a <=( (not A201)  and  A166 );
 a59925a <=( a59924a  and  a59921a );
 a59928a <=( (not A203)  and  (not A202) );
 a59931a <=( (not A233)  and  (not A232) );
 a59932a <=( a59931a  and  a59928a );
 a59933a <=( a59932a  and  a59925a );
 a59936a <=( A265  and  (not A235) );
 a59939a <=( (not A267)  and  A266 );
 a59940a <=( a59939a  and  a59936a );
 a59943a <=( A298  and  (not A268) );
 a59946a <=( A302  and  (not A299) );
 a59947a <=( a59946a  and  a59943a );
 a59948a <=( a59947a  and  a59940a );
 a59951a <=( (not A167)  and  A170 );
 a59954a <=( (not A201)  and  A166 );
 a59955a <=( a59954a  and  a59951a );
 a59958a <=( (not A203)  and  (not A202) );
 a59961a <=( (not A233)  and  (not A232) );
 a59962a <=( a59961a  and  a59958a );
 a59963a <=( a59962a  and  a59955a );
 a59966a <=( A265  and  (not A235) );
 a59969a <=( (not A267)  and  A266 );
 a59970a <=( a59969a  and  a59966a );
 a59973a <=( (not A298)  and  (not A268) );
 a59976a <=( A302  and  A299 );
 a59977a <=( a59976a  and  a59973a );
 a59978a <=( a59977a  and  a59970a );
 a59981a <=( (not A167)  and  A170 );
 a59984a <=( A199  and  A166 );
 a59985a <=( a59984a  and  a59981a );
 a59988a <=( (not A201)  and  A200 );
 a59991a <=( (not A234)  and  (not A202) );
 a59992a <=( a59991a  and  a59988a );
 a59993a <=( a59992a  and  a59985a );
 a59996a <=( (not A236)  and  (not A235) );
 a59999a <=( (not A268)  and  (not A267) );
 a60000a <=( a59999a  and  a59996a );
 a60003a <=( A298  and  (not A269) );
 a60006a <=( A302  and  (not A299) );
 a60007a <=( a60006a  and  a60003a );
 a60008a <=( a60007a  and  a60000a );
 a60011a <=( (not A167)  and  A170 );
 a60014a <=( A199  and  A166 );
 a60015a <=( a60014a  and  a60011a );
 a60018a <=( (not A201)  and  A200 );
 a60021a <=( (not A234)  and  (not A202) );
 a60022a <=( a60021a  and  a60018a );
 a60023a <=( a60022a  and  a60015a );
 a60026a <=( (not A236)  and  (not A235) );
 a60029a <=( (not A268)  and  (not A267) );
 a60030a <=( a60029a  and  a60026a );
 a60033a <=( (not A298)  and  (not A269) );
 a60036a <=( A302  and  A299 );
 a60037a <=( a60036a  and  a60033a );
 a60038a <=( a60037a  and  a60030a );
 a60041a <=( (not A167)  and  A170 );
 a60044a <=( A199  and  A166 );
 a60045a <=( a60044a  and  a60041a );
 a60048a <=( (not A201)  and  A200 );
 a60051a <=( (not A234)  and  (not A202) );
 a60052a <=( a60051a  and  a60048a );
 a60053a <=( a60052a  and  a60045a );
 a60056a <=( (not A236)  and  (not A235) );
 a60059a <=( A266  and  A265 );
 a60060a <=( a60059a  and  a60056a );
 a60063a <=( (not A268)  and  (not A267) );
 a60066a <=( A300  and  A299 );
 a60067a <=( a60066a  and  a60063a );
 a60068a <=( a60067a  and  a60060a );
 a60071a <=( (not A167)  and  A170 );
 a60074a <=( A199  and  A166 );
 a60075a <=( a60074a  and  a60071a );
 a60078a <=( (not A201)  and  A200 );
 a60081a <=( (not A234)  and  (not A202) );
 a60082a <=( a60081a  and  a60078a );
 a60083a <=( a60082a  and  a60075a );
 a60086a <=( (not A236)  and  (not A235) );
 a60089a <=( A266  and  A265 );
 a60090a <=( a60089a  and  a60086a );
 a60093a <=( (not A268)  and  (not A267) );
 a60096a <=( A300  and  A298 );
 a60097a <=( a60096a  and  a60093a );
 a60098a <=( a60097a  and  a60090a );
 a60101a <=( (not A167)  and  A170 );
 a60104a <=( A199  and  A166 );
 a60105a <=( a60104a  and  a60101a );
 a60108a <=( (not A201)  and  A200 );
 a60111a <=( (not A234)  and  (not A202) );
 a60112a <=( a60111a  and  a60108a );
 a60113a <=( a60112a  and  a60105a );
 a60116a <=( (not A236)  and  (not A235) );
 a60119a <=( (not A266)  and  (not A265) );
 a60120a <=( a60119a  and  a60116a );
 a60123a <=( A298  and  (not A268) );
 a60126a <=( A302  and  (not A299) );
 a60127a <=( a60126a  and  a60123a );
 a60128a <=( a60127a  and  a60120a );
 a60131a <=( (not A167)  and  A170 );
 a60134a <=( A199  and  A166 );
 a60135a <=( a60134a  and  a60131a );
 a60138a <=( (not A201)  and  A200 );
 a60141a <=( (not A234)  and  (not A202) );
 a60142a <=( a60141a  and  a60138a );
 a60143a <=( a60142a  and  a60135a );
 a60146a <=( (not A236)  and  (not A235) );
 a60149a <=( (not A266)  and  (not A265) );
 a60150a <=( a60149a  and  a60146a );
 a60153a <=( (not A298)  and  (not A268) );
 a60156a <=( A302  and  A299 );
 a60157a <=( a60156a  and  a60153a );
 a60158a <=( a60157a  and  a60150a );
 a60161a <=( (not A167)  and  A170 );
 a60164a <=( A199  and  A166 );
 a60165a <=( a60164a  and  a60161a );
 a60168a <=( (not A201)  and  A200 );
 a60171a <=( A232  and  (not A202) );
 a60172a <=( a60171a  and  a60168a );
 a60173a <=( a60172a  and  a60165a );
 a60176a <=( (not A234)  and  A233 );
 a60179a <=( (not A267)  and  (not A235) );
 a60180a <=( a60179a  and  a60176a );
 a60183a <=( (not A269)  and  (not A268) );
 a60186a <=( A300  and  A299 );
 a60187a <=( a60186a  and  a60183a );
 a60188a <=( a60187a  and  a60180a );
 a60191a <=( (not A167)  and  A170 );
 a60194a <=( A199  and  A166 );
 a60195a <=( a60194a  and  a60191a );
 a60198a <=( (not A201)  and  A200 );
 a60201a <=( A232  and  (not A202) );
 a60202a <=( a60201a  and  a60198a );
 a60203a <=( a60202a  and  a60195a );
 a60206a <=( (not A234)  and  A233 );
 a60209a <=( (not A267)  and  (not A235) );
 a60210a <=( a60209a  and  a60206a );
 a60213a <=( (not A269)  and  (not A268) );
 a60216a <=( A300  and  A298 );
 a60217a <=( a60216a  and  a60213a );
 a60218a <=( a60217a  and  a60210a );
 a60221a <=( (not A167)  and  A170 );
 a60224a <=( A199  and  A166 );
 a60225a <=( a60224a  and  a60221a );
 a60228a <=( (not A201)  and  A200 );
 a60231a <=( A232  and  (not A202) );
 a60232a <=( a60231a  and  a60228a );
 a60233a <=( a60232a  and  a60225a );
 a60236a <=( (not A234)  and  A233 );
 a60239a <=( A265  and  (not A235) );
 a60240a <=( a60239a  and  a60236a );
 a60243a <=( (not A267)  and  A266 );
 a60246a <=( A301  and  (not A268) );
 a60247a <=( a60246a  and  a60243a );
 a60248a <=( a60247a  and  a60240a );
 a60251a <=( (not A167)  and  A170 );
 a60254a <=( A199  and  A166 );
 a60255a <=( a60254a  and  a60251a );
 a60258a <=( (not A201)  and  A200 );
 a60261a <=( A232  and  (not A202) );
 a60262a <=( a60261a  and  a60258a );
 a60263a <=( a60262a  and  a60255a );
 a60266a <=( (not A234)  and  A233 );
 a60269a <=( (not A265)  and  (not A235) );
 a60270a <=( a60269a  and  a60266a );
 a60273a <=( (not A268)  and  (not A266) );
 a60276a <=( A300  and  A299 );
 a60277a <=( a60276a  and  a60273a );
 a60278a <=( a60277a  and  a60270a );
 a60281a <=( (not A167)  and  A170 );
 a60284a <=( A199  and  A166 );
 a60285a <=( a60284a  and  a60281a );
 a60288a <=( (not A201)  and  A200 );
 a60291a <=( A232  and  (not A202) );
 a60292a <=( a60291a  and  a60288a );
 a60293a <=( a60292a  and  a60285a );
 a60296a <=( (not A234)  and  A233 );
 a60299a <=( (not A265)  and  (not A235) );
 a60300a <=( a60299a  and  a60296a );
 a60303a <=( (not A268)  and  (not A266) );
 a60306a <=( A300  and  A298 );
 a60307a <=( a60306a  and  a60303a );
 a60308a <=( a60307a  and  a60300a );
 a60311a <=( (not A167)  and  A170 );
 a60314a <=( A199  and  A166 );
 a60315a <=( a60314a  and  a60311a );
 a60318a <=( (not A201)  and  A200 );
 a60321a <=( (not A232)  and  (not A202) );
 a60322a <=( a60321a  and  a60318a );
 a60323a <=( a60322a  and  a60315a );
 a60326a <=( (not A235)  and  (not A233) );
 a60329a <=( (not A268)  and  (not A267) );
 a60330a <=( a60329a  and  a60326a );
 a60333a <=( A298  and  (not A269) );
 a60336a <=( A302  and  (not A299) );
 a60337a <=( a60336a  and  a60333a );
 a60338a <=( a60337a  and  a60330a );
 a60341a <=( (not A167)  and  A170 );
 a60344a <=( A199  and  A166 );
 a60345a <=( a60344a  and  a60341a );
 a60348a <=( (not A201)  and  A200 );
 a60351a <=( (not A232)  and  (not A202) );
 a60352a <=( a60351a  and  a60348a );
 a60353a <=( a60352a  and  a60345a );
 a60356a <=( (not A235)  and  (not A233) );
 a60359a <=( (not A268)  and  (not A267) );
 a60360a <=( a60359a  and  a60356a );
 a60363a <=( (not A298)  and  (not A269) );
 a60366a <=( A302  and  A299 );
 a60367a <=( a60366a  and  a60363a );
 a60368a <=( a60367a  and  a60360a );
 a60371a <=( (not A167)  and  A170 );
 a60374a <=( A199  and  A166 );
 a60375a <=( a60374a  and  a60371a );
 a60378a <=( (not A201)  and  A200 );
 a60381a <=( (not A232)  and  (not A202) );
 a60382a <=( a60381a  and  a60378a );
 a60383a <=( a60382a  and  a60375a );
 a60386a <=( (not A235)  and  (not A233) );
 a60389a <=( A266  and  A265 );
 a60390a <=( a60389a  and  a60386a );
 a60393a <=( (not A268)  and  (not A267) );
 a60396a <=( A300  and  A299 );
 a60397a <=( a60396a  and  a60393a );
 a60398a <=( a60397a  and  a60390a );
 a60401a <=( (not A167)  and  A170 );
 a60404a <=( A199  and  A166 );
 a60405a <=( a60404a  and  a60401a );
 a60408a <=( (not A201)  and  A200 );
 a60411a <=( (not A232)  and  (not A202) );
 a60412a <=( a60411a  and  a60408a );
 a60413a <=( a60412a  and  a60405a );
 a60416a <=( (not A235)  and  (not A233) );
 a60419a <=( A266  and  A265 );
 a60420a <=( a60419a  and  a60416a );
 a60423a <=( (not A268)  and  (not A267) );
 a60426a <=( A300  and  A298 );
 a60427a <=( a60426a  and  a60423a );
 a60428a <=( a60427a  and  a60420a );
 a60431a <=( (not A167)  and  A170 );
 a60434a <=( A199  and  A166 );
 a60435a <=( a60434a  and  a60431a );
 a60438a <=( (not A201)  and  A200 );
 a60441a <=( (not A232)  and  (not A202) );
 a60442a <=( a60441a  and  a60438a );
 a60443a <=( a60442a  and  a60435a );
 a60446a <=( (not A235)  and  (not A233) );
 a60449a <=( (not A266)  and  (not A265) );
 a60450a <=( a60449a  and  a60446a );
 a60453a <=( A298  and  (not A268) );
 a60456a <=( A302  and  (not A299) );
 a60457a <=( a60456a  and  a60453a );
 a60458a <=( a60457a  and  a60450a );
 a60461a <=( (not A167)  and  A170 );
 a60464a <=( A199  and  A166 );
 a60465a <=( a60464a  and  a60461a );
 a60468a <=( (not A201)  and  A200 );
 a60471a <=( (not A232)  and  (not A202) );
 a60472a <=( a60471a  and  a60468a );
 a60473a <=( a60472a  and  a60465a );
 a60476a <=( (not A235)  and  (not A233) );
 a60479a <=( (not A266)  and  (not A265) );
 a60480a <=( a60479a  and  a60476a );
 a60483a <=( (not A298)  and  (not A268) );
 a60486a <=( A302  and  A299 );
 a60487a <=( a60486a  and  a60483a );
 a60488a <=( a60487a  and  a60480a );
 a60491a <=( (not A167)  and  A170 );
 a60494a <=( (not A199)  and  A166 );
 a60495a <=( a60494a  and  a60491a );
 a60498a <=( (not A202)  and  (not A200) );
 a60501a <=( (not A235)  and  (not A234) );
 a60502a <=( a60501a  and  a60498a );
 a60503a <=( a60502a  and  a60495a );
 a60506a <=( A265  and  (not A236) );
 a60509a <=( (not A267)  and  A266 );
 a60510a <=( a60509a  and  a60506a );
 a60513a <=( A298  and  (not A268) );
 a60516a <=( A302  and  (not A299) );
 a60517a <=( a60516a  and  a60513a );
 a60518a <=( a60517a  and  a60510a );
 a60521a <=( (not A167)  and  A170 );
 a60524a <=( (not A199)  and  A166 );
 a60525a <=( a60524a  and  a60521a );
 a60528a <=( (not A202)  and  (not A200) );
 a60531a <=( (not A235)  and  (not A234) );
 a60532a <=( a60531a  and  a60528a );
 a60533a <=( a60532a  and  a60525a );
 a60536a <=( A265  and  (not A236) );
 a60539a <=( (not A267)  and  A266 );
 a60540a <=( a60539a  and  a60536a );
 a60543a <=( (not A298)  and  (not A268) );
 a60546a <=( A302  and  A299 );
 a60547a <=( a60546a  and  a60543a );
 a60548a <=( a60547a  and  a60540a );
 a60551a <=( (not A167)  and  A170 );
 a60554a <=( (not A199)  and  A166 );
 a60555a <=( a60554a  and  a60551a );
 a60558a <=( (not A202)  and  (not A200) );
 a60561a <=( A233  and  A232 );
 a60562a <=( a60561a  and  a60558a );
 a60563a <=( a60562a  and  a60555a );
 a60566a <=( (not A235)  and  (not A234) );
 a60569a <=( (not A268)  and  (not A267) );
 a60570a <=( a60569a  and  a60566a );
 a60573a <=( A298  and  (not A269) );
 a60576a <=( A302  and  (not A299) );
 a60577a <=( a60576a  and  a60573a );
 a60578a <=( a60577a  and  a60570a );
 a60581a <=( (not A167)  and  A170 );
 a60584a <=( (not A199)  and  A166 );
 a60585a <=( a60584a  and  a60581a );
 a60588a <=( (not A202)  and  (not A200) );
 a60591a <=( A233  and  A232 );
 a60592a <=( a60591a  and  a60588a );
 a60593a <=( a60592a  and  a60585a );
 a60596a <=( (not A235)  and  (not A234) );
 a60599a <=( (not A268)  and  (not A267) );
 a60600a <=( a60599a  and  a60596a );
 a60603a <=( (not A298)  and  (not A269) );
 a60606a <=( A302  and  A299 );
 a60607a <=( a60606a  and  a60603a );
 a60608a <=( a60607a  and  a60600a );
 a60611a <=( (not A167)  and  A170 );
 a60614a <=( (not A199)  and  A166 );
 a60615a <=( a60614a  and  a60611a );
 a60618a <=( (not A202)  and  (not A200) );
 a60621a <=( A233  and  A232 );
 a60622a <=( a60621a  and  a60618a );
 a60623a <=( a60622a  and  a60615a );
 a60626a <=( (not A235)  and  (not A234) );
 a60629a <=( A266  and  A265 );
 a60630a <=( a60629a  and  a60626a );
 a60633a <=( (not A268)  and  (not A267) );
 a60636a <=( A300  and  A299 );
 a60637a <=( a60636a  and  a60633a );
 a60638a <=( a60637a  and  a60630a );
 a60641a <=( (not A167)  and  A170 );
 a60644a <=( (not A199)  and  A166 );
 a60645a <=( a60644a  and  a60641a );
 a60648a <=( (not A202)  and  (not A200) );
 a60651a <=( A233  and  A232 );
 a60652a <=( a60651a  and  a60648a );
 a60653a <=( a60652a  and  a60645a );
 a60656a <=( (not A235)  and  (not A234) );
 a60659a <=( A266  and  A265 );
 a60660a <=( a60659a  and  a60656a );
 a60663a <=( (not A268)  and  (not A267) );
 a60666a <=( A300  and  A298 );
 a60667a <=( a60666a  and  a60663a );
 a60668a <=( a60667a  and  a60660a );
 a60671a <=( (not A167)  and  A170 );
 a60674a <=( (not A199)  and  A166 );
 a60675a <=( a60674a  and  a60671a );
 a60678a <=( (not A202)  and  (not A200) );
 a60681a <=( A233  and  A232 );
 a60682a <=( a60681a  and  a60678a );
 a60683a <=( a60682a  and  a60675a );
 a60686a <=( (not A235)  and  (not A234) );
 a60689a <=( (not A266)  and  (not A265) );
 a60690a <=( a60689a  and  a60686a );
 a60693a <=( A298  and  (not A268) );
 a60696a <=( A302  and  (not A299) );
 a60697a <=( a60696a  and  a60693a );
 a60698a <=( a60697a  and  a60690a );
 a60701a <=( (not A167)  and  A170 );
 a60704a <=( (not A199)  and  A166 );
 a60705a <=( a60704a  and  a60701a );
 a60708a <=( (not A202)  and  (not A200) );
 a60711a <=( A233  and  A232 );
 a60712a <=( a60711a  and  a60708a );
 a60713a <=( a60712a  and  a60705a );
 a60716a <=( (not A235)  and  (not A234) );
 a60719a <=( (not A266)  and  (not A265) );
 a60720a <=( a60719a  and  a60716a );
 a60723a <=( (not A298)  and  (not A268) );
 a60726a <=( A302  and  A299 );
 a60727a <=( a60726a  and  a60723a );
 a60728a <=( a60727a  and  a60720a );
 a60731a <=( (not A167)  and  A170 );
 a60734a <=( (not A199)  and  A166 );
 a60735a <=( a60734a  and  a60731a );
 a60738a <=( (not A202)  and  (not A200) );
 a60741a <=( (not A233)  and  (not A232) );
 a60742a <=( a60741a  and  a60738a );
 a60743a <=( a60742a  and  a60735a );
 a60746a <=( A265  and  (not A235) );
 a60749a <=( (not A267)  and  A266 );
 a60750a <=( a60749a  and  a60746a );
 a60753a <=( A298  and  (not A268) );
 a60756a <=( A302  and  (not A299) );
 a60757a <=( a60756a  and  a60753a );
 a60758a <=( a60757a  and  a60750a );
 a60761a <=( (not A167)  and  A170 );
 a60764a <=( (not A199)  and  A166 );
 a60765a <=( a60764a  and  a60761a );
 a60768a <=( (not A202)  and  (not A200) );
 a60771a <=( (not A233)  and  (not A232) );
 a60772a <=( a60771a  and  a60768a );
 a60773a <=( a60772a  and  a60765a );
 a60776a <=( A265  and  (not A235) );
 a60779a <=( (not A267)  and  A266 );
 a60780a <=( a60779a  and  a60776a );
 a60783a <=( (not A298)  and  (not A268) );
 a60786a <=( A302  and  A299 );
 a60787a <=( a60786a  and  a60783a );
 a60788a <=( a60787a  and  a60780a );
 a60791a <=( A199  and  A169 );
 a60794a <=( (not A201)  and  A200 );
 a60795a <=( a60794a  and  a60791a );
 a60798a <=( A232  and  (not A202) );
 a60801a <=( (not A234)  and  A233 );
 a60802a <=( a60801a  and  a60798a );
 a60803a <=( a60802a  and  a60795a );
 a60806a <=( A265  and  (not A235) );
 a60809a <=( (not A267)  and  A266 );
 a60810a <=( a60809a  and  a60806a );
 a60813a <=( A298  and  (not A268) );
 a60816a <=( A302  and  (not A299) );
 a60817a <=( a60816a  and  a60813a );
 a60818a <=( a60817a  and  a60810a );
 a60821a <=( A199  and  A169 );
 a60824a <=( (not A201)  and  A200 );
 a60825a <=( a60824a  and  a60821a );
 a60828a <=( A232  and  (not A202) );
 a60831a <=( (not A234)  and  A233 );
 a60832a <=( a60831a  and  a60828a );
 a60833a <=( a60832a  and  a60825a );
 a60836a <=( A265  and  (not A235) );
 a60839a <=( (not A267)  and  A266 );
 a60840a <=( a60839a  and  a60836a );
 a60843a <=( (not A298)  and  (not A268) );
 a60846a <=( A302  and  A299 );
 a60847a <=( a60846a  and  a60843a );
 a60848a <=( a60847a  and  a60840a );
 a60851a <=( (not A167)  and  (not A169) );
 a60854a <=( A199  and  (not A166) );
 a60855a <=( a60854a  and  a60851a );
 a60858a <=( A232  and  A201 );
 a60861a <=( (not A234)  and  A233 );
 a60862a <=( a60861a  and  a60858a );
 a60863a <=( a60862a  and  a60855a );
 a60866a <=( A265  and  (not A235) );
 a60869a <=( (not A267)  and  A266 );
 a60870a <=( a60869a  and  a60866a );
 a60873a <=( A298  and  (not A268) );
 a60876a <=( A302  and  (not A299) );
 a60877a <=( a60876a  and  a60873a );
 a60878a <=( a60877a  and  a60870a );
 a60881a <=( (not A167)  and  (not A169) );
 a60884a <=( A199  and  (not A166) );
 a60885a <=( a60884a  and  a60881a );
 a60888a <=( A232  and  A201 );
 a60891a <=( (not A234)  and  A233 );
 a60892a <=( a60891a  and  a60888a );
 a60893a <=( a60892a  and  a60885a );
 a60896a <=( A265  and  (not A235) );
 a60899a <=( (not A267)  and  A266 );
 a60900a <=( a60899a  and  a60896a );
 a60903a <=( (not A298)  and  (not A268) );
 a60906a <=( A302  and  A299 );
 a60907a <=( a60906a  and  a60903a );
 a60908a <=( a60907a  and  a60900a );
 a60911a <=( (not A167)  and  (not A169) );
 a60914a <=( A200  and  (not A166) );
 a60915a <=( a60914a  and  a60911a );
 a60918a <=( A232  and  A201 );
 a60921a <=( (not A234)  and  A233 );
 a60922a <=( a60921a  and  a60918a );
 a60923a <=( a60922a  and  a60915a );
 a60926a <=( A265  and  (not A235) );
 a60929a <=( (not A267)  and  A266 );
 a60930a <=( a60929a  and  a60926a );
 a60933a <=( A298  and  (not A268) );
 a60936a <=( A302  and  (not A299) );
 a60937a <=( a60936a  and  a60933a );
 a60938a <=( a60937a  and  a60930a );
 a60941a <=( (not A167)  and  (not A169) );
 a60944a <=( A200  and  (not A166) );
 a60945a <=( a60944a  and  a60941a );
 a60948a <=( A232  and  A201 );
 a60951a <=( (not A234)  and  A233 );
 a60952a <=( a60951a  and  a60948a );
 a60953a <=( a60952a  and  a60945a );
 a60956a <=( A265  and  (not A235) );
 a60959a <=( (not A267)  and  A266 );
 a60960a <=( a60959a  and  a60956a );
 a60963a <=( (not A298)  and  (not A268) );
 a60966a <=( A302  and  A299 );
 a60967a <=( a60966a  and  a60963a );
 a60968a <=( a60967a  and  a60960a );
 a60971a <=( (not A167)  and  (not A169) );
 a60974a <=( (not A199)  and  (not A166) );
 a60975a <=( a60974a  and  a60971a );
 a60978a <=( A203  and  A200 );
 a60981a <=( (not A235)  and  (not A234) );
 a60982a <=( a60981a  and  a60978a );
 a60983a <=( a60982a  and  a60975a );
 a60986a <=( A265  and  (not A236) );
 a60989a <=( (not A267)  and  A266 );
 a60990a <=( a60989a  and  a60986a );
 a60993a <=( A298  and  (not A268) );
 a60996a <=( A302  and  (not A299) );
 a60997a <=( a60996a  and  a60993a );
 a60998a <=( a60997a  and  a60990a );
 a61001a <=( (not A167)  and  (not A169) );
 a61004a <=( (not A199)  and  (not A166) );
 a61005a <=( a61004a  and  a61001a );
 a61008a <=( A203  and  A200 );
 a61011a <=( (not A235)  and  (not A234) );
 a61012a <=( a61011a  and  a61008a );
 a61013a <=( a61012a  and  a61005a );
 a61016a <=( A265  and  (not A236) );
 a61019a <=( (not A267)  and  A266 );
 a61020a <=( a61019a  and  a61016a );
 a61023a <=( (not A298)  and  (not A268) );
 a61026a <=( A302  and  A299 );
 a61027a <=( a61026a  and  a61023a );
 a61028a <=( a61027a  and  a61020a );
 a61031a <=( (not A167)  and  (not A169) );
 a61034a <=( (not A199)  and  (not A166) );
 a61035a <=( a61034a  and  a61031a );
 a61038a <=( A203  and  A200 );
 a61041a <=( A233  and  A232 );
 a61042a <=( a61041a  and  a61038a );
 a61043a <=( a61042a  and  a61035a );
 a61046a <=( (not A235)  and  (not A234) );
 a61049a <=( (not A268)  and  (not A267) );
 a61050a <=( a61049a  and  a61046a );
 a61053a <=( A298  and  (not A269) );
 a61056a <=( A302  and  (not A299) );
 a61057a <=( a61056a  and  a61053a );
 a61058a <=( a61057a  and  a61050a );
 a61061a <=( (not A167)  and  (not A169) );
 a61064a <=( (not A199)  and  (not A166) );
 a61065a <=( a61064a  and  a61061a );
 a61068a <=( A203  and  A200 );
 a61071a <=( A233  and  A232 );
 a61072a <=( a61071a  and  a61068a );
 a61073a <=( a61072a  and  a61065a );
 a61076a <=( (not A235)  and  (not A234) );
 a61079a <=( (not A268)  and  (not A267) );
 a61080a <=( a61079a  and  a61076a );
 a61083a <=( (not A298)  and  (not A269) );
 a61086a <=( A302  and  A299 );
 a61087a <=( a61086a  and  a61083a );
 a61088a <=( a61087a  and  a61080a );
 a61091a <=( (not A167)  and  (not A169) );
 a61094a <=( (not A199)  and  (not A166) );
 a61095a <=( a61094a  and  a61091a );
 a61098a <=( A203  and  A200 );
 a61101a <=( A233  and  A232 );
 a61102a <=( a61101a  and  a61098a );
 a61103a <=( a61102a  and  a61095a );
 a61106a <=( (not A235)  and  (not A234) );
 a61109a <=( A266  and  A265 );
 a61110a <=( a61109a  and  a61106a );
 a61113a <=( (not A268)  and  (not A267) );
 a61116a <=( A300  and  A299 );
 a61117a <=( a61116a  and  a61113a );
 a61118a <=( a61117a  and  a61110a );
 a61121a <=( (not A167)  and  (not A169) );
 a61124a <=( (not A199)  and  (not A166) );
 a61125a <=( a61124a  and  a61121a );
 a61128a <=( A203  and  A200 );
 a61131a <=( A233  and  A232 );
 a61132a <=( a61131a  and  a61128a );
 a61133a <=( a61132a  and  a61125a );
 a61136a <=( (not A235)  and  (not A234) );
 a61139a <=( A266  and  A265 );
 a61140a <=( a61139a  and  a61136a );
 a61143a <=( (not A268)  and  (not A267) );
 a61146a <=( A300  and  A298 );
 a61147a <=( a61146a  and  a61143a );
 a61148a <=( a61147a  and  a61140a );
 a61151a <=( (not A167)  and  (not A169) );
 a61154a <=( (not A199)  and  (not A166) );
 a61155a <=( a61154a  and  a61151a );
 a61158a <=( A203  and  A200 );
 a61161a <=( A233  and  A232 );
 a61162a <=( a61161a  and  a61158a );
 a61163a <=( a61162a  and  a61155a );
 a61166a <=( (not A235)  and  (not A234) );
 a61169a <=( (not A266)  and  (not A265) );
 a61170a <=( a61169a  and  a61166a );
 a61173a <=( A298  and  (not A268) );
 a61176a <=( A302  and  (not A299) );
 a61177a <=( a61176a  and  a61173a );
 a61178a <=( a61177a  and  a61170a );
 a61181a <=( (not A167)  and  (not A169) );
 a61184a <=( (not A199)  and  (not A166) );
 a61185a <=( a61184a  and  a61181a );
 a61188a <=( A203  and  A200 );
 a61191a <=( A233  and  A232 );
 a61192a <=( a61191a  and  a61188a );
 a61193a <=( a61192a  and  a61185a );
 a61196a <=( (not A235)  and  (not A234) );
 a61199a <=( (not A266)  and  (not A265) );
 a61200a <=( a61199a  and  a61196a );
 a61203a <=( (not A298)  and  (not A268) );
 a61206a <=( A302  and  A299 );
 a61207a <=( a61206a  and  a61203a );
 a61208a <=( a61207a  and  a61200a );
 a61211a <=( (not A167)  and  (not A169) );
 a61214a <=( (not A199)  and  (not A166) );
 a61215a <=( a61214a  and  a61211a );
 a61218a <=( A203  and  A200 );
 a61221a <=( (not A233)  and  (not A232) );
 a61222a <=( a61221a  and  a61218a );
 a61223a <=( a61222a  and  a61215a );
 a61226a <=( A265  and  (not A235) );
 a61229a <=( (not A267)  and  A266 );
 a61230a <=( a61229a  and  a61226a );
 a61233a <=( A298  and  (not A268) );
 a61236a <=( A302  and  (not A299) );
 a61237a <=( a61236a  and  a61233a );
 a61238a <=( a61237a  and  a61230a );
 a61241a <=( (not A167)  and  (not A169) );
 a61244a <=( (not A199)  and  (not A166) );
 a61245a <=( a61244a  and  a61241a );
 a61248a <=( A203  and  A200 );
 a61251a <=( (not A233)  and  (not A232) );
 a61252a <=( a61251a  and  a61248a );
 a61253a <=( a61252a  and  a61245a );
 a61256a <=( A265  and  (not A235) );
 a61259a <=( (not A267)  and  A266 );
 a61260a <=( a61259a  and  a61256a );
 a61263a <=( (not A298)  and  (not A268) );
 a61266a <=( A302  and  A299 );
 a61267a <=( a61266a  and  a61263a );
 a61268a <=( a61267a  and  a61260a );
 a61271a <=( (not A167)  and  (not A169) );
 a61274a <=( A199  and  (not A166) );
 a61275a <=( a61274a  and  a61271a );
 a61278a <=( A203  and  (not A200) );
 a61281a <=( (not A235)  and  (not A234) );
 a61282a <=( a61281a  and  a61278a );
 a61283a <=( a61282a  and  a61275a );
 a61286a <=( A265  and  (not A236) );
 a61289a <=( (not A267)  and  A266 );
 a61290a <=( a61289a  and  a61286a );
 a61293a <=( A298  and  (not A268) );
 a61296a <=( A302  and  (not A299) );
 a61297a <=( a61296a  and  a61293a );
 a61298a <=( a61297a  and  a61290a );
 a61301a <=( (not A167)  and  (not A169) );
 a61304a <=( A199  and  (not A166) );
 a61305a <=( a61304a  and  a61301a );
 a61308a <=( A203  and  (not A200) );
 a61311a <=( (not A235)  and  (not A234) );
 a61312a <=( a61311a  and  a61308a );
 a61313a <=( a61312a  and  a61305a );
 a61316a <=( A265  and  (not A236) );
 a61319a <=( (not A267)  and  A266 );
 a61320a <=( a61319a  and  a61316a );
 a61323a <=( (not A298)  and  (not A268) );
 a61326a <=( A302  and  A299 );
 a61327a <=( a61326a  and  a61323a );
 a61328a <=( a61327a  and  a61320a );
 a61331a <=( (not A167)  and  (not A169) );
 a61334a <=( A199  and  (not A166) );
 a61335a <=( a61334a  and  a61331a );
 a61338a <=( A203  and  (not A200) );
 a61341a <=( A233  and  A232 );
 a61342a <=( a61341a  and  a61338a );
 a61343a <=( a61342a  and  a61335a );
 a61346a <=( (not A235)  and  (not A234) );
 a61349a <=( (not A268)  and  (not A267) );
 a61350a <=( a61349a  and  a61346a );
 a61353a <=( A298  and  (not A269) );
 a61356a <=( A302  and  (not A299) );
 a61357a <=( a61356a  and  a61353a );
 a61358a <=( a61357a  and  a61350a );
 a61361a <=( (not A167)  and  (not A169) );
 a61364a <=( A199  and  (not A166) );
 a61365a <=( a61364a  and  a61361a );
 a61368a <=( A203  and  (not A200) );
 a61371a <=( A233  and  A232 );
 a61372a <=( a61371a  and  a61368a );
 a61373a <=( a61372a  and  a61365a );
 a61376a <=( (not A235)  and  (not A234) );
 a61379a <=( (not A268)  and  (not A267) );
 a61380a <=( a61379a  and  a61376a );
 a61383a <=( (not A298)  and  (not A269) );
 a61386a <=( A302  and  A299 );
 a61387a <=( a61386a  and  a61383a );
 a61388a <=( a61387a  and  a61380a );
 a61391a <=( (not A167)  and  (not A169) );
 a61394a <=( A199  and  (not A166) );
 a61395a <=( a61394a  and  a61391a );
 a61398a <=( A203  and  (not A200) );
 a61401a <=( A233  and  A232 );
 a61402a <=( a61401a  and  a61398a );
 a61403a <=( a61402a  and  a61395a );
 a61406a <=( (not A235)  and  (not A234) );
 a61409a <=( A266  and  A265 );
 a61410a <=( a61409a  and  a61406a );
 a61413a <=( (not A268)  and  (not A267) );
 a61416a <=( A300  and  A299 );
 a61417a <=( a61416a  and  a61413a );
 a61418a <=( a61417a  and  a61410a );
 a61421a <=( (not A167)  and  (not A169) );
 a61424a <=( A199  and  (not A166) );
 a61425a <=( a61424a  and  a61421a );
 a61428a <=( A203  and  (not A200) );
 a61431a <=( A233  and  A232 );
 a61432a <=( a61431a  and  a61428a );
 a61433a <=( a61432a  and  a61425a );
 a61436a <=( (not A235)  and  (not A234) );
 a61439a <=( A266  and  A265 );
 a61440a <=( a61439a  and  a61436a );
 a61443a <=( (not A268)  and  (not A267) );
 a61446a <=( A300  and  A298 );
 a61447a <=( a61446a  and  a61443a );
 a61448a <=( a61447a  and  a61440a );
 a61451a <=( (not A167)  and  (not A169) );
 a61454a <=( A199  and  (not A166) );
 a61455a <=( a61454a  and  a61451a );
 a61458a <=( A203  and  (not A200) );
 a61461a <=( A233  and  A232 );
 a61462a <=( a61461a  and  a61458a );
 a61463a <=( a61462a  and  a61455a );
 a61466a <=( (not A235)  and  (not A234) );
 a61469a <=( (not A266)  and  (not A265) );
 a61470a <=( a61469a  and  a61466a );
 a61473a <=( A298  and  (not A268) );
 a61476a <=( A302  and  (not A299) );
 a61477a <=( a61476a  and  a61473a );
 a61478a <=( a61477a  and  a61470a );
 a61481a <=( (not A167)  and  (not A169) );
 a61484a <=( A199  and  (not A166) );
 a61485a <=( a61484a  and  a61481a );
 a61488a <=( A203  and  (not A200) );
 a61491a <=( A233  and  A232 );
 a61492a <=( a61491a  and  a61488a );
 a61493a <=( a61492a  and  a61485a );
 a61496a <=( (not A235)  and  (not A234) );
 a61499a <=( (not A266)  and  (not A265) );
 a61500a <=( a61499a  and  a61496a );
 a61503a <=( (not A298)  and  (not A268) );
 a61506a <=( A302  and  A299 );
 a61507a <=( a61506a  and  a61503a );
 a61508a <=( a61507a  and  a61500a );
 a61511a <=( (not A167)  and  (not A169) );
 a61514a <=( A199  and  (not A166) );
 a61515a <=( a61514a  and  a61511a );
 a61518a <=( A203  and  (not A200) );
 a61521a <=( (not A233)  and  (not A232) );
 a61522a <=( a61521a  and  a61518a );
 a61523a <=( a61522a  and  a61515a );
 a61526a <=( A265  and  (not A235) );
 a61529a <=( (not A267)  and  A266 );
 a61530a <=( a61529a  and  a61526a );
 a61533a <=( A298  and  (not A268) );
 a61536a <=( A302  and  (not A299) );
 a61537a <=( a61536a  and  a61533a );
 a61538a <=( a61537a  and  a61530a );
 a61541a <=( (not A167)  and  (not A169) );
 a61544a <=( A199  and  (not A166) );
 a61545a <=( a61544a  and  a61541a );
 a61548a <=( A203  and  (not A200) );
 a61551a <=( (not A233)  and  (not A232) );
 a61552a <=( a61551a  and  a61548a );
 a61553a <=( a61552a  and  a61545a );
 a61556a <=( A265  and  (not A235) );
 a61559a <=( (not A267)  and  A266 );
 a61560a <=( a61559a  and  a61556a );
 a61563a <=( (not A298)  and  (not A268) );
 a61566a <=( A302  and  A299 );
 a61567a <=( a61566a  and  a61563a );
 a61568a <=( a61567a  and  a61560a );
 a61571a <=( (not A168)  and  (not A169) );
 a61574a <=( A166  and  A167 );
 a61575a <=( a61574a  and  a61571a );
 a61578a <=( A232  and  A202 );
 a61581a <=( (not A234)  and  A233 );
 a61582a <=( a61581a  and  a61578a );
 a61583a <=( a61582a  and  a61575a );
 a61586a <=( A265  and  (not A235) );
 a61589a <=( (not A267)  and  A266 );
 a61590a <=( a61589a  and  a61586a );
 a61593a <=( A298  and  (not A268) );
 a61596a <=( A302  and  (not A299) );
 a61597a <=( a61596a  and  a61593a );
 a61598a <=( a61597a  and  a61590a );
 a61601a <=( (not A168)  and  (not A169) );
 a61604a <=( A166  and  A167 );
 a61605a <=( a61604a  and  a61601a );
 a61608a <=( A232  and  A202 );
 a61611a <=( (not A234)  and  A233 );
 a61612a <=( a61611a  and  a61608a );
 a61613a <=( a61612a  and  a61605a );
 a61616a <=( A265  and  (not A235) );
 a61619a <=( (not A267)  and  A266 );
 a61620a <=( a61619a  and  a61616a );
 a61623a <=( (not A298)  and  (not A268) );
 a61626a <=( A302  and  A299 );
 a61627a <=( a61626a  and  a61623a );
 a61628a <=( a61627a  and  a61620a );
 a61631a <=( (not A168)  and  (not A169) );
 a61634a <=( A166  and  A167 );
 a61635a <=( a61634a  and  a61631a );
 a61638a <=( A201  and  A199 );
 a61641a <=( (not A235)  and  (not A234) );
 a61642a <=( a61641a  and  a61638a );
 a61643a <=( a61642a  and  a61635a );
 a61646a <=( A265  and  (not A236) );
 a61649a <=( (not A267)  and  A266 );
 a61650a <=( a61649a  and  a61646a );
 a61653a <=( A298  and  (not A268) );
 a61656a <=( A302  and  (not A299) );
 a61657a <=( a61656a  and  a61653a );
 a61658a <=( a61657a  and  a61650a );
 a61661a <=( (not A168)  and  (not A169) );
 a61664a <=( A166  and  A167 );
 a61665a <=( a61664a  and  a61661a );
 a61668a <=( A201  and  A199 );
 a61671a <=( (not A235)  and  (not A234) );
 a61672a <=( a61671a  and  a61668a );
 a61673a <=( a61672a  and  a61665a );
 a61676a <=( A265  and  (not A236) );
 a61679a <=( (not A267)  and  A266 );
 a61680a <=( a61679a  and  a61676a );
 a61683a <=( (not A298)  and  (not A268) );
 a61686a <=( A302  and  A299 );
 a61687a <=( a61686a  and  a61683a );
 a61688a <=( a61687a  and  a61680a );
 a61691a <=( (not A168)  and  (not A169) );
 a61694a <=( A166  and  A167 );
 a61695a <=( a61694a  and  a61691a );
 a61698a <=( A201  and  A199 );
 a61701a <=( A233  and  A232 );
 a61702a <=( a61701a  and  a61698a );
 a61703a <=( a61702a  and  a61695a );
 a61706a <=( (not A235)  and  (not A234) );
 a61709a <=( (not A268)  and  (not A267) );
 a61710a <=( a61709a  and  a61706a );
 a61713a <=( A298  and  (not A269) );
 a61716a <=( A302  and  (not A299) );
 a61717a <=( a61716a  and  a61713a );
 a61718a <=( a61717a  and  a61710a );
 a61721a <=( (not A168)  and  (not A169) );
 a61724a <=( A166  and  A167 );
 a61725a <=( a61724a  and  a61721a );
 a61728a <=( A201  and  A199 );
 a61731a <=( A233  and  A232 );
 a61732a <=( a61731a  and  a61728a );
 a61733a <=( a61732a  and  a61725a );
 a61736a <=( (not A235)  and  (not A234) );
 a61739a <=( (not A268)  and  (not A267) );
 a61740a <=( a61739a  and  a61736a );
 a61743a <=( (not A298)  and  (not A269) );
 a61746a <=( A302  and  A299 );
 a61747a <=( a61746a  and  a61743a );
 a61748a <=( a61747a  and  a61740a );
 a61751a <=( (not A168)  and  (not A169) );
 a61754a <=( A166  and  A167 );
 a61755a <=( a61754a  and  a61751a );
 a61758a <=( A201  and  A199 );
 a61761a <=( A233  and  A232 );
 a61762a <=( a61761a  and  a61758a );
 a61763a <=( a61762a  and  a61755a );
 a61766a <=( (not A235)  and  (not A234) );
 a61769a <=( A266  and  A265 );
 a61770a <=( a61769a  and  a61766a );
 a61773a <=( (not A268)  and  (not A267) );
 a61776a <=( A300  and  A299 );
 a61777a <=( a61776a  and  a61773a );
 a61778a <=( a61777a  and  a61770a );
 a61781a <=( (not A168)  and  (not A169) );
 a61784a <=( A166  and  A167 );
 a61785a <=( a61784a  and  a61781a );
 a61788a <=( A201  and  A199 );
 a61791a <=( A233  and  A232 );
 a61792a <=( a61791a  and  a61788a );
 a61793a <=( a61792a  and  a61785a );
 a61796a <=( (not A235)  and  (not A234) );
 a61799a <=( A266  and  A265 );
 a61800a <=( a61799a  and  a61796a );
 a61803a <=( (not A268)  and  (not A267) );
 a61806a <=( A300  and  A298 );
 a61807a <=( a61806a  and  a61803a );
 a61808a <=( a61807a  and  a61800a );
 a61811a <=( (not A168)  and  (not A169) );
 a61814a <=( A166  and  A167 );
 a61815a <=( a61814a  and  a61811a );
 a61818a <=( A201  and  A199 );
 a61821a <=( A233  and  A232 );
 a61822a <=( a61821a  and  a61818a );
 a61823a <=( a61822a  and  a61815a );
 a61826a <=( (not A235)  and  (not A234) );
 a61829a <=( (not A266)  and  (not A265) );
 a61830a <=( a61829a  and  a61826a );
 a61833a <=( A298  and  (not A268) );
 a61836a <=( A302  and  (not A299) );
 a61837a <=( a61836a  and  a61833a );
 a61838a <=( a61837a  and  a61830a );
 a61841a <=( (not A168)  and  (not A169) );
 a61844a <=( A166  and  A167 );
 a61845a <=( a61844a  and  a61841a );
 a61848a <=( A201  and  A199 );
 a61851a <=( A233  and  A232 );
 a61852a <=( a61851a  and  a61848a );
 a61853a <=( a61852a  and  a61845a );
 a61856a <=( (not A235)  and  (not A234) );
 a61859a <=( (not A266)  and  (not A265) );
 a61860a <=( a61859a  and  a61856a );
 a61863a <=( (not A298)  and  (not A268) );
 a61866a <=( A302  and  A299 );
 a61867a <=( a61866a  and  a61863a );
 a61868a <=( a61867a  and  a61860a );
 a61871a <=( (not A168)  and  (not A169) );
 a61874a <=( A166  and  A167 );
 a61875a <=( a61874a  and  a61871a );
 a61878a <=( A201  and  A199 );
 a61881a <=( (not A233)  and  (not A232) );
 a61882a <=( a61881a  and  a61878a );
 a61883a <=( a61882a  and  a61875a );
 a61886a <=( A265  and  (not A235) );
 a61889a <=( (not A267)  and  A266 );
 a61890a <=( a61889a  and  a61886a );
 a61893a <=( A298  and  (not A268) );
 a61896a <=( A302  and  (not A299) );
 a61897a <=( a61896a  and  a61893a );
 a61898a <=( a61897a  and  a61890a );
 a61901a <=( (not A168)  and  (not A169) );
 a61904a <=( A166  and  A167 );
 a61905a <=( a61904a  and  a61901a );
 a61908a <=( A201  and  A199 );
 a61911a <=( (not A233)  and  (not A232) );
 a61912a <=( a61911a  and  a61908a );
 a61913a <=( a61912a  and  a61905a );
 a61916a <=( A265  and  (not A235) );
 a61919a <=( (not A267)  and  A266 );
 a61920a <=( a61919a  and  a61916a );
 a61923a <=( (not A298)  and  (not A268) );
 a61926a <=( A302  and  A299 );
 a61927a <=( a61926a  and  a61923a );
 a61928a <=( a61927a  and  a61920a );
 a61931a <=( (not A168)  and  (not A169) );
 a61934a <=( A166  and  A167 );
 a61935a <=( a61934a  and  a61931a );
 a61938a <=( A201  and  A200 );
 a61941a <=( (not A235)  and  (not A234) );
 a61942a <=( a61941a  and  a61938a );
 a61943a <=( a61942a  and  a61935a );
 a61946a <=( A265  and  (not A236) );
 a61949a <=( (not A267)  and  A266 );
 a61950a <=( a61949a  and  a61946a );
 a61953a <=( A298  and  (not A268) );
 a61956a <=( A302  and  (not A299) );
 a61957a <=( a61956a  and  a61953a );
 a61958a <=( a61957a  and  a61950a );
 a61961a <=( (not A168)  and  (not A169) );
 a61964a <=( A166  and  A167 );
 a61965a <=( a61964a  and  a61961a );
 a61968a <=( A201  and  A200 );
 a61971a <=( (not A235)  and  (not A234) );
 a61972a <=( a61971a  and  a61968a );
 a61973a <=( a61972a  and  a61965a );
 a61976a <=( A265  and  (not A236) );
 a61979a <=( (not A267)  and  A266 );
 a61980a <=( a61979a  and  a61976a );
 a61983a <=( (not A298)  and  (not A268) );
 a61986a <=( A302  and  A299 );
 a61987a <=( a61986a  and  a61983a );
 a61988a <=( a61987a  and  a61980a );
 a61991a <=( (not A168)  and  (not A169) );
 a61994a <=( A166  and  A167 );
 a61995a <=( a61994a  and  a61991a );
 a61998a <=( A201  and  A200 );
 a62001a <=( A233  and  A232 );
 a62002a <=( a62001a  and  a61998a );
 a62003a <=( a62002a  and  a61995a );
 a62006a <=( (not A235)  and  (not A234) );
 a62009a <=( (not A268)  and  (not A267) );
 a62010a <=( a62009a  and  a62006a );
 a62013a <=( A298  and  (not A269) );
 a62016a <=( A302  and  (not A299) );
 a62017a <=( a62016a  and  a62013a );
 a62018a <=( a62017a  and  a62010a );
 a62021a <=( (not A168)  and  (not A169) );
 a62024a <=( A166  and  A167 );
 a62025a <=( a62024a  and  a62021a );
 a62028a <=( A201  and  A200 );
 a62031a <=( A233  and  A232 );
 a62032a <=( a62031a  and  a62028a );
 a62033a <=( a62032a  and  a62025a );
 a62036a <=( (not A235)  and  (not A234) );
 a62039a <=( (not A268)  and  (not A267) );
 a62040a <=( a62039a  and  a62036a );
 a62043a <=( (not A298)  and  (not A269) );
 a62046a <=( A302  and  A299 );
 a62047a <=( a62046a  and  a62043a );
 a62048a <=( a62047a  and  a62040a );
 a62051a <=( (not A168)  and  (not A169) );
 a62054a <=( A166  and  A167 );
 a62055a <=( a62054a  and  a62051a );
 a62058a <=( A201  and  A200 );
 a62061a <=( A233  and  A232 );
 a62062a <=( a62061a  and  a62058a );
 a62063a <=( a62062a  and  a62055a );
 a62066a <=( (not A235)  and  (not A234) );
 a62069a <=( A266  and  A265 );
 a62070a <=( a62069a  and  a62066a );
 a62073a <=( (not A268)  and  (not A267) );
 a62076a <=( A300  and  A299 );
 a62077a <=( a62076a  and  a62073a );
 a62078a <=( a62077a  and  a62070a );
 a62081a <=( (not A168)  and  (not A169) );
 a62084a <=( A166  and  A167 );
 a62085a <=( a62084a  and  a62081a );
 a62088a <=( A201  and  A200 );
 a62091a <=( A233  and  A232 );
 a62092a <=( a62091a  and  a62088a );
 a62093a <=( a62092a  and  a62085a );
 a62096a <=( (not A235)  and  (not A234) );
 a62099a <=( A266  and  A265 );
 a62100a <=( a62099a  and  a62096a );
 a62103a <=( (not A268)  and  (not A267) );
 a62106a <=( A300  and  A298 );
 a62107a <=( a62106a  and  a62103a );
 a62108a <=( a62107a  and  a62100a );
 a62111a <=( (not A168)  and  (not A169) );
 a62114a <=( A166  and  A167 );
 a62115a <=( a62114a  and  a62111a );
 a62118a <=( A201  and  A200 );
 a62121a <=( A233  and  A232 );
 a62122a <=( a62121a  and  a62118a );
 a62123a <=( a62122a  and  a62115a );
 a62126a <=( (not A235)  and  (not A234) );
 a62129a <=( (not A266)  and  (not A265) );
 a62130a <=( a62129a  and  a62126a );
 a62133a <=( A298  and  (not A268) );
 a62136a <=( A302  and  (not A299) );
 a62137a <=( a62136a  and  a62133a );
 a62138a <=( a62137a  and  a62130a );
 a62141a <=( (not A168)  and  (not A169) );
 a62144a <=( A166  and  A167 );
 a62145a <=( a62144a  and  a62141a );
 a62148a <=( A201  and  A200 );
 a62151a <=( A233  and  A232 );
 a62152a <=( a62151a  and  a62148a );
 a62153a <=( a62152a  and  a62145a );
 a62156a <=( (not A235)  and  (not A234) );
 a62159a <=( (not A266)  and  (not A265) );
 a62160a <=( a62159a  and  a62156a );
 a62163a <=( (not A298)  and  (not A268) );
 a62166a <=( A302  and  A299 );
 a62167a <=( a62166a  and  a62163a );
 a62168a <=( a62167a  and  a62160a );
 a62171a <=( (not A168)  and  (not A169) );
 a62174a <=( A166  and  A167 );
 a62175a <=( a62174a  and  a62171a );
 a62178a <=( A201  and  A200 );
 a62181a <=( (not A233)  and  (not A232) );
 a62182a <=( a62181a  and  a62178a );
 a62183a <=( a62182a  and  a62175a );
 a62186a <=( A265  and  (not A235) );
 a62189a <=( (not A267)  and  A266 );
 a62190a <=( a62189a  and  a62186a );
 a62193a <=( A298  and  (not A268) );
 a62196a <=( A302  and  (not A299) );
 a62197a <=( a62196a  and  a62193a );
 a62198a <=( a62197a  and  a62190a );
 a62201a <=( (not A168)  and  (not A169) );
 a62204a <=( A166  and  A167 );
 a62205a <=( a62204a  and  a62201a );
 a62208a <=( A201  and  A200 );
 a62211a <=( (not A233)  and  (not A232) );
 a62212a <=( a62211a  and  a62208a );
 a62213a <=( a62212a  and  a62205a );
 a62216a <=( A265  and  (not A235) );
 a62219a <=( (not A267)  and  A266 );
 a62220a <=( a62219a  and  a62216a );
 a62223a <=( (not A298)  and  (not A268) );
 a62226a <=( A302  and  A299 );
 a62227a <=( a62226a  and  a62223a );
 a62228a <=( a62227a  and  a62220a );
 a62231a <=( (not A168)  and  (not A169) );
 a62234a <=( A166  and  A167 );
 a62235a <=( a62234a  and  a62231a );
 a62238a <=( A200  and  (not A199) );
 a62241a <=( (not A234)  and  A203 );
 a62242a <=( a62241a  and  a62238a );
 a62243a <=( a62242a  and  a62235a );
 a62246a <=( (not A236)  and  (not A235) );
 a62249a <=( (not A268)  and  (not A267) );
 a62250a <=( a62249a  and  a62246a );
 a62253a <=( A298  and  (not A269) );
 a62256a <=( A302  and  (not A299) );
 a62257a <=( a62256a  and  a62253a );
 a62258a <=( a62257a  and  a62250a );
 a62261a <=( (not A168)  and  (not A169) );
 a62264a <=( A166  and  A167 );
 a62265a <=( a62264a  and  a62261a );
 a62268a <=( A200  and  (not A199) );
 a62271a <=( (not A234)  and  A203 );
 a62272a <=( a62271a  and  a62268a );
 a62273a <=( a62272a  and  a62265a );
 a62276a <=( (not A236)  and  (not A235) );
 a62279a <=( (not A268)  and  (not A267) );
 a62280a <=( a62279a  and  a62276a );
 a62283a <=( (not A298)  and  (not A269) );
 a62286a <=( A302  and  A299 );
 a62287a <=( a62286a  and  a62283a );
 a62288a <=( a62287a  and  a62280a );
 a62291a <=( (not A168)  and  (not A169) );
 a62294a <=( A166  and  A167 );
 a62295a <=( a62294a  and  a62291a );
 a62298a <=( A200  and  (not A199) );
 a62301a <=( (not A234)  and  A203 );
 a62302a <=( a62301a  and  a62298a );
 a62303a <=( a62302a  and  a62295a );
 a62306a <=( (not A236)  and  (not A235) );
 a62309a <=( A266  and  A265 );
 a62310a <=( a62309a  and  a62306a );
 a62313a <=( (not A268)  and  (not A267) );
 a62316a <=( A300  and  A299 );
 a62317a <=( a62316a  and  a62313a );
 a62318a <=( a62317a  and  a62310a );
 a62321a <=( (not A168)  and  (not A169) );
 a62324a <=( A166  and  A167 );
 a62325a <=( a62324a  and  a62321a );
 a62328a <=( A200  and  (not A199) );
 a62331a <=( (not A234)  and  A203 );
 a62332a <=( a62331a  and  a62328a );
 a62333a <=( a62332a  and  a62325a );
 a62336a <=( (not A236)  and  (not A235) );
 a62339a <=( A266  and  A265 );
 a62340a <=( a62339a  and  a62336a );
 a62343a <=( (not A268)  and  (not A267) );
 a62346a <=( A300  and  A298 );
 a62347a <=( a62346a  and  a62343a );
 a62348a <=( a62347a  and  a62340a );
 a62351a <=( (not A168)  and  (not A169) );
 a62354a <=( A166  and  A167 );
 a62355a <=( a62354a  and  a62351a );
 a62358a <=( A200  and  (not A199) );
 a62361a <=( (not A234)  and  A203 );
 a62362a <=( a62361a  and  a62358a );
 a62363a <=( a62362a  and  a62355a );
 a62366a <=( (not A236)  and  (not A235) );
 a62369a <=( (not A266)  and  (not A265) );
 a62370a <=( a62369a  and  a62366a );
 a62373a <=( A298  and  (not A268) );
 a62376a <=( A302  and  (not A299) );
 a62377a <=( a62376a  and  a62373a );
 a62378a <=( a62377a  and  a62370a );
 a62381a <=( (not A168)  and  (not A169) );
 a62384a <=( A166  and  A167 );
 a62385a <=( a62384a  and  a62381a );
 a62388a <=( A200  and  (not A199) );
 a62391a <=( (not A234)  and  A203 );
 a62392a <=( a62391a  and  a62388a );
 a62393a <=( a62392a  and  a62385a );
 a62396a <=( (not A236)  and  (not A235) );
 a62399a <=( (not A266)  and  (not A265) );
 a62400a <=( a62399a  and  a62396a );
 a62403a <=( (not A298)  and  (not A268) );
 a62406a <=( A302  and  A299 );
 a62407a <=( a62406a  and  a62403a );
 a62408a <=( a62407a  and  a62400a );
 a62411a <=( (not A168)  and  (not A169) );
 a62414a <=( A166  and  A167 );
 a62415a <=( a62414a  and  a62411a );
 a62418a <=( A200  and  (not A199) );
 a62421a <=( A232  and  A203 );
 a62422a <=( a62421a  and  a62418a );
 a62423a <=( a62422a  and  a62415a );
 a62426a <=( (not A234)  and  A233 );
 a62429a <=( (not A267)  and  (not A235) );
 a62430a <=( a62429a  and  a62426a );
 a62433a <=( (not A269)  and  (not A268) );
 a62436a <=( A300  and  A299 );
 a62437a <=( a62436a  and  a62433a );
 a62438a <=( a62437a  and  a62430a );
 a62441a <=( (not A168)  and  (not A169) );
 a62444a <=( A166  and  A167 );
 a62445a <=( a62444a  and  a62441a );
 a62448a <=( A200  and  (not A199) );
 a62451a <=( A232  and  A203 );
 a62452a <=( a62451a  and  a62448a );
 a62453a <=( a62452a  and  a62445a );
 a62456a <=( (not A234)  and  A233 );
 a62459a <=( (not A267)  and  (not A235) );
 a62460a <=( a62459a  and  a62456a );
 a62463a <=( (not A269)  and  (not A268) );
 a62466a <=( A300  and  A298 );
 a62467a <=( a62466a  and  a62463a );
 a62468a <=( a62467a  and  a62460a );
 a62471a <=( (not A168)  and  (not A169) );
 a62474a <=( A166  and  A167 );
 a62475a <=( a62474a  and  a62471a );
 a62478a <=( A200  and  (not A199) );
 a62481a <=( A232  and  A203 );
 a62482a <=( a62481a  and  a62478a );
 a62483a <=( a62482a  and  a62475a );
 a62486a <=( (not A234)  and  A233 );
 a62489a <=( A265  and  (not A235) );
 a62490a <=( a62489a  and  a62486a );
 a62493a <=( (not A267)  and  A266 );
 a62496a <=( A301  and  (not A268) );
 a62497a <=( a62496a  and  a62493a );
 a62498a <=( a62497a  and  a62490a );
 a62501a <=( (not A168)  and  (not A169) );
 a62504a <=( A166  and  A167 );
 a62505a <=( a62504a  and  a62501a );
 a62508a <=( A200  and  (not A199) );
 a62511a <=( A232  and  A203 );
 a62512a <=( a62511a  and  a62508a );
 a62513a <=( a62512a  and  a62505a );
 a62516a <=( (not A234)  and  A233 );
 a62519a <=( (not A265)  and  (not A235) );
 a62520a <=( a62519a  and  a62516a );
 a62523a <=( (not A268)  and  (not A266) );
 a62526a <=( A300  and  A299 );
 a62527a <=( a62526a  and  a62523a );
 a62528a <=( a62527a  and  a62520a );
 a62531a <=( (not A168)  and  (not A169) );
 a62534a <=( A166  and  A167 );
 a62535a <=( a62534a  and  a62531a );
 a62538a <=( A200  and  (not A199) );
 a62541a <=( A232  and  A203 );
 a62542a <=( a62541a  and  a62538a );
 a62543a <=( a62542a  and  a62535a );
 a62546a <=( (not A234)  and  A233 );
 a62549a <=( (not A265)  and  (not A235) );
 a62550a <=( a62549a  and  a62546a );
 a62553a <=( (not A268)  and  (not A266) );
 a62556a <=( A300  and  A298 );
 a62557a <=( a62556a  and  a62553a );
 a62558a <=( a62557a  and  a62550a );
 a62561a <=( (not A168)  and  (not A169) );
 a62564a <=( A166  and  A167 );
 a62565a <=( a62564a  and  a62561a );
 a62568a <=( A200  and  (not A199) );
 a62571a <=( (not A232)  and  A203 );
 a62572a <=( a62571a  and  a62568a );
 a62573a <=( a62572a  and  a62565a );
 a62576a <=( (not A235)  and  (not A233) );
 a62579a <=( (not A268)  and  (not A267) );
 a62580a <=( a62579a  and  a62576a );
 a62583a <=( A298  and  (not A269) );
 a62586a <=( A302  and  (not A299) );
 a62587a <=( a62586a  and  a62583a );
 a62588a <=( a62587a  and  a62580a );
 a62591a <=( (not A168)  and  (not A169) );
 a62594a <=( A166  and  A167 );
 a62595a <=( a62594a  and  a62591a );
 a62598a <=( A200  and  (not A199) );
 a62601a <=( (not A232)  and  A203 );
 a62602a <=( a62601a  and  a62598a );
 a62603a <=( a62602a  and  a62595a );
 a62606a <=( (not A235)  and  (not A233) );
 a62609a <=( (not A268)  and  (not A267) );
 a62610a <=( a62609a  and  a62606a );
 a62613a <=( (not A298)  and  (not A269) );
 a62616a <=( A302  and  A299 );
 a62617a <=( a62616a  and  a62613a );
 a62618a <=( a62617a  and  a62610a );
 a62621a <=( (not A168)  and  (not A169) );
 a62624a <=( A166  and  A167 );
 a62625a <=( a62624a  and  a62621a );
 a62628a <=( A200  and  (not A199) );
 a62631a <=( (not A232)  and  A203 );
 a62632a <=( a62631a  and  a62628a );
 a62633a <=( a62632a  and  a62625a );
 a62636a <=( (not A235)  and  (not A233) );
 a62639a <=( A266  and  A265 );
 a62640a <=( a62639a  and  a62636a );
 a62643a <=( (not A268)  and  (not A267) );
 a62646a <=( A300  and  A299 );
 a62647a <=( a62646a  and  a62643a );
 a62648a <=( a62647a  and  a62640a );
 a62651a <=( (not A168)  and  (not A169) );
 a62654a <=( A166  and  A167 );
 a62655a <=( a62654a  and  a62651a );
 a62658a <=( A200  and  (not A199) );
 a62661a <=( (not A232)  and  A203 );
 a62662a <=( a62661a  and  a62658a );
 a62663a <=( a62662a  and  a62655a );
 a62666a <=( (not A235)  and  (not A233) );
 a62669a <=( A266  and  A265 );
 a62670a <=( a62669a  and  a62666a );
 a62673a <=( (not A268)  and  (not A267) );
 a62676a <=( A300  and  A298 );
 a62677a <=( a62676a  and  a62673a );
 a62678a <=( a62677a  and  a62670a );
 a62681a <=( (not A168)  and  (not A169) );
 a62684a <=( A166  and  A167 );
 a62685a <=( a62684a  and  a62681a );
 a62688a <=( A200  and  (not A199) );
 a62691a <=( (not A232)  and  A203 );
 a62692a <=( a62691a  and  a62688a );
 a62693a <=( a62692a  and  a62685a );
 a62696a <=( (not A235)  and  (not A233) );
 a62699a <=( (not A266)  and  (not A265) );
 a62700a <=( a62699a  and  a62696a );
 a62703a <=( A298  and  (not A268) );
 a62706a <=( A302  and  (not A299) );
 a62707a <=( a62706a  and  a62703a );
 a62708a <=( a62707a  and  a62700a );
 a62711a <=( (not A168)  and  (not A169) );
 a62714a <=( A166  and  A167 );
 a62715a <=( a62714a  and  a62711a );
 a62718a <=( A200  and  (not A199) );
 a62721a <=( (not A232)  and  A203 );
 a62722a <=( a62721a  and  a62718a );
 a62723a <=( a62722a  and  a62715a );
 a62726a <=( (not A235)  and  (not A233) );
 a62729a <=( (not A266)  and  (not A265) );
 a62730a <=( a62729a  and  a62726a );
 a62733a <=( (not A298)  and  (not A268) );
 a62736a <=( A302  and  A299 );
 a62737a <=( a62736a  and  a62733a );
 a62738a <=( a62737a  and  a62730a );
 a62741a <=( (not A168)  and  (not A169) );
 a62744a <=( A166  and  A167 );
 a62745a <=( a62744a  and  a62741a );
 a62748a <=( (not A200)  and  A199 );
 a62751a <=( (not A234)  and  A203 );
 a62752a <=( a62751a  and  a62748a );
 a62753a <=( a62752a  and  a62745a );
 a62756a <=( (not A236)  and  (not A235) );
 a62759a <=( (not A268)  and  (not A267) );
 a62760a <=( a62759a  and  a62756a );
 a62763a <=( A298  and  (not A269) );
 a62766a <=( A302  and  (not A299) );
 a62767a <=( a62766a  and  a62763a );
 a62768a <=( a62767a  and  a62760a );
 a62771a <=( (not A168)  and  (not A169) );
 a62774a <=( A166  and  A167 );
 a62775a <=( a62774a  and  a62771a );
 a62778a <=( (not A200)  and  A199 );
 a62781a <=( (not A234)  and  A203 );
 a62782a <=( a62781a  and  a62778a );
 a62783a <=( a62782a  and  a62775a );
 a62786a <=( (not A236)  and  (not A235) );
 a62789a <=( (not A268)  and  (not A267) );
 a62790a <=( a62789a  and  a62786a );
 a62793a <=( (not A298)  and  (not A269) );
 a62796a <=( A302  and  A299 );
 a62797a <=( a62796a  and  a62793a );
 a62798a <=( a62797a  and  a62790a );
 a62801a <=( (not A168)  and  (not A169) );
 a62804a <=( A166  and  A167 );
 a62805a <=( a62804a  and  a62801a );
 a62808a <=( (not A200)  and  A199 );
 a62811a <=( (not A234)  and  A203 );
 a62812a <=( a62811a  and  a62808a );
 a62813a <=( a62812a  and  a62805a );
 a62816a <=( (not A236)  and  (not A235) );
 a62819a <=( A266  and  A265 );
 a62820a <=( a62819a  and  a62816a );
 a62823a <=( (not A268)  and  (not A267) );
 a62826a <=( A300  and  A299 );
 a62827a <=( a62826a  and  a62823a );
 a62828a <=( a62827a  and  a62820a );
 a62831a <=( (not A168)  and  (not A169) );
 a62834a <=( A166  and  A167 );
 a62835a <=( a62834a  and  a62831a );
 a62838a <=( (not A200)  and  A199 );
 a62841a <=( (not A234)  and  A203 );
 a62842a <=( a62841a  and  a62838a );
 a62843a <=( a62842a  and  a62835a );
 a62846a <=( (not A236)  and  (not A235) );
 a62849a <=( A266  and  A265 );
 a62850a <=( a62849a  and  a62846a );
 a62853a <=( (not A268)  and  (not A267) );
 a62856a <=( A300  and  A298 );
 a62857a <=( a62856a  and  a62853a );
 a62858a <=( a62857a  and  a62850a );
 a62861a <=( (not A168)  and  (not A169) );
 a62864a <=( A166  and  A167 );
 a62865a <=( a62864a  and  a62861a );
 a62868a <=( (not A200)  and  A199 );
 a62871a <=( (not A234)  and  A203 );
 a62872a <=( a62871a  and  a62868a );
 a62873a <=( a62872a  and  a62865a );
 a62876a <=( (not A236)  and  (not A235) );
 a62879a <=( (not A266)  and  (not A265) );
 a62880a <=( a62879a  and  a62876a );
 a62883a <=( A298  and  (not A268) );
 a62886a <=( A302  and  (not A299) );
 a62887a <=( a62886a  and  a62883a );
 a62888a <=( a62887a  and  a62880a );
 a62891a <=( (not A168)  and  (not A169) );
 a62894a <=( A166  and  A167 );
 a62895a <=( a62894a  and  a62891a );
 a62898a <=( (not A200)  and  A199 );
 a62901a <=( (not A234)  and  A203 );
 a62902a <=( a62901a  and  a62898a );
 a62903a <=( a62902a  and  a62895a );
 a62906a <=( (not A236)  and  (not A235) );
 a62909a <=( (not A266)  and  (not A265) );
 a62910a <=( a62909a  and  a62906a );
 a62913a <=( (not A298)  and  (not A268) );
 a62916a <=( A302  and  A299 );
 a62917a <=( a62916a  and  a62913a );
 a62918a <=( a62917a  and  a62910a );
 a62921a <=( (not A168)  and  (not A169) );
 a62924a <=( A166  and  A167 );
 a62925a <=( a62924a  and  a62921a );
 a62928a <=( (not A200)  and  A199 );
 a62931a <=( A232  and  A203 );
 a62932a <=( a62931a  and  a62928a );
 a62933a <=( a62932a  and  a62925a );
 a62936a <=( (not A234)  and  A233 );
 a62939a <=( (not A267)  and  (not A235) );
 a62940a <=( a62939a  and  a62936a );
 a62943a <=( (not A269)  and  (not A268) );
 a62946a <=( A300  and  A299 );
 a62947a <=( a62946a  and  a62943a );
 a62948a <=( a62947a  and  a62940a );
 a62951a <=( (not A168)  and  (not A169) );
 a62954a <=( A166  and  A167 );
 a62955a <=( a62954a  and  a62951a );
 a62958a <=( (not A200)  and  A199 );
 a62961a <=( A232  and  A203 );
 a62962a <=( a62961a  and  a62958a );
 a62963a <=( a62962a  and  a62955a );
 a62966a <=( (not A234)  and  A233 );
 a62969a <=( (not A267)  and  (not A235) );
 a62970a <=( a62969a  and  a62966a );
 a62973a <=( (not A269)  and  (not A268) );
 a62976a <=( A300  and  A298 );
 a62977a <=( a62976a  and  a62973a );
 a62978a <=( a62977a  and  a62970a );
 a62981a <=( (not A168)  and  (not A169) );
 a62984a <=( A166  and  A167 );
 a62985a <=( a62984a  and  a62981a );
 a62988a <=( (not A200)  and  A199 );
 a62991a <=( A232  and  A203 );
 a62992a <=( a62991a  and  a62988a );
 a62993a <=( a62992a  and  a62985a );
 a62996a <=( (not A234)  and  A233 );
 a62999a <=( A265  and  (not A235) );
 a63000a <=( a62999a  and  a62996a );
 a63003a <=( (not A267)  and  A266 );
 a63006a <=( A301  and  (not A268) );
 a63007a <=( a63006a  and  a63003a );
 a63008a <=( a63007a  and  a63000a );
 a63011a <=( (not A168)  and  (not A169) );
 a63014a <=( A166  and  A167 );
 a63015a <=( a63014a  and  a63011a );
 a63018a <=( (not A200)  and  A199 );
 a63021a <=( A232  and  A203 );
 a63022a <=( a63021a  and  a63018a );
 a63023a <=( a63022a  and  a63015a );
 a63026a <=( (not A234)  and  A233 );
 a63029a <=( (not A265)  and  (not A235) );
 a63030a <=( a63029a  and  a63026a );
 a63033a <=( (not A268)  and  (not A266) );
 a63036a <=( A300  and  A299 );
 a63037a <=( a63036a  and  a63033a );
 a63038a <=( a63037a  and  a63030a );
 a63041a <=( (not A168)  and  (not A169) );
 a63044a <=( A166  and  A167 );
 a63045a <=( a63044a  and  a63041a );
 a63048a <=( (not A200)  and  A199 );
 a63051a <=( A232  and  A203 );
 a63052a <=( a63051a  and  a63048a );
 a63053a <=( a63052a  and  a63045a );
 a63056a <=( (not A234)  and  A233 );
 a63059a <=( (not A265)  and  (not A235) );
 a63060a <=( a63059a  and  a63056a );
 a63063a <=( (not A268)  and  (not A266) );
 a63066a <=( A300  and  A298 );
 a63067a <=( a63066a  and  a63063a );
 a63068a <=( a63067a  and  a63060a );
 a63071a <=( (not A168)  and  (not A169) );
 a63074a <=( A166  and  A167 );
 a63075a <=( a63074a  and  a63071a );
 a63078a <=( (not A200)  and  A199 );
 a63081a <=( (not A232)  and  A203 );
 a63082a <=( a63081a  and  a63078a );
 a63083a <=( a63082a  and  a63075a );
 a63086a <=( (not A235)  and  (not A233) );
 a63089a <=( (not A268)  and  (not A267) );
 a63090a <=( a63089a  and  a63086a );
 a63093a <=( A298  and  (not A269) );
 a63096a <=( A302  and  (not A299) );
 a63097a <=( a63096a  and  a63093a );
 a63098a <=( a63097a  and  a63090a );
 a63101a <=( (not A168)  and  (not A169) );
 a63104a <=( A166  and  A167 );
 a63105a <=( a63104a  and  a63101a );
 a63108a <=( (not A200)  and  A199 );
 a63111a <=( (not A232)  and  A203 );
 a63112a <=( a63111a  and  a63108a );
 a63113a <=( a63112a  and  a63105a );
 a63116a <=( (not A235)  and  (not A233) );
 a63119a <=( (not A268)  and  (not A267) );
 a63120a <=( a63119a  and  a63116a );
 a63123a <=( (not A298)  and  (not A269) );
 a63126a <=( A302  and  A299 );
 a63127a <=( a63126a  and  a63123a );
 a63128a <=( a63127a  and  a63120a );
 a63131a <=( (not A168)  and  (not A169) );
 a63134a <=( A166  and  A167 );
 a63135a <=( a63134a  and  a63131a );
 a63138a <=( (not A200)  and  A199 );
 a63141a <=( (not A232)  and  A203 );
 a63142a <=( a63141a  and  a63138a );
 a63143a <=( a63142a  and  a63135a );
 a63146a <=( (not A235)  and  (not A233) );
 a63149a <=( A266  and  A265 );
 a63150a <=( a63149a  and  a63146a );
 a63153a <=( (not A268)  and  (not A267) );
 a63156a <=( A300  and  A299 );
 a63157a <=( a63156a  and  a63153a );
 a63158a <=( a63157a  and  a63150a );
 a63161a <=( (not A168)  and  (not A169) );
 a63164a <=( A166  and  A167 );
 a63165a <=( a63164a  and  a63161a );
 a63168a <=( (not A200)  and  A199 );
 a63171a <=( (not A232)  and  A203 );
 a63172a <=( a63171a  and  a63168a );
 a63173a <=( a63172a  and  a63165a );
 a63176a <=( (not A235)  and  (not A233) );
 a63179a <=( A266  and  A265 );
 a63180a <=( a63179a  and  a63176a );
 a63183a <=( (not A268)  and  (not A267) );
 a63186a <=( A300  and  A298 );
 a63187a <=( a63186a  and  a63183a );
 a63188a <=( a63187a  and  a63180a );
 a63191a <=( (not A168)  and  (not A169) );
 a63194a <=( A166  and  A167 );
 a63195a <=( a63194a  and  a63191a );
 a63198a <=( (not A200)  and  A199 );
 a63201a <=( (not A232)  and  A203 );
 a63202a <=( a63201a  and  a63198a );
 a63203a <=( a63202a  and  a63195a );
 a63206a <=( (not A235)  and  (not A233) );
 a63209a <=( (not A266)  and  (not A265) );
 a63210a <=( a63209a  and  a63206a );
 a63213a <=( A298  and  (not A268) );
 a63216a <=( A302  and  (not A299) );
 a63217a <=( a63216a  and  a63213a );
 a63218a <=( a63217a  and  a63210a );
 a63221a <=( (not A168)  and  (not A169) );
 a63224a <=( A166  and  A167 );
 a63225a <=( a63224a  and  a63221a );
 a63228a <=( (not A200)  and  A199 );
 a63231a <=( (not A232)  and  A203 );
 a63232a <=( a63231a  and  a63228a );
 a63233a <=( a63232a  and  a63225a );
 a63236a <=( (not A235)  and  (not A233) );
 a63239a <=( (not A266)  and  (not A265) );
 a63240a <=( a63239a  and  a63236a );
 a63243a <=( (not A298)  and  (not A268) );
 a63246a <=( A302  and  A299 );
 a63247a <=( a63246a  and  a63243a );
 a63248a <=( a63247a  and  a63240a );
 a63251a <=( (not A169)  and  (not A170) );
 a63254a <=( A199  and  (not A168) );
 a63255a <=( a63254a  and  a63251a );
 a63258a <=( A232  and  A201 );
 a63261a <=( (not A234)  and  A233 );
 a63262a <=( a63261a  and  a63258a );
 a63263a <=( a63262a  and  a63255a );
 a63266a <=( A265  and  (not A235) );
 a63269a <=( (not A267)  and  A266 );
 a63270a <=( a63269a  and  a63266a );
 a63273a <=( A298  and  (not A268) );
 a63276a <=( A302  and  (not A299) );
 a63277a <=( a63276a  and  a63273a );
 a63278a <=( a63277a  and  a63270a );
 a63281a <=( (not A169)  and  (not A170) );
 a63284a <=( A199  and  (not A168) );
 a63285a <=( a63284a  and  a63281a );
 a63288a <=( A232  and  A201 );
 a63291a <=( (not A234)  and  A233 );
 a63292a <=( a63291a  and  a63288a );
 a63293a <=( a63292a  and  a63285a );
 a63296a <=( A265  and  (not A235) );
 a63299a <=( (not A267)  and  A266 );
 a63300a <=( a63299a  and  a63296a );
 a63303a <=( (not A298)  and  (not A268) );
 a63306a <=( A302  and  A299 );
 a63307a <=( a63306a  and  a63303a );
 a63308a <=( a63307a  and  a63300a );
 a63311a <=( (not A169)  and  (not A170) );
 a63314a <=( A200  and  (not A168) );
 a63315a <=( a63314a  and  a63311a );
 a63318a <=( A232  and  A201 );
 a63321a <=( (not A234)  and  A233 );
 a63322a <=( a63321a  and  a63318a );
 a63323a <=( a63322a  and  a63315a );
 a63326a <=( A265  and  (not A235) );
 a63329a <=( (not A267)  and  A266 );
 a63330a <=( a63329a  and  a63326a );
 a63333a <=( A298  and  (not A268) );
 a63336a <=( A302  and  (not A299) );
 a63337a <=( a63336a  and  a63333a );
 a63338a <=( a63337a  and  a63330a );
 a63341a <=( (not A169)  and  (not A170) );
 a63344a <=( A200  and  (not A168) );
 a63345a <=( a63344a  and  a63341a );
 a63348a <=( A232  and  A201 );
 a63351a <=( (not A234)  and  A233 );
 a63352a <=( a63351a  and  a63348a );
 a63353a <=( a63352a  and  a63345a );
 a63356a <=( A265  and  (not A235) );
 a63359a <=( (not A267)  and  A266 );
 a63360a <=( a63359a  and  a63356a );
 a63363a <=( (not A298)  and  (not A268) );
 a63366a <=( A302  and  A299 );
 a63367a <=( a63366a  and  a63363a );
 a63368a <=( a63367a  and  a63360a );
 a63371a <=( (not A169)  and  (not A170) );
 a63374a <=( (not A199)  and  (not A168) );
 a63375a <=( a63374a  and  a63371a );
 a63378a <=( A203  and  A200 );
 a63381a <=( (not A235)  and  (not A234) );
 a63382a <=( a63381a  and  a63378a );
 a63383a <=( a63382a  and  a63375a );
 a63386a <=( A265  and  (not A236) );
 a63389a <=( (not A267)  and  A266 );
 a63390a <=( a63389a  and  a63386a );
 a63393a <=( A298  and  (not A268) );
 a63396a <=( A302  and  (not A299) );
 a63397a <=( a63396a  and  a63393a );
 a63398a <=( a63397a  and  a63390a );
 a63401a <=( (not A169)  and  (not A170) );
 a63404a <=( (not A199)  and  (not A168) );
 a63405a <=( a63404a  and  a63401a );
 a63408a <=( A203  and  A200 );
 a63411a <=( (not A235)  and  (not A234) );
 a63412a <=( a63411a  and  a63408a );
 a63413a <=( a63412a  and  a63405a );
 a63416a <=( A265  and  (not A236) );
 a63419a <=( (not A267)  and  A266 );
 a63420a <=( a63419a  and  a63416a );
 a63423a <=( (not A298)  and  (not A268) );
 a63426a <=( A302  and  A299 );
 a63427a <=( a63426a  and  a63423a );
 a63428a <=( a63427a  and  a63420a );
 a63431a <=( (not A169)  and  (not A170) );
 a63434a <=( (not A199)  and  (not A168) );
 a63435a <=( a63434a  and  a63431a );
 a63438a <=( A203  and  A200 );
 a63441a <=( A233  and  A232 );
 a63442a <=( a63441a  and  a63438a );
 a63443a <=( a63442a  and  a63435a );
 a63446a <=( (not A235)  and  (not A234) );
 a63449a <=( (not A268)  and  (not A267) );
 a63450a <=( a63449a  and  a63446a );
 a63453a <=( A298  and  (not A269) );
 a63456a <=( A302  and  (not A299) );
 a63457a <=( a63456a  and  a63453a );
 a63458a <=( a63457a  and  a63450a );
 a63461a <=( (not A169)  and  (not A170) );
 a63464a <=( (not A199)  and  (not A168) );
 a63465a <=( a63464a  and  a63461a );
 a63468a <=( A203  and  A200 );
 a63471a <=( A233  and  A232 );
 a63472a <=( a63471a  and  a63468a );
 a63473a <=( a63472a  and  a63465a );
 a63476a <=( (not A235)  and  (not A234) );
 a63479a <=( (not A268)  and  (not A267) );
 a63480a <=( a63479a  and  a63476a );
 a63483a <=( (not A298)  and  (not A269) );
 a63486a <=( A302  and  A299 );
 a63487a <=( a63486a  and  a63483a );
 a63488a <=( a63487a  and  a63480a );
 a63491a <=( (not A169)  and  (not A170) );
 a63494a <=( (not A199)  and  (not A168) );
 a63495a <=( a63494a  and  a63491a );
 a63498a <=( A203  and  A200 );
 a63501a <=( A233  and  A232 );
 a63502a <=( a63501a  and  a63498a );
 a63503a <=( a63502a  and  a63495a );
 a63506a <=( (not A235)  and  (not A234) );
 a63509a <=( A266  and  A265 );
 a63510a <=( a63509a  and  a63506a );
 a63513a <=( (not A268)  and  (not A267) );
 a63516a <=( A300  and  A299 );
 a63517a <=( a63516a  and  a63513a );
 a63518a <=( a63517a  and  a63510a );
 a63521a <=( (not A169)  and  (not A170) );
 a63524a <=( (not A199)  and  (not A168) );
 a63525a <=( a63524a  and  a63521a );
 a63528a <=( A203  and  A200 );
 a63531a <=( A233  and  A232 );
 a63532a <=( a63531a  and  a63528a );
 a63533a <=( a63532a  and  a63525a );
 a63536a <=( (not A235)  and  (not A234) );
 a63539a <=( A266  and  A265 );
 a63540a <=( a63539a  and  a63536a );
 a63543a <=( (not A268)  and  (not A267) );
 a63546a <=( A300  and  A298 );
 a63547a <=( a63546a  and  a63543a );
 a63548a <=( a63547a  and  a63540a );
 a63551a <=( (not A169)  and  (not A170) );
 a63554a <=( (not A199)  and  (not A168) );
 a63555a <=( a63554a  and  a63551a );
 a63558a <=( A203  and  A200 );
 a63561a <=( A233  and  A232 );
 a63562a <=( a63561a  and  a63558a );
 a63563a <=( a63562a  and  a63555a );
 a63566a <=( (not A235)  and  (not A234) );
 a63569a <=( (not A266)  and  (not A265) );
 a63570a <=( a63569a  and  a63566a );
 a63573a <=( A298  and  (not A268) );
 a63576a <=( A302  and  (not A299) );
 a63577a <=( a63576a  and  a63573a );
 a63578a <=( a63577a  and  a63570a );
 a63581a <=( (not A169)  and  (not A170) );
 a63584a <=( (not A199)  and  (not A168) );
 a63585a <=( a63584a  and  a63581a );
 a63588a <=( A203  and  A200 );
 a63591a <=( A233  and  A232 );
 a63592a <=( a63591a  and  a63588a );
 a63593a <=( a63592a  and  a63585a );
 a63596a <=( (not A235)  and  (not A234) );
 a63599a <=( (not A266)  and  (not A265) );
 a63600a <=( a63599a  and  a63596a );
 a63603a <=( (not A298)  and  (not A268) );
 a63606a <=( A302  and  A299 );
 a63607a <=( a63606a  and  a63603a );
 a63608a <=( a63607a  and  a63600a );
 a63611a <=( (not A169)  and  (not A170) );
 a63614a <=( (not A199)  and  (not A168) );
 a63615a <=( a63614a  and  a63611a );
 a63618a <=( A203  and  A200 );
 a63621a <=( (not A233)  and  (not A232) );
 a63622a <=( a63621a  and  a63618a );
 a63623a <=( a63622a  and  a63615a );
 a63626a <=( A265  and  (not A235) );
 a63629a <=( (not A267)  and  A266 );
 a63630a <=( a63629a  and  a63626a );
 a63633a <=( A298  and  (not A268) );
 a63636a <=( A302  and  (not A299) );
 a63637a <=( a63636a  and  a63633a );
 a63638a <=( a63637a  and  a63630a );
 a63641a <=( (not A169)  and  (not A170) );
 a63644a <=( (not A199)  and  (not A168) );
 a63645a <=( a63644a  and  a63641a );
 a63648a <=( A203  and  A200 );
 a63651a <=( (not A233)  and  (not A232) );
 a63652a <=( a63651a  and  a63648a );
 a63653a <=( a63652a  and  a63645a );
 a63656a <=( A265  and  (not A235) );
 a63659a <=( (not A267)  and  A266 );
 a63660a <=( a63659a  and  a63656a );
 a63663a <=( (not A298)  and  (not A268) );
 a63666a <=( A302  and  A299 );
 a63667a <=( a63666a  and  a63663a );
 a63668a <=( a63667a  and  a63660a );
 a63671a <=( (not A169)  and  (not A170) );
 a63674a <=( A199  and  (not A168) );
 a63675a <=( a63674a  and  a63671a );
 a63678a <=( A203  and  (not A200) );
 a63681a <=( (not A235)  and  (not A234) );
 a63682a <=( a63681a  and  a63678a );
 a63683a <=( a63682a  and  a63675a );
 a63686a <=( A265  and  (not A236) );
 a63689a <=( (not A267)  and  A266 );
 a63690a <=( a63689a  and  a63686a );
 a63693a <=( A298  and  (not A268) );
 a63696a <=( A302  and  (not A299) );
 a63697a <=( a63696a  and  a63693a );
 a63698a <=( a63697a  and  a63690a );
 a63701a <=( (not A169)  and  (not A170) );
 a63704a <=( A199  and  (not A168) );
 a63705a <=( a63704a  and  a63701a );
 a63708a <=( A203  and  (not A200) );
 a63711a <=( (not A235)  and  (not A234) );
 a63712a <=( a63711a  and  a63708a );
 a63713a <=( a63712a  and  a63705a );
 a63716a <=( A265  and  (not A236) );
 a63719a <=( (not A267)  and  A266 );
 a63720a <=( a63719a  and  a63716a );
 a63723a <=( (not A298)  and  (not A268) );
 a63726a <=( A302  and  A299 );
 a63727a <=( a63726a  and  a63723a );
 a63728a <=( a63727a  and  a63720a );
 a63731a <=( (not A169)  and  (not A170) );
 a63734a <=( A199  and  (not A168) );
 a63735a <=( a63734a  and  a63731a );
 a63738a <=( A203  and  (not A200) );
 a63741a <=( A233  and  A232 );
 a63742a <=( a63741a  and  a63738a );
 a63743a <=( a63742a  and  a63735a );
 a63746a <=( (not A235)  and  (not A234) );
 a63749a <=( (not A268)  and  (not A267) );
 a63750a <=( a63749a  and  a63746a );
 a63753a <=( A298  and  (not A269) );
 a63756a <=( A302  and  (not A299) );
 a63757a <=( a63756a  and  a63753a );
 a63758a <=( a63757a  and  a63750a );
 a63761a <=( (not A169)  and  (not A170) );
 a63764a <=( A199  and  (not A168) );
 a63765a <=( a63764a  and  a63761a );
 a63768a <=( A203  and  (not A200) );
 a63771a <=( A233  and  A232 );
 a63772a <=( a63771a  and  a63768a );
 a63773a <=( a63772a  and  a63765a );
 a63776a <=( (not A235)  and  (not A234) );
 a63779a <=( (not A268)  and  (not A267) );
 a63780a <=( a63779a  and  a63776a );
 a63783a <=( (not A298)  and  (not A269) );
 a63786a <=( A302  and  A299 );
 a63787a <=( a63786a  and  a63783a );
 a63788a <=( a63787a  and  a63780a );
 a63791a <=( (not A169)  and  (not A170) );
 a63794a <=( A199  and  (not A168) );
 a63795a <=( a63794a  and  a63791a );
 a63798a <=( A203  and  (not A200) );
 a63801a <=( A233  and  A232 );
 a63802a <=( a63801a  and  a63798a );
 a63803a <=( a63802a  and  a63795a );
 a63806a <=( (not A235)  and  (not A234) );
 a63809a <=( A266  and  A265 );
 a63810a <=( a63809a  and  a63806a );
 a63813a <=( (not A268)  and  (not A267) );
 a63816a <=( A300  and  A299 );
 a63817a <=( a63816a  and  a63813a );
 a63818a <=( a63817a  and  a63810a );
 a63821a <=( (not A169)  and  (not A170) );
 a63824a <=( A199  and  (not A168) );
 a63825a <=( a63824a  and  a63821a );
 a63828a <=( A203  and  (not A200) );
 a63831a <=( A233  and  A232 );
 a63832a <=( a63831a  and  a63828a );
 a63833a <=( a63832a  and  a63825a );
 a63836a <=( (not A235)  and  (not A234) );
 a63839a <=( A266  and  A265 );
 a63840a <=( a63839a  and  a63836a );
 a63843a <=( (not A268)  and  (not A267) );
 a63846a <=( A300  and  A298 );
 a63847a <=( a63846a  and  a63843a );
 a63848a <=( a63847a  and  a63840a );
 a63851a <=( (not A169)  and  (not A170) );
 a63854a <=( A199  and  (not A168) );
 a63855a <=( a63854a  and  a63851a );
 a63858a <=( A203  and  (not A200) );
 a63861a <=( A233  and  A232 );
 a63862a <=( a63861a  and  a63858a );
 a63863a <=( a63862a  and  a63855a );
 a63866a <=( (not A235)  and  (not A234) );
 a63869a <=( (not A266)  and  (not A265) );
 a63870a <=( a63869a  and  a63866a );
 a63873a <=( A298  and  (not A268) );
 a63876a <=( A302  and  (not A299) );
 a63877a <=( a63876a  and  a63873a );
 a63878a <=( a63877a  and  a63870a );
 a63881a <=( (not A169)  and  (not A170) );
 a63884a <=( A199  and  (not A168) );
 a63885a <=( a63884a  and  a63881a );
 a63888a <=( A203  and  (not A200) );
 a63891a <=( A233  and  A232 );
 a63892a <=( a63891a  and  a63888a );
 a63893a <=( a63892a  and  a63885a );
 a63896a <=( (not A235)  and  (not A234) );
 a63899a <=( (not A266)  and  (not A265) );
 a63900a <=( a63899a  and  a63896a );
 a63903a <=( (not A298)  and  (not A268) );
 a63906a <=( A302  and  A299 );
 a63907a <=( a63906a  and  a63903a );
 a63908a <=( a63907a  and  a63900a );
 a63911a <=( (not A169)  and  (not A170) );
 a63914a <=( A199  and  (not A168) );
 a63915a <=( a63914a  and  a63911a );
 a63918a <=( A203  and  (not A200) );
 a63921a <=( (not A233)  and  (not A232) );
 a63922a <=( a63921a  and  a63918a );
 a63923a <=( a63922a  and  a63915a );
 a63926a <=( A265  and  (not A235) );
 a63929a <=( (not A267)  and  A266 );
 a63930a <=( a63929a  and  a63926a );
 a63933a <=( A298  and  (not A268) );
 a63936a <=( A302  and  (not A299) );
 a63937a <=( a63936a  and  a63933a );
 a63938a <=( a63937a  and  a63930a );
 a63941a <=( (not A169)  and  (not A170) );
 a63944a <=( A199  and  (not A168) );
 a63945a <=( a63944a  and  a63941a );
 a63948a <=( A203  and  (not A200) );
 a63951a <=( (not A233)  and  (not A232) );
 a63952a <=( a63951a  and  a63948a );
 a63953a <=( a63952a  and  a63945a );
 a63956a <=( A265  and  (not A235) );
 a63959a <=( (not A267)  and  A266 );
 a63960a <=( a63959a  and  a63956a );
 a63963a <=( (not A298)  and  (not A268) );
 a63966a <=( A302  and  A299 );
 a63967a <=( a63966a  and  a63963a );
 a63968a <=( a63967a  and  a63960a );
 a63971a <=( A166  and  A168 );
 a63974a <=( A200  and  A199 );
 a63975a <=( a63974a  and  a63971a );
 a63978a <=( (not A202)  and  (not A201) );
 a63981a <=( A233  and  A232 );
 a63982a <=( a63981a  and  a63978a );
 a63983a <=( a63982a  and  a63975a );
 a63986a <=( (not A235)  and  (not A234) );
 a63989a <=( A266  and  A265 );
 a63990a <=( a63989a  and  a63986a );
 a63993a <=( (not A268)  and  (not A267) );
 a63997a <=( A302  and  (not A299) );
 a63998a <=( A298  and  a63997a );
 a63999a <=( a63998a  and  a63993a );
 a64000a <=( a63999a  and  a63990a );
 a64003a <=( A166  and  A168 );
 a64006a <=( A200  and  A199 );
 a64007a <=( a64006a  and  a64003a );
 a64010a <=( (not A202)  and  (not A201) );
 a64013a <=( A233  and  A232 );
 a64014a <=( a64013a  and  a64010a );
 a64015a <=( a64014a  and  a64007a );
 a64018a <=( (not A235)  and  (not A234) );
 a64021a <=( A266  and  A265 );
 a64022a <=( a64021a  and  a64018a );
 a64025a <=( (not A268)  and  (not A267) );
 a64029a <=( A302  and  A299 );
 a64030a <=( (not A298)  and  a64029a );
 a64031a <=( a64030a  and  a64025a );
 a64032a <=( a64031a  and  a64022a );
 a64035a <=( A167  and  A168 );
 a64038a <=( A200  and  A199 );
 a64039a <=( a64038a  and  a64035a );
 a64042a <=( (not A202)  and  (not A201) );
 a64045a <=( A233  and  A232 );
 a64046a <=( a64045a  and  a64042a );
 a64047a <=( a64046a  and  a64039a );
 a64050a <=( (not A235)  and  (not A234) );
 a64053a <=( A266  and  A265 );
 a64054a <=( a64053a  and  a64050a );
 a64057a <=( (not A268)  and  (not A267) );
 a64061a <=( A302  and  (not A299) );
 a64062a <=( A298  and  a64061a );
 a64063a <=( a64062a  and  a64057a );
 a64064a <=( a64063a  and  a64054a );
 a64067a <=( A167  and  A168 );
 a64070a <=( A200  and  A199 );
 a64071a <=( a64070a  and  a64067a );
 a64074a <=( (not A202)  and  (not A201) );
 a64077a <=( A233  and  A232 );
 a64078a <=( a64077a  and  a64074a );
 a64079a <=( a64078a  and  a64071a );
 a64082a <=( (not A235)  and  (not A234) );
 a64085a <=( A266  and  A265 );
 a64086a <=( a64085a  and  a64082a );
 a64089a <=( (not A268)  and  (not A267) );
 a64093a <=( A302  and  A299 );
 a64094a <=( (not A298)  and  a64093a );
 a64095a <=( a64094a  and  a64089a );
 a64096a <=( a64095a  and  a64086a );
 a64099a <=( A167  and  A170 );
 a64102a <=( (not A201)  and  (not A166) );
 a64103a <=( a64102a  and  a64099a );
 a64106a <=( (not A203)  and  (not A202) );
 a64109a <=( A233  and  A232 );
 a64110a <=( a64109a  and  a64106a );
 a64111a <=( a64110a  and  a64103a );
 a64114a <=( (not A235)  and  (not A234) );
 a64117a <=( A266  and  A265 );
 a64118a <=( a64117a  and  a64114a );
 a64121a <=( (not A268)  and  (not A267) );
 a64125a <=( A302  and  (not A299) );
 a64126a <=( A298  and  a64125a );
 a64127a <=( a64126a  and  a64121a );
 a64128a <=( a64127a  and  a64118a );
 a64131a <=( A167  and  A170 );
 a64134a <=( (not A201)  and  (not A166) );
 a64135a <=( a64134a  and  a64131a );
 a64138a <=( (not A203)  and  (not A202) );
 a64141a <=( A233  and  A232 );
 a64142a <=( a64141a  and  a64138a );
 a64143a <=( a64142a  and  a64135a );
 a64146a <=( (not A235)  and  (not A234) );
 a64149a <=( A266  and  A265 );
 a64150a <=( a64149a  and  a64146a );
 a64153a <=( (not A268)  and  (not A267) );
 a64157a <=( A302  and  A299 );
 a64158a <=( (not A298)  and  a64157a );
 a64159a <=( a64158a  and  a64153a );
 a64160a <=( a64159a  and  a64150a );
 a64163a <=( A167  and  A170 );
 a64166a <=( A199  and  (not A166) );
 a64167a <=( a64166a  and  a64163a );
 a64170a <=( (not A201)  and  A200 );
 a64173a <=( (not A234)  and  (not A202) );
 a64174a <=( a64173a  and  a64170a );
 a64175a <=( a64174a  and  a64167a );
 a64178a <=( (not A236)  and  (not A235) );
 a64181a <=( A266  and  A265 );
 a64182a <=( a64181a  and  a64178a );
 a64185a <=( (not A268)  and  (not A267) );
 a64189a <=( A302  and  (not A299) );
 a64190a <=( A298  and  a64189a );
 a64191a <=( a64190a  and  a64185a );
 a64192a <=( a64191a  and  a64182a );
 a64195a <=( A167  and  A170 );
 a64198a <=( A199  and  (not A166) );
 a64199a <=( a64198a  and  a64195a );
 a64202a <=( (not A201)  and  A200 );
 a64205a <=( (not A234)  and  (not A202) );
 a64206a <=( a64205a  and  a64202a );
 a64207a <=( a64206a  and  a64199a );
 a64210a <=( (not A236)  and  (not A235) );
 a64213a <=( A266  and  A265 );
 a64214a <=( a64213a  and  a64210a );
 a64217a <=( (not A268)  and  (not A267) );
 a64221a <=( A302  and  A299 );
 a64222a <=( (not A298)  and  a64221a );
 a64223a <=( a64222a  and  a64217a );
 a64224a <=( a64223a  and  a64214a );
 a64227a <=( A167  and  A170 );
 a64230a <=( A199  and  (not A166) );
 a64231a <=( a64230a  and  a64227a );
 a64234a <=( (not A201)  and  A200 );
 a64237a <=( A232  and  (not A202) );
 a64238a <=( a64237a  and  a64234a );
 a64239a <=( a64238a  and  a64231a );
 a64242a <=( (not A234)  and  A233 );
 a64245a <=( (not A267)  and  (not A235) );
 a64246a <=( a64245a  and  a64242a );
 a64249a <=( (not A269)  and  (not A268) );
 a64253a <=( A302  and  (not A299) );
 a64254a <=( A298  and  a64253a );
 a64255a <=( a64254a  and  a64249a );
 a64256a <=( a64255a  and  a64246a );
 a64259a <=( A167  and  A170 );
 a64262a <=( A199  and  (not A166) );
 a64263a <=( a64262a  and  a64259a );
 a64266a <=( (not A201)  and  A200 );
 a64269a <=( A232  and  (not A202) );
 a64270a <=( a64269a  and  a64266a );
 a64271a <=( a64270a  and  a64263a );
 a64274a <=( (not A234)  and  A233 );
 a64277a <=( (not A267)  and  (not A235) );
 a64278a <=( a64277a  and  a64274a );
 a64281a <=( (not A269)  and  (not A268) );
 a64285a <=( A302  and  A299 );
 a64286a <=( (not A298)  and  a64285a );
 a64287a <=( a64286a  and  a64281a );
 a64288a <=( a64287a  and  a64278a );
 a64291a <=( A167  and  A170 );
 a64294a <=( A199  and  (not A166) );
 a64295a <=( a64294a  and  a64291a );
 a64298a <=( (not A201)  and  A200 );
 a64301a <=( A232  and  (not A202) );
 a64302a <=( a64301a  and  a64298a );
 a64303a <=( a64302a  and  a64295a );
 a64306a <=( (not A234)  and  A233 );
 a64309a <=( A265  and  (not A235) );
 a64310a <=( a64309a  and  a64306a );
 a64313a <=( (not A267)  and  A266 );
 a64317a <=( A300  and  A299 );
 a64318a <=( (not A268)  and  a64317a );
 a64319a <=( a64318a  and  a64313a );
 a64320a <=( a64319a  and  a64310a );
 a64323a <=( A167  and  A170 );
 a64326a <=( A199  and  (not A166) );
 a64327a <=( a64326a  and  a64323a );
 a64330a <=( (not A201)  and  A200 );
 a64333a <=( A232  and  (not A202) );
 a64334a <=( a64333a  and  a64330a );
 a64335a <=( a64334a  and  a64327a );
 a64338a <=( (not A234)  and  A233 );
 a64341a <=( A265  and  (not A235) );
 a64342a <=( a64341a  and  a64338a );
 a64345a <=( (not A267)  and  A266 );
 a64349a <=( A300  and  A298 );
 a64350a <=( (not A268)  and  a64349a );
 a64351a <=( a64350a  and  a64345a );
 a64352a <=( a64351a  and  a64342a );
 a64355a <=( A167  and  A170 );
 a64358a <=( A199  and  (not A166) );
 a64359a <=( a64358a  and  a64355a );
 a64362a <=( (not A201)  and  A200 );
 a64365a <=( A232  and  (not A202) );
 a64366a <=( a64365a  and  a64362a );
 a64367a <=( a64366a  and  a64359a );
 a64370a <=( (not A234)  and  A233 );
 a64373a <=( (not A265)  and  (not A235) );
 a64374a <=( a64373a  and  a64370a );
 a64377a <=( (not A268)  and  (not A266) );
 a64381a <=( A302  and  (not A299) );
 a64382a <=( A298  and  a64381a );
 a64383a <=( a64382a  and  a64377a );
 a64384a <=( a64383a  and  a64374a );
 a64387a <=( A167  and  A170 );
 a64390a <=( A199  and  (not A166) );
 a64391a <=( a64390a  and  a64387a );
 a64394a <=( (not A201)  and  A200 );
 a64397a <=( A232  and  (not A202) );
 a64398a <=( a64397a  and  a64394a );
 a64399a <=( a64398a  and  a64391a );
 a64402a <=( (not A234)  and  A233 );
 a64405a <=( (not A265)  and  (not A235) );
 a64406a <=( a64405a  and  a64402a );
 a64409a <=( (not A268)  and  (not A266) );
 a64413a <=( A302  and  A299 );
 a64414a <=( (not A298)  and  a64413a );
 a64415a <=( a64414a  and  a64409a );
 a64416a <=( a64415a  and  a64406a );
 a64419a <=( A167  and  A170 );
 a64422a <=( A199  and  (not A166) );
 a64423a <=( a64422a  and  a64419a );
 a64426a <=( (not A201)  and  A200 );
 a64429a <=( (not A232)  and  (not A202) );
 a64430a <=( a64429a  and  a64426a );
 a64431a <=( a64430a  and  a64423a );
 a64434a <=( (not A235)  and  (not A233) );
 a64437a <=( A266  and  A265 );
 a64438a <=( a64437a  and  a64434a );
 a64441a <=( (not A268)  and  (not A267) );
 a64445a <=( A302  and  (not A299) );
 a64446a <=( A298  and  a64445a );
 a64447a <=( a64446a  and  a64441a );
 a64448a <=( a64447a  and  a64438a );
 a64451a <=( A167  and  A170 );
 a64454a <=( A199  and  (not A166) );
 a64455a <=( a64454a  and  a64451a );
 a64458a <=( (not A201)  and  A200 );
 a64461a <=( (not A232)  and  (not A202) );
 a64462a <=( a64461a  and  a64458a );
 a64463a <=( a64462a  and  a64455a );
 a64466a <=( (not A235)  and  (not A233) );
 a64469a <=( A266  and  A265 );
 a64470a <=( a64469a  and  a64466a );
 a64473a <=( (not A268)  and  (not A267) );
 a64477a <=( A302  and  A299 );
 a64478a <=( (not A298)  and  a64477a );
 a64479a <=( a64478a  and  a64473a );
 a64480a <=( a64479a  and  a64470a );
 a64483a <=( A167  and  A170 );
 a64486a <=( (not A199)  and  (not A166) );
 a64487a <=( a64486a  and  a64483a );
 a64490a <=( (not A202)  and  (not A200) );
 a64493a <=( A233  and  A232 );
 a64494a <=( a64493a  and  a64490a );
 a64495a <=( a64494a  and  a64487a );
 a64498a <=( (not A235)  and  (not A234) );
 a64501a <=( A266  and  A265 );
 a64502a <=( a64501a  and  a64498a );
 a64505a <=( (not A268)  and  (not A267) );
 a64509a <=( A302  and  (not A299) );
 a64510a <=( A298  and  a64509a );
 a64511a <=( a64510a  and  a64505a );
 a64512a <=( a64511a  and  a64502a );
 a64515a <=( A167  and  A170 );
 a64518a <=( (not A199)  and  (not A166) );
 a64519a <=( a64518a  and  a64515a );
 a64522a <=( (not A202)  and  (not A200) );
 a64525a <=( A233  and  A232 );
 a64526a <=( a64525a  and  a64522a );
 a64527a <=( a64526a  and  a64519a );
 a64530a <=( (not A235)  and  (not A234) );
 a64533a <=( A266  and  A265 );
 a64534a <=( a64533a  and  a64530a );
 a64537a <=( (not A268)  and  (not A267) );
 a64541a <=( A302  and  A299 );
 a64542a <=( (not A298)  and  a64541a );
 a64543a <=( a64542a  and  a64537a );
 a64544a <=( a64543a  and  a64534a );
 a64547a <=( (not A167)  and  A170 );
 a64550a <=( (not A201)  and  A166 );
 a64551a <=( a64550a  and  a64547a );
 a64554a <=( (not A203)  and  (not A202) );
 a64557a <=( A233  and  A232 );
 a64558a <=( a64557a  and  a64554a );
 a64559a <=( a64558a  and  a64551a );
 a64562a <=( (not A235)  and  (not A234) );
 a64565a <=( A266  and  A265 );
 a64566a <=( a64565a  and  a64562a );
 a64569a <=( (not A268)  and  (not A267) );
 a64573a <=( A302  and  (not A299) );
 a64574a <=( A298  and  a64573a );
 a64575a <=( a64574a  and  a64569a );
 a64576a <=( a64575a  and  a64566a );
 a64579a <=( (not A167)  and  A170 );
 a64582a <=( (not A201)  and  A166 );
 a64583a <=( a64582a  and  a64579a );
 a64586a <=( (not A203)  and  (not A202) );
 a64589a <=( A233  and  A232 );
 a64590a <=( a64589a  and  a64586a );
 a64591a <=( a64590a  and  a64583a );
 a64594a <=( (not A235)  and  (not A234) );
 a64597a <=( A266  and  A265 );
 a64598a <=( a64597a  and  a64594a );
 a64601a <=( (not A268)  and  (not A267) );
 a64605a <=( A302  and  A299 );
 a64606a <=( (not A298)  and  a64605a );
 a64607a <=( a64606a  and  a64601a );
 a64608a <=( a64607a  and  a64598a );
 a64611a <=( (not A167)  and  A170 );
 a64614a <=( A199  and  A166 );
 a64615a <=( a64614a  and  a64611a );
 a64618a <=( (not A201)  and  A200 );
 a64621a <=( (not A234)  and  (not A202) );
 a64622a <=( a64621a  and  a64618a );
 a64623a <=( a64622a  and  a64615a );
 a64626a <=( (not A236)  and  (not A235) );
 a64629a <=( A266  and  A265 );
 a64630a <=( a64629a  and  a64626a );
 a64633a <=( (not A268)  and  (not A267) );
 a64637a <=( A302  and  (not A299) );
 a64638a <=( A298  and  a64637a );
 a64639a <=( a64638a  and  a64633a );
 a64640a <=( a64639a  and  a64630a );
 a64643a <=( (not A167)  and  A170 );
 a64646a <=( A199  and  A166 );
 a64647a <=( a64646a  and  a64643a );
 a64650a <=( (not A201)  and  A200 );
 a64653a <=( (not A234)  and  (not A202) );
 a64654a <=( a64653a  and  a64650a );
 a64655a <=( a64654a  and  a64647a );
 a64658a <=( (not A236)  and  (not A235) );
 a64661a <=( A266  and  A265 );
 a64662a <=( a64661a  and  a64658a );
 a64665a <=( (not A268)  and  (not A267) );
 a64669a <=( A302  and  A299 );
 a64670a <=( (not A298)  and  a64669a );
 a64671a <=( a64670a  and  a64665a );
 a64672a <=( a64671a  and  a64662a );
 a64675a <=( (not A167)  and  A170 );
 a64678a <=( A199  and  A166 );
 a64679a <=( a64678a  and  a64675a );
 a64682a <=( (not A201)  and  A200 );
 a64685a <=( A232  and  (not A202) );
 a64686a <=( a64685a  and  a64682a );
 a64687a <=( a64686a  and  a64679a );
 a64690a <=( (not A234)  and  A233 );
 a64693a <=( (not A267)  and  (not A235) );
 a64694a <=( a64693a  and  a64690a );
 a64697a <=( (not A269)  and  (not A268) );
 a64701a <=( A302  and  (not A299) );
 a64702a <=( A298  and  a64701a );
 a64703a <=( a64702a  and  a64697a );
 a64704a <=( a64703a  and  a64694a );
 a64707a <=( (not A167)  and  A170 );
 a64710a <=( A199  and  A166 );
 a64711a <=( a64710a  and  a64707a );
 a64714a <=( (not A201)  and  A200 );
 a64717a <=( A232  and  (not A202) );
 a64718a <=( a64717a  and  a64714a );
 a64719a <=( a64718a  and  a64711a );
 a64722a <=( (not A234)  and  A233 );
 a64725a <=( (not A267)  and  (not A235) );
 a64726a <=( a64725a  and  a64722a );
 a64729a <=( (not A269)  and  (not A268) );
 a64733a <=( A302  and  A299 );
 a64734a <=( (not A298)  and  a64733a );
 a64735a <=( a64734a  and  a64729a );
 a64736a <=( a64735a  and  a64726a );
 a64739a <=( (not A167)  and  A170 );
 a64742a <=( A199  and  A166 );
 a64743a <=( a64742a  and  a64739a );
 a64746a <=( (not A201)  and  A200 );
 a64749a <=( A232  and  (not A202) );
 a64750a <=( a64749a  and  a64746a );
 a64751a <=( a64750a  and  a64743a );
 a64754a <=( (not A234)  and  A233 );
 a64757a <=( A265  and  (not A235) );
 a64758a <=( a64757a  and  a64754a );
 a64761a <=( (not A267)  and  A266 );
 a64765a <=( A300  and  A299 );
 a64766a <=( (not A268)  and  a64765a );
 a64767a <=( a64766a  and  a64761a );
 a64768a <=( a64767a  and  a64758a );
 a64771a <=( (not A167)  and  A170 );
 a64774a <=( A199  and  A166 );
 a64775a <=( a64774a  and  a64771a );
 a64778a <=( (not A201)  and  A200 );
 a64781a <=( A232  and  (not A202) );
 a64782a <=( a64781a  and  a64778a );
 a64783a <=( a64782a  and  a64775a );
 a64786a <=( (not A234)  and  A233 );
 a64789a <=( A265  and  (not A235) );
 a64790a <=( a64789a  and  a64786a );
 a64793a <=( (not A267)  and  A266 );
 a64797a <=( A300  and  A298 );
 a64798a <=( (not A268)  and  a64797a );
 a64799a <=( a64798a  and  a64793a );
 a64800a <=( a64799a  and  a64790a );
 a64803a <=( (not A167)  and  A170 );
 a64806a <=( A199  and  A166 );
 a64807a <=( a64806a  and  a64803a );
 a64810a <=( (not A201)  and  A200 );
 a64813a <=( A232  and  (not A202) );
 a64814a <=( a64813a  and  a64810a );
 a64815a <=( a64814a  and  a64807a );
 a64818a <=( (not A234)  and  A233 );
 a64821a <=( (not A265)  and  (not A235) );
 a64822a <=( a64821a  and  a64818a );
 a64825a <=( (not A268)  and  (not A266) );
 a64829a <=( A302  and  (not A299) );
 a64830a <=( A298  and  a64829a );
 a64831a <=( a64830a  and  a64825a );
 a64832a <=( a64831a  and  a64822a );
 a64835a <=( (not A167)  and  A170 );
 a64838a <=( A199  and  A166 );
 a64839a <=( a64838a  and  a64835a );
 a64842a <=( (not A201)  and  A200 );
 a64845a <=( A232  and  (not A202) );
 a64846a <=( a64845a  and  a64842a );
 a64847a <=( a64846a  and  a64839a );
 a64850a <=( (not A234)  and  A233 );
 a64853a <=( (not A265)  and  (not A235) );
 a64854a <=( a64853a  and  a64850a );
 a64857a <=( (not A268)  and  (not A266) );
 a64861a <=( A302  and  A299 );
 a64862a <=( (not A298)  and  a64861a );
 a64863a <=( a64862a  and  a64857a );
 a64864a <=( a64863a  and  a64854a );
 a64867a <=( (not A167)  and  A170 );
 a64870a <=( A199  and  A166 );
 a64871a <=( a64870a  and  a64867a );
 a64874a <=( (not A201)  and  A200 );
 a64877a <=( (not A232)  and  (not A202) );
 a64878a <=( a64877a  and  a64874a );
 a64879a <=( a64878a  and  a64871a );
 a64882a <=( (not A235)  and  (not A233) );
 a64885a <=( A266  and  A265 );
 a64886a <=( a64885a  and  a64882a );
 a64889a <=( (not A268)  and  (not A267) );
 a64893a <=( A302  and  (not A299) );
 a64894a <=( A298  and  a64893a );
 a64895a <=( a64894a  and  a64889a );
 a64896a <=( a64895a  and  a64886a );
 a64899a <=( (not A167)  and  A170 );
 a64902a <=( A199  and  A166 );
 a64903a <=( a64902a  and  a64899a );
 a64906a <=( (not A201)  and  A200 );
 a64909a <=( (not A232)  and  (not A202) );
 a64910a <=( a64909a  and  a64906a );
 a64911a <=( a64910a  and  a64903a );
 a64914a <=( (not A235)  and  (not A233) );
 a64917a <=( A266  and  A265 );
 a64918a <=( a64917a  and  a64914a );
 a64921a <=( (not A268)  and  (not A267) );
 a64925a <=( A302  and  A299 );
 a64926a <=( (not A298)  and  a64925a );
 a64927a <=( a64926a  and  a64921a );
 a64928a <=( a64927a  and  a64918a );
 a64931a <=( (not A167)  and  A170 );
 a64934a <=( (not A199)  and  A166 );
 a64935a <=( a64934a  and  a64931a );
 a64938a <=( (not A202)  and  (not A200) );
 a64941a <=( A233  and  A232 );
 a64942a <=( a64941a  and  a64938a );
 a64943a <=( a64942a  and  a64935a );
 a64946a <=( (not A235)  and  (not A234) );
 a64949a <=( A266  and  A265 );
 a64950a <=( a64949a  and  a64946a );
 a64953a <=( (not A268)  and  (not A267) );
 a64957a <=( A302  and  (not A299) );
 a64958a <=( A298  and  a64957a );
 a64959a <=( a64958a  and  a64953a );
 a64960a <=( a64959a  and  a64950a );
 a64963a <=( (not A167)  and  A170 );
 a64966a <=( (not A199)  and  A166 );
 a64967a <=( a64966a  and  a64963a );
 a64970a <=( (not A202)  and  (not A200) );
 a64973a <=( A233  and  A232 );
 a64974a <=( a64973a  and  a64970a );
 a64975a <=( a64974a  and  a64967a );
 a64978a <=( (not A235)  and  (not A234) );
 a64981a <=( A266  and  A265 );
 a64982a <=( a64981a  and  a64978a );
 a64985a <=( (not A268)  and  (not A267) );
 a64989a <=( A302  and  A299 );
 a64990a <=( (not A298)  and  a64989a );
 a64991a <=( a64990a  and  a64985a );
 a64992a <=( a64991a  and  a64982a );
 a64995a <=( (not A167)  and  (not A169) );
 a64998a <=( (not A199)  and  (not A166) );
 a64999a <=( a64998a  and  a64995a );
 a65002a <=( A203  and  A200 );
 a65005a <=( A233  and  A232 );
 a65006a <=( a65005a  and  a65002a );
 a65007a <=( a65006a  and  a64999a );
 a65010a <=( (not A235)  and  (not A234) );
 a65013a <=( A266  and  A265 );
 a65014a <=( a65013a  and  a65010a );
 a65017a <=( (not A268)  and  (not A267) );
 a65021a <=( A302  and  (not A299) );
 a65022a <=( A298  and  a65021a );
 a65023a <=( a65022a  and  a65017a );
 a65024a <=( a65023a  and  a65014a );
 a65027a <=( (not A167)  and  (not A169) );
 a65030a <=( (not A199)  and  (not A166) );
 a65031a <=( a65030a  and  a65027a );
 a65034a <=( A203  and  A200 );
 a65037a <=( A233  and  A232 );
 a65038a <=( a65037a  and  a65034a );
 a65039a <=( a65038a  and  a65031a );
 a65042a <=( (not A235)  and  (not A234) );
 a65045a <=( A266  and  A265 );
 a65046a <=( a65045a  and  a65042a );
 a65049a <=( (not A268)  and  (not A267) );
 a65053a <=( A302  and  A299 );
 a65054a <=( (not A298)  and  a65053a );
 a65055a <=( a65054a  and  a65049a );
 a65056a <=( a65055a  and  a65046a );
 a65059a <=( (not A167)  and  (not A169) );
 a65062a <=( A199  and  (not A166) );
 a65063a <=( a65062a  and  a65059a );
 a65066a <=( A203  and  (not A200) );
 a65069a <=( A233  and  A232 );
 a65070a <=( a65069a  and  a65066a );
 a65071a <=( a65070a  and  a65063a );
 a65074a <=( (not A235)  and  (not A234) );
 a65077a <=( A266  and  A265 );
 a65078a <=( a65077a  and  a65074a );
 a65081a <=( (not A268)  and  (not A267) );
 a65085a <=( A302  and  (not A299) );
 a65086a <=( A298  and  a65085a );
 a65087a <=( a65086a  and  a65081a );
 a65088a <=( a65087a  and  a65078a );
 a65091a <=( (not A167)  and  (not A169) );
 a65094a <=( A199  and  (not A166) );
 a65095a <=( a65094a  and  a65091a );
 a65098a <=( A203  and  (not A200) );
 a65101a <=( A233  and  A232 );
 a65102a <=( a65101a  and  a65098a );
 a65103a <=( a65102a  and  a65095a );
 a65106a <=( (not A235)  and  (not A234) );
 a65109a <=( A266  and  A265 );
 a65110a <=( a65109a  and  a65106a );
 a65113a <=( (not A268)  and  (not A267) );
 a65117a <=( A302  and  A299 );
 a65118a <=( (not A298)  and  a65117a );
 a65119a <=( a65118a  and  a65113a );
 a65120a <=( a65119a  and  a65110a );
 a65123a <=( (not A168)  and  (not A169) );
 a65126a <=( A166  and  A167 );
 a65127a <=( a65126a  and  a65123a );
 a65130a <=( A201  and  A199 );
 a65133a <=( A233  and  A232 );
 a65134a <=( a65133a  and  a65130a );
 a65135a <=( a65134a  and  a65127a );
 a65138a <=( (not A235)  and  (not A234) );
 a65141a <=( A266  and  A265 );
 a65142a <=( a65141a  and  a65138a );
 a65145a <=( (not A268)  and  (not A267) );
 a65149a <=( A302  and  (not A299) );
 a65150a <=( A298  and  a65149a );
 a65151a <=( a65150a  and  a65145a );
 a65152a <=( a65151a  and  a65142a );
 a65155a <=( (not A168)  and  (not A169) );
 a65158a <=( A166  and  A167 );
 a65159a <=( a65158a  and  a65155a );
 a65162a <=( A201  and  A199 );
 a65165a <=( A233  and  A232 );
 a65166a <=( a65165a  and  a65162a );
 a65167a <=( a65166a  and  a65159a );
 a65170a <=( (not A235)  and  (not A234) );
 a65173a <=( A266  and  A265 );
 a65174a <=( a65173a  and  a65170a );
 a65177a <=( (not A268)  and  (not A267) );
 a65181a <=( A302  and  A299 );
 a65182a <=( (not A298)  and  a65181a );
 a65183a <=( a65182a  and  a65177a );
 a65184a <=( a65183a  and  a65174a );
 a65187a <=( (not A168)  and  (not A169) );
 a65190a <=( A166  and  A167 );
 a65191a <=( a65190a  and  a65187a );
 a65194a <=( A201  and  A200 );
 a65197a <=( A233  and  A232 );
 a65198a <=( a65197a  and  a65194a );
 a65199a <=( a65198a  and  a65191a );
 a65202a <=( (not A235)  and  (not A234) );
 a65205a <=( A266  and  A265 );
 a65206a <=( a65205a  and  a65202a );
 a65209a <=( (not A268)  and  (not A267) );
 a65213a <=( A302  and  (not A299) );
 a65214a <=( A298  and  a65213a );
 a65215a <=( a65214a  and  a65209a );
 a65216a <=( a65215a  and  a65206a );
 a65219a <=( (not A168)  and  (not A169) );
 a65222a <=( A166  and  A167 );
 a65223a <=( a65222a  and  a65219a );
 a65226a <=( A201  and  A200 );
 a65229a <=( A233  and  A232 );
 a65230a <=( a65229a  and  a65226a );
 a65231a <=( a65230a  and  a65223a );
 a65234a <=( (not A235)  and  (not A234) );
 a65237a <=( A266  and  A265 );
 a65238a <=( a65237a  and  a65234a );
 a65241a <=( (not A268)  and  (not A267) );
 a65245a <=( A302  and  A299 );
 a65246a <=( (not A298)  and  a65245a );
 a65247a <=( a65246a  and  a65241a );
 a65248a <=( a65247a  and  a65238a );
 a65251a <=( (not A168)  and  (not A169) );
 a65254a <=( A166  and  A167 );
 a65255a <=( a65254a  and  a65251a );
 a65258a <=( A200  and  (not A199) );
 a65261a <=( (not A234)  and  A203 );
 a65262a <=( a65261a  and  a65258a );
 a65263a <=( a65262a  and  a65255a );
 a65266a <=( (not A236)  and  (not A235) );
 a65269a <=( A266  and  A265 );
 a65270a <=( a65269a  and  a65266a );
 a65273a <=( (not A268)  and  (not A267) );
 a65277a <=( A302  and  (not A299) );
 a65278a <=( A298  and  a65277a );
 a65279a <=( a65278a  and  a65273a );
 a65280a <=( a65279a  and  a65270a );
 a65283a <=( (not A168)  and  (not A169) );
 a65286a <=( A166  and  A167 );
 a65287a <=( a65286a  and  a65283a );
 a65290a <=( A200  and  (not A199) );
 a65293a <=( (not A234)  and  A203 );
 a65294a <=( a65293a  and  a65290a );
 a65295a <=( a65294a  and  a65287a );
 a65298a <=( (not A236)  and  (not A235) );
 a65301a <=( A266  and  A265 );
 a65302a <=( a65301a  and  a65298a );
 a65305a <=( (not A268)  and  (not A267) );
 a65309a <=( A302  and  A299 );
 a65310a <=( (not A298)  and  a65309a );
 a65311a <=( a65310a  and  a65305a );
 a65312a <=( a65311a  and  a65302a );
 a65315a <=( (not A168)  and  (not A169) );
 a65318a <=( A166  and  A167 );
 a65319a <=( a65318a  and  a65315a );
 a65322a <=( A200  and  (not A199) );
 a65325a <=( A232  and  A203 );
 a65326a <=( a65325a  and  a65322a );
 a65327a <=( a65326a  and  a65319a );
 a65330a <=( (not A234)  and  A233 );
 a65333a <=( (not A267)  and  (not A235) );
 a65334a <=( a65333a  and  a65330a );
 a65337a <=( (not A269)  and  (not A268) );
 a65341a <=( A302  and  (not A299) );
 a65342a <=( A298  and  a65341a );
 a65343a <=( a65342a  and  a65337a );
 a65344a <=( a65343a  and  a65334a );
 a65347a <=( (not A168)  and  (not A169) );
 a65350a <=( A166  and  A167 );
 a65351a <=( a65350a  and  a65347a );
 a65354a <=( A200  and  (not A199) );
 a65357a <=( A232  and  A203 );
 a65358a <=( a65357a  and  a65354a );
 a65359a <=( a65358a  and  a65351a );
 a65362a <=( (not A234)  and  A233 );
 a65365a <=( (not A267)  and  (not A235) );
 a65366a <=( a65365a  and  a65362a );
 a65369a <=( (not A269)  and  (not A268) );
 a65373a <=( A302  and  A299 );
 a65374a <=( (not A298)  and  a65373a );
 a65375a <=( a65374a  and  a65369a );
 a65376a <=( a65375a  and  a65366a );
 a65379a <=( (not A168)  and  (not A169) );
 a65382a <=( A166  and  A167 );
 a65383a <=( a65382a  and  a65379a );
 a65386a <=( A200  and  (not A199) );
 a65389a <=( A232  and  A203 );
 a65390a <=( a65389a  and  a65386a );
 a65391a <=( a65390a  and  a65383a );
 a65394a <=( (not A234)  and  A233 );
 a65397a <=( A265  and  (not A235) );
 a65398a <=( a65397a  and  a65394a );
 a65401a <=( (not A267)  and  A266 );
 a65405a <=( A300  and  A299 );
 a65406a <=( (not A268)  and  a65405a );
 a65407a <=( a65406a  and  a65401a );
 a65408a <=( a65407a  and  a65398a );
 a65411a <=( (not A168)  and  (not A169) );
 a65414a <=( A166  and  A167 );
 a65415a <=( a65414a  and  a65411a );
 a65418a <=( A200  and  (not A199) );
 a65421a <=( A232  and  A203 );
 a65422a <=( a65421a  and  a65418a );
 a65423a <=( a65422a  and  a65415a );
 a65426a <=( (not A234)  and  A233 );
 a65429a <=( A265  and  (not A235) );
 a65430a <=( a65429a  and  a65426a );
 a65433a <=( (not A267)  and  A266 );
 a65437a <=( A300  and  A298 );
 a65438a <=( (not A268)  and  a65437a );
 a65439a <=( a65438a  and  a65433a );
 a65440a <=( a65439a  and  a65430a );
 a65443a <=( (not A168)  and  (not A169) );
 a65446a <=( A166  and  A167 );
 a65447a <=( a65446a  and  a65443a );
 a65450a <=( A200  and  (not A199) );
 a65453a <=( A232  and  A203 );
 a65454a <=( a65453a  and  a65450a );
 a65455a <=( a65454a  and  a65447a );
 a65458a <=( (not A234)  and  A233 );
 a65461a <=( (not A265)  and  (not A235) );
 a65462a <=( a65461a  and  a65458a );
 a65465a <=( (not A268)  and  (not A266) );
 a65469a <=( A302  and  (not A299) );
 a65470a <=( A298  and  a65469a );
 a65471a <=( a65470a  and  a65465a );
 a65472a <=( a65471a  and  a65462a );
 a65475a <=( (not A168)  and  (not A169) );
 a65478a <=( A166  and  A167 );
 a65479a <=( a65478a  and  a65475a );
 a65482a <=( A200  and  (not A199) );
 a65485a <=( A232  and  A203 );
 a65486a <=( a65485a  and  a65482a );
 a65487a <=( a65486a  and  a65479a );
 a65490a <=( (not A234)  and  A233 );
 a65493a <=( (not A265)  and  (not A235) );
 a65494a <=( a65493a  and  a65490a );
 a65497a <=( (not A268)  and  (not A266) );
 a65501a <=( A302  and  A299 );
 a65502a <=( (not A298)  and  a65501a );
 a65503a <=( a65502a  and  a65497a );
 a65504a <=( a65503a  and  a65494a );
 a65507a <=( (not A168)  and  (not A169) );
 a65510a <=( A166  and  A167 );
 a65511a <=( a65510a  and  a65507a );
 a65514a <=( A200  and  (not A199) );
 a65517a <=( (not A232)  and  A203 );
 a65518a <=( a65517a  and  a65514a );
 a65519a <=( a65518a  and  a65511a );
 a65522a <=( (not A235)  and  (not A233) );
 a65525a <=( A266  and  A265 );
 a65526a <=( a65525a  and  a65522a );
 a65529a <=( (not A268)  and  (not A267) );
 a65533a <=( A302  and  (not A299) );
 a65534a <=( A298  and  a65533a );
 a65535a <=( a65534a  and  a65529a );
 a65536a <=( a65535a  and  a65526a );
 a65539a <=( (not A168)  and  (not A169) );
 a65542a <=( A166  and  A167 );
 a65543a <=( a65542a  and  a65539a );
 a65546a <=( A200  and  (not A199) );
 a65549a <=( (not A232)  and  A203 );
 a65550a <=( a65549a  and  a65546a );
 a65551a <=( a65550a  and  a65543a );
 a65554a <=( (not A235)  and  (not A233) );
 a65557a <=( A266  and  A265 );
 a65558a <=( a65557a  and  a65554a );
 a65561a <=( (not A268)  and  (not A267) );
 a65565a <=( A302  and  A299 );
 a65566a <=( (not A298)  and  a65565a );
 a65567a <=( a65566a  and  a65561a );
 a65568a <=( a65567a  and  a65558a );
 a65571a <=( (not A168)  and  (not A169) );
 a65574a <=( A166  and  A167 );
 a65575a <=( a65574a  and  a65571a );
 a65578a <=( (not A200)  and  A199 );
 a65581a <=( (not A234)  and  A203 );
 a65582a <=( a65581a  and  a65578a );
 a65583a <=( a65582a  and  a65575a );
 a65586a <=( (not A236)  and  (not A235) );
 a65589a <=( A266  and  A265 );
 a65590a <=( a65589a  and  a65586a );
 a65593a <=( (not A268)  and  (not A267) );
 a65597a <=( A302  and  (not A299) );
 a65598a <=( A298  and  a65597a );
 a65599a <=( a65598a  and  a65593a );
 a65600a <=( a65599a  and  a65590a );
 a65603a <=( (not A168)  and  (not A169) );
 a65606a <=( A166  and  A167 );
 a65607a <=( a65606a  and  a65603a );
 a65610a <=( (not A200)  and  A199 );
 a65613a <=( (not A234)  and  A203 );
 a65614a <=( a65613a  and  a65610a );
 a65615a <=( a65614a  and  a65607a );
 a65618a <=( (not A236)  and  (not A235) );
 a65621a <=( A266  and  A265 );
 a65622a <=( a65621a  and  a65618a );
 a65625a <=( (not A268)  and  (not A267) );
 a65629a <=( A302  and  A299 );
 a65630a <=( (not A298)  and  a65629a );
 a65631a <=( a65630a  and  a65625a );
 a65632a <=( a65631a  and  a65622a );
 a65635a <=( (not A168)  and  (not A169) );
 a65638a <=( A166  and  A167 );
 a65639a <=( a65638a  and  a65635a );
 a65642a <=( (not A200)  and  A199 );
 a65645a <=( A232  and  A203 );
 a65646a <=( a65645a  and  a65642a );
 a65647a <=( a65646a  and  a65639a );
 a65650a <=( (not A234)  and  A233 );
 a65653a <=( (not A267)  and  (not A235) );
 a65654a <=( a65653a  and  a65650a );
 a65657a <=( (not A269)  and  (not A268) );
 a65661a <=( A302  and  (not A299) );
 a65662a <=( A298  and  a65661a );
 a65663a <=( a65662a  and  a65657a );
 a65664a <=( a65663a  and  a65654a );
 a65667a <=( (not A168)  and  (not A169) );
 a65670a <=( A166  and  A167 );
 a65671a <=( a65670a  and  a65667a );
 a65674a <=( (not A200)  and  A199 );
 a65677a <=( A232  and  A203 );
 a65678a <=( a65677a  and  a65674a );
 a65679a <=( a65678a  and  a65671a );
 a65682a <=( (not A234)  and  A233 );
 a65685a <=( (not A267)  and  (not A235) );
 a65686a <=( a65685a  and  a65682a );
 a65689a <=( (not A269)  and  (not A268) );
 a65693a <=( A302  and  A299 );
 a65694a <=( (not A298)  and  a65693a );
 a65695a <=( a65694a  and  a65689a );
 a65696a <=( a65695a  and  a65686a );
 a65699a <=( (not A168)  and  (not A169) );
 a65702a <=( A166  and  A167 );
 a65703a <=( a65702a  and  a65699a );
 a65706a <=( (not A200)  and  A199 );
 a65709a <=( A232  and  A203 );
 a65710a <=( a65709a  and  a65706a );
 a65711a <=( a65710a  and  a65703a );
 a65714a <=( (not A234)  and  A233 );
 a65717a <=( A265  and  (not A235) );
 a65718a <=( a65717a  and  a65714a );
 a65721a <=( (not A267)  and  A266 );
 a65725a <=( A300  and  A299 );
 a65726a <=( (not A268)  and  a65725a );
 a65727a <=( a65726a  and  a65721a );
 a65728a <=( a65727a  and  a65718a );
 a65731a <=( (not A168)  and  (not A169) );
 a65734a <=( A166  and  A167 );
 a65735a <=( a65734a  and  a65731a );
 a65738a <=( (not A200)  and  A199 );
 a65741a <=( A232  and  A203 );
 a65742a <=( a65741a  and  a65738a );
 a65743a <=( a65742a  and  a65735a );
 a65746a <=( (not A234)  and  A233 );
 a65749a <=( A265  and  (not A235) );
 a65750a <=( a65749a  and  a65746a );
 a65753a <=( (not A267)  and  A266 );
 a65757a <=( A300  and  A298 );
 a65758a <=( (not A268)  and  a65757a );
 a65759a <=( a65758a  and  a65753a );
 a65760a <=( a65759a  and  a65750a );
 a65763a <=( (not A168)  and  (not A169) );
 a65766a <=( A166  and  A167 );
 a65767a <=( a65766a  and  a65763a );
 a65770a <=( (not A200)  and  A199 );
 a65773a <=( A232  and  A203 );
 a65774a <=( a65773a  and  a65770a );
 a65775a <=( a65774a  and  a65767a );
 a65778a <=( (not A234)  and  A233 );
 a65781a <=( (not A265)  and  (not A235) );
 a65782a <=( a65781a  and  a65778a );
 a65785a <=( (not A268)  and  (not A266) );
 a65789a <=( A302  and  (not A299) );
 a65790a <=( A298  and  a65789a );
 a65791a <=( a65790a  and  a65785a );
 a65792a <=( a65791a  and  a65782a );
 a65795a <=( (not A168)  and  (not A169) );
 a65798a <=( A166  and  A167 );
 a65799a <=( a65798a  and  a65795a );
 a65802a <=( (not A200)  and  A199 );
 a65805a <=( A232  and  A203 );
 a65806a <=( a65805a  and  a65802a );
 a65807a <=( a65806a  and  a65799a );
 a65810a <=( (not A234)  and  A233 );
 a65813a <=( (not A265)  and  (not A235) );
 a65814a <=( a65813a  and  a65810a );
 a65817a <=( (not A268)  and  (not A266) );
 a65821a <=( A302  and  A299 );
 a65822a <=( (not A298)  and  a65821a );
 a65823a <=( a65822a  and  a65817a );
 a65824a <=( a65823a  and  a65814a );
 a65827a <=( (not A168)  and  (not A169) );
 a65830a <=( A166  and  A167 );
 a65831a <=( a65830a  and  a65827a );
 a65834a <=( (not A200)  and  A199 );
 a65837a <=( (not A232)  and  A203 );
 a65838a <=( a65837a  and  a65834a );
 a65839a <=( a65838a  and  a65831a );
 a65842a <=( (not A235)  and  (not A233) );
 a65845a <=( A266  and  A265 );
 a65846a <=( a65845a  and  a65842a );
 a65849a <=( (not A268)  and  (not A267) );
 a65853a <=( A302  and  (not A299) );
 a65854a <=( A298  and  a65853a );
 a65855a <=( a65854a  and  a65849a );
 a65856a <=( a65855a  and  a65846a );
 a65859a <=( (not A168)  and  (not A169) );
 a65862a <=( A166  and  A167 );
 a65863a <=( a65862a  and  a65859a );
 a65866a <=( (not A200)  and  A199 );
 a65869a <=( (not A232)  and  A203 );
 a65870a <=( a65869a  and  a65866a );
 a65871a <=( a65870a  and  a65863a );
 a65874a <=( (not A235)  and  (not A233) );
 a65877a <=( A266  and  A265 );
 a65878a <=( a65877a  and  a65874a );
 a65881a <=( (not A268)  and  (not A267) );
 a65885a <=( A302  and  A299 );
 a65886a <=( (not A298)  and  a65885a );
 a65887a <=( a65886a  and  a65881a );
 a65888a <=( a65887a  and  a65878a );
 a65891a <=( (not A169)  and  (not A170) );
 a65894a <=( (not A199)  and  (not A168) );
 a65895a <=( a65894a  and  a65891a );
 a65898a <=( A203  and  A200 );
 a65901a <=( A233  and  A232 );
 a65902a <=( a65901a  and  a65898a );
 a65903a <=( a65902a  and  a65895a );
 a65906a <=( (not A235)  and  (not A234) );
 a65909a <=( A266  and  A265 );
 a65910a <=( a65909a  and  a65906a );
 a65913a <=( (not A268)  and  (not A267) );
 a65917a <=( A302  and  (not A299) );
 a65918a <=( A298  and  a65917a );
 a65919a <=( a65918a  and  a65913a );
 a65920a <=( a65919a  and  a65910a );
 a65923a <=( (not A169)  and  (not A170) );
 a65926a <=( (not A199)  and  (not A168) );
 a65927a <=( a65926a  and  a65923a );
 a65930a <=( A203  and  A200 );
 a65933a <=( A233  and  A232 );
 a65934a <=( a65933a  and  a65930a );
 a65935a <=( a65934a  and  a65927a );
 a65938a <=( (not A235)  and  (not A234) );
 a65941a <=( A266  and  A265 );
 a65942a <=( a65941a  and  a65938a );
 a65945a <=( (not A268)  and  (not A267) );
 a65949a <=( A302  and  A299 );
 a65950a <=( (not A298)  and  a65949a );
 a65951a <=( a65950a  and  a65945a );
 a65952a <=( a65951a  and  a65942a );
 a65955a <=( (not A169)  and  (not A170) );
 a65958a <=( A199  and  (not A168) );
 a65959a <=( a65958a  and  a65955a );
 a65962a <=( A203  and  (not A200) );
 a65965a <=( A233  and  A232 );
 a65966a <=( a65965a  and  a65962a );
 a65967a <=( a65966a  and  a65959a );
 a65970a <=( (not A235)  and  (not A234) );
 a65973a <=( A266  and  A265 );
 a65974a <=( a65973a  and  a65970a );
 a65977a <=( (not A268)  and  (not A267) );
 a65981a <=( A302  and  (not A299) );
 a65982a <=( A298  and  a65981a );
 a65983a <=( a65982a  and  a65977a );
 a65984a <=( a65983a  and  a65974a );
 a65987a <=( (not A169)  and  (not A170) );
 a65990a <=( A199  and  (not A168) );
 a65991a <=( a65990a  and  a65987a );
 a65994a <=( A203  and  (not A200) );
 a65997a <=( A233  and  A232 );
 a65998a <=( a65997a  and  a65994a );
 a65999a <=( a65998a  and  a65991a );
 a66002a <=( (not A235)  and  (not A234) );
 a66005a <=( A266  and  A265 );
 a66006a <=( a66005a  and  a66002a );
 a66009a <=( (not A268)  and  (not A267) );
 a66013a <=( A302  and  A299 );
 a66014a <=( (not A298)  and  a66013a );
 a66015a <=( a66014a  and  a66009a );
 a66016a <=( a66015a  and  a66006a );
 a66019a <=( A167  and  A170 );
 a66022a <=( A199  and  (not A166) );
 a66023a <=( a66022a  and  a66019a );
 a66026a <=( (not A201)  and  A200 );
 a66030a <=( A233  and  A232 );
 a66031a <=( (not A202)  and  a66030a );
 a66032a <=( a66031a  and  a66026a );
 a66033a <=( a66032a  and  a66023a );
 a66036a <=( (not A235)  and  (not A234) );
 a66039a <=( A266  and  A265 );
 a66040a <=( a66039a  and  a66036a );
 a66043a <=( (not A268)  and  (not A267) );
 a66047a <=( A302  and  (not A299) );
 a66048a <=( A298  and  a66047a );
 a66049a <=( a66048a  and  a66043a );
 a66050a <=( a66049a  and  a66040a );
 a66053a <=( A167  and  A170 );
 a66056a <=( A199  and  (not A166) );
 a66057a <=( a66056a  and  a66053a );
 a66060a <=( (not A201)  and  A200 );
 a66064a <=( A233  and  A232 );
 a66065a <=( (not A202)  and  a66064a );
 a66066a <=( a66065a  and  a66060a );
 a66067a <=( a66066a  and  a66057a );
 a66070a <=( (not A235)  and  (not A234) );
 a66073a <=( A266  and  A265 );
 a66074a <=( a66073a  and  a66070a );
 a66077a <=( (not A268)  and  (not A267) );
 a66081a <=( A302  and  A299 );
 a66082a <=( (not A298)  and  a66081a );
 a66083a <=( a66082a  and  a66077a );
 a66084a <=( a66083a  and  a66074a );
 a66087a <=( (not A167)  and  A170 );
 a66090a <=( A199  and  A166 );
 a66091a <=( a66090a  and  a66087a );
 a66094a <=( (not A201)  and  A200 );
 a66098a <=( A233  and  A232 );
 a66099a <=( (not A202)  and  a66098a );
 a66100a <=( a66099a  and  a66094a );
 a66101a <=( a66100a  and  a66091a );
 a66104a <=( (not A235)  and  (not A234) );
 a66107a <=( A266  and  A265 );
 a66108a <=( a66107a  and  a66104a );
 a66111a <=( (not A268)  and  (not A267) );
 a66115a <=( A302  and  (not A299) );
 a66116a <=( A298  and  a66115a );
 a66117a <=( a66116a  and  a66111a );
 a66118a <=( a66117a  and  a66108a );
 a66121a <=( (not A167)  and  A170 );
 a66124a <=( A199  and  A166 );
 a66125a <=( a66124a  and  a66121a );
 a66128a <=( (not A201)  and  A200 );
 a66132a <=( A233  and  A232 );
 a66133a <=( (not A202)  and  a66132a );
 a66134a <=( a66133a  and  a66128a );
 a66135a <=( a66134a  and  a66125a );
 a66138a <=( (not A235)  and  (not A234) );
 a66141a <=( A266  and  A265 );
 a66142a <=( a66141a  and  a66138a );
 a66145a <=( (not A268)  and  (not A267) );
 a66149a <=( A302  and  A299 );
 a66150a <=( (not A298)  and  a66149a );
 a66151a <=( a66150a  and  a66145a );
 a66152a <=( a66151a  and  a66142a );
 a66155a <=( (not A168)  and  (not A169) );
 a66158a <=( A166  and  A167 );
 a66159a <=( a66158a  and  a66155a );
 a66162a <=( A200  and  (not A199) );
 a66166a <=( A233  and  A232 );
 a66167a <=( A203  and  a66166a );
 a66168a <=( a66167a  and  a66162a );
 a66169a <=( a66168a  and  a66159a );
 a66172a <=( (not A235)  and  (not A234) );
 a66175a <=( A266  and  A265 );
 a66176a <=( a66175a  and  a66172a );
 a66179a <=( (not A268)  and  (not A267) );
 a66183a <=( A302  and  (not A299) );
 a66184a <=( A298  and  a66183a );
 a66185a <=( a66184a  and  a66179a );
 a66186a <=( a66185a  and  a66176a );
 a66189a <=( (not A168)  and  (not A169) );
 a66192a <=( A166  and  A167 );
 a66193a <=( a66192a  and  a66189a );
 a66196a <=( A200  and  (not A199) );
 a66200a <=( A233  and  A232 );
 a66201a <=( A203  and  a66200a );
 a66202a <=( a66201a  and  a66196a );
 a66203a <=( a66202a  and  a66193a );
 a66206a <=( (not A235)  and  (not A234) );
 a66209a <=( A266  and  A265 );
 a66210a <=( a66209a  and  a66206a );
 a66213a <=( (not A268)  and  (not A267) );
 a66217a <=( A302  and  A299 );
 a66218a <=( (not A298)  and  a66217a );
 a66219a <=( a66218a  and  a66213a );
 a66220a <=( a66219a  and  a66210a );
 a66223a <=( (not A168)  and  (not A169) );
 a66226a <=( A166  and  A167 );
 a66227a <=( a66226a  and  a66223a );
 a66230a <=( (not A200)  and  A199 );
 a66234a <=( A233  and  A232 );
 a66235a <=( A203  and  a66234a );
 a66236a <=( a66235a  and  a66230a );
 a66237a <=( a66236a  and  a66227a );
 a66240a <=( (not A235)  and  (not A234) );
 a66243a <=( A266  and  A265 );
 a66244a <=( a66243a  and  a66240a );
 a66247a <=( (not A268)  and  (not A267) );
 a66251a <=( A302  and  (not A299) );
 a66252a <=( A298  and  a66251a );
 a66253a <=( a66252a  and  a66247a );
 a66254a <=( a66253a  and  a66244a );
 a66257a <=( (not A168)  and  (not A169) );
 a66260a <=( A166  and  A167 );
 a66261a <=( a66260a  and  a66257a );
 a66264a <=( (not A200)  and  A199 );
 a66268a <=( A233  and  A232 );
 a66269a <=( A203  and  a66268a );
 a66270a <=( a66269a  and  a66264a );
 a66271a <=( a66270a  and  a66261a );
 a66274a <=( (not A235)  and  (not A234) );
 a66277a <=( A266  and  A265 );
 a66278a <=( a66277a  and  a66274a );
 a66281a <=( (not A268)  and  (not A267) );
 a66285a <=( A302  and  A299 );
 a66286a <=( (not A298)  and  a66285a );
 a66287a <=( a66286a  and  a66281a );
 a66288a <=( a66287a  and  a66278a );


end x25_15x_behav;
