Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_13x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A74: buffer std_logic
);
end x25_13x;

architecture x25_13x_behav of x25_13x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a209a,a210a,a214a,a215a,a216a,a220a,a221a,a225a,a226a,a227a,a228a,a232a,a233a,a237a,a238a,a239a,a243a,a244a,a247a,a250a,a251a,a252a,a253a,a254a,a258a,a259a,a263a,a264a,a265a,a269a,a270a,a273a,a276a,a277a,a278a,a279a,a283a,a284a,a288a,a289a,a290a,a294a,a295a,a298a,a301a,a302a,a303a,a304a,a305a,a306a,a310a,a311a,a315a,a316a,a317a,a321a,a322a,a326a,a327a,a328a,a329a,a333a,a334a,a338a,a339a,a340a,a344a,a345a,a348a,a351a,a352a,a353a,a354a,a355a,a359a,a360a,a364a,a365a,a366a,a370a,a371a,a374a,a377a,a378a,a379a,a380a,a384a,a385a,a389a,a390a,a391a,a395a,a396a,a399a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a412a,a413a,a417a,a418a,a419a,a423a,a424a,a428a,a429a,a430a,a431a,a435a,a436a,a440a,a441a,a442a,a446a,a447a,a450a,a453a,a454a,a455a,a456a,a457a,a461a,a462a,a466a,a467a,a468a,a472a,a473a,a476a,a479a,a480a,a481a,a482a,a486a,a487a,a491a,a492a,a493a,a497a,a498a,a501a,a504a,a505a,a506a,a507a,a508a,a509a,a513a,a514a,a518a,a519a,a520a,a524a,a525a,a528a,a531a,a532a,a533a,a534a,a538a,a539a,a543a,a544a,a545a,a549a,a550a,a553a,a556a,a557a,a558a,a559a,a560a,a564a,a565a,a569a,a570a,a571a,a575a,a576a,a579a,a582a,a583a,a584a,a585a,a589a,a590a,a594a,a595a,a596a,a600a,a601a,a604a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a625a,a629a,a633a,a637a,a641a,a645a,a649a,a653a,a657a,a661a,a664a,a667a,a670a,a673a,a676a,a679a,a682a,a685a,a688a,a691a,a694a,a697a,a700a,a703a,a706a,a709a,a712a,a715a,a718a,a721a,a724a,a727a,a730a,a733a,a736a,a739a,a742a,a745a,a748a,a751a,a754a,a757a,a760a,a764a,a765a,a768a,a772a,a773a,a776a,a780a,a781a,a784a,a788a,a789a,a792a,a796a,a797a,a800a,a804a,a805a,a808a,a812a,a813a,a816a,a820a,a821a,a824a,a828a,a829a,a832a,a836a,a837a,a840a,a844a,a845a,a848a,a852a,a853a,a856a,a860a,a861a,a864a,a868a,a869a,a872a,a876a,a877a,a880a,a884a,a885a,a888a,a892a,a893a,a896a,a900a,a901a,a904a,a908a,a909a,a912a,a916a,a917a,a921a,a922a,a926a,a927a,a931a,a932a,a936a,a937a,a941a,a942a,a946a,a947a,a951a,a952a,a956a,a957a,a961a,a962a,a966a,a967a,a971a,a972a,a976a,a977a,a981a,a982a,a986a,a987a,a991a,a992a,a996a,a997a,a1001a,a1002a,a1006a,a1007a,a1011a,a1012a,a1016a,a1017a,a1021a,a1022a,a1026a,a1027a,a1031a,a1032a,a1036a,a1037a,a1041a,a1042a,a1046a,a1047a,a1051a,a1052a,a1056a,a1057a,a1061a,a1062a,a1066a,a1067a,a1071a,a1072a,a1076a,a1077a,a1081a,a1082a,a1086a,a1087a,a1091a,a1092a,a1096a,a1097a,a1101a,a1102a,a1106a,a1107a,a1111a,a1112a,a1116a,a1117a,a1121a,a1122a,a1126a,a1127a,a1131a,a1132a,a1136a,a1137a,a1141a,a1142a,a1146a,a1147a,a1151a,a1152a,a1156a,a1157a,a1161a,a1162a,a1166a,a1167a,a1171a,a1172a,a1176a,a1177a,a1181a,a1182a,a1185a,a1188a,a1189a,a1193a,a1194a,a1197a,a1200a,a1201a,a1205a,a1206a,a1209a,a1212a,a1213a,a1217a,a1218a,a1221a,a1224a,a1225a,a1229a,a1230a,a1233a,a1236a,a1237a,a1241a,a1242a,a1245a,a1248a,a1249a,a1253a,a1254a,a1257a,a1260a,a1261a,a1265a,a1266a,a1269a,a1272a,a1273a,a1277a,a1278a,a1281a,a1284a,a1285a,a1289a,a1290a,a1293a,a1296a,a1297a,a1301a,a1302a,a1305a,a1308a,a1309a,a1313a,a1314a,a1317a,a1320a,a1321a,a1325a,a1326a,a1329a,a1332a,a1333a,a1337a,a1338a,a1341a,a1344a,a1345a,a1349a,a1350a,a1353a,a1356a,a1357a,a1361a,a1362a,a1365a,a1368a,a1369a,a1373a,a1374a,a1377a,a1380a,a1381a,a1385a,a1386a,a1389a,a1392a,a1393a,a1397a,a1398a,a1401a,a1404a,a1405a,a1409a,a1410a,a1413a,a1416a,a1417a,a1421a,a1422a,a1425a,a1428a,a1429a,a1433a,a1434a,a1437a,a1440a,a1441a,a1445a,a1446a,a1449a,a1452a,a1453a,a1457a,a1458a,a1461a,a1464a,a1465a,a1469a,a1470a,a1473a,a1476a,a1477a,a1481a,a1482a,a1485a,a1488a,a1489a,a1493a,a1494a,a1497a,a1500a,a1501a,a1505a,a1506a,a1509a,a1512a,a1513a,a1517a,a1518a,a1521a,a1524a,a1525a,a1529a,a1530a,a1533a,a1536a,a1537a,a1541a,a1542a,a1545a,a1548a,a1549a,a1553a,a1554a,a1557a,a1560a,a1561a,a1565a,a1566a,a1569a,a1572a,a1573a,a1577a,a1578a,a1581a,a1584a,a1585a,a1589a,a1590a,a1593a,a1596a,a1597a,a1601a,a1602a,a1605a,a1608a,a1609a,a1613a,a1614a,a1617a,a1620a,a1621a,a1625a,a1626a,a1629a,a1632a,a1633a,a1637a,a1638a,a1641a,a1644a,a1645a,a1649a,a1650a,a1653a,a1656a,a1657a,a1660a,a1663a,a1664a,a1667a,a1670a,a1671a,a1674a,a1677a,a1678a,a1681a,a1684a,a1685a,a1688a,a1691a,a1692a,a1695a,a1698a,a1699a,a1702a,a1705a,a1706a,a1709a,a1712a,a1713a,a1716a,a1719a,a1720a,a1723a,a1726a,a1727a,a1730a,a1733a,a1734a,a1737a,a1740a,a1741a,a1744a,a1747a,a1748a,a1751a,a1754a,a1755a,a1758a,a1761a,a1762a,a1765a,a1768a,a1769a,a1772a,a1775a,a1776a,a1779a,a1782a,a1783a,a1786a,a1789a,a1790a,a1793a,a1796a,a1797a,a1800a,a1803a,a1804a,a1807a,a1810a,a1811a,a1814a,a1817a,a1818a,a1821a,a1824a,a1825a,a1828a,a1831a,a1832a,a1835a,a1838a,a1839a,a1842a,a1845a,a1846a,a1849a,a1852a,a1853a,a1856a,a1859a,a1860a,a1863a,a1866a,a1867a,a1870a,a1873a,a1874a,a1877a,a1880a,a1881a,a1884a,a1887a,a1888a,a1891a,a1894a,a1895a,a1898a,a1901a,a1902a,a1905a,a1908a,a1909a,a1912a,a1915a,a1916a,a1919a,a1922a,a1923a,a1926a,a1929a,a1930a,a1933a,a1936a,a1937a,a1940a,a1943a,a1944a,a1947a,a1950a,a1951a,a1954a,a1957a,a1958a,a1961a,a1964a,a1965a,a1968a,a1971a,a1972a,a1975a,a1978a,a1979a,a1982a,a1985a,a1986a,a1989a,a1992a,a1993a,a1996a,a1999a,a2000a,a2003a,a2006a,a2007a,a2010a,a2013a,a2014a,a2017a,a2020a,a2021a,a2024a,a2027a,a2028a,a2031a,a2034a,a2035a,a2038a,a2041a,a2042a,a2045a,a2048a,a2049a,a2052a,a2055a,a2056a,a2059a,a2062a,a2063a,a2066a,a2069a,a2070a,a2073a,a2076a,a2077a,a2080a,a2083a,a2084a,a2087a,a2090a,a2091a,a2094a,a2097a,a2098a,a2101a,a2104a,a2105a,a2108a,a2111a,a2112a,a2115a,a2118a,a2119a,a2122a,a2125a,a2126a,a2129a,a2132a,a2133a,a2136a,a2139a,a2140a,a2143a,a2146a,a2147a,a2150a,a2153a,a2154a,a2157a,a2160a,a2161a,a2164a,a2167a,a2168a,a2171a,a2174a,a2175a,a2178a,a2181a,a2182a,a2185a,a2188a,a2189a,a2192a,a2195a,a2196a,a2199a,a2202a,a2203a,a2206a,a2209a,a2210a,a2213a,a2216a,a2217a,a2220a,a2223a,a2224a,a2227a,a2230a,a2231a,a2234a,a2237a,a2238a,a2241a,a2244a,a2245a,a2248a,a2251a,a2252a,a2255a,a2258a,a2259a,a2262a,a2265a,a2266a,a2269a,a2272a,a2273a,a2276a,a2279a,a2280a,a2283a,a2286a,a2287a,a2290a,a2293a,a2294a,a2297a,a2300a,a2301a,a2304a,a2307a,a2308a,a2311a,a2314a,a2315a,a2318a,a2321a,a2322a,a2325a,a2328a,a2329a,a2332a,a2335a,a2336a,a2339a,a2343a,a2344a,a2345a,a2348a,a2351a,a2352a,a2355a,a2359a,a2360a,a2361a,a2364a,a2367a,a2368a,a2371a,a2375a,a2376a,a2377a,a2380a,a2383a,a2384a,a2387a,a2391a,a2392a,a2393a,a2396a,a2399a,a2400a,a2403a,a2407a,a2408a,a2409a,a2412a,a2415a,a2416a,a2419a,a2423a,a2424a,a2425a,a2428a,a2431a,a2432a,a2435a,a2439a,a2440a,a2441a,a2444a,a2447a,a2448a,a2451a,a2455a,a2456a,a2457a,a2460a,a2463a,a2464a,a2467a,a2471a,a2472a,a2473a,a2476a,a2479a,a2480a,a2483a,a2487a,a2488a,a2489a,a2492a,a2495a,a2496a,a2499a,a2503a,a2504a,a2505a,a2508a,a2511a,a2512a,a2515a,a2519a,a2520a,a2521a,a2524a,a2527a,a2528a,a2531a,a2535a,a2536a,a2537a,a2540a,a2543a,a2544a,a2547a,a2551a,a2552a,a2553a,a2556a,a2559a,a2560a,a2563a,a2567a,a2568a,a2569a,a2572a,a2575a,a2576a,a2579a,a2583a,a2584a,a2585a,a2588a,a2591a,a2592a,a2595a,a2599a,a2600a,a2601a,a2604a,a2607a,a2608a,a2611a,a2615a,a2616a,a2617a,a2620a,a2623a,a2624a,a2627a,a2631a,a2632a,a2633a,a2636a,a2639a,a2640a,a2643a,a2647a,a2648a,a2649a,a2652a,a2655a,a2656a,a2659a,a2663a,a2664a,a2665a,a2668a,a2671a,a2672a,a2675a,a2679a,a2680a,a2681a,a2684a,a2687a,a2688a,a2691a,a2695a,a2696a,a2697a,a2700a,a2703a,a2704a,a2707a,a2711a,a2712a,a2713a,a2716a,a2719a,a2720a,a2723a,a2727a,a2728a,a2729a,a2732a,a2735a,a2736a,a2739a,a2743a,a2744a,a2745a,a2748a,a2751a,a2752a,a2755a,a2759a,a2760a,a2761a,a2764a,a2767a,a2768a,a2771a,a2775a,a2776a,a2777a,a2780a,a2783a,a2784a,a2787a,a2791a,a2792a,a2793a,a2796a,a2799a,a2800a,a2803a,a2807a,a2808a,a2809a,a2812a,a2815a,a2816a,a2819a,a2823a,a2824a,a2825a,a2828a,a2831a,a2832a,a2835a,a2839a,a2840a,a2841a,a2844a,a2848a,a2849a,a2850a,a2853a,a2857a,a2858a,a2859a,a2862a,a2866a,a2867a,a2868a,a2871a,a2875a,a2876a,a2877a,a2880a,a2884a,a2885a,a2886a,a2889a,a2893a,a2894a,a2895a,a2898a,a2902a,a2903a,a2904a,a2907a,a2911a,a2912a,a2913a,a2916a,a2920a,a2921a,a2922a,a2925a,a2929a,a2930a,a2931a,a2934a,a2938a,a2939a,a2940a,a2943a,a2947a,a2948a,a2949a,a2952a,a2956a,a2957a,a2958a,a2961a,a2965a,a2966a,a2967a,a2970a,a2974a,a2975a,a2976a,a2979a,a2983a,a2984a,a2985a: std_logic;
begin

A74 <=( a613a ) or ( a408a );
 a1a <=( a2985a  and  a2976a );
 a2a <=( a2967a  and  a2958a );
 a3a <=( a2949a  and  a2940a );
 a4a <=( a2931a  and  a2922a );
 a5a <=( a2913a  and  a2904a );
 a6a <=( a2895a  and  a2886a );
 a7a <=( a2877a  and  a2868a );
 a8a <=( a2859a  and  a2850a );
 a9a <=( a2841a  and  a2832a );
 a10a <=( a2825a  and  a2816a );
 a11a <=( a2809a  and  a2800a );
 a12a <=( a2793a  and  a2784a );
 a13a <=( a2777a  and  a2768a );
 a14a <=( a2761a  and  a2752a );
 a15a <=( a2745a  and  a2736a );
 a16a <=( a2729a  and  a2720a );
 a17a <=( a2713a  and  a2704a );
 a18a <=( a2697a  and  a2688a );
 a19a <=( a2681a  and  a2672a );
 a20a <=( a2665a  and  a2656a );
 a21a <=( a2649a  and  a2640a );
 a22a <=( a2633a  and  a2624a );
 a23a <=( a2617a  and  a2608a );
 a24a <=( a2601a  and  a2592a );
 a25a <=( a2585a  and  a2576a );
 a26a <=( a2569a  and  a2560a );
 a27a <=( a2553a  and  a2544a );
 a28a <=( a2537a  and  a2528a );
 a29a <=( a2521a  and  a2512a );
 a30a <=( a2505a  and  a2496a );
 a31a <=( a2489a  and  a2480a );
 a32a <=( a2473a  and  a2464a );
 a33a <=( a2457a  and  a2448a );
 a34a <=( a2441a  and  a2432a );
 a35a <=( a2425a  and  a2416a );
 a36a <=( a2409a  and  a2400a );
 a37a <=( a2393a  and  a2384a );
 a38a <=( a2377a  and  a2368a );
 a39a <=( a2361a  and  a2352a );
 a40a <=( a2345a  and  a2336a );
 a41a <=( a2329a  and  a2322a );
 a42a <=( a2315a  and  a2308a );
 a43a <=( a2301a  and  a2294a );
 a44a <=( a2287a  and  a2280a );
 a45a <=( a2273a  and  a2266a );
 a46a <=( a2259a  and  a2252a );
 a47a <=( a2245a  and  a2238a );
 a48a <=( a2231a  and  a2224a );
 a49a <=( a2217a  and  a2210a );
 a50a <=( a2203a  and  a2196a );
 a51a <=( a2189a  and  a2182a );
 a52a <=( a2175a  and  a2168a );
 a53a <=( a2161a  and  a2154a );
 a54a <=( a2147a  and  a2140a );
 a55a <=( a2133a  and  a2126a );
 a56a <=( a2119a  and  a2112a );
 a57a <=( a2105a  and  a2098a );
 a58a <=( a2091a  and  a2084a );
 a59a <=( a2077a  and  a2070a );
 a60a <=( a2063a  and  a2056a );
 a61a <=( a2049a  and  a2042a );
 a62a <=( a2035a  and  a2028a );
 a63a <=( a2021a  and  a2014a );
 a64a <=( a2007a  and  a2000a );
 a65a <=( a1993a  and  a1986a );
 a66a <=( a1979a  and  a1972a );
 a67a <=( a1965a  and  a1958a );
 a68a <=( a1951a  and  a1944a );
 a69a <=( a1937a  and  a1930a );
 a70a <=( a1923a  and  a1916a );
 a71a <=( a1909a  and  a1902a );
 a72a <=( a1895a  and  a1888a );
 a73a <=( a1881a  and  a1874a );
 a74a <=( a1867a  and  a1860a );
 a75a <=( a1853a  and  a1846a );
 a76a <=( a1839a  and  a1832a );
 a77a <=( a1825a  and  a1818a );
 a78a <=( a1811a  and  a1804a );
 a79a <=( a1797a  and  a1790a );
 a80a <=( a1783a  and  a1776a );
 a81a <=( a1769a  and  a1762a );
 a82a <=( a1755a  and  a1748a );
 a83a <=( a1741a  and  a1734a );
 a84a <=( a1727a  and  a1720a );
 a85a <=( a1713a  and  a1706a );
 a86a <=( a1699a  and  a1692a );
 a87a <=( a1685a  and  a1678a );
 a88a <=( a1671a  and  a1664a );
 a89a <=( a1657a  and  a1650a );
 a90a <=( a1645a  and  a1638a );
 a91a <=( a1633a  and  a1626a );
 a92a <=( a1621a  and  a1614a );
 a93a <=( a1609a  and  a1602a );
 a94a <=( a1597a  and  a1590a );
 a95a <=( a1585a  and  a1578a );
 a96a <=( a1573a  and  a1566a );
 a97a <=( a1561a  and  a1554a );
 a98a <=( a1549a  and  a1542a );
 a99a <=( a1537a  and  a1530a );
 a100a <=( a1525a  and  a1518a );
 a101a <=( a1513a  and  a1506a );
 a102a <=( a1501a  and  a1494a );
 a103a <=( a1489a  and  a1482a );
 a104a <=( a1477a  and  a1470a );
 a105a <=( a1465a  and  a1458a );
 a106a <=( a1453a  and  a1446a );
 a107a <=( a1441a  and  a1434a );
 a108a <=( a1429a  and  a1422a );
 a109a <=( a1417a  and  a1410a );
 a110a <=( a1405a  and  a1398a );
 a111a <=( a1393a  and  a1386a );
 a112a <=( a1381a  and  a1374a );
 a113a <=( a1369a  and  a1362a );
 a114a <=( a1357a  and  a1350a );
 a115a <=( a1345a  and  a1338a );
 a116a <=( a1333a  and  a1326a );
 a117a <=( a1321a  and  a1314a );
 a118a <=( a1309a  and  a1302a );
 a119a <=( a1297a  and  a1290a );
 a120a <=( a1285a  and  a1278a );
 a121a <=( a1273a  and  a1266a );
 a122a <=( a1261a  and  a1254a );
 a123a <=( a1249a  and  a1242a );
 a124a <=( a1237a  and  a1230a );
 a125a <=( a1225a  and  a1218a );
 a126a <=( a1213a  and  a1206a );
 a127a <=( a1201a  and  a1194a );
 a128a <=( a1189a  and  a1182a );
 a129a <=( a1177a  and  a1172a );
 a130a <=( a1167a  and  a1162a );
 a131a <=( a1157a  and  a1152a );
 a132a <=( a1147a  and  a1142a );
 a133a <=( a1137a  and  a1132a );
 a134a <=( a1127a  and  a1122a );
 a135a <=( a1117a  and  a1112a );
 a136a <=( a1107a  and  a1102a );
 a137a <=( a1097a  and  a1092a );
 a138a <=( a1087a  and  a1082a );
 a139a <=( a1077a  and  a1072a );
 a140a <=( a1067a  and  a1062a );
 a141a <=( a1057a  and  a1052a );
 a142a <=( a1047a  and  a1042a );
 a143a <=( a1037a  and  a1032a );
 a144a <=( a1027a  and  a1022a );
 a145a <=( a1017a  and  a1012a );
 a146a <=( a1007a  and  a1002a );
 a147a <=( a997a  and  a992a );
 a148a <=( a987a  and  a982a );
 a149a <=( a977a  and  a972a );
 a150a <=( a967a  and  a962a );
 a151a <=( a957a  and  a952a );
 a152a <=( a947a  and  a942a );
 a153a <=( a937a  and  a932a );
 a154a <=( a927a  and  a922a );
 a155a <=( a917a  and  a912a );
 a156a <=( a909a  and  a904a );
 a157a <=( a901a  and  a896a );
 a158a <=( a893a  and  a888a );
 a159a <=( a885a  and  a880a );
 a160a <=( a877a  and  a872a );
 a161a <=( a869a  and  a864a );
 a162a <=( a861a  and  a856a );
 a163a <=( a853a  and  a848a );
 a164a <=( a845a  and  a840a );
 a165a <=( a837a  and  a832a );
 a166a <=( a829a  and  a824a );
 a167a <=( a821a  and  a816a );
 a168a <=( a813a  and  a808a );
 a169a <=( a805a  and  a800a );
 a170a <=( a797a  and  a792a );
 a171a <=( a789a  and  a784a );
 a172a <=( a781a  and  a776a );
 a173a <=( a773a  and  a768a );
 a174a <=( a765a  and  a760a );
 a175a <=( a757a  and  a754a );
 a176a <=( a751a  and  a748a );
 a177a <=( a745a  and  a742a );
 a178a <=( a739a  and  a736a );
 a179a <=( a733a  and  a730a );
 a180a <=( a727a  and  a724a );
 a181a <=( a721a  and  a718a );
 a182a <=( a715a  and  a712a );
 a183a <=( a709a  and  a706a );
 a184a <=( a703a  and  a700a );
 a185a <=( a697a  and  a694a );
 a186a <=( a691a  and  a688a );
 a187a <=( a685a  and  a682a );
 a188a <=( a679a  and  a676a );
 a189a <=( a673a  and  a670a );
 a190a <=( a667a  and  a664a );
 a191a <=( A169  and  a661a );
 a192a <=( A169  and  a657a );
 a193a <=( A168  and  a653a );
 a194a <=( A168  and  a649a );
 a195a <=( A200  and  a645a );
 a196a <=( A199  and  a641a );
 a197a <=( A202  and  a637a );
 a198a <=( A202  and  a633a );
 a199a <=( A265  and  a629a );
 a200a <=( (not A265)  and  a625a );
 a201a <=( A235  and  A169 );
 a202a <=( A235  and  A202 );
 a203a <=( A267  and  A266 );
 a204a <=( A267  and  A265 );
 a209a <=( a203a ) or ( a204a );
 a210a <=( A268 ) or ( a209a );
 a214a <=( a200a ) or ( a201a );
 a215a <=( a202a ) or ( a214a );
 a216a <=( a215a ) or ( a210a );
 a220a <=( a197a ) or ( a198a );
 a221a <=( a199a ) or ( a220a );
 a225a <=( a194a ) or ( a195a );
 a226a <=( a196a ) or ( a225a );
 a227a <=( a226a ) or ( a221a );
 a228a <=( a227a ) or ( a216a );
 a232a <=( a191a ) or ( a192a );
 a233a <=( a193a ) or ( a232a );
 a237a <=( a188a ) or ( a189a );
 a238a <=( a190a ) or ( a237a );
 a239a <=( a238a ) or ( a233a );
 a243a <=( a185a ) or ( a186a );
 a244a <=( a187a ) or ( a243a );
 a247a <=( a183a ) or ( a184a );
 a250a <=( a181a ) or ( a182a );
 a251a <=( a250a ) or ( a247a );
 a252a <=( a251a ) or ( a244a );
 a253a <=( a252a ) or ( a239a );
 a254a <=( a253a ) or ( a228a );
 a258a <=( a178a ) or ( a179a );
 a259a <=( a180a ) or ( a258a );
 a263a <=( a175a ) or ( a176a );
 a264a <=( a177a ) or ( a263a );
 a265a <=( a264a ) or ( a259a );
 a269a <=( a172a ) or ( a173a );
 a270a <=( a174a ) or ( a269a );
 a273a <=( a170a ) or ( a171a );
 a276a <=( a168a ) or ( a169a );
 a277a <=( a276a ) or ( a273a );
 a278a <=( a277a ) or ( a270a );
 a279a <=( a278a ) or ( a265a );
 a283a <=( a165a ) or ( a166a );
 a284a <=( a167a ) or ( a283a );
 a288a <=( a162a ) or ( a163a );
 a289a <=( a164a ) or ( a288a );
 a290a <=( a289a ) or ( a284a );
 a294a <=( a159a ) or ( a160a );
 a295a <=( a161a ) or ( a294a );
 a298a <=( a157a ) or ( a158a );
 a301a <=( a155a ) or ( a156a );
 a302a <=( a301a ) or ( a298a );
 a303a <=( a302a ) or ( a295a );
 a304a <=( a303a ) or ( a290a );
 a305a <=( a304a ) or ( a279a );
 a306a <=( a305a ) or ( a254a );
 a310a <=( a152a ) or ( a153a );
 a311a <=( a154a ) or ( a310a );
 a315a <=( a149a ) or ( a150a );
 a316a <=( a151a ) or ( a315a );
 a317a <=( a316a ) or ( a311a );
 a321a <=( a146a ) or ( a147a );
 a322a <=( a148a ) or ( a321a );
 a326a <=( a143a ) or ( a144a );
 a327a <=( a145a ) or ( a326a );
 a328a <=( a327a ) or ( a322a );
 a329a <=( a328a ) or ( a317a );
 a333a <=( a140a ) or ( a141a );
 a334a <=( a142a ) or ( a333a );
 a338a <=( a137a ) or ( a138a );
 a339a <=( a139a ) or ( a338a );
 a340a <=( a339a ) or ( a334a );
 a344a <=( a134a ) or ( a135a );
 a345a <=( a136a ) or ( a344a );
 a348a <=( a132a ) or ( a133a );
 a351a <=( a130a ) or ( a131a );
 a352a <=( a351a ) or ( a348a );
 a353a <=( a352a ) or ( a345a );
 a354a <=( a353a ) or ( a340a );
 a355a <=( a354a ) or ( a329a );
 a359a <=( a127a ) or ( a128a );
 a360a <=( a129a ) or ( a359a );
 a364a <=( a124a ) or ( a125a );
 a365a <=( a126a ) or ( a364a );
 a366a <=( a365a ) or ( a360a );
 a370a <=( a121a ) or ( a122a );
 a371a <=( a123a ) or ( a370a );
 a374a <=( a119a ) or ( a120a );
 a377a <=( a117a ) or ( a118a );
 a378a <=( a377a ) or ( a374a );
 a379a <=( a378a ) or ( a371a );
 a380a <=( a379a ) or ( a366a );
 a384a <=( a114a ) or ( a115a );
 a385a <=( a116a ) or ( a384a );
 a389a <=( a111a ) or ( a112a );
 a390a <=( a113a ) or ( a389a );
 a391a <=( a390a ) or ( a385a );
 a395a <=( a108a ) or ( a109a );
 a396a <=( a110a ) or ( a395a );
 a399a <=( a106a ) or ( a107a );
 a402a <=( a104a ) or ( a105a );
 a403a <=( a402a ) or ( a399a );
 a404a <=( a403a ) or ( a396a );
 a405a <=( a404a ) or ( a391a );
 a406a <=( a405a ) or ( a380a );
 a407a <=( a406a ) or ( a355a );
 a408a <=( a407a ) or ( a306a );
 a412a <=( a101a ) or ( a102a );
 a413a <=( a103a ) or ( a412a );
 a417a <=( a98a ) or ( a99a );
 a418a <=( a100a ) or ( a417a );
 a419a <=( a418a ) or ( a413a );
 a423a <=( a95a ) or ( a96a );
 a424a <=( a97a ) or ( a423a );
 a428a <=( a92a ) or ( a93a );
 a429a <=( a94a ) or ( a428a );
 a430a <=( a429a ) or ( a424a );
 a431a <=( a430a ) or ( a419a );
 a435a <=( a89a ) or ( a90a );
 a436a <=( a91a ) or ( a435a );
 a440a <=( a86a ) or ( a87a );
 a441a <=( a88a ) or ( a440a );
 a442a <=( a441a ) or ( a436a );
 a446a <=( a83a ) or ( a84a );
 a447a <=( a85a ) or ( a446a );
 a450a <=( a81a ) or ( a82a );
 a453a <=( a79a ) or ( a80a );
 a454a <=( a453a ) or ( a450a );
 a455a <=( a454a ) or ( a447a );
 a456a <=( a455a ) or ( a442a );
 a457a <=( a456a ) or ( a431a );
 a461a <=( a76a ) or ( a77a );
 a462a <=( a78a ) or ( a461a );
 a466a <=( a73a ) or ( a74a );
 a467a <=( a75a ) or ( a466a );
 a468a <=( a467a ) or ( a462a );
 a472a <=( a70a ) or ( a71a );
 a473a <=( a72a ) or ( a472a );
 a476a <=( a68a ) or ( a69a );
 a479a <=( a66a ) or ( a67a );
 a480a <=( a479a ) or ( a476a );
 a481a <=( a480a ) or ( a473a );
 a482a <=( a481a ) or ( a468a );
 a486a <=( a63a ) or ( a64a );
 a487a <=( a65a ) or ( a486a );
 a491a <=( a60a ) or ( a61a );
 a492a <=( a62a ) or ( a491a );
 a493a <=( a492a ) or ( a487a );
 a497a <=( a57a ) or ( a58a );
 a498a <=( a59a ) or ( a497a );
 a501a <=( a55a ) or ( a56a );
 a504a <=( a53a ) or ( a54a );
 a505a <=( a504a ) or ( a501a );
 a506a <=( a505a ) or ( a498a );
 a507a <=( a506a ) or ( a493a );
 a508a <=( a507a ) or ( a482a );
 a509a <=( a508a ) or ( a457a );
 a513a <=( a50a ) or ( a51a );
 a514a <=( a52a ) or ( a513a );
 a518a <=( a47a ) or ( a48a );
 a519a <=( a49a ) or ( a518a );
 a520a <=( a519a ) or ( a514a );
 a524a <=( a44a ) or ( a45a );
 a525a <=( a46a ) or ( a524a );
 a528a <=( a42a ) or ( a43a );
 a531a <=( a40a ) or ( a41a );
 a532a <=( a531a ) or ( a528a );
 a533a <=( a532a ) or ( a525a );
 a534a <=( a533a ) or ( a520a );
 a538a <=( a37a ) or ( a38a );
 a539a <=( a39a ) or ( a538a );
 a543a <=( a34a ) or ( a35a );
 a544a <=( a36a ) or ( a543a );
 a545a <=( a544a ) or ( a539a );
 a549a <=( a31a ) or ( a32a );
 a550a <=( a33a ) or ( a549a );
 a553a <=( a29a ) or ( a30a );
 a556a <=( a27a ) or ( a28a );
 a557a <=( a556a ) or ( a553a );
 a558a <=( a557a ) or ( a550a );
 a559a <=( a558a ) or ( a545a );
 a560a <=( a559a ) or ( a534a );
 a564a <=( a24a ) or ( a25a );
 a565a <=( a26a ) or ( a564a );
 a569a <=( a21a ) or ( a22a );
 a570a <=( a23a ) or ( a569a );
 a571a <=( a570a ) or ( a565a );
 a575a <=( a18a ) or ( a19a );
 a576a <=( a20a ) or ( a575a );
 a579a <=( a16a ) or ( a17a );
 a582a <=( a14a ) or ( a15a );
 a583a <=( a582a ) or ( a579a );
 a584a <=( a583a ) or ( a576a );
 a585a <=( a584a ) or ( a571a );
 a589a <=( a11a ) or ( a12a );
 a590a <=( a13a ) or ( a589a );
 a594a <=( a8a ) or ( a9a );
 a595a <=( a10a ) or ( a594a );
 a596a <=( a595a ) or ( a590a );
 a600a <=( a5a ) or ( a6a );
 a601a <=( a7a ) or ( a600a );
 a604a <=( a3a ) or ( a4a );
 a607a <=( a1a ) or ( a2a );
 a608a <=( a607a ) or ( a604a );
 a609a <=( a608a ) or ( a601a );
 a610a <=( a609a ) or ( a596a );
 a611a <=( a610a ) or ( a585a );
 a612a <=( a611a ) or ( a560a );
 a613a <=( a612a ) or ( a509a );
 a625a <=( A269  and  A266 );
 a629a <=( A269  and  (not A266) );
 a633a <=( A234  and  A232 );
 a637a <=( A234  and  A233 );
 a641a <=( A235  and  A201 );
 a645a <=( A235  and  A201 );
 a649a <=( A235  and  A166 );
 a653a <=( A235  and  A167 );
 a657a <=( A234  and  A232 );
 a661a <=( A234  and  A233 );
 a664a <=( (not A232)  and  A202 );
 a667a <=( A236  and  A233 );
 a670a <=( A232  and  A202 );
 a673a <=( A236  and  (not A233) );
 a676a <=( A201  and  A199 );
 a679a <=( A234  and  A232 );
 a682a <=( A201  and  A199 );
 a685a <=( A234  and  A233 );
 a688a <=( A201  and  A200 );
 a691a <=( A234  and  A232 );
 a694a <=( A201  and  A200 );
 a697a <=( A234  and  A233 );
 a700a <=( A200  and  (not A199) );
 a703a <=( A235  and  A203 );
 a706a <=( (not A200)  and  A199 );
 a709a <=( A235  and  A203 );
 a712a <=( A166  and  A168 );
 a715a <=( A234  and  A232 );
 a718a <=( A166  and  A168 );
 a721a <=( A234  and  A233 );
 a724a <=( A167  and  A168 );
 a727a <=( A234  and  A232 );
 a730a <=( A167  and  A168 );
 a733a <=( A234  and  A233 );
 a736a <=( A167  and  A170 );
 a739a <=( A235  and  (not A166) );
 a742a <=( (not A167)  and  A170 );
 a745a <=( A235  and  A166 );
 a748a <=( (not A232)  and  A169 );
 a751a <=( A236  and  A233 );
 a754a <=( A232  and  A169 );
 a757a <=( A236  and  (not A233) );
 a760a <=( A201  and  A199 );
 a764a <=( A236  and  A233 );
 a765a <=( (not A232)  and  a764a );
 a768a <=( A201  and  A199 );
 a772a <=( A236  and  (not A233) );
 a773a <=( A232  and  a772a );
 a776a <=( A201  and  A200 );
 a780a <=( A236  and  A233 );
 a781a <=( (not A232)  and  a780a );
 a784a <=( A201  and  A200 );
 a788a <=( A236  and  (not A233) );
 a789a <=( A232  and  a788a );
 a792a <=( A200  and  (not A199) );
 a796a <=( A234  and  A232 );
 a797a <=( A203  and  a796a );
 a800a <=( A200  and  (not A199) );
 a804a <=( A234  and  A233 );
 a805a <=( A203  and  a804a );
 a808a <=( (not A200)  and  A199 );
 a812a <=( A234  and  A232 );
 a813a <=( A203  and  a812a );
 a816a <=( (not A200)  and  A199 );
 a820a <=( A234  and  A233 );
 a821a <=( A203  and  a820a );
 a824a <=( A166  and  A168 );
 a828a <=( A236  and  A233 );
 a829a <=( (not A232)  and  a828a );
 a832a <=( A166  and  A168 );
 a836a <=( A236  and  (not A233) );
 a837a <=( A232  and  a836a );
 a840a <=( A167  and  A168 );
 a844a <=( A236  and  A233 );
 a845a <=( (not A232)  and  a844a );
 a848a <=( A167  and  A168 );
 a852a <=( A236  and  (not A233) );
 a853a <=( A232  and  a852a );
 a856a <=( A167  and  A170 );
 a860a <=( A234  and  A232 );
 a861a <=( (not A166)  and  a860a );
 a864a <=( A167  and  A170 );
 a868a <=( A234  and  A233 );
 a869a <=( (not A166)  and  a868a );
 a872a <=( (not A167)  and  A170 );
 a876a <=( A234  and  A232 );
 a877a <=( A166  and  a876a );
 a880a <=( (not A167)  and  A170 );
 a884a <=( A234  and  A233 );
 a885a <=( A166  and  a884a );
 a888a <=( (not A201)  and  A169 );
 a892a <=( A301  and  (not A203) );
 a893a <=( (not A202)  and  a892a );
 a896a <=( (not A199)  and  A169 );
 a900a <=( A301  and  (not A202) );
 a901a <=( (not A200)  and  a900a );
 a904a <=( (not A167)  and  (not A169) );
 a908a <=( A301  and  A202 );
 a909a <=( (not A166)  and  a908a );
 a912a <=( (not A169)  and  (not A170) );
 a916a <=( A301  and  A202 );
 a917a <=( (not A168)  and  a916a );
 a921a <=( A203  and  A200 );
 a922a <=( (not A199)  and  a921a );
 a926a <=( A236  and  A233 );
 a927a <=( (not A232)  and  a926a );
 a931a <=( A203  and  A200 );
 a932a <=( (not A199)  and  a931a );
 a936a <=( A236  and  (not A233) );
 a937a <=( A232  and  a936a );
 a941a <=( A203  and  (not A200) );
 a942a <=( A199  and  a941a );
 a946a <=( A236  and  A233 );
 a947a <=( (not A232)  and  a946a );
 a951a <=( A203  and  (not A200) );
 a952a <=( A199  and  a951a );
 a956a <=( A236  and  (not A233) );
 a957a <=( A232  and  a956a );
 a961a <=( (not A201)  and  A166 );
 a962a <=( A168  and  a961a );
 a966a <=( A301  and  (not A203) );
 a967a <=( (not A202)  and  a966a );
 a971a <=( (not A199)  and  A166 );
 a972a <=( A168  and  a971a );
 a976a <=( A301  and  (not A202) );
 a977a <=( (not A200)  and  a976a );
 a981a <=( (not A201)  and  A167 );
 a982a <=( A168  and  a981a );
 a986a <=( A301  and  (not A203) );
 a987a <=( (not A202)  and  a986a );
 a991a <=( (not A199)  and  A167 );
 a992a <=( A168  and  a991a );
 a996a <=( A301  and  (not A202) );
 a997a <=( (not A200)  and  a996a );
 a1001a <=( (not A166)  and  A167 );
 a1002a <=( A170  and  a1001a );
 a1006a <=( A236  and  A233 );
 a1007a <=( (not A232)  and  a1006a );
 a1011a <=( (not A166)  and  A167 );
 a1012a <=( A170  and  a1011a );
 a1016a <=( A236  and  (not A233) );
 a1017a <=( A232  and  a1016a );
 a1021a <=( A166  and  (not A167) );
 a1022a <=( A170  and  a1021a );
 a1026a <=( A236  and  A233 );
 a1027a <=( (not A232)  and  a1026a );
 a1031a <=( A166  and  (not A167) );
 a1032a <=( A170  and  a1031a );
 a1036a <=( A236  and  (not A233) );
 a1037a <=( A232  and  a1036a );
 a1041a <=( (not A202)  and  (not A201) );
 a1042a <=( A169  and  a1041a );
 a1046a <=( A300  and  A299 );
 a1047a <=( (not A203)  and  a1046a );
 a1051a <=( (not A202)  and  (not A201) );
 a1052a <=( A169  and  a1051a );
 a1056a <=( A300  and  A298 );
 a1057a <=( (not A203)  and  a1056a );
 a1061a <=( A200  and  A199 );
 a1062a <=( A169  and  a1061a );
 a1066a <=( A301  and  (not A202) );
 a1067a <=( (not A201)  and  a1066a );
 a1071a <=( (not A200)  and  (not A199) );
 a1072a <=( A169  and  a1071a );
 a1076a <=( A300  and  A299 );
 a1077a <=( (not A202)  and  a1076a );
 a1081a <=( (not A200)  and  (not A199) );
 a1082a <=( A169  and  a1081a );
 a1086a <=( A300  and  A298 );
 a1087a <=( (not A202)  and  a1086a );
 a1091a <=( (not A166)  and  (not A167) );
 a1092a <=( (not A169)  and  a1091a );
 a1096a <=( A300  and  A299 );
 a1097a <=( A202  and  a1096a );
 a1101a <=( (not A166)  and  (not A167) );
 a1102a <=( (not A169)  and  a1101a );
 a1106a <=( A300  and  A298 );
 a1107a <=( A202  and  a1106a );
 a1111a <=( (not A166)  and  (not A167) );
 a1112a <=( (not A169)  and  a1111a );
 a1116a <=( A301  and  A201 );
 a1117a <=( A199  and  a1116a );
 a1121a <=( (not A166)  and  (not A167) );
 a1122a <=( (not A169)  and  a1121a );
 a1126a <=( A301  and  A201 );
 a1127a <=( A200  and  a1126a );
 a1131a <=( A167  and  (not A168) );
 a1132a <=( (not A169)  and  a1131a );
 a1136a <=( A301  and  A202 );
 a1137a <=( A166  and  a1136a );
 a1141a <=( (not A168)  and  (not A169) );
 a1142a <=( (not A170)  and  a1141a );
 a1146a <=( A300  and  A299 );
 a1147a <=( A202  and  a1146a );
 a1151a <=( (not A168)  and  (not A169) );
 a1152a <=( (not A170)  and  a1151a );
 a1156a <=( A300  and  A298 );
 a1157a <=( A202  and  a1156a );
 a1161a <=( (not A168)  and  (not A169) );
 a1162a <=( (not A170)  and  a1161a );
 a1166a <=( A301  and  A201 );
 a1167a <=( A199  and  a1166a );
 a1171a <=( (not A168)  and  (not A169) );
 a1172a <=( (not A170)  and  a1171a );
 a1176a <=( A301  and  A201 );
 a1177a <=( A200  and  a1176a );
 a1181a <=( (not A201)  and  A166 );
 a1182a <=( A168  and  a1181a );
 a1185a <=( (not A203)  and  (not A202) );
 a1188a <=( A300  and  A299 );
 a1189a <=( a1188a  and  a1185a );
 a1193a <=( (not A201)  and  A166 );
 a1194a <=( A168  and  a1193a );
 a1197a <=( (not A203)  and  (not A202) );
 a1200a <=( A300  and  A298 );
 a1201a <=( a1200a  and  a1197a );
 a1205a <=( A199  and  A166 );
 a1206a <=( A168  and  a1205a );
 a1209a <=( (not A201)  and  A200 );
 a1212a <=( A301  and  (not A202) );
 a1213a <=( a1212a  and  a1209a );
 a1217a <=( (not A199)  and  A166 );
 a1218a <=( A168  and  a1217a );
 a1221a <=( (not A202)  and  (not A200) );
 a1224a <=( A300  and  A299 );
 a1225a <=( a1224a  and  a1221a );
 a1229a <=( (not A199)  and  A166 );
 a1230a <=( A168  and  a1229a );
 a1233a <=( (not A202)  and  (not A200) );
 a1236a <=( A300  and  A298 );
 a1237a <=( a1236a  and  a1233a );
 a1241a <=( (not A201)  and  A167 );
 a1242a <=( A168  and  a1241a );
 a1245a <=( (not A203)  and  (not A202) );
 a1248a <=( A300  and  A299 );
 a1249a <=( a1248a  and  a1245a );
 a1253a <=( (not A201)  and  A167 );
 a1254a <=( A168  and  a1253a );
 a1257a <=( (not A203)  and  (not A202) );
 a1260a <=( A300  and  A298 );
 a1261a <=( a1260a  and  a1257a );
 a1265a <=( A199  and  A167 );
 a1266a <=( A168  and  a1265a );
 a1269a <=( (not A201)  and  A200 );
 a1272a <=( A301  and  (not A202) );
 a1273a <=( a1272a  and  a1269a );
 a1277a <=( (not A199)  and  A167 );
 a1278a <=( A168  and  a1277a );
 a1281a <=( (not A202)  and  (not A200) );
 a1284a <=( A300  and  A299 );
 a1285a <=( a1284a  and  a1281a );
 a1289a <=( (not A199)  and  A167 );
 a1290a <=( A168  and  a1289a );
 a1293a <=( (not A202)  and  (not A200) );
 a1296a <=( A300  and  A298 );
 a1297a <=( a1296a  and  a1293a );
 a1301a <=( (not A166)  and  A167 );
 a1302a <=( A170  and  a1301a );
 a1305a <=( (not A202)  and  (not A201) );
 a1308a <=( A301  and  (not A203) );
 a1309a <=( a1308a  and  a1305a );
 a1313a <=( (not A166)  and  A167 );
 a1314a <=( A170  and  a1313a );
 a1317a <=( (not A200)  and  (not A199) );
 a1320a <=( A301  and  (not A202) );
 a1321a <=( a1320a  and  a1317a );
 a1325a <=( A166  and  (not A167) );
 a1326a <=( A170  and  a1325a );
 a1329a <=( (not A202)  and  (not A201) );
 a1332a <=( A301  and  (not A203) );
 a1333a <=( a1332a  and  a1329a );
 a1337a <=( A166  and  (not A167) );
 a1338a <=( A170  and  a1337a );
 a1341a <=( (not A200)  and  (not A199) );
 a1344a <=( A301  and  (not A202) );
 a1345a <=( a1344a  and  a1341a );
 a1349a <=( (not A202)  and  (not A201) );
 a1350a <=( A169  and  a1349a );
 a1353a <=( A298  and  (not A203) );
 a1356a <=( A302  and  (not A299) );
 a1357a <=( a1356a  and  a1353a );
 a1361a <=( (not A202)  and  (not A201) );
 a1362a <=( A169  and  a1361a );
 a1365a <=( (not A298)  and  (not A203) );
 a1368a <=( A302  and  A299 );
 a1369a <=( a1368a  and  a1365a );
 a1373a <=( A200  and  A199 );
 a1374a <=( A169  and  a1373a );
 a1377a <=( (not A202)  and  (not A201) );
 a1380a <=( A300  and  A299 );
 a1381a <=( a1380a  and  a1377a );
 a1385a <=( A200  and  A199 );
 a1386a <=( A169  and  a1385a );
 a1389a <=( (not A202)  and  (not A201) );
 a1392a <=( A300  and  A298 );
 a1393a <=( a1392a  and  a1389a );
 a1397a <=( (not A200)  and  (not A199) );
 a1398a <=( A169  and  a1397a );
 a1401a <=( A298  and  (not A202) );
 a1404a <=( A302  and  (not A299) );
 a1405a <=( a1404a  and  a1401a );
 a1409a <=( (not A200)  and  (not A199) );
 a1410a <=( A169  and  a1409a );
 a1413a <=( (not A298)  and  (not A202) );
 a1416a <=( A302  and  A299 );
 a1417a <=( a1416a  and  a1413a );
 a1421a <=( (not A166)  and  (not A167) );
 a1422a <=( (not A169)  and  a1421a );
 a1425a <=( A298  and  A202 );
 a1428a <=( A302  and  (not A299) );
 a1429a <=( a1428a  and  a1425a );
 a1433a <=( (not A166)  and  (not A167) );
 a1434a <=( (not A169)  and  a1433a );
 a1437a <=( (not A298)  and  A202 );
 a1440a <=( A302  and  A299 );
 a1441a <=( a1440a  and  a1437a );
 a1445a <=( (not A166)  and  (not A167) );
 a1446a <=( (not A169)  and  a1445a );
 a1449a <=( A201  and  A199 );
 a1452a <=( A300  and  A299 );
 a1453a <=( a1452a  and  a1449a );
 a1457a <=( (not A166)  and  (not A167) );
 a1458a <=( (not A169)  and  a1457a );
 a1461a <=( A201  and  A199 );
 a1464a <=( A300  and  A298 );
 a1465a <=( a1464a  and  a1461a );
 a1469a <=( (not A166)  and  (not A167) );
 a1470a <=( (not A169)  and  a1469a );
 a1473a <=( A201  and  A200 );
 a1476a <=( A300  and  A299 );
 a1477a <=( a1476a  and  a1473a );
 a1481a <=( (not A166)  and  (not A167) );
 a1482a <=( (not A169)  and  a1481a );
 a1485a <=( A201  and  A200 );
 a1488a <=( A300  and  A298 );
 a1489a <=( a1488a  and  a1485a );
 a1493a <=( (not A166)  and  (not A167) );
 a1494a <=( (not A169)  and  a1493a );
 a1497a <=( A200  and  (not A199) );
 a1500a <=( A301  and  A203 );
 a1501a <=( a1500a  and  a1497a );
 a1505a <=( (not A166)  and  (not A167) );
 a1506a <=( (not A169)  and  a1505a );
 a1509a <=( (not A200)  and  A199 );
 a1512a <=( A301  and  A203 );
 a1513a <=( a1512a  and  a1509a );
 a1517a <=( A167  and  (not A168) );
 a1518a <=( (not A169)  and  a1517a );
 a1521a <=( A202  and  A166 );
 a1524a <=( A300  and  A299 );
 a1525a <=( a1524a  and  a1521a );
 a1529a <=( A167  and  (not A168) );
 a1530a <=( (not A169)  and  a1529a );
 a1533a <=( A202  and  A166 );
 a1536a <=( A300  and  A298 );
 a1537a <=( a1536a  and  a1533a );
 a1541a <=( A167  and  (not A168) );
 a1542a <=( (not A169)  and  a1541a );
 a1545a <=( A199  and  A166 );
 a1548a <=( A301  and  A201 );
 a1549a <=( a1548a  and  a1545a );
 a1553a <=( A167  and  (not A168) );
 a1554a <=( (not A169)  and  a1553a );
 a1557a <=( A200  and  A166 );
 a1560a <=( A301  and  A201 );
 a1561a <=( a1560a  and  a1557a );
 a1565a <=( (not A168)  and  (not A169) );
 a1566a <=( (not A170)  and  a1565a );
 a1569a <=( A298  and  A202 );
 a1572a <=( A302  and  (not A299) );
 a1573a <=( a1572a  and  a1569a );
 a1577a <=( (not A168)  and  (not A169) );
 a1578a <=( (not A170)  and  a1577a );
 a1581a <=( (not A298)  and  A202 );
 a1584a <=( A302  and  A299 );
 a1585a <=( a1584a  and  a1581a );
 a1589a <=( (not A168)  and  (not A169) );
 a1590a <=( (not A170)  and  a1589a );
 a1593a <=( A201  and  A199 );
 a1596a <=( A300  and  A299 );
 a1597a <=( a1596a  and  a1593a );
 a1601a <=( (not A168)  and  (not A169) );
 a1602a <=( (not A170)  and  a1601a );
 a1605a <=( A201  and  A199 );
 a1608a <=( A300  and  A298 );
 a1609a <=( a1608a  and  a1605a );
 a1613a <=( (not A168)  and  (not A169) );
 a1614a <=( (not A170)  and  a1613a );
 a1617a <=( A201  and  A200 );
 a1620a <=( A300  and  A299 );
 a1621a <=( a1620a  and  a1617a );
 a1625a <=( (not A168)  and  (not A169) );
 a1626a <=( (not A170)  and  a1625a );
 a1629a <=( A201  and  A200 );
 a1632a <=( A300  and  A298 );
 a1633a <=( a1632a  and  a1629a );
 a1637a <=( (not A168)  and  (not A169) );
 a1638a <=( (not A170)  and  a1637a );
 a1641a <=( A200  and  (not A199) );
 a1644a <=( A301  and  A203 );
 a1645a <=( a1644a  and  a1641a );
 a1649a <=( (not A168)  and  (not A169) );
 a1650a <=( (not A170)  and  a1649a );
 a1653a <=( (not A200)  and  A199 );
 a1656a <=( A301  and  A203 );
 a1657a <=( a1656a  and  a1653a );
 a1660a <=( A166  and  A168 );
 a1663a <=( (not A202)  and  (not A201) );
 a1664a <=( a1663a  and  a1660a );
 a1667a <=( A298  and  (not A203) );
 a1670a <=( A302  and  (not A299) );
 a1671a <=( a1670a  and  a1667a );
 a1674a <=( A166  and  A168 );
 a1677a <=( (not A202)  and  (not A201) );
 a1678a <=( a1677a  and  a1674a );
 a1681a <=( (not A298)  and  (not A203) );
 a1684a <=( A302  and  A299 );
 a1685a <=( a1684a  and  a1681a );
 a1688a <=( A166  and  A168 );
 a1691a <=( A200  and  A199 );
 a1692a <=( a1691a  and  a1688a );
 a1695a <=( (not A202)  and  (not A201) );
 a1698a <=( A300  and  A299 );
 a1699a <=( a1698a  and  a1695a );
 a1702a <=( A166  and  A168 );
 a1705a <=( A200  and  A199 );
 a1706a <=( a1705a  and  a1702a );
 a1709a <=( (not A202)  and  (not A201) );
 a1712a <=( A300  and  A298 );
 a1713a <=( a1712a  and  a1709a );
 a1716a <=( A166  and  A168 );
 a1719a <=( (not A200)  and  (not A199) );
 a1720a <=( a1719a  and  a1716a );
 a1723a <=( A298  and  (not A202) );
 a1726a <=( A302  and  (not A299) );
 a1727a <=( a1726a  and  a1723a );
 a1730a <=( A166  and  A168 );
 a1733a <=( (not A200)  and  (not A199) );
 a1734a <=( a1733a  and  a1730a );
 a1737a <=( (not A298)  and  (not A202) );
 a1740a <=( A302  and  A299 );
 a1741a <=( a1740a  and  a1737a );
 a1744a <=( A167  and  A168 );
 a1747a <=( (not A202)  and  (not A201) );
 a1748a <=( a1747a  and  a1744a );
 a1751a <=( A298  and  (not A203) );
 a1754a <=( A302  and  (not A299) );
 a1755a <=( a1754a  and  a1751a );
 a1758a <=( A167  and  A168 );
 a1761a <=( (not A202)  and  (not A201) );
 a1762a <=( a1761a  and  a1758a );
 a1765a <=( (not A298)  and  (not A203) );
 a1768a <=( A302  and  A299 );
 a1769a <=( a1768a  and  a1765a );
 a1772a <=( A167  and  A168 );
 a1775a <=( A200  and  A199 );
 a1776a <=( a1775a  and  a1772a );
 a1779a <=( (not A202)  and  (not A201) );
 a1782a <=( A300  and  A299 );
 a1783a <=( a1782a  and  a1779a );
 a1786a <=( A167  and  A168 );
 a1789a <=( A200  and  A199 );
 a1790a <=( a1789a  and  a1786a );
 a1793a <=( (not A202)  and  (not A201) );
 a1796a <=( A300  and  A298 );
 a1797a <=( a1796a  and  a1793a );
 a1800a <=( A167  and  A168 );
 a1803a <=( (not A200)  and  (not A199) );
 a1804a <=( a1803a  and  a1800a );
 a1807a <=( A298  and  (not A202) );
 a1810a <=( A302  and  (not A299) );
 a1811a <=( a1810a  and  a1807a );
 a1814a <=( A167  and  A168 );
 a1817a <=( (not A200)  and  (not A199) );
 a1818a <=( a1817a  and  a1814a );
 a1821a <=( (not A298)  and  (not A202) );
 a1824a <=( A302  and  A299 );
 a1825a <=( a1824a  and  a1821a );
 a1828a <=( A167  and  A170 );
 a1831a <=( (not A201)  and  (not A166) );
 a1832a <=( a1831a  and  a1828a );
 a1835a <=( (not A203)  and  (not A202) );
 a1838a <=( A300  and  A299 );
 a1839a <=( a1838a  and  a1835a );
 a1842a <=( A167  and  A170 );
 a1845a <=( (not A201)  and  (not A166) );
 a1846a <=( a1845a  and  a1842a );
 a1849a <=( (not A203)  and  (not A202) );
 a1852a <=( A300  and  A298 );
 a1853a <=( a1852a  and  a1849a );
 a1856a <=( A167  and  A170 );
 a1859a <=( A199  and  (not A166) );
 a1860a <=( a1859a  and  a1856a );
 a1863a <=( (not A201)  and  A200 );
 a1866a <=( A301  and  (not A202) );
 a1867a <=( a1866a  and  a1863a );
 a1870a <=( A167  and  A170 );
 a1873a <=( (not A199)  and  (not A166) );
 a1874a <=( a1873a  and  a1870a );
 a1877a <=( (not A202)  and  (not A200) );
 a1880a <=( A300  and  A299 );
 a1881a <=( a1880a  and  a1877a );
 a1884a <=( A167  and  A170 );
 a1887a <=( (not A199)  and  (not A166) );
 a1888a <=( a1887a  and  a1884a );
 a1891a <=( (not A202)  and  (not A200) );
 a1894a <=( A300  and  A298 );
 a1895a <=( a1894a  and  a1891a );
 a1898a <=( (not A167)  and  A170 );
 a1901a <=( (not A201)  and  A166 );
 a1902a <=( a1901a  and  a1898a );
 a1905a <=( (not A203)  and  (not A202) );
 a1908a <=( A300  and  A299 );
 a1909a <=( a1908a  and  a1905a );
 a1912a <=( (not A167)  and  A170 );
 a1915a <=( (not A201)  and  A166 );
 a1916a <=( a1915a  and  a1912a );
 a1919a <=( (not A203)  and  (not A202) );
 a1922a <=( A300  and  A298 );
 a1923a <=( a1922a  and  a1919a );
 a1926a <=( (not A167)  and  A170 );
 a1929a <=( A199  and  A166 );
 a1930a <=( a1929a  and  a1926a );
 a1933a <=( (not A201)  and  A200 );
 a1936a <=( A301  and  (not A202) );
 a1937a <=( a1936a  and  a1933a );
 a1940a <=( (not A167)  and  A170 );
 a1943a <=( (not A199)  and  A166 );
 a1944a <=( a1943a  and  a1940a );
 a1947a <=( (not A202)  and  (not A200) );
 a1950a <=( A300  and  A299 );
 a1951a <=( a1950a  and  a1947a );
 a1954a <=( (not A167)  and  A170 );
 a1957a <=( (not A199)  and  A166 );
 a1958a <=( a1957a  and  a1954a );
 a1961a <=( (not A202)  and  (not A200) );
 a1964a <=( A300  and  A298 );
 a1965a <=( a1964a  and  a1961a );
 a1968a <=( A199  and  A169 );
 a1971a <=( (not A201)  and  A200 );
 a1972a <=( a1971a  and  a1968a );
 a1975a <=( A298  and  (not A202) );
 a1978a <=( A302  and  (not A299) );
 a1979a <=( a1978a  and  a1975a );
 a1982a <=( A199  and  A169 );
 a1985a <=( (not A201)  and  A200 );
 a1986a <=( a1985a  and  a1982a );
 a1989a <=( (not A298)  and  (not A202) );
 a1992a <=( A302  and  A299 );
 a1993a <=( a1992a  and  a1989a );
 a1996a <=( (not A167)  and  (not A169) );
 a1999a <=( A199  and  (not A166) );
 a2000a <=( a1999a  and  a1996a );
 a2003a <=( A298  and  A201 );
 a2006a <=( A302  and  (not A299) );
 a2007a <=( a2006a  and  a2003a );
 a2010a <=( (not A167)  and  (not A169) );
 a2013a <=( A199  and  (not A166) );
 a2014a <=( a2013a  and  a2010a );
 a2017a <=( (not A298)  and  A201 );
 a2020a <=( A302  and  A299 );
 a2021a <=( a2020a  and  a2017a );
 a2024a <=( (not A167)  and  (not A169) );
 a2027a <=( A200  and  (not A166) );
 a2028a <=( a2027a  and  a2024a );
 a2031a <=( A298  and  A201 );
 a2034a <=( A302  and  (not A299) );
 a2035a <=( a2034a  and  a2031a );
 a2038a <=( (not A167)  and  (not A169) );
 a2041a <=( A200  and  (not A166) );
 a2042a <=( a2041a  and  a2038a );
 a2045a <=( (not A298)  and  A201 );
 a2048a <=( A302  and  A299 );
 a2049a <=( a2048a  and  a2045a );
 a2052a <=( (not A167)  and  (not A169) );
 a2055a <=( (not A199)  and  (not A166) );
 a2056a <=( a2055a  and  a2052a );
 a2059a <=( A203  and  A200 );
 a2062a <=( A300  and  A299 );
 a2063a <=( a2062a  and  a2059a );
 a2066a <=( (not A167)  and  (not A169) );
 a2069a <=( (not A199)  and  (not A166) );
 a2070a <=( a2069a  and  a2066a );
 a2073a <=( A203  and  A200 );
 a2076a <=( A300  and  A298 );
 a2077a <=( a2076a  and  a2073a );
 a2080a <=( (not A167)  and  (not A169) );
 a2083a <=( A199  and  (not A166) );
 a2084a <=( a2083a  and  a2080a );
 a2087a <=( A203  and  (not A200) );
 a2090a <=( A300  and  A299 );
 a2091a <=( a2090a  and  a2087a );
 a2094a <=( (not A167)  and  (not A169) );
 a2097a <=( A199  and  (not A166) );
 a2098a <=( a2097a  and  a2094a );
 a2101a <=( A203  and  (not A200) );
 a2104a <=( A300  and  A298 );
 a2105a <=( a2104a  and  a2101a );
 a2108a <=( (not A168)  and  (not A169) );
 a2111a <=( A166  and  A167 );
 a2112a <=( a2111a  and  a2108a );
 a2115a <=( A298  and  A202 );
 a2118a <=( A302  and  (not A299) );
 a2119a <=( a2118a  and  a2115a );
 a2122a <=( (not A168)  and  (not A169) );
 a2125a <=( A166  and  A167 );
 a2126a <=( a2125a  and  a2122a );
 a2129a <=( (not A298)  and  A202 );
 a2132a <=( A302  and  A299 );
 a2133a <=( a2132a  and  a2129a );
 a2136a <=( (not A168)  and  (not A169) );
 a2139a <=( A166  and  A167 );
 a2140a <=( a2139a  and  a2136a );
 a2143a <=( A201  and  A199 );
 a2146a <=( A300  and  A299 );
 a2147a <=( a2146a  and  a2143a );
 a2150a <=( (not A168)  and  (not A169) );
 a2153a <=( A166  and  A167 );
 a2154a <=( a2153a  and  a2150a );
 a2157a <=( A201  and  A199 );
 a2160a <=( A300  and  A298 );
 a2161a <=( a2160a  and  a2157a );
 a2164a <=( (not A168)  and  (not A169) );
 a2167a <=( A166  and  A167 );
 a2168a <=( a2167a  and  a2164a );
 a2171a <=( A201  and  A200 );
 a2174a <=( A300  and  A299 );
 a2175a <=( a2174a  and  a2171a );
 a2178a <=( (not A168)  and  (not A169) );
 a2181a <=( A166  and  A167 );
 a2182a <=( a2181a  and  a2178a );
 a2185a <=( A201  and  A200 );
 a2188a <=( A300  and  A298 );
 a2189a <=( a2188a  and  a2185a );
 a2192a <=( (not A168)  and  (not A169) );
 a2195a <=( A166  and  A167 );
 a2196a <=( a2195a  and  a2192a );
 a2199a <=( A200  and  (not A199) );
 a2202a <=( A301  and  A203 );
 a2203a <=( a2202a  and  a2199a );
 a2206a <=( (not A168)  and  (not A169) );
 a2209a <=( A166  and  A167 );
 a2210a <=( a2209a  and  a2206a );
 a2213a <=( (not A200)  and  A199 );
 a2216a <=( A301  and  A203 );
 a2217a <=( a2216a  and  a2213a );
 a2220a <=( (not A169)  and  (not A170) );
 a2223a <=( A199  and  (not A168) );
 a2224a <=( a2223a  and  a2220a );
 a2227a <=( A298  and  A201 );
 a2230a <=( A302  and  (not A299) );
 a2231a <=( a2230a  and  a2227a );
 a2234a <=( (not A169)  and  (not A170) );
 a2237a <=( A199  and  (not A168) );
 a2238a <=( a2237a  and  a2234a );
 a2241a <=( (not A298)  and  A201 );
 a2244a <=( A302  and  A299 );
 a2245a <=( a2244a  and  a2241a );
 a2248a <=( (not A169)  and  (not A170) );
 a2251a <=( A200  and  (not A168) );
 a2252a <=( a2251a  and  a2248a );
 a2255a <=( A298  and  A201 );
 a2258a <=( A302  and  (not A299) );
 a2259a <=( a2258a  and  a2255a );
 a2262a <=( (not A169)  and  (not A170) );
 a2265a <=( A200  and  (not A168) );
 a2266a <=( a2265a  and  a2262a );
 a2269a <=( (not A298)  and  A201 );
 a2272a <=( A302  and  A299 );
 a2273a <=( a2272a  and  a2269a );
 a2276a <=( (not A169)  and  (not A170) );
 a2279a <=( (not A199)  and  (not A168) );
 a2280a <=( a2279a  and  a2276a );
 a2283a <=( A203  and  A200 );
 a2286a <=( A300  and  A299 );
 a2287a <=( a2286a  and  a2283a );
 a2290a <=( (not A169)  and  (not A170) );
 a2293a <=( (not A199)  and  (not A168) );
 a2294a <=( a2293a  and  a2290a );
 a2297a <=( A203  and  A200 );
 a2300a <=( A300  and  A298 );
 a2301a <=( a2300a  and  a2297a );
 a2304a <=( (not A169)  and  (not A170) );
 a2307a <=( A199  and  (not A168) );
 a2308a <=( a2307a  and  a2304a );
 a2311a <=( A203  and  (not A200) );
 a2314a <=( A300  and  A299 );
 a2315a <=( a2314a  and  a2311a );
 a2318a <=( (not A169)  and  (not A170) );
 a2321a <=( A199  and  (not A168) );
 a2322a <=( a2321a  and  a2318a );
 a2325a <=( A203  and  (not A200) );
 a2328a <=( A300  and  A298 );
 a2329a <=( a2328a  and  a2325a );
 a2332a <=( A166  and  A168 );
 a2335a <=( A200  and  A199 );
 a2336a <=( a2335a  and  a2332a );
 a2339a <=( (not A202)  and  (not A201) );
 a2343a <=( A302  and  (not A299) );
 a2344a <=( A298  and  a2343a );
 a2345a <=( a2344a  and  a2339a );
 a2348a <=( A166  and  A168 );
 a2351a <=( A200  and  A199 );
 a2352a <=( a2351a  and  a2348a );
 a2355a <=( (not A202)  and  (not A201) );
 a2359a <=( A302  and  A299 );
 a2360a <=( (not A298)  and  a2359a );
 a2361a <=( a2360a  and  a2355a );
 a2364a <=( A167  and  A168 );
 a2367a <=( A200  and  A199 );
 a2368a <=( a2367a  and  a2364a );
 a2371a <=( (not A202)  and  (not A201) );
 a2375a <=( A302  and  (not A299) );
 a2376a <=( A298  and  a2375a );
 a2377a <=( a2376a  and  a2371a );
 a2380a <=( A167  and  A168 );
 a2383a <=( A200  and  A199 );
 a2384a <=( a2383a  and  a2380a );
 a2387a <=( (not A202)  and  (not A201) );
 a2391a <=( A302  and  A299 );
 a2392a <=( (not A298)  and  a2391a );
 a2393a <=( a2392a  and  a2387a );
 a2396a <=( A167  and  A170 );
 a2399a <=( (not A201)  and  (not A166) );
 a2400a <=( a2399a  and  a2396a );
 a2403a <=( (not A203)  and  (not A202) );
 a2407a <=( A302  and  (not A299) );
 a2408a <=( A298  and  a2407a );
 a2409a <=( a2408a  and  a2403a );
 a2412a <=( A167  and  A170 );
 a2415a <=( (not A201)  and  (not A166) );
 a2416a <=( a2415a  and  a2412a );
 a2419a <=( (not A203)  and  (not A202) );
 a2423a <=( A302  and  A299 );
 a2424a <=( (not A298)  and  a2423a );
 a2425a <=( a2424a  and  a2419a );
 a2428a <=( A167  and  A170 );
 a2431a <=( A199  and  (not A166) );
 a2432a <=( a2431a  and  a2428a );
 a2435a <=( (not A201)  and  A200 );
 a2439a <=( A300  and  A299 );
 a2440a <=( (not A202)  and  a2439a );
 a2441a <=( a2440a  and  a2435a );
 a2444a <=( A167  and  A170 );
 a2447a <=( A199  and  (not A166) );
 a2448a <=( a2447a  and  a2444a );
 a2451a <=( (not A201)  and  A200 );
 a2455a <=( A300  and  A298 );
 a2456a <=( (not A202)  and  a2455a );
 a2457a <=( a2456a  and  a2451a );
 a2460a <=( A167  and  A170 );
 a2463a <=( (not A199)  and  (not A166) );
 a2464a <=( a2463a  and  a2460a );
 a2467a <=( (not A202)  and  (not A200) );
 a2471a <=( A302  and  (not A299) );
 a2472a <=( A298  and  a2471a );
 a2473a <=( a2472a  and  a2467a );
 a2476a <=( A167  and  A170 );
 a2479a <=( (not A199)  and  (not A166) );
 a2480a <=( a2479a  and  a2476a );
 a2483a <=( (not A202)  and  (not A200) );
 a2487a <=( A302  and  A299 );
 a2488a <=( (not A298)  and  a2487a );
 a2489a <=( a2488a  and  a2483a );
 a2492a <=( (not A167)  and  A170 );
 a2495a <=( (not A201)  and  A166 );
 a2496a <=( a2495a  and  a2492a );
 a2499a <=( (not A203)  and  (not A202) );
 a2503a <=( A302  and  (not A299) );
 a2504a <=( A298  and  a2503a );
 a2505a <=( a2504a  and  a2499a );
 a2508a <=( (not A167)  and  A170 );
 a2511a <=( (not A201)  and  A166 );
 a2512a <=( a2511a  and  a2508a );
 a2515a <=( (not A203)  and  (not A202) );
 a2519a <=( A302  and  A299 );
 a2520a <=( (not A298)  and  a2519a );
 a2521a <=( a2520a  and  a2515a );
 a2524a <=( (not A167)  and  A170 );
 a2527a <=( A199  and  A166 );
 a2528a <=( a2527a  and  a2524a );
 a2531a <=( (not A201)  and  A200 );
 a2535a <=( A300  and  A299 );
 a2536a <=( (not A202)  and  a2535a );
 a2537a <=( a2536a  and  a2531a );
 a2540a <=( (not A167)  and  A170 );
 a2543a <=( A199  and  A166 );
 a2544a <=( a2543a  and  a2540a );
 a2547a <=( (not A201)  and  A200 );
 a2551a <=( A300  and  A298 );
 a2552a <=( (not A202)  and  a2551a );
 a2553a <=( a2552a  and  a2547a );
 a2556a <=( (not A167)  and  A170 );
 a2559a <=( (not A199)  and  A166 );
 a2560a <=( a2559a  and  a2556a );
 a2563a <=( (not A202)  and  (not A200) );
 a2567a <=( A302  and  (not A299) );
 a2568a <=( A298  and  a2567a );
 a2569a <=( a2568a  and  a2563a );
 a2572a <=( (not A167)  and  A170 );
 a2575a <=( (not A199)  and  A166 );
 a2576a <=( a2575a  and  a2572a );
 a2579a <=( (not A202)  and  (not A200) );
 a2583a <=( A302  and  A299 );
 a2584a <=( (not A298)  and  a2583a );
 a2585a <=( a2584a  and  a2579a );
 a2588a <=( (not A167)  and  (not A169) );
 a2591a <=( (not A199)  and  (not A166) );
 a2592a <=( a2591a  and  a2588a );
 a2595a <=( A203  and  A200 );
 a2599a <=( A302  and  (not A299) );
 a2600a <=( A298  and  a2599a );
 a2601a <=( a2600a  and  a2595a );
 a2604a <=( (not A167)  and  (not A169) );
 a2607a <=( (not A199)  and  (not A166) );
 a2608a <=( a2607a  and  a2604a );
 a2611a <=( A203  and  A200 );
 a2615a <=( A302  and  A299 );
 a2616a <=( (not A298)  and  a2615a );
 a2617a <=( a2616a  and  a2611a );
 a2620a <=( (not A167)  and  (not A169) );
 a2623a <=( A199  and  (not A166) );
 a2624a <=( a2623a  and  a2620a );
 a2627a <=( A203  and  (not A200) );
 a2631a <=( A302  and  (not A299) );
 a2632a <=( A298  and  a2631a );
 a2633a <=( a2632a  and  a2627a );
 a2636a <=( (not A167)  and  (not A169) );
 a2639a <=( A199  and  (not A166) );
 a2640a <=( a2639a  and  a2636a );
 a2643a <=( A203  and  (not A200) );
 a2647a <=( A302  and  A299 );
 a2648a <=( (not A298)  and  a2647a );
 a2649a <=( a2648a  and  a2643a );
 a2652a <=( (not A168)  and  (not A169) );
 a2655a <=( A166  and  A167 );
 a2656a <=( a2655a  and  a2652a );
 a2659a <=( A201  and  A199 );
 a2663a <=( A302  and  (not A299) );
 a2664a <=( A298  and  a2663a );
 a2665a <=( a2664a  and  a2659a );
 a2668a <=( (not A168)  and  (not A169) );
 a2671a <=( A166  and  A167 );
 a2672a <=( a2671a  and  a2668a );
 a2675a <=( A201  and  A199 );
 a2679a <=( A302  and  A299 );
 a2680a <=( (not A298)  and  a2679a );
 a2681a <=( a2680a  and  a2675a );
 a2684a <=( (not A168)  and  (not A169) );
 a2687a <=( A166  and  A167 );
 a2688a <=( a2687a  and  a2684a );
 a2691a <=( A201  and  A200 );
 a2695a <=( A302  and  (not A299) );
 a2696a <=( A298  and  a2695a );
 a2697a <=( a2696a  and  a2691a );
 a2700a <=( (not A168)  and  (not A169) );
 a2703a <=( A166  and  A167 );
 a2704a <=( a2703a  and  a2700a );
 a2707a <=( A201  and  A200 );
 a2711a <=( A302  and  A299 );
 a2712a <=( (not A298)  and  a2711a );
 a2713a <=( a2712a  and  a2707a );
 a2716a <=( (not A168)  and  (not A169) );
 a2719a <=( A166  and  A167 );
 a2720a <=( a2719a  and  a2716a );
 a2723a <=( A200  and  (not A199) );
 a2727a <=( A300  and  A299 );
 a2728a <=( A203  and  a2727a );
 a2729a <=( a2728a  and  a2723a );
 a2732a <=( (not A168)  and  (not A169) );
 a2735a <=( A166  and  A167 );
 a2736a <=( a2735a  and  a2732a );
 a2739a <=( A200  and  (not A199) );
 a2743a <=( A300  and  A298 );
 a2744a <=( A203  and  a2743a );
 a2745a <=( a2744a  and  a2739a );
 a2748a <=( (not A168)  and  (not A169) );
 a2751a <=( A166  and  A167 );
 a2752a <=( a2751a  and  a2748a );
 a2755a <=( (not A200)  and  A199 );
 a2759a <=( A300  and  A299 );
 a2760a <=( A203  and  a2759a );
 a2761a <=( a2760a  and  a2755a );
 a2764a <=( (not A168)  and  (not A169) );
 a2767a <=( A166  and  A167 );
 a2768a <=( a2767a  and  a2764a );
 a2771a <=( (not A200)  and  A199 );
 a2775a <=( A300  and  A298 );
 a2776a <=( A203  and  a2775a );
 a2777a <=( a2776a  and  a2771a );
 a2780a <=( (not A169)  and  (not A170) );
 a2783a <=( (not A199)  and  (not A168) );
 a2784a <=( a2783a  and  a2780a );
 a2787a <=( A203  and  A200 );
 a2791a <=( A302  and  (not A299) );
 a2792a <=( A298  and  a2791a );
 a2793a <=( a2792a  and  a2787a );
 a2796a <=( (not A169)  and  (not A170) );
 a2799a <=( (not A199)  and  (not A168) );
 a2800a <=( a2799a  and  a2796a );
 a2803a <=( A203  and  A200 );
 a2807a <=( A302  and  A299 );
 a2808a <=( (not A298)  and  a2807a );
 a2809a <=( a2808a  and  a2803a );
 a2812a <=( (not A169)  and  (not A170) );
 a2815a <=( A199  and  (not A168) );
 a2816a <=( a2815a  and  a2812a );
 a2819a <=( A203  and  (not A200) );
 a2823a <=( A302  and  (not A299) );
 a2824a <=( A298  and  a2823a );
 a2825a <=( a2824a  and  a2819a );
 a2828a <=( (not A169)  and  (not A170) );
 a2831a <=( A199  and  (not A168) );
 a2832a <=( a2831a  and  a2828a );
 a2835a <=( A203  and  (not A200) );
 a2839a <=( A302  and  A299 );
 a2840a <=( (not A298)  and  a2839a );
 a2841a <=( a2840a  and  a2835a );
 a2844a <=( A167  and  A170 );
 a2848a <=( A200  and  A199 );
 a2849a <=( (not A166)  and  a2848a );
 a2850a <=( a2849a  and  a2844a );
 a2853a <=( (not A202)  and  (not A201) );
 a2857a <=( A302  and  (not A299) );
 a2858a <=( A298  and  a2857a );
 a2859a <=( a2858a  and  a2853a );
 a2862a <=( A167  and  A170 );
 a2866a <=( A200  and  A199 );
 a2867a <=( (not A166)  and  a2866a );
 a2868a <=( a2867a  and  a2862a );
 a2871a <=( (not A202)  and  (not A201) );
 a2875a <=( A302  and  A299 );
 a2876a <=( (not A298)  and  a2875a );
 a2877a <=( a2876a  and  a2871a );
 a2880a <=( (not A167)  and  A170 );
 a2884a <=( A200  and  A199 );
 a2885a <=( A166  and  a2884a );
 a2886a <=( a2885a  and  a2880a );
 a2889a <=( (not A202)  and  (not A201) );
 a2893a <=( A302  and  (not A299) );
 a2894a <=( A298  and  a2893a );
 a2895a <=( a2894a  and  a2889a );
 a2898a <=( (not A167)  and  A170 );
 a2902a <=( A200  and  A199 );
 a2903a <=( A166  and  a2902a );
 a2904a <=( a2903a  and  a2898a );
 a2907a <=( (not A202)  and  (not A201) );
 a2911a <=( A302  and  A299 );
 a2912a <=( (not A298)  and  a2911a );
 a2913a <=( a2912a  and  a2907a );
 a2916a <=( (not A168)  and  (not A169) );
 a2920a <=( (not A199)  and  A166 );
 a2921a <=( A167  and  a2920a );
 a2922a <=( a2921a  and  a2916a );
 a2925a <=( A203  and  A200 );
 a2929a <=( A302  and  (not A299) );
 a2930a <=( A298  and  a2929a );
 a2931a <=( a2930a  and  a2925a );
 a2934a <=( (not A168)  and  (not A169) );
 a2938a <=( (not A199)  and  A166 );
 a2939a <=( A167  and  a2938a );
 a2940a <=( a2939a  and  a2934a );
 a2943a <=( A203  and  A200 );
 a2947a <=( A302  and  A299 );
 a2948a <=( (not A298)  and  a2947a );
 a2949a <=( a2948a  and  a2943a );
 a2952a <=( (not A168)  and  (not A169) );
 a2956a <=( A199  and  A166 );
 a2957a <=( A167  and  a2956a );
 a2958a <=( a2957a  and  a2952a );
 a2961a <=( A203  and  (not A200) );
 a2965a <=( A302  and  (not A299) );
 a2966a <=( A298  and  a2965a );
 a2967a <=( a2966a  and  a2961a );
 a2970a <=( (not A168)  and  (not A169) );
 a2974a <=( A199  and  A166 );
 a2975a <=( A167  and  a2974a );
 a2976a <=( a2975a  and  a2970a );
 a2979a <=( A203  and  (not A200) );
 a2983a <=( A302  and  A299 );
 a2984a <=( (not A298)  and  a2983a );
 a2985a <=( a2984a  and  a2979a );


end x25_13x_behav;
